module fake_jpeg_10870_n_590 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_590);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_590;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_0),
.B(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_62),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g152 ( 
.A(n_63),
.Y(n_152)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_64),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_32),
.A2(n_11),
.B1(n_1),
.B2(n_2),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_65),
.A2(n_89),
.B1(n_92),
.B2(n_41),
.Y(n_150)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx5_ASAP7_75t_SL g160 ( 
.A(n_66),
.Y(n_160)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_67),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_68),
.Y(n_178)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_55),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g163 ( 
.A(n_72),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_32),
.B(n_11),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_73),
.B(n_74),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_23),
.B(n_11),
.C(n_1),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_75),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_77),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_78),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g202 ( 
.A(n_79),
.Y(n_202)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_80),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_81),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_82),
.Y(n_198)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_83),
.Y(n_153)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_84),
.Y(n_183)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_85),
.Y(n_180)
);

BUFx16f_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx6_ASAP7_75t_SL g140 ( 
.A(n_86),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_87),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_31),
.Y(n_88)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_88),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_37),
.A2(n_18),
.B1(n_4),
.B2(n_5),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_21),
.B(n_12),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_90),
.B(n_125),
.Y(n_135)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_91),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_21),
.B(n_14),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_92),
.B(n_98),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_94),
.Y(n_199)
);

INVx6_ASAP7_75t_SL g95 ( 
.A(n_55),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_95),
.B(n_122),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_96),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_SL g98 ( 
.A1(n_55),
.A2(n_14),
.B(n_4),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_100),
.Y(n_162)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_102),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_103),
.Y(n_151)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_27),
.Y(n_104)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_104),
.Y(n_154)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_30),
.Y(n_105)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_30),
.Y(n_106)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_107),
.Y(n_185)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_33),
.Y(n_108)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_108),
.Y(n_190)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_33),
.Y(n_109)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_109),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_26),
.B(n_29),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_110),
.B(n_50),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_111),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_112),
.Y(n_197)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_37),
.Y(n_113)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_113),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_43),
.Y(n_114)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_114),
.Y(n_189)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_35),
.Y(n_115)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_115),
.Y(n_172)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_116),
.Y(n_204)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_117),
.Y(n_205)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_35),
.Y(n_118)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_118),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_37),
.Y(n_119)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_119),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_31),
.Y(n_120)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_120),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_31),
.Y(n_121)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_121),
.Y(n_192)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_44),
.Y(n_122)
);

BUFx12f_ASAP7_75t_SL g123 ( 
.A(n_59),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_123),
.B(n_124),
.Y(n_173)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_44),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_26),
.B(n_14),
.Y(n_125)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_59),
.Y(n_126)
);

BUFx4f_ASAP7_75t_L g203 ( 
.A(n_126),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_46),
.Y(n_127)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_127),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_62),
.A2(n_59),
.B1(n_49),
.B2(n_53),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_131),
.A2(n_133),
.B1(n_142),
.B2(n_147),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_76),
.A2(n_59),
.B1(n_49),
.B2(n_53),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_134),
.B(n_164),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_73),
.B(n_50),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_138),
.B(n_159),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_93),
.A2(n_59),
.B1(n_46),
.B2(n_49),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_78),
.A2(n_53),
.B1(n_49),
.B2(n_46),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_68),
.A2(n_57),
.B1(n_56),
.B2(n_45),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_148),
.A2(n_150),
.B1(n_184),
.B2(n_99),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_36),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_88),
.B(n_36),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_161),
.B(n_166),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_72),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_103),
.B(n_41),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_86),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_167),
.B(n_193),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_78),
.A2(n_46),
.B1(n_53),
.B2(n_56),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_168),
.A2(n_176),
.B1(n_179),
.B2(n_48),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_127),
.B(n_29),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_175),
.B(n_182),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_64),
.A2(n_52),
.B1(n_45),
.B2(n_57),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_117),
.A2(n_52),
.B1(n_28),
.B2(n_42),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_113),
.B(n_28),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_70),
.A2(n_34),
.B1(n_30),
.B2(n_42),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_120),
.B(n_34),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_77),
.A2(n_42),
.B1(n_51),
.B2(n_34),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_200),
.A2(n_206),
.B1(n_97),
.B2(n_96),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_81),
.A2(n_51),
.B1(n_34),
.B2(n_0),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_121),
.B(n_15),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_207),
.B(n_210),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_126),
.B(n_16),
.Y(n_210)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_212),
.Y(n_284)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_140),
.Y(n_213)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_213),
.Y(n_315)
);

INVx3_ASAP7_75t_SL g214 ( 
.A(n_160),
.Y(n_214)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_214),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_132),
.B(n_119),
.C(n_112),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_215),
.B(n_218),
.C(n_256),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_144),
.B(n_17),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_216),
.B(n_238),
.Y(n_319)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_178),
.Y(n_217)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_217),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_130),
.B(n_111),
.C(n_102),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_171),
.Y(n_220)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_220),
.Y(n_288)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_151),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_221),
.Y(n_295)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_183),
.Y(n_222)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_222),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_223),
.B(n_224),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_128),
.A2(n_94),
.B1(n_87),
.B2(n_82),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_226),
.A2(n_267),
.B(n_195),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_149),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_227),
.Y(n_287)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_190),
.Y(n_228)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_228),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_173),
.A2(n_51),
.B(n_54),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_229),
.B(n_277),
.Y(n_294)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_155),
.Y(n_230)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_230),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_135),
.A2(n_54),
.B1(n_48),
.B2(n_6),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_231),
.A2(n_233),
.B1(n_249),
.B2(n_269),
.Y(n_306)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_155),
.Y(n_232)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_232),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_206),
.A2(n_54),
.B1(n_48),
.B2(n_6),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_163),
.B(n_188),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_234),
.B(n_247),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

INVx11_ASAP7_75t_L g286 ( 
.A(n_235),
.Y(n_286)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_203),
.Y(n_236)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_236),
.Y(n_298)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_203),
.Y(n_237)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_237),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_160),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_239),
.Y(n_303)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_197),
.Y(n_242)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_242),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_156),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_243),
.B(n_248),
.Y(n_289)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_154),
.Y(n_244)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_244),
.Y(n_313)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_197),
.Y(n_245)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_245),
.Y(n_322)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_172),
.Y(n_246)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_246),
.Y(n_323)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_163),
.Y(n_247)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_162),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_131),
.A2(n_54),
.B1(n_48),
.B2(n_6),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_141),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_250),
.B(n_251),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_200),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_252),
.Y(n_308)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_146),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_253),
.B(n_257),
.Y(n_302)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_170),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_254),
.B(n_255),
.Y(n_334)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_186),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_137),
.B(n_4),
.C(n_7),
.Y(n_256)
);

CKINVDCx6p67_ASAP7_75t_R g257 ( 
.A(n_202),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_174),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_258),
.B(n_259),
.Y(n_310)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_165),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_192),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_260),
.B(n_261),
.Y(n_317)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_194),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_148),
.A2(n_17),
.B1(n_7),
.B2(n_15),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_262),
.A2(n_179),
.B1(n_181),
.B2(n_158),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_202),
.B(n_7),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_263),
.B(n_266),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_139),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_264),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_168),
.Y(n_265)
);

NAND3xp33_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_274),
.C(n_278),
.Y(n_292)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_136),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_145),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_133),
.A2(n_0),
.B1(n_16),
.B2(n_142),
.Y(n_269)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_170),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_271),
.B(n_273),
.Y(n_330)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_157),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_272),
.Y(n_300)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_153),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_187),
.B(n_0),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_143),
.A2(n_0),
.B1(n_191),
.B2(n_181),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_275),
.A2(n_199),
.B1(n_196),
.B2(n_169),
.Y(n_314)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_162),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_276),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_176),
.B(n_143),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_208),
.Y(n_278)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_185),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_279),
.Y(n_327)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_180),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_280),
.Y(n_333)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_158),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_282),
.Y(n_285)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_185),
.Y(n_282)
);

AND2x2_ASAP7_75t_SL g283 ( 
.A(n_215),
.B(n_189),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_283),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_147),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_291),
.B(n_324),
.C(n_328),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_293),
.A2(n_314),
.B1(n_331),
.B2(n_235),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_268),
.B(n_191),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_304),
.B(n_305),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_256),
.B(n_129),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_311),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_265),
.A2(n_129),
.B1(n_198),
.B2(n_169),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_320),
.A2(n_329),
.B1(n_332),
.B2(n_307),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_241),
.B(n_152),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_218),
.B(n_177),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_325),
.B(n_335),
.Y(n_349)
);

MAJx2_ASAP7_75t_L g328 ( 
.A(n_234),
.B(n_204),
.C(n_180),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_252),
.A2(n_177),
.B1(n_198),
.B2(n_209),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_219),
.A2(n_209),
.B1(n_199),
.B2(n_205),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_219),
.A2(n_195),
.B1(n_240),
.B2(n_255),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_221),
.B(n_247),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_338),
.A2(n_245),
.B1(n_272),
.B2(n_237),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g416 ( 
.A1(n_340),
.A2(n_363),
.B1(n_373),
.B2(n_376),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_308),
.A2(n_275),
.B1(n_212),
.B2(n_217),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_344),
.A2(n_345),
.B1(n_352),
.B2(n_375),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_308),
.A2(n_225),
.B1(n_214),
.B2(n_271),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_294),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_346),
.B(n_350),
.Y(n_406)
);

OA21x2_ASAP7_75t_L g347 ( 
.A1(n_293),
.A2(n_282),
.B(n_276),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_347),
.A2(n_356),
.B(n_334),
.Y(n_392)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_285),
.Y(n_348)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_348),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_318),
.B(n_211),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_319),
.B(n_304),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_351),
.B(n_369),
.Y(n_405)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_285),
.Y(n_353)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_353),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_305),
.B(n_279),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_354),
.B(n_357),
.Y(n_394)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_335),
.Y(n_355)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_355),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_294),
.A2(n_257),
.B(n_213),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_312),
.B(n_254),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_312),
.B(n_236),
.C(n_227),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_358),
.B(n_359),
.C(n_374),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_283),
.B(n_257),
.C(n_248),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_360),
.A2(n_368),
.B1(n_287),
.B2(n_309),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_283),
.B(n_325),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_361),
.B(n_366),
.Y(n_398)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_313),
.Y(n_362)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_362),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_L g363 ( 
.A1(n_338),
.A2(n_230),
.B1(n_232),
.B2(n_242),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_313),
.Y(n_364)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_364),
.Y(n_397)
);

INVx2_ASAP7_75t_SL g365 ( 
.A(n_326),
.Y(n_365)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_365),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_324),
.B(n_291),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_310),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_367),
.B(n_370),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_338),
.A2(n_331),
.B1(n_311),
.B2(n_314),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_332),
.B(n_316),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_333),
.B(n_290),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_323),
.Y(n_371)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_371),
.Y(n_402)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_323),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_372),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_307),
.A2(n_315),
.B1(n_300),
.B2(n_298),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_328),
.B(n_316),
.C(n_288),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_306),
.A2(n_329),
.B1(n_299),
.B2(n_320),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_315),
.A2(n_300),
.B1(n_301),
.B2(n_298),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_288),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_377),
.B(n_378),
.Y(n_413)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_290),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_289),
.B(n_333),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_379),
.B(n_380),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_296),
.B(n_327),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_316),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_381),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_342),
.A2(n_292),
.B(n_302),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_383),
.A2(n_389),
.B(n_407),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_368),
.A2(n_306),
.B1(n_330),
.B2(n_326),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_385),
.A2(n_386),
.B1(n_410),
.B2(n_396),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_349),
.A2(n_317),
.B1(n_296),
.B2(n_284),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_375),
.A2(n_321),
.B1(n_334),
.B2(n_327),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_388),
.A2(n_390),
.B1(n_414),
.B2(n_417),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_356),
.A2(n_321),
.B(n_334),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_347),
.A2(n_352),
.B1(n_369),
.B2(n_355),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_392),
.A2(n_408),
.B(n_359),
.Y(n_424)
);

OA21x2_ASAP7_75t_L g396 ( 
.A1(n_360),
.A2(n_301),
.B(n_297),
.Y(n_396)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_396),
.Y(n_439)
);

A2O1A1Ixp33_ASAP7_75t_L g404 ( 
.A1(n_361),
.A2(n_297),
.B(n_303),
.C(n_322),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_404),
.B(n_412),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_356),
.A2(n_303),
.B(n_286),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_341),
.A2(n_287),
.B(n_337),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_SL g409 ( 
.A(n_366),
.B(n_322),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_409),
.B(n_339),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_380),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_347),
.A2(n_284),
.B1(n_309),
.B2(n_337),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_339),
.B(n_286),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_415),
.B(n_379),
.C(n_345),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_347),
.A2(n_284),
.B1(n_336),
.B2(n_295),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_413),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_418),
.B(n_420),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_419),
.B(n_415),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_413),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_395),
.B(n_357),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_421),
.B(n_437),
.C(n_440),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_400),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_422),
.B(n_427),
.Y(n_458)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_393),
.Y(n_423)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_423),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_424),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_390),
.A2(n_349),
.B1(n_343),
.B2(n_341),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_426),
.A2(n_428),
.B1(n_434),
.B2(n_445),
.Y(n_460)
);

OA22x2_ASAP7_75t_L g427 ( 
.A1(n_382),
.A2(n_341),
.B1(n_353),
.B2(n_348),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_382),
.A2(n_343),
.B1(n_354),
.B2(n_358),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_393),
.Y(n_429)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_429),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_406),
.B(n_350),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_431),
.B(n_432),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_406),
.B(n_351),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_407),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_433),
.B(n_392),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_412),
.A2(n_374),
.B1(n_381),
.B2(n_367),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_400),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_435),
.B(n_447),
.Y(n_478)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_397),
.Y(n_436)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_436),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_394),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_438),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_395),
.B(n_378),
.C(n_377),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_397),
.Y(n_441)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_441),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_442),
.A2(n_446),
.B1(n_394),
.B2(n_398),
.Y(n_451)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_402),
.Y(n_444)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_444),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_388),
.A2(n_391),
.B1(n_384),
.B2(n_387),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_410),
.A2(n_385),
.B1(n_396),
.B2(n_386),
.Y(n_446)
);

INVxp33_ASAP7_75t_L g447 ( 
.A(n_405),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_405),
.A2(n_370),
.B1(n_344),
.B2(n_372),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_448),
.A2(n_403),
.B1(n_408),
.B2(n_399),
.Y(n_476)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_402),
.Y(n_449)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_449),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_442),
.A2(n_391),
.B1(n_387),
.B2(n_384),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_450),
.A2(n_451),
.B1(n_455),
.B2(n_467),
.Y(n_481)
);

OAI22xp33_ASAP7_75t_SL g452 ( 
.A1(n_446),
.A2(n_414),
.B1(n_417),
.B2(n_416),
.Y(n_452)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_452),
.Y(n_492)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_445),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_453),
.B(n_474),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_439),
.A2(n_416),
.B1(n_389),
.B2(n_398),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_457),
.B(n_473),
.Y(n_480)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_464),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_421),
.B(n_409),
.C(n_411),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_466),
.B(n_437),
.C(n_440),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_439),
.A2(n_396),
.B1(n_404),
.B2(n_411),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_422),
.B(n_401),
.Y(n_470)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_470),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_418),
.B(n_404),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_471),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_419),
.B(n_409),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_443),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_439),
.A2(n_403),
.B1(n_383),
.B2(n_399),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_475),
.A2(n_423),
.B1(n_441),
.B2(n_436),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_476),
.A2(n_424),
.B1(n_433),
.B2(n_420),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_482),
.B(n_470),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_483),
.A2(n_485),
.B1(n_487),
.B2(n_491),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_455),
.B(n_430),
.Y(n_484)
);

CKINVDCx14_ASAP7_75t_R g517 ( 
.A(n_484),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_453),
.A2(n_443),
.B1(n_430),
.B2(n_426),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_460),
.A2(n_425),
.B1(n_427),
.B2(n_428),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_459),
.B(n_434),
.C(n_427),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_488),
.B(n_499),
.C(n_501),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_457),
.B(n_448),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_489),
.B(n_502),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_463),
.B(n_371),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_490),
.B(n_493),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_460),
.A2(n_425),
.B1(n_427),
.B2(n_449),
.Y(n_491)
);

INVxp33_ASAP7_75t_L g494 ( 
.A(n_478),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_494),
.B(n_496),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_474),
.B(n_429),
.Y(n_495)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_495),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_451),
.A2(n_444),
.B1(n_365),
.B2(n_362),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_459),
.B(n_364),
.C(n_365),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_454),
.Y(n_500)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_500),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_473),
.B(n_336),
.C(n_295),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_466),
.B(n_462),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_471),
.B(n_456),
.Y(n_503)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_503),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_475),
.B(n_464),
.C(n_450),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_504),
.B(n_468),
.C(n_458),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_509),
.B(n_521),
.C(n_523),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_482),
.B(n_476),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_514),
.B(n_520),
.Y(n_542)
);

BUFx24_ASAP7_75t_SL g515 ( 
.A(n_497),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_515),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_484),
.A2(n_488),
.B(n_499),
.Y(n_516)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_516),
.Y(n_539)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_500),
.Y(n_518)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_518),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_480),
.B(n_458),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_519),
.B(n_522),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_489),
.B(n_502),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_485),
.B(n_467),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_SL g523 ( 
.A(n_480),
.B(n_456),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_495),
.Y(n_524)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_524),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_504),
.B(n_468),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_525),
.A2(n_483),
.B1(n_487),
.B2(n_498),
.Y(n_538)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_506),
.Y(n_526)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_526),
.Y(n_543)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_507),
.Y(n_527)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_527),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_508),
.A2(n_492),
.B1(n_481),
.B2(n_505),
.Y(n_528)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_528),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_508),
.A2(n_481),
.B1(n_479),
.B2(n_493),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_529),
.B(n_531),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_509),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_530),
.B(n_538),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_517),
.A2(n_484),
.B(n_486),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_521),
.B(n_486),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_532),
.B(n_519),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_522),
.A2(n_503),
.B(n_498),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_534),
.B(n_491),
.Y(n_545)
);

INVxp33_ASAP7_75t_L g535 ( 
.A(n_512),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_535),
.A2(n_513),
.B1(n_510),
.B2(n_501),
.Y(n_546)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_544),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_545),
.B(n_546),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_533),
.B(n_510),
.C(n_514),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_547),
.B(n_549),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_535),
.A2(n_511),
.B1(n_461),
.B2(n_465),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_536),
.B(n_523),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_SL g558 ( 
.A(n_551),
.B(n_556),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_534),
.A2(n_496),
.B1(n_461),
.B2(n_465),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_552),
.B(n_527),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_533),
.B(n_511),
.C(n_520),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_554),
.B(n_542),
.C(n_539),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_530),
.B(n_454),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_557),
.B(n_559),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_SL g559 ( 
.A1(n_547),
.A2(n_532),
.B(n_541),
.Y(n_559)
);

OAI21xp5_ASAP7_75t_L g560 ( 
.A1(n_553),
.A2(n_531),
.B(n_532),
.Y(n_560)
);

AOI21x1_ASAP7_75t_L g571 ( 
.A1(n_560),
.A2(n_544),
.B(n_545),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_562),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_553),
.B(n_542),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_SL g570 ( 
.A(n_564),
.B(n_565),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_555),
.B(n_540),
.Y(n_565)
);

INVx6_ASAP7_75t_L g567 ( 
.A(n_548),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_567),
.B(n_549),
.Y(n_575)
);

NOR2xp67_ASAP7_75t_L g568 ( 
.A(n_558),
.B(n_554),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_568),
.B(n_566),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_557),
.B(n_546),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g576 ( 
.A(n_569),
.B(n_571),
.Y(n_576)
);

A2O1A1Ixp33_ASAP7_75t_SL g573 ( 
.A1(n_560),
.A2(n_550),
.B(n_552),
.C(n_544),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_573),
.Y(n_578)
);

CKINVDCx16_ASAP7_75t_R g580 ( 
.A(n_575),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_SL g583 ( 
.A1(n_577),
.A2(n_561),
.B(n_563),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_570),
.B(n_574),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_579),
.B(n_581),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_SL g581 ( 
.A(n_572),
.B(n_561),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_583),
.B(n_584),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_576),
.B(n_573),
.C(n_526),
.Y(n_584)
);

AOI321xp33_ASAP7_75t_L g586 ( 
.A1(n_582),
.A2(n_577),
.A3(n_578),
.B1(n_580),
.B2(n_543),
.C(n_567),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_586),
.B(n_469),
.C(n_472),
.Y(n_587)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_587),
.B(n_585),
.Y(n_588)
);

OAI22xp33_ASAP7_75t_L g589 ( 
.A1(n_588),
.A2(n_469),
.B1(n_472),
.B2(n_477),
.Y(n_589)
);

AOI31xp33_ASAP7_75t_L g590 ( 
.A1(n_589),
.A2(n_477),
.A3(n_537),
.B(n_579),
.Y(n_590)
);


endmodule