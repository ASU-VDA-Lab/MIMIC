module real_aes_639_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_798, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_798;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_503;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_769;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_753;
wire n_314;
wire n_252;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_0), .B(n_119), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_1), .A2(n_128), .B(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_2), .B(n_765), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_3), .B(n_119), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_4), .B(n_135), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_5), .B(n_135), .Y(n_198) );
INVx1_ASAP7_75t_L g126 ( .A(n_6), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_7), .B(n_135), .Y(n_173) );
CKINVDCx16_ASAP7_75t_R g765 ( .A(n_8), .Y(n_765) );
NAND2xp33_ASAP7_75t_L g136 ( .A(n_9), .B(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g460 ( .A(n_10), .B(n_145), .Y(n_460) );
AND2x2_ASAP7_75t_L g520 ( .A(n_11), .B(n_114), .Y(n_520) );
INVx2_ASAP7_75t_L g116 ( .A(n_12), .Y(n_116) );
AOI221x1_ASAP7_75t_L g214 ( .A1(n_13), .A2(n_24), .B1(n_119), .B2(n_128), .C(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_14), .B(n_135), .Y(n_494) );
CKINVDCx16_ASAP7_75t_R g432 ( .A(n_15), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g118 ( .A(n_16), .B(n_119), .Y(n_118) );
AO21x2_ASAP7_75t_L g113 ( .A1(n_17), .A2(n_114), .B(n_117), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_18), .B(n_153), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_19), .B(n_135), .Y(n_162) );
AO21x1_ASAP7_75t_L g193 ( .A1(n_20), .A2(n_119), .B(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_21), .B(n_119), .Y(n_525) );
INVx1_ASAP7_75t_L g436 ( .A(n_22), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_23), .A2(n_89), .B1(n_119), .B2(n_465), .Y(n_464) );
NAND2x1_ASAP7_75t_L g184 ( .A(n_25), .B(n_135), .Y(n_184) );
NAND2x1_ASAP7_75t_L g172 ( .A(n_26), .B(n_137), .Y(n_172) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_27), .A2(n_86), .B(n_116), .Y(n_115) );
OR2x2_ASAP7_75t_L g140 ( .A(n_27), .B(n_86), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_28), .B(n_137), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_29), .B(n_135), .Y(n_134) );
AO21x2_ASAP7_75t_L g489 ( .A1(n_30), .A2(n_145), .B(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_31), .B(n_137), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_32), .A2(n_128), .B(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_33), .B(n_135), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_34), .A2(n_128), .B(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g125 ( .A(n_35), .B(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g129 ( .A(n_35), .B(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g473 ( .A(n_35), .Y(n_473) );
OR2x6_ASAP7_75t_L g434 ( .A(n_36), .B(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_37), .B(n_119), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_38), .B(n_119), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_39), .B(n_135), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_40), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_41), .B(n_137), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_42), .B(n_119), .Y(n_446) );
XNOR2xp5_ASAP7_75t_L g746 ( .A(n_43), .B(n_747), .Y(n_746) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_44), .A2(n_128), .B(n_456), .Y(n_455) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_45), .A2(n_103), .B1(n_758), .B2(n_769), .C1(n_786), .C2(n_790), .Y(n_102) );
OAI22xp5_ASAP7_75t_SL g774 ( .A1(n_45), .A2(n_775), .B1(n_776), .B2(n_777), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_45), .Y(n_775) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_46), .A2(n_128), .B(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_47), .B(n_137), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_48), .B(n_137), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_49), .B(n_119), .Y(n_491) );
INVx1_ASAP7_75t_L g122 ( .A(n_50), .Y(n_122) );
INVx1_ASAP7_75t_L g132 ( .A(n_50), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_51), .B(n_135), .Y(n_458) );
AND2x2_ASAP7_75t_L g480 ( .A(n_52), .B(n_153), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_53), .B(n_137), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_54), .B(n_135), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_55), .B(n_137), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_56), .A2(n_128), .B(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_57), .B(n_119), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_58), .B(n_119), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_59), .A2(n_128), .B(n_499), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_60), .A2(n_99), .B1(n_748), .B2(n_749), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_60), .Y(n_749) );
AO21x1_ASAP7_75t_L g195 ( .A1(n_61), .A2(n_128), .B(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g531 ( .A(n_62), .B(n_154), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_63), .B(n_119), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_64), .B(n_137), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_65), .B(n_119), .Y(n_174) );
AOI22xp5_ASAP7_75t_L g777 ( .A1(n_66), .A2(n_79), .B1(n_778), .B2(n_779), .Y(n_777) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_66), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_67), .B(n_137), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_68), .A2(n_93), .B1(n_128), .B2(n_471), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_69), .Y(n_755) );
AND2x2_ASAP7_75t_L g208 ( .A(n_70), .B(n_154), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_71), .B(n_135), .Y(n_528) );
INVx1_ASAP7_75t_L g124 ( .A(n_72), .Y(n_124) );
INVx1_ASAP7_75t_L g130 ( .A(n_72), .Y(n_130) );
AND2x2_ASAP7_75t_L g176 ( .A(n_73), .B(n_145), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_74), .B(n_137), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_75), .A2(n_128), .B(n_484), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g447 ( .A1(n_76), .A2(n_128), .B(n_448), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_77), .A2(n_128), .B(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g503 ( .A(n_78), .B(n_154), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_79), .Y(n_778) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_80), .B(n_153), .Y(n_462) );
INVx1_ASAP7_75t_L g437 ( .A(n_81), .Y(n_437) );
AND2x2_ASAP7_75t_L g144 ( .A(n_82), .B(n_145), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_83), .B(n_119), .Y(n_164) );
AND2x2_ASAP7_75t_L g451 ( .A(n_84), .B(n_114), .Y(n_451) );
AND2x2_ASAP7_75t_L g194 ( .A(n_85), .B(n_139), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_87), .B(n_137), .Y(n_163) );
AND2x2_ASAP7_75t_L g188 ( .A(n_88), .B(n_145), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_90), .B(n_135), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_91), .A2(n_128), .B(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_92), .B(n_137), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_94), .A2(n_128), .B(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_95), .B(n_135), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_96), .B(n_135), .Y(n_151) );
BUFx2_ASAP7_75t_L g530 ( .A(n_97), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_98), .Y(n_785) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_99), .Y(n_748) );
BUFx2_ASAP7_75t_L g766 ( .A(n_100), .Y(n_766) );
BUFx2_ASAP7_75t_SL g794 ( .A(n_100), .Y(n_794) );
AOI21xp5_ASAP7_75t_L g127 ( .A1(n_101), .A2(n_128), .B(n_133), .Y(n_127) );
OAI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_746), .B(n_750), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OAI22x1_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_429), .B1(n_438), .B2(n_742), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_107), .A2(n_439), .B1(n_752), .B2(n_753), .Y(n_751) );
AND2x4_ASAP7_75t_L g107 ( .A(n_108), .B(n_350), .Y(n_107) );
NOR3xp33_ASAP7_75t_SL g108 ( .A(n_109), .B(n_262), .C(n_302), .Y(n_108) );
OAI221xp5_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_177), .B1(n_226), .B2(n_241), .C(n_244), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_141), .Y(n_111) );
INVx2_ASAP7_75t_L g259 ( .A(n_112), .Y(n_259) );
AND2x2_ASAP7_75t_L g289 ( .A(n_112), .B(n_290), .Y(n_289) );
BUFx3_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_L g227 ( .A(n_113), .B(n_228), .Y(n_227) );
OR2x2_ASAP7_75t_L g234 ( .A(n_113), .B(n_167), .Y(n_234) );
INVx2_ASAP7_75t_L g240 ( .A(n_113), .Y(n_240) );
AND2x2_ASAP7_75t_L g249 ( .A(n_113), .B(n_143), .Y(n_249) );
INVx1_ASAP7_75t_L g265 ( .A(n_113), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_113), .B(n_311), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_114), .A2(n_525), .B(n_526), .Y(n_524) );
BUFx4f_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx3_ASAP7_75t_L g146 ( .A(n_115), .Y(n_146) );
AND2x4_ASAP7_75t_L g139 ( .A(n_116), .B(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_SL g154 ( .A(n_116), .B(n_140), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_127), .B(n_139), .Y(n_117) );
AND2x4_ASAP7_75t_L g119 ( .A(n_120), .B(n_125), .Y(n_119) );
AND2x4_ASAP7_75t_L g120 ( .A(n_121), .B(n_123), .Y(n_120) );
AND2x6_ASAP7_75t_L g137 ( .A(n_121), .B(n_130), .Y(n_137) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x4_ASAP7_75t_L g135 ( .A(n_123), .B(n_132), .Y(n_135) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx5_ASAP7_75t_L g138 ( .A(n_125), .Y(n_138) );
AND2x2_ASAP7_75t_L g131 ( .A(n_126), .B(n_132), .Y(n_131) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_126), .Y(n_468) );
AND2x6_ASAP7_75t_L g128 ( .A(n_129), .B(n_131), .Y(n_128) );
BUFx3_ASAP7_75t_L g469 ( .A(n_129), .Y(n_469) );
INVx2_ASAP7_75t_L g475 ( .A(n_130), .Y(n_475) );
AND2x4_ASAP7_75t_L g471 ( .A(n_131), .B(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g467 ( .A(n_132), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_136), .B(n_138), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_137), .B(n_530), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_138), .A2(n_151), .B(n_152), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_138), .A2(n_162), .B(n_163), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_138), .A2(n_172), .B(n_173), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_138), .A2(n_184), .B(n_185), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_138), .A2(n_197), .B(n_198), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_138), .A2(n_205), .B(n_206), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_138), .A2(n_216), .B(n_217), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_138), .A2(n_449), .B(n_450), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_138), .A2(n_457), .B(n_458), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_138), .A2(n_485), .B(n_486), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_138), .A2(n_494), .B(n_495), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_138), .A2(n_500), .B(n_501), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_138), .A2(n_517), .B(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_138), .A2(n_528), .B(n_529), .Y(n_527) );
INVx1_ASAP7_75t_SL g158 ( .A(n_139), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_139), .B(n_200), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_139), .A2(n_482), .B(n_483), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_139), .A2(n_491), .B(n_492), .Y(n_490) );
AND2x2_ASAP7_75t_SL g141 ( .A(n_142), .B(n_155), .Y(n_141) );
INVx4_ASAP7_75t_L g230 ( .A(n_142), .Y(n_230) );
AND2x2_ASAP7_75t_L g261 ( .A(n_142), .B(n_168), .Y(n_261) );
AND2x2_ASAP7_75t_L g337 ( .A(n_142), .B(n_311), .Y(n_337) );
NAND2x1p5_ASAP7_75t_L g379 ( .A(n_142), .B(n_167), .Y(n_379) );
INVx5_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_143), .B(n_167), .Y(n_266) );
AND2x2_ASAP7_75t_L g290 ( .A(n_143), .B(n_168), .Y(n_290) );
BUFx2_ASAP7_75t_L g306 ( .A(n_143), .Y(n_306) );
NOR2x1_ASAP7_75t_SL g409 ( .A(n_143), .B(n_311), .Y(n_409) );
OR2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_147), .Y(n_143) );
INVx3_ASAP7_75t_L g187 ( .A(n_145), .Y(n_187) );
INVx4_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AO21x2_ASAP7_75t_L g453 ( .A1(n_146), .A2(n_454), .B(n_460), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_149), .B(n_153), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_153), .Y(n_175) );
OA21x2_ASAP7_75t_L g213 ( .A1(n_153), .A2(n_214), .B(n_218), .Y(n_213) );
OA21x2_ASAP7_75t_L g276 ( .A1(n_153), .A2(n_214), .B(n_218), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_153), .A2(n_446), .B(n_447), .Y(n_445) );
AO21x2_ASAP7_75t_L g463 ( .A1(n_153), .A2(n_464), .B(n_470), .Y(n_463) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g286 ( .A(n_155), .Y(n_286) );
AOI221xp5_ASAP7_75t_L g352 ( .A1(n_155), .A2(n_353), .B1(n_355), .B2(n_357), .C(n_362), .Y(n_352) );
AND2x2_ASAP7_75t_L g372 ( .A(n_155), .B(n_265), .Y(n_372) );
AND2x4_ASAP7_75t_L g155 ( .A(n_156), .B(n_167), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g228 ( .A(n_157), .Y(n_228) );
INVx1_ASAP7_75t_L g281 ( .A(n_157), .Y(n_281) );
AO21x2_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B(n_165), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_158), .B(n_166), .Y(n_165) );
AO21x2_ASAP7_75t_L g311 ( .A1(n_158), .A2(n_159), .B(n_165), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_164), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_167), .B(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g250 ( .A(n_167), .B(n_238), .Y(n_250) );
INVx2_ASAP7_75t_L g292 ( .A(n_167), .Y(n_292) );
AND2x2_ASAP7_75t_L g425 ( .A(n_167), .B(n_240), .Y(n_425) );
INVx4_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_168), .Y(n_282) );
AO21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_175), .B(n_176), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_170), .B(n_174), .Y(n_169) );
AOI21x1_ASAP7_75t_L g513 ( .A1(n_175), .A2(n_514), .B(n_520), .Y(n_513) );
NOR3xp33_ASAP7_75t_L g177 ( .A(n_178), .B(n_209), .C(n_224), .Y(n_177) );
AND2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_189), .Y(n_178) );
INVx2_ASAP7_75t_L g339 ( .A(n_179), .Y(n_339) );
AND2x2_ASAP7_75t_L g384 ( .A(n_179), .B(n_261), .Y(n_384) );
BUFx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g329 ( .A(n_180), .Y(n_329) );
AND2x4_ASAP7_75t_SL g344 ( .A(n_180), .B(n_256), .Y(n_344) );
AO21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_187), .B(n_188), .Y(n_180) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_181), .A2(n_187), .B(n_188), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_182), .B(n_186), .Y(n_181) );
AO21x2_ASAP7_75t_L g201 ( .A1(n_187), .A2(n_202), .B(n_208), .Y(n_201) );
AO21x2_ASAP7_75t_L g221 ( .A1(n_187), .A2(n_202), .B(n_208), .Y(n_221) );
AO21x1_ASAP7_75t_SL g496 ( .A1(n_187), .A2(n_497), .B(n_503), .Y(n_496) );
AO21x2_ASAP7_75t_L g554 ( .A1(n_187), .A2(n_497), .B(n_503), .Y(n_554) );
INVx2_ASAP7_75t_L g298 ( .A(n_189), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_189), .B(n_328), .Y(n_354) );
AND2x4_ASAP7_75t_L g387 ( .A(n_189), .B(n_334), .Y(n_387) );
AND2x4_ASAP7_75t_L g189 ( .A(n_190), .B(n_201), .Y(n_189) );
AND2x2_ASAP7_75t_L g225 ( .A(n_190), .B(n_220), .Y(n_225) );
OR2x2_ASAP7_75t_L g255 ( .A(n_190), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_SL g324 ( .A(n_190), .B(n_276), .Y(n_324) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
BUFx2_ASAP7_75t_L g269 ( .A(n_191), .Y(n_269) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g243 ( .A(n_192), .Y(n_243) );
OAI21x1_ASAP7_75t_SL g192 ( .A1(n_193), .A2(n_195), .B(n_199), .Y(n_192) );
INVx1_ASAP7_75t_L g200 ( .A(n_194), .Y(n_200) );
INVx2_ASAP7_75t_L g256 ( .A(n_201), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_203), .B(n_207), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_209), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_211), .B(n_219), .Y(n_210) );
AND2x2_ASAP7_75t_L g224 ( .A(n_211), .B(n_225), .Y(n_224) );
OR2x2_ASAP7_75t_L g297 ( .A(n_211), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g382 ( .A(n_211), .Y(n_382) );
BUFx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x4_ASAP7_75t_L g242 ( .A(n_212), .B(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g361 ( .A(n_212), .B(n_221), .Y(n_361) );
AND2x2_ASAP7_75t_L g365 ( .A(n_212), .B(n_231), .Y(n_365) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g334 ( .A(n_213), .Y(n_334) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_213), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_219), .B(n_242), .Y(n_318) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_222), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_220), .B(n_243), .Y(n_428) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g232 ( .A(n_221), .B(n_223), .Y(n_232) );
AND2x2_ASAP7_75t_L g314 ( .A(n_221), .B(n_276), .Y(n_314) );
AND2x2_ASAP7_75t_L g333 ( .A(n_221), .B(n_222), .Y(n_333) );
BUFx2_ASAP7_75t_L g254 ( .A(n_222), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_222), .B(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
BUFx3_ASAP7_75t_L g231 ( .A(n_223), .Y(n_231) );
INVxp67_ASAP7_75t_L g274 ( .A(n_223), .Y(n_274) );
INVx1_ASAP7_75t_L g247 ( .A(n_225), .Y(n_247) );
AND2x2_ASAP7_75t_L g283 ( .A(n_225), .B(n_254), .Y(n_283) );
NAND2xp33_ASAP7_75t_L g364 ( .A(n_225), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g401 ( .A(n_225), .B(n_402), .Y(n_401) );
AOI221xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_229), .B1(n_232), .B2(n_233), .C(n_235), .Y(n_226) );
AND2x2_ASAP7_75t_L g330 ( .A(n_227), .B(n_230), .Y(n_330) );
AND2x2_ASAP7_75t_SL g349 ( .A(n_227), .B(n_290), .Y(n_349) );
AND2x2_ASAP7_75t_L g367 ( .A(n_227), .B(n_292), .Y(n_367) );
AND2x2_ASAP7_75t_L g422 ( .A(n_227), .B(n_261), .Y(n_422) );
INVx1_ASAP7_75t_L g238 ( .A(n_228), .Y(n_238) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_228), .Y(n_294) );
CKINVDCx16_ASAP7_75t_R g374 ( .A(n_229), .Y(n_374) );
AND2x4_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_230), .B(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_230), .B(n_281), .Y(n_356) );
AND2x2_ASAP7_75t_L g323 ( .A(n_231), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_SL g359 ( .A(n_231), .Y(n_359) );
AND2x2_ASAP7_75t_L g268 ( .A(n_232), .B(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_232), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g410 ( .A(n_232), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_232), .B(n_334), .Y(n_420) );
AND2x4_ASAP7_75t_L g336 ( .A(n_233), .B(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
OR2x2_ASAP7_75t_L g407 ( .A(n_234), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
OR2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_239), .Y(n_236) );
OR2x2_ASAP7_75t_L g278 ( .A(n_239), .B(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g285 ( .A(n_240), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g316 ( .A(n_240), .B(n_290), .Y(n_316) );
AND2x2_ASAP7_75t_L g390 ( .A(n_240), .B(n_311), .Y(n_390) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g338 ( .A(n_242), .B(n_339), .Y(n_338) );
OAI32xp33_ASAP7_75t_L g403 ( .A1(n_242), .A2(n_404), .A3(n_406), .B1(n_407), .B2(n_410), .Y(n_403) );
AND2x4_ASAP7_75t_L g275 ( .A(n_243), .B(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g373 ( .A(n_243), .B(n_276), .Y(n_373) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_248), .B1(n_251), .B2(n_257), .Y(n_244) );
INVxp67_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_SL g362 ( .A1(n_246), .A2(n_260), .B(n_363), .C(n_364), .Y(n_362) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g346 ( .A(n_247), .B(n_274), .Y(n_346) );
INVx1_ASAP7_75t_SL g417 ( .A(n_248), .Y(n_417) );
AND2x4_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
AND2x4_ASAP7_75t_L g320 ( .A(n_250), .B(n_259), .Y(n_320) );
AOI221xp5_ASAP7_75t_L g398 ( .A1(n_250), .A2(n_399), .B1(n_400), .B2(n_401), .C(n_403), .Y(n_398) );
INVx1_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_255), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_255), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OAI22xp33_ASAP7_75t_L g340 ( .A1(n_258), .A2(n_288), .B1(n_341), .B2(n_342), .Y(n_340) );
OR2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
OAI211xp5_ASAP7_75t_SL g376 ( .A1(n_259), .A2(n_377), .B(n_385), .C(n_398), .Y(n_376) );
INVx2_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g296 ( .A(n_261), .B(n_265), .Y(n_296) );
OAI211xp5_ASAP7_75t_SL g262 ( .A1(n_263), .A2(n_267), .B(n_270), .C(n_299), .Y(n_262) );
OR2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g293 ( .A(n_265), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g413 ( .A(n_265), .B(n_409), .Y(n_413) );
OAI32xp33_ASAP7_75t_L g370 ( .A1(n_266), .A2(n_371), .A3(n_373), .B1(n_374), .B2(n_375), .Y(n_370) );
INVx1_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_SL g360 ( .A(n_269), .B(n_361), .Y(n_360) );
AOI221xp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_277), .B1(n_283), .B2(n_284), .C(n_287), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_273), .B(n_275), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g427 ( .A(n_274), .B(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_SL g341 ( .A(n_275), .B(n_339), .Y(n_341) );
A2O1A1O1Ixp25_ASAP7_75t_L g412 ( .A1(n_275), .A2(n_344), .B(n_360), .C(n_406), .D(n_413), .Y(n_412) );
AOI31xp33_ASAP7_75t_L g414 ( .A1(n_275), .A2(n_296), .A3(n_406), .B(n_413), .Y(n_414) );
AND2x2_ASAP7_75t_L g328 ( .A(n_276), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_278), .B(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
INVx2_ASAP7_75t_L g405 ( .A(n_280), .Y(n_405) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g400 ( .A(n_281), .B(n_292), .Y(n_400) );
INVx1_ASAP7_75t_L g315 ( .A(n_283), .Y(n_315) );
AND2x2_ASAP7_75t_L g300 ( .A(n_284), .B(n_301), .Y(n_300) );
INVx2_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
AOI31xp33_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_291), .A3(n_295), .B(n_297), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_290), .B(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g423 ( .A(n_290), .B(n_369), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
AND2x2_ASAP7_75t_L g368 ( .A(n_292), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g394 ( .A(n_292), .Y(n_394) );
INVxp67_ASAP7_75t_L g363 ( .A(n_293), .Y(n_363) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g301 ( .A(n_297), .Y(n_301) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND3xp33_ASAP7_75t_SL g302 ( .A(n_303), .B(n_319), .C(n_335), .Y(n_302) );
AOI22xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_312), .B1(n_316), .B2(n_317), .Y(n_303) );
INVxp67_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx2_ASAP7_75t_L g389 ( .A(n_306), .Y(n_389) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVxp67_ASAP7_75t_SL g369 ( .A(n_310), .Y(n_369) );
INVxp67_ASAP7_75t_SL g395 ( .A(n_310), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_310), .B(n_379), .Y(n_396) );
NAND2xp33_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
INVx1_ASAP7_75t_L g347 ( .A(n_314), .Y(n_347) );
INVx1_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_321), .B1(n_330), .B2(n_331), .Y(n_319) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_322), .B(n_325), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
AOI221xp5_ASAP7_75t_L g366 ( .A1(n_328), .A2(n_333), .B1(n_367), .B2(n_368), .C(n_370), .Y(n_366) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2x1_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx1_ASAP7_75t_L g406 ( .A(n_333), .Y(n_406) );
AND2x2_ASAP7_75t_L g343 ( .A(n_334), .B(n_344), .Y(n_343) );
O2A1O1Ixp33_ASAP7_75t_SL g391 ( .A1(n_334), .A2(n_392), .B(n_396), .C(n_397), .Y(n_391) );
AOI211xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_338), .B(n_340), .C(n_345), .Y(n_335) );
AND2x2_ASAP7_75t_L g386 ( .A(n_339), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g397 ( .A(n_344), .Y(n_397) );
AOI21xp33_ASAP7_75t_SL g345 ( .A1(n_346), .A2(n_347), .B(n_348), .Y(n_345) );
INVx2_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
NOR3xp33_ASAP7_75t_L g350 ( .A(n_351), .B(n_376), .C(n_411), .Y(n_350) );
NAND2xp5_ASAP7_75t_SL g351 ( .A(n_352), .B(n_366), .Y(n_351) );
INVx1_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
INVxp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx1_ASAP7_75t_L g375 ( .A(n_360), .Y(n_375) );
INVxp67_ASAP7_75t_L g399 ( .A(n_364), .Y(n_399) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_SL g383 ( .A(n_373), .Y(n_383) );
AOI22xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_380), .B1(n_383), .B2(n_384), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AOI21xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_388), .B(n_391), .Y(n_385) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g424 ( .A(n_409), .B(n_425), .Y(n_424) );
OAI221xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_414), .B1(n_415), .B2(n_418), .C(n_421), .Y(n_411) );
INVxp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OAI31xp33_ASAP7_75t_SL g421 ( .A1(n_422), .A2(n_423), .A3(n_424), .B(n_426), .Y(n_421) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx4f_ASAP7_75t_SL g752 ( .A(n_429), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_430), .Y(n_429) );
CKINVDCx11_ASAP7_75t_R g430 ( .A(n_431), .Y(n_430) );
OR2x6_ASAP7_75t_SL g431 ( .A(n_432), .B(n_433), .Y(n_431) );
AND2x6_ASAP7_75t_SL g745 ( .A(n_432), .B(n_434), .Y(n_745) );
OR2x2_ASAP7_75t_L g757 ( .A(n_432), .B(n_434), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_432), .B(n_433), .Y(n_768) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
INVx3_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
XNOR2xp5_ASAP7_75t_L g773 ( .A(n_439), .B(n_774), .Y(n_773) );
AND2x4_ASAP7_75t_SL g439 ( .A(n_440), .B(n_638), .Y(n_439) );
NOR3xp33_ASAP7_75t_SL g440 ( .A(n_441), .B(n_547), .C(n_579), .Y(n_440) );
OAI221xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_476), .B1(n_504), .B2(n_521), .C(n_532), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_452), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g510 ( .A(n_444), .B(n_453), .Y(n_510) );
INVx4_ASAP7_75t_L g538 ( .A(n_444), .Y(n_538) );
AND2x4_ASAP7_75t_SL g578 ( .A(n_444), .B(n_512), .Y(n_578) );
BUFx2_ASAP7_75t_L g588 ( .A(n_444), .Y(n_588) );
NOR2x1_ASAP7_75t_L g654 ( .A(n_444), .B(n_593), .Y(n_654) );
AND2x2_ASAP7_75t_L g663 ( .A(n_444), .B(n_591), .Y(n_663) );
OR2x2_ASAP7_75t_L g671 ( .A(n_444), .B(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g697 ( .A(n_444), .B(n_536), .Y(n_697) );
AND2x4_ASAP7_75t_L g716 ( .A(n_444), .B(n_717), .Y(n_716) );
OR2x6_ASAP7_75t_L g444 ( .A(n_445), .B(n_451), .Y(n_444) );
INVx2_ASAP7_75t_SL g629 ( .A(n_452), .Y(n_629) );
OR2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_461), .Y(n_452) );
AND2x2_ASAP7_75t_L g536 ( .A(n_453), .B(n_513), .Y(n_536) );
INVx2_ASAP7_75t_L g563 ( .A(n_453), .Y(n_563) );
INVx2_ASAP7_75t_L g593 ( .A(n_453), .Y(n_593) );
AND2x2_ASAP7_75t_L g607 ( .A(n_453), .B(n_512), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_459), .Y(n_454) );
AND2x2_ASAP7_75t_L g537 ( .A(n_461), .B(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g560 ( .A(n_461), .Y(n_560) );
BUFx3_ASAP7_75t_L g574 ( .A(n_461), .Y(n_574) );
AND2x2_ASAP7_75t_L g603 ( .A(n_461), .B(n_604), .Y(n_603) );
AND2x4_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
AND2x4_ASAP7_75t_L g508 ( .A(n_462), .B(n_463), .Y(n_508) );
AND2x4_ASAP7_75t_L g465 ( .A(n_466), .B(n_469), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
NOR2x1p5_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
INVx3_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g609 ( .A(n_476), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_487), .Y(n_476) );
OR2x2_ASAP7_75t_L g720 ( .A(n_477), .B(n_521), .Y(n_720) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g576 ( .A(n_478), .B(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_478), .B(n_487), .Y(n_637) );
OR2x2_ASAP7_75t_L g735 ( .A(n_478), .B(n_657), .Y(n_735) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g546 ( .A(n_479), .B(n_522), .Y(n_546) );
OR2x2_ASAP7_75t_SL g556 ( .A(n_479), .B(n_557), .Y(n_556) );
INVx4_ASAP7_75t_L g567 ( .A(n_479), .Y(n_567) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_479), .Y(n_618) );
NAND2x1_ASAP7_75t_L g624 ( .A(n_479), .B(n_523), .Y(n_624) );
AND2x2_ASAP7_75t_L g649 ( .A(n_479), .B(n_489), .Y(n_649) );
OR2x2_ASAP7_75t_L g670 ( .A(n_479), .B(n_553), .Y(n_670) );
OR2x6_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
INVx1_ASAP7_75t_L g565 ( .A(n_487), .Y(n_565) );
O2A1O1Ixp33_ASAP7_75t_L g658 ( .A1(n_487), .A2(n_659), .B(n_662), .C(n_664), .Y(n_658) );
AND2x2_ASAP7_75t_L g731 ( .A(n_487), .B(n_507), .Y(n_731) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_496), .Y(n_487) );
INVx1_ASAP7_75t_L g598 ( .A(n_488), .Y(n_598) );
AND2x2_ASAP7_75t_L g668 ( .A(n_488), .B(n_523), .Y(n_668) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g542 ( .A(n_489), .Y(n_542) );
OR2x2_ASAP7_75t_L g557 ( .A(n_489), .B(n_523), .Y(n_557) );
INVx1_ASAP7_75t_L g573 ( .A(n_489), .Y(n_573) );
AND2x2_ASAP7_75t_L g585 ( .A(n_489), .B(n_496), .Y(n_585) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_489), .Y(n_691) );
NOR2x1_ASAP7_75t_SL g522 ( .A(n_496), .B(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_502), .Y(n_497) );
INVxp67_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_509), .Y(n_505) );
OR2x2_ASAP7_75t_L g655 ( .A(n_506), .B(n_590), .Y(n_655) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_507), .B(n_673), .Y(n_672) );
OR2x2_ASAP7_75t_L g737 ( .A(n_507), .B(n_634), .Y(n_737) );
INVx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g582 ( .A(n_508), .B(n_563), .Y(n_582) );
AND2x2_ASAP7_75t_L g678 ( .A(n_508), .B(n_591), .Y(n_678) );
INVx1_ASAP7_75t_L g595 ( .A(n_509), .Y(n_595) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
INVx1_ASAP7_75t_L g645 ( .A(n_510), .Y(n_645) );
INVx2_ASAP7_75t_L g612 ( .A(n_511), .Y(n_612) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g562 ( .A(n_512), .B(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g592 ( .A(n_512), .Y(n_592) );
INVx1_ASAP7_75t_L g717 ( .A(n_512), .Y(n_717) );
INVx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_513), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_519), .Y(n_514) );
OR2x2_ASAP7_75t_L g688 ( .A(n_521), .B(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_SL g543 ( .A(n_523), .Y(n_543) );
OR2x2_ASAP7_75t_L g566 ( .A(n_523), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g577 ( .A(n_523), .B(n_553), .Y(n_577) );
AND2x2_ASAP7_75t_L g651 ( .A(n_523), .B(n_567), .Y(n_651) );
BUFx2_ASAP7_75t_L g734 ( .A(n_523), .Y(n_734) );
OR2x6_ASAP7_75t_L g523 ( .A(n_524), .B(n_531), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_539), .B(n_544), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_537), .Y(n_534) );
AND2x2_ASAP7_75t_L g686 ( .A(n_535), .B(n_608), .Y(n_686) );
BUFx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g545 ( .A(n_536), .B(n_538), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_537), .B(n_607), .Y(n_708) );
INVx1_ASAP7_75t_L g738 ( .A(n_537), .Y(n_738) );
NAND2x1p5_ASAP7_75t_L g634 ( .A(n_538), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_538), .B(n_674), .Y(n_711) );
INVxp67_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
AND2x4_ASAP7_75t_SL g575 ( .A(n_541), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_541), .B(n_569), .Y(n_722) );
INVx3_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_542), .B(n_624), .Y(n_680) );
AND2x2_ASAP7_75t_L g698 ( .A(n_542), .B(n_651), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_543), .B(n_585), .Y(n_601) );
A2O1A1Ixp33_ASAP7_75t_L g630 ( .A1(n_543), .A2(n_589), .B(n_631), .C(n_636), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_543), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
AOI221xp5_ASAP7_75t_L g725 ( .A1(n_545), .A2(n_618), .B1(n_726), .B2(n_732), .C(n_736), .Y(n_725) );
INVx1_ASAP7_75t_SL g713 ( .A(n_546), .Y(n_713) );
OAI221xp5_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_558), .B1(n_564), .B2(n_568), .C(n_798), .Y(n_547) );
INVx2_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
AND2x4_ASAP7_75t_L g549 ( .A(n_550), .B(n_555), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g623 ( .A(n_552), .Y(n_623) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g597 ( .A(n_553), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g628 ( .A(n_553), .B(n_573), .Y(n_628) );
INVx2_ASAP7_75t_L g661 ( .A(n_553), .Y(n_661) );
INVx3_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OAI32xp33_ASAP7_75t_L g712 ( .A1(n_556), .A2(n_603), .A3(n_634), .B1(n_713), .B2(n_714), .Y(n_712) );
OR2x2_ASAP7_75t_L g683 ( .A(n_557), .B(n_670), .Y(n_683) );
INVx1_ASAP7_75t_L g693 ( .A(n_558), .Y(n_693) );
OR2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
INVx2_ASAP7_75t_L g608 ( .A(n_559), .Y(n_608) );
AND2x2_ASAP7_75t_L g679 ( .A(n_559), .B(n_654), .Y(n_679) );
OR2x2_ASAP7_75t_L g710 ( .A(n_559), .B(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_560), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g604 ( .A(n_563), .Y(n_604) );
OR2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
INVx2_ASAP7_75t_SL g569 ( .A(n_566), .Y(n_569) );
OR2x2_ASAP7_75t_L g656 ( .A(n_566), .B(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_567), .B(n_585), .Y(n_584) );
NOR2xp67_ASAP7_75t_L g690 ( .A(n_567), .B(n_691), .Y(n_690) );
BUFx2_ASAP7_75t_L g703 ( .A(n_567), .Y(n_703) );
A2O1A1Ixp33_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_570), .B(n_575), .C(n_578), .Y(n_568) );
AND2x2_ASAP7_75t_L g718 ( .A(n_570), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
BUFx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g644 ( .A(n_574), .B(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_574), .B(n_578), .Y(n_665) );
AND2x2_ASAP7_75t_L g696 ( .A(n_574), .B(n_697), .Y(n_696) );
O2A1O1Ixp33_ASAP7_75t_L g706 ( .A1(n_576), .A2(n_707), .B(n_709), .C(n_712), .Y(n_706) );
AOI222xp33_ASAP7_75t_L g580 ( .A1(n_577), .A2(n_581), .B1(n_583), .B2(n_586), .C1(n_594), .C2(n_596), .Y(n_580) );
AND2x2_ASAP7_75t_L g648 ( .A(n_577), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g581 ( .A(n_578), .B(n_582), .Y(n_581) );
INVx2_ASAP7_75t_SL g602 ( .A(n_578), .Y(n_602) );
NAND4xp25_ASAP7_75t_L g579 ( .A(n_580), .B(n_599), .C(n_620), .D(n_630), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_582), .B(n_588), .Y(n_642) );
INVx1_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g650 ( .A(n_585), .B(n_651), .Y(n_650) );
INVx2_ASAP7_75t_SL g657 ( .A(n_585), .Y(n_657) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
A2O1A1Ixp33_ASAP7_75t_L g620 ( .A1(n_587), .A2(n_621), .B(n_625), .C(n_629), .Y(n_620) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_588), .B(n_603), .Y(n_724) );
OR2x2_ASAP7_75t_L g728 ( .A(n_588), .B(n_614), .Y(n_728) );
INVx1_ASAP7_75t_L g701 ( .A(n_589), .Y(n_701) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVx1_ASAP7_75t_SL g635 ( .A(n_592), .Y(n_635) );
INVx1_ASAP7_75t_L g615 ( .A(n_593), .Y(n_615) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_595), .B(n_632), .Y(n_631) );
BUFx2_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g619 ( .A(n_597), .Y(n_619) );
AOI322xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_602), .A3(n_603), .B1(n_605), .B2(n_609), .C1(n_610), .C2(n_616), .Y(n_599) );
INVxp67_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
O2A1O1Ixp33_ASAP7_75t_SL g681 ( .A1(n_602), .A2(n_682), .B(n_683), .C(n_684), .Y(n_681) );
INVx1_ASAP7_75t_L g704 ( .A(n_603), .Y(n_704) );
NOR2xp67_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g662 ( .A(n_608), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_614), .Y(n_684) );
INVx2_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
INVx3_ASAP7_75t_L g627 ( .A(n_624), .Y(n_627) );
OR2x2_ASAP7_75t_L g695 ( .A(n_624), .B(n_657), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_624), .B(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
INVx1_ASAP7_75t_SL g727 ( .A(n_628), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_629), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND3xp33_ASAP7_75t_SL g732 ( .A(n_637), .B(n_733), .C(n_735), .Y(n_732) );
NOR3xp33_ASAP7_75t_SL g638 ( .A(n_639), .B(n_676), .C(n_705), .Y(n_638) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_640), .B(n_658), .Y(n_639) );
O2A1O1Ixp33_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_643), .B(n_646), .C(n_652), .Y(n_640) );
OAI31xp33_ASAP7_75t_L g685 ( .A1(n_641), .A2(n_663), .A3(n_686), .B(n_687), .Y(n_685) );
INVx1_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .Y(n_647) );
INVx2_ASAP7_75t_L g700 ( .A(n_648), .Y(n_700) );
INVx1_ASAP7_75t_L g675 ( .A(n_650), .Y(n_675) );
AOI21xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_655), .B(n_656), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OR2x2_ASAP7_75t_L g702 ( .A(n_660), .B(n_703), .Y(n_702) );
INVxp67_ASAP7_75t_L g741 ( .A(n_661), .Y(n_741) );
OAI22xp33_ASAP7_75t_SL g664 ( .A1(n_665), .A2(n_666), .B1(n_671), .B2(n_675), .Y(n_664) );
INVx3_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AND2x4_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_670), .Y(n_682) );
OR2x2_ASAP7_75t_L g733 ( .A(n_670), .B(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
NAND3xp33_ASAP7_75t_SL g676 ( .A(n_677), .B(n_685), .C(n_692), .Y(n_676) );
O2A1O1Ixp33_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B(n_680), .C(n_681), .Y(n_677) );
INVx2_ASAP7_75t_L g714 ( .A(n_678), .Y(n_714) );
INVx1_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AOI221xp5_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_694), .B1(n_696), .B2(n_698), .C(n_699), .Y(n_692) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OAI22xp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_701), .B1(n_702), .B2(n_704), .Y(n_699) );
NAND3xp33_ASAP7_75t_SL g705 ( .A(n_706), .B(n_715), .C(n_725), .Y(n_705) );
INVxp33_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_718), .B1(n_721), .B2(n_723), .Y(n_715) );
INVx2_ASAP7_75t_L g729 ( .A(n_716), .Y(n_729) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_728), .B1(n_729), .B2(n_730), .Y(n_726) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
OAI22xp33_ASAP7_75t_SL g736 ( .A1(n_735), .A2(n_737), .B1(n_738), .B2(n_739), .Y(n_736) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
CKINVDCx6p67_ASAP7_75t_R g742 ( .A(n_743), .Y(n_742) );
INVx4_ASAP7_75t_SL g753 ( .A(n_743), .Y(n_753) );
INVx3_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
CKINVDCx5p33_ASAP7_75t_R g744 ( .A(n_745), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g750 ( .A1(n_746), .A2(n_751), .B(n_754), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
BUFx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_761), .B(n_767), .Y(n_760) );
INVxp67_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
NAND2xp5_ASAP7_75t_SL g762 ( .A(n_763), .B(n_766), .Y(n_762) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
OR2x2_ASAP7_75t_SL g789 ( .A(n_764), .B(n_766), .Y(n_789) );
AOI21xp5_ASAP7_75t_L g791 ( .A1(n_764), .A2(n_792), .B(n_795), .Y(n_791) );
INVx1_ASAP7_75t_SL g772 ( .A(n_767), .Y(n_772) );
BUFx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
BUFx3_ASAP7_75t_L g784 ( .A(n_768), .Y(n_784) );
BUFx2_ASAP7_75t_L g796 ( .A(n_768), .Y(n_796) );
INVxp67_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
AOI21xp33_ASAP7_75t_SL g770 ( .A1(n_771), .A2(n_773), .B(n_780), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
CKINVDCx16_ASAP7_75t_R g776 ( .A(n_777), .Y(n_776) );
NOR2xp33_ASAP7_75t_SL g780 ( .A(n_781), .B(n_785), .Y(n_780) );
INVx1_ASAP7_75t_SL g781 ( .A(n_782), .Y(n_781) );
BUFx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_784), .Y(n_783) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_SL g790 ( .A(n_791), .Y(n_790) );
CKINVDCx11_ASAP7_75t_R g792 ( .A(n_793), .Y(n_792) );
CKINVDCx8_ASAP7_75t_R g793 ( .A(n_794), .Y(n_793) );
INVx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
endmodule