module fake_jpeg_26124_n_299 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_299);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_299;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_265;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

HAxp5_ASAP7_75t_SL g42 ( 
.A(n_39),
.B(n_24),
.CON(n_42),
.SN(n_42)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_42),
.B(n_34),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_38),
.A2(n_21),
.B1(n_25),
.B2(n_32),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_25),
.B1(n_32),
.B2(n_20),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_36),
.B(n_26),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_50),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_30),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_57),
.Y(n_67)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_26),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_54),
.Y(n_69)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_37),
.Y(n_61)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_33),
.B1(n_21),
.B2(n_25),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_65),
.A2(n_73),
.B1(n_35),
.B2(n_59),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_68),
.A2(n_33),
.B1(n_34),
.B2(n_56),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_39),
.B1(n_33),
.B2(n_20),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_70),
.A2(n_78),
.B1(n_81),
.B2(n_35),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_34),
.C(n_40),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_35),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_42),
.A2(n_20),
.B1(n_32),
.B2(n_17),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_43),
.B(n_41),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_55),
.Y(n_88)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_46),
.A2(n_17),
.B1(n_23),
.B2(n_28),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_51),
.A2(n_39),
.B1(n_33),
.B2(n_34),
.Y(n_81)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_61),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_83),
.B(n_85),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_90),
.Y(n_135)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_103),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_46),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_75),
.Y(n_114)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_94),
.B(n_99),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_69),
.A2(n_85),
.B1(n_78),
.B2(n_65),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_95),
.A2(n_102),
.B1(n_86),
.B2(n_76),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_98),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_23),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_39),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_75),
.C(n_81),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_71),
.A2(n_35),
.B1(n_59),
.B2(n_40),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_104),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_109),
.Y(n_126)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_76),
.B1(n_63),
.B2(n_77),
.Y(n_129)
);

NAND2x1_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_37),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_31),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_31),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_111),
.Y(n_131)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_88),
.B1(n_111),
.B2(n_108),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_136),
.B1(n_138),
.B2(n_96),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_118),
.Y(n_145)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_115),
.B(n_116),
.Y(n_146)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_85),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_37),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_75),
.C(n_64),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_122),
.C(n_133),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_74),
.C(n_70),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_125),
.B(n_132),
.Y(n_157)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_129),
.A2(n_91),
.B1(n_80),
.B2(n_106),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_97),
.B(n_24),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_130),
.B(n_22),
.Y(n_166)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_93),
.B(n_74),
.C(n_86),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_134),
.B(n_80),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_96),
.A2(n_79),
.B1(n_82),
.B2(n_83),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_139),
.A2(n_149),
.B1(n_166),
.B2(n_128),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_140),
.B(n_153),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_89),
.B(n_1),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_141),
.Y(n_172)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_144),
.Y(n_177)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_101),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_148),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_101),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_137),
.A2(n_28),
.B(n_16),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_150),
.A2(n_151),
.B(n_162),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_137),
.A2(n_16),
.B(n_19),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_154),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_40),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_104),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_135),
.B(n_30),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_122),
.Y(n_169)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_13),
.C(n_15),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_156),
.B(n_160),
.Y(n_171)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_123),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_125),
.Y(n_161)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_119),
.A2(n_19),
.B(n_30),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_163),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_134),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_132),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_167),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_146),
.A2(n_124),
.B1(n_116),
.B2(n_115),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_168),
.A2(n_173),
.B1(n_185),
.B2(n_187),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_178),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_139),
.A2(n_121),
.B1(n_136),
.B2(n_120),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_113),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_179),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_126),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_190),
.C(n_193),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_143),
.A2(n_152),
.B1(n_141),
.B2(n_144),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_147),
.A2(n_112),
.B1(n_130),
.B2(n_31),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_148),
.A2(n_154),
.B1(n_145),
.B2(n_155),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_140),
.B(n_112),
.C(n_40),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_157),
.A2(n_27),
.B1(n_22),
.B2(n_53),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_192),
.A2(n_29),
.B1(n_1),
.B2(n_2),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_153),
.B(n_145),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_172),
.A2(n_162),
.B(n_161),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_194),
.A2(n_200),
.B(n_211),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_197),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_171),
.B(n_163),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_159),
.Y(n_198)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_198),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_172),
.A2(n_150),
.B(n_151),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_186),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_208),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_173),
.A2(n_158),
.B1(n_27),
.B2(n_22),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_206),
.A2(n_210),
.B1(n_212),
.B2(n_215),
.Y(n_226)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_168),
.Y(n_209)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_187),
.A2(n_27),
.B1(n_53),
.B2(n_40),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_175),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_40),
.C(n_29),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_176),
.C(n_207),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_214),
.A2(n_191),
.B1(n_181),
.B2(n_174),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_191),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_170),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_183),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_194),
.Y(n_218)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_219),
.B(n_235),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_204),
.B(n_169),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_210),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_234),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_180),
.C(n_176),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_228),
.C(n_229),
.Y(n_238)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_227),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_190),
.C(n_193),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_29),
.C(n_8),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_29),
.C(n_9),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_232),
.C(n_214),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_7),
.C(n_14),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_7),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_199),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_195),
.Y(n_237)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_237),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_249),
.Y(n_259)
);

NOR2xp67_ASAP7_75t_SL g240 ( 
.A(n_222),
.B(n_199),
.Y(n_240)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_240),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_206),
.C(n_201),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_246),
.C(n_232),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_245),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_230),
.A2(n_196),
.B(n_215),
.Y(n_244)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_244),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_223),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_215),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_211),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_247),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_6),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_246),
.Y(n_251)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_251),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_3),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_250),
.A2(n_233),
.B1(n_231),
.B2(n_226),
.Y(n_254)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_254),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_241),
.A2(n_239),
.B(n_243),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_255),
.A2(n_258),
.B(n_263),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_236),
.A2(n_229),
.B(n_6),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_242),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_262)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_262),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_10),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_259),
.B(n_238),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_272),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_256),
.A2(n_238),
.B(n_245),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_266),
.B(n_269),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_10),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_261),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_271),
.A2(n_251),
.B1(n_255),
.B2(n_252),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_263),
.B(n_11),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_11),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_258),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_262),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_279),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_277),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_274),
.B(n_253),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_270),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_269),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_281),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_257),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_267),
.A2(n_257),
.B1(n_4),
.B2(n_5),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_283),
.B(n_268),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_288),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_282),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_289),
.B(n_276),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_291),
.B(n_292),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_265),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_290),
.A2(n_282),
.B(n_287),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_294),
.A2(n_286),
.B(n_271),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_293),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_12),
.C(n_14),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_12),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_2),
.B1(n_15),
.B2(n_287),
.Y(n_299)
);


endmodule