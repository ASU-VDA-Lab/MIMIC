module real_aes_17718_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_453;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_815;
wire n_638;
wire n_564;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_756;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g832 ( .A(n_0), .B(n_833), .Y(n_832) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_1), .A2(n_4), .B1(n_201), .B2(n_586), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g138 ( .A1(n_2), .A2(n_45), .B1(n_139), .B2(n_141), .Y(n_138) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_3), .A2(n_26), .B1(n_141), .B2(n_165), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_5), .A2(n_16), .B1(n_182), .B2(n_219), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_6), .A2(n_62), .B1(n_167), .B2(n_239), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_7), .A2(n_17), .B1(n_139), .B2(n_186), .Y(n_509) );
INVx1_ASAP7_75t_L g833 ( .A(n_8), .Y(n_833) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_9), .Y(n_571) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_10), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_11), .A2(n_18), .B1(n_184), .B2(n_238), .Y(n_237) );
AOI22xp5_ASAP7_75t_L g810 ( .A1(n_12), .A2(n_66), .B1(n_811), .B2(n_812), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_12), .Y(n_811) );
OR2x2_ASAP7_75t_L g120 ( .A(n_13), .B(n_40), .Y(n_120) );
BUFx2_ASAP7_75t_L g836 ( .A(n_13), .Y(n_836) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_14), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_15), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_19), .A2(n_104), .B1(n_823), .B2(n_839), .Y(n_103) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_20), .A2(n_101), .B1(n_182), .B2(n_201), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g815 ( .A1(n_21), .A2(n_475), .B(n_816), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_22), .A2(n_41), .B1(n_215), .B2(n_216), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_23), .B(n_183), .Y(n_256) );
OAI22x1_ASAP7_75t_SL g808 ( .A1(n_24), .A2(n_809), .B1(n_810), .B2(n_813), .Y(n_808) );
CKINVDCx5p33_ASAP7_75t_R g813 ( .A(n_24), .Y(n_813) );
OAI21x1_ASAP7_75t_L g155 ( .A1(n_25), .A2(n_60), .B(n_156), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_27), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g579 ( .A(n_28), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_29), .B(n_145), .Y(n_533) );
INVx4_ASAP7_75t_R g522 ( .A(n_30), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g146 ( .A1(n_31), .A2(n_49), .B1(n_147), .B2(n_149), .Y(n_146) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_32), .A2(n_56), .B1(n_149), .B2(n_182), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_33), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_34), .B(n_215), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_35), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_36), .B(n_141), .Y(n_540) );
INVx1_ASAP7_75t_L g588 ( .A(n_37), .Y(n_588) );
A2O1A1Ixp33_ASAP7_75t_SL g569 ( .A1(n_38), .A2(n_139), .B(n_151), .C(n_570), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_39), .A2(n_57), .B1(n_139), .B2(n_149), .Y(n_577) );
HB1xp67_ASAP7_75t_L g838 ( .A(n_40), .Y(n_838) );
AOI22xp5_ASAP7_75t_L g163 ( .A1(n_42), .A2(n_89), .B1(n_139), .B2(n_164), .Y(n_163) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_43), .A2(n_55), .B1(n_124), .B2(n_125), .Y(n_123) );
INVx1_ASAP7_75t_L g125 ( .A(n_43), .Y(n_125) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_44), .A2(n_48), .B1(n_139), .B2(n_186), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g567 ( .A(n_46), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_47), .A2(n_61), .B1(n_182), .B2(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g537 ( .A(n_50), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_51), .B(n_139), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_52), .Y(n_550) );
INVx2_ASAP7_75t_L g108 ( .A(n_53), .Y(n_108) );
INVx1_ASAP7_75t_L g118 ( .A(n_54), .Y(n_118) );
BUFx3_ASAP7_75t_L g485 ( .A(n_54), .Y(n_485) );
INVx1_ASAP7_75t_L g124 ( .A(n_55), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g523 ( .A(n_58), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_59), .A2(n_90), .B1(n_139), .B2(n_149), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_63), .A2(n_78), .B1(n_147), .B2(n_204), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g512 ( .A(n_64), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g185 ( .A1(n_65), .A2(n_80), .B1(n_139), .B2(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g812 ( .A(n_66), .Y(n_812) );
CKINVDCx5p33_ASAP7_75t_R g476 ( .A(n_67), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_68), .A2(n_100), .B1(n_182), .B2(n_184), .Y(n_181) );
AND2x4_ASAP7_75t_L g135 ( .A(n_69), .B(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g156 ( .A(n_70), .Y(n_156) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_71), .A2(n_92), .B1(n_147), .B2(n_149), .Y(n_584) );
AO22x1_ASAP7_75t_L g498 ( .A1(n_72), .A2(n_79), .B1(n_216), .B2(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g136 ( .A(n_73), .Y(n_136) );
AND2x2_ASAP7_75t_L g572 ( .A(n_74), .B(n_153), .Y(n_572) );
CKINVDCx14_ASAP7_75t_R g112 ( .A(n_75), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_75), .B(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_76), .B(n_167), .Y(n_556) );
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_77), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_81), .B(n_141), .Y(n_551) );
INVx2_ASAP7_75t_L g145 ( .A(n_82), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_83), .B(n_153), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g519 ( .A(n_84), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g166 ( .A1(n_85), .A2(n_99), .B1(n_149), .B2(n_167), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_86), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_87), .B(n_174), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_88), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_91), .B(n_153), .Y(n_261) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_93), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_94), .B(n_153), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_95), .B(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g806 ( .A(n_95), .Y(n_806) );
NAND2xp33_ASAP7_75t_L g259 ( .A(n_96), .B(n_183), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_97), .A2(n_167), .B(n_169), .C(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g524 ( .A(n_98), .B(n_525), .Y(n_524) );
NAND2xp33_ASAP7_75t_L g555 ( .A(n_102), .B(n_148), .Y(n_555) );
OR2x6_ASAP7_75t_L g104 ( .A(n_105), .B(n_478), .Y(n_104) );
NOR2x1_ASAP7_75t_L g105 ( .A(n_106), .B(n_109), .Y(n_105) );
BUFx8_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVx3_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g482 ( .A(n_108), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_108), .B(n_820), .Y(n_819) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_470), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_121), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
INVx3_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
CKINVDCx8_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
INVx4_ASAP7_75t_L g474 ( .A(n_115), .Y(n_474) );
INVx5_ASAP7_75t_L g477 ( .A(n_115), .Y(n_477) );
AND2x6_ASAP7_75t_SL g115 ( .A(n_116), .B(n_119), .Y(n_115) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
HB1xp67_ASAP7_75t_L g829 ( .A(n_118), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_119), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NOR2x1_ASAP7_75t_L g822 ( .A(n_120), .B(n_485), .Y(n_822) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AOI21xp33_ASAP7_75t_SL g470 ( .A1(n_122), .A2(n_471), .B(n_475), .Y(n_470) );
XNOR2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_126), .Y(n_122) );
OAI22x1_ASAP7_75t_L g488 ( .A1(n_126), .A2(n_489), .B1(n_803), .B2(n_807), .Y(n_488) );
NOR2x1p5_ASAP7_75t_L g126 ( .A(n_127), .B(n_380), .Y(n_126) );
NAND4xp75_ASAP7_75t_L g127 ( .A(n_128), .B(n_325), .C(n_345), .D(n_361), .Y(n_127) );
NOR2x1p5_ASAP7_75t_SL g128 ( .A(n_129), .B(n_295), .Y(n_128) );
NAND4xp75_ASAP7_75t_L g129 ( .A(n_130), .B(n_231), .C(n_272), .D(n_281), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_192), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_159), .Y(n_131) );
AND2x4_ASAP7_75t_L g405 ( .A(n_132), .B(n_332), .Y(n_405) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_133), .Y(n_248) );
INVx2_ASAP7_75t_L g266 ( .A(n_133), .Y(n_266) );
AND2x2_ASAP7_75t_L g289 ( .A(n_133), .B(n_251), .Y(n_289) );
OR2x2_ASAP7_75t_L g344 ( .A(n_133), .B(n_160), .Y(n_344) );
AO31x2_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_137), .A3(n_152), .B(n_157), .Y(n_133) );
INVx2_ASAP7_75t_L g189 ( .A(n_134), .Y(n_189) );
AO31x2_ASAP7_75t_L g212 ( .A1(n_134), .A2(n_161), .A3(n_213), .B(n_221), .Y(n_212) );
AO31x2_ASAP7_75t_L g235 ( .A1(n_134), .A2(n_178), .A3(n_236), .B(n_242), .Y(n_235) );
AO31x2_ASAP7_75t_L g507 ( .A1(n_134), .A2(n_209), .A3(n_508), .B(n_511), .Y(n_507) );
BUFx10_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g171 ( .A(n_135), .Y(n_171) );
INVx1_ASAP7_75t_L g505 ( .A(n_135), .Y(n_505) );
BUFx10_ASAP7_75t_L g542 ( .A(n_135), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_142), .B1(n_146), .B2(n_150), .Y(n_137) );
INVx1_ASAP7_75t_L g184 ( .A(n_139), .Y(n_184) );
INVx4_ASAP7_75t_L g186 ( .A(n_139), .Y(n_186) );
INVx1_ASAP7_75t_L g204 ( .A(n_139), .Y(n_204) );
INVx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_140), .Y(n_141) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_140), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_140), .Y(n_149) );
INVx2_ASAP7_75t_L g165 ( .A(n_140), .Y(n_165) );
INVx1_ASAP7_75t_L g167 ( .A(n_140), .Y(n_167) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_140), .Y(n_183) );
INVx1_ASAP7_75t_L g202 ( .A(n_140), .Y(n_202) );
INVx1_ASAP7_75t_L g217 ( .A(n_140), .Y(n_217) );
INVx1_ASAP7_75t_L g220 ( .A(n_140), .Y(n_220) );
INVx1_ASAP7_75t_L g240 ( .A(n_140), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_141), .B(n_565), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_142), .A2(n_150), .B1(n_200), .B2(n_203), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g213 ( .A1(n_142), .A2(n_150), .B1(n_214), .B2(n_218), .Y(n_213) );
OAI22xp5_ASAP7_75t_L g226 ( .A1(n_142), .A2(n_150), .B1(n_227), .B2(n_228), .Y(n_226) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g501 ( .A(n_143), .Y(n_501) );
BUFx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g553 ( .A(n_144), .Y(n_553) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
BUFx8_ASAP7_75t_L g151 ( .A(n_145), .Y(n_151) );
INVx1_ASAP7_75t_L g169 ( .A(n_145), .Y(n_169) );
INVx1_ASAP7_75t_L g536 ( .A(n_145), .Y(n_536) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g215 ( .A(n_148), .Y(n_215) );
OAI22xp33_ASAP7_75t_L g521 ( .A1(n_148), .A2(n_220), .B1(n_522), .B2(n_523), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_149), .B(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g586 ( .A(n_149), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g162 ( .A1(n_150), .A2(n_163), .B1(n_166), .B2(n_168), .Y(n_162) );
OAI22xp5_ASAP7_75t_L g180 ( .A1(n_150), .A2(n_181), .B1(n_185), .B2(n_187), .Y(n_180) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_150), .A2(n_187), .B1(n_237), .B2(n_241), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_150), .A2(n_258), .B(n_259), .Y(n_257) );
OAI22x1_ASAP7_75t_L g508 ( .A1(n_150), .A2(n_168), .B1(n_509), .B2(n_510), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_150), .A2(n_501), .B1(n_576), .B2(n_577), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_150), .A2(n_168), .B1(n_584), .B2(n_585), .Y(n_583) );
INVx6_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
O2A1O1Ixp5_ASAP7_75t_L g254 ( .A1(n_151), .A2(n_186), .B(n_255), .C(n_256), .Y(n_254) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_151), .A2(n_498), .B(n_500), .C(n_504), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_151), .A2(n_555), .B(n_556), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_151), .B(n_498), .Y(n_600) );
AO31x2_ASAP7_75t_L g574 ( .A1(n_152), .A2(n_542), .A3(n_575), .B(n_578), .Y(n_574) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NOR2x1_ASAP7_75t_L g557 ( .A(n_153), .B(n_558), .Y(n_557) );
INVx4_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_154), .B(n_158), .Y(n_157) );
BUFx3_ASAP7_75t_L g161 ( .A(n_154), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_154), .B(n_191), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_154), .B(n_222), .Y(n_221) );
INVx2_ASAP7_75t_SL g252 ( .A(n_154), .Y(n_252) );
AND2x2_ASAP7_75t_L g541 ( .A(n_154), .B(n_542), .Y(n_541) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g174 ( .A(n_155), .Y(n_174) );
AND2x2_ASAP7_75t_L g262 ( .A(n_159), .B(n_263), .Y(n_262) );
AND2x4_ASAP7_75t_L g412 ( .A(n_159), .B(n_289), .Y(n_412) );
AND2x4_ASAP7_75t_L g159 ( .A(n_160), .B(n_176), .Y(n_159) );
OR2x2_ASAP7_75t_L g249 ( .A(n_160), .B(n_250), .Y(n_249) );
BUFx2_ASAP7_75t_L g280 ( .A(n_160), .Y(n_280) );
AND2x2_ASAP7_75t_L g286 ( .A(n_160), .B(n_177), .Y(n_286) );
INVx1_ASAP7_75t_L g304 ( .A(n_160), .Y(n_304) );
INVx2_ASAP7_75t_L g333 ( .A(n_160), .Y(n_333) );
AO31x2_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_162), .A3(n_170), .B(n_172), .Y(n_160) );
INVx2_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_165), .B(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_168), .B(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_SL g187 ( .A(n_169), .Y(n_187) );
AO31x2_ASAP7_75t_L g225 ( .A1(n_170), .A2(n_205), .A3(n_226), .B(n_229), .Y(n_225) );
AO31x2_ASAP7_75t_L g582 ( .A1(n_170), .A2(n_178), .A3(n_583), .B(n_587), .Y(n_582) );
INVx2_ASAP7_75t_SL g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_SL g260 ( .A(n_171), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_173), .B(n_175), .Y(n_172) );
INVx2_ASAP7_75t_L g206 ( .A(n_173), .Y(n_206) );
NOR2xp33_ASAP7_75t_SL g242 ( .A(n_173), .B(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g179 ( .A(n_174), .Y(n_179) );
INVx2_ASAP7_75t_L g209 ( .A(n_174), .Y(n_209) );
OAI21xp33_ASAP7_75t_L g504 ( .A1(n_174), .A2(n_503), .B(n_505), .Y(n_504) );
INVx3_ASAP7_75t_L g309 ( .A(n_176), .Y(n_309) );
INVx2_ASAP7_75t_L g314 ( .A(n_176), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_176), .B(n_265), .Y(n_319) );
AND2x2_ASAP7_75t_L g342 ( .A(n_176), .B(n_321), .Y(n_342) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_176), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_176), .B(n_397), .Y(n_396) );
INVx3_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
BUFx2_ASAP7_75t_L g331 ( .A(n_177), .Y(n_331) );
AND2x2_ASAP7_75t_L g379 ( .A(n_177), .B(n_333), .Y(n_379) );
AO31x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_180), .A3(n_188), .B(n_190), .Y(n_177) );
AOI21x1_ASAP7_75t_L g561 ( .A1(n_178), .A2(n_562), .B(n_572), .Y(n_561) );
BUFx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_179), .B(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g525 ( .A(n_179), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_179), .B(n_579), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_179), .B(n_588), .Y(n_587) );
INVx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVxp67_ASAP7_75t_SL g499 ( .A(n_183), .Y(n_499) );
O2A1O1Ixp33_ASAP7_75t_L g549 ( .A1(n_186), .A2(n_550), .B(n_551), .C(n_552), .Y(n_549) );
AO31x2_ASAP7_75t_L g198 ( .A1(n_188), .A2(n_199), .A3(n_205), .B(n_207), .Y(n_198) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_189), .A2(n_517), .B(n_520), .Y(n_516) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_194), .B(n_210), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_194), .B(n_323), .Y(n_370) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NAND2x1p5_ASAP7_75t_L g367 ( .A(n_195), .B(n_323), .Y(n_367) );
INVx1_ASAP7_75t_L g468 ( .A(n_195), .Y(n_468) );
INVx3_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g418 ( .A(n_196), .B(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g271 ( .A(n_197), .Y(n_271) );
OR2x2_ASAP7_75t_L g352 ( .A(n_197), .B(n_224), .Y(n_352) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g294 ( .A(n_198), .Y(n_294) );
AND2x4_ASAP7_75t_L g300 ( .A(n_198), .B(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_202), .B(n_567), .Y(n_566) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_205), .A2(n_516), .B(n_524), .Y(n_515) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_209), .B(n_230), .Y(n_229) );
AOI32xp33_ASAP7_75t_L g438 ( .A1(n_210), .A2(n_341), .A3(n_439), .B1(n_441), .B2(n_442), .Y(n_438) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
OR2x2_ASAP7_75t_L g387 ( .A(n_211), .B(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_212), .B(n_223), .Y(n_211) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_212), .Y(n_233) );
OR2x2_ASAP7_75t_L g269 ( .A(n_212), .B(n_225), .Y(n_269) );
INVx1_ASAP7_75t_L g284 ( .A(n_212), .Y(n_284) );
AND2x2_ASAP7_75t_L g293 ( .A(n_212), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g299 ( .A(n_212), .Y(n_299) );
INVx2_ASAP7_75t_L g324 ( .A(n_212), .Y(n_324) );
AND2x2_ASAP7_75t_L g443 ( .A(n_212), .B(n_235), .Y(n_443) );
OAI21xp33_ASAP7_75t_SL g532 ( .A1(n_216), .A2(n_533), .B(n_534), .Y(n_532) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_223), .B(n_276), .Y(n_363) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g234 ( .A(n_225), .B(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g292 ( .A(n_225), .Y(n_292) );
INVx2_ASAP7_75t_L g301 ( .A(n_225), .Y(n_301) );
AND2x4_ASAP7_75t_L g323 ( .A(n_225), .B(n_324), .Y(n_323) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_225), .Y(n_415) );
AOI22x1_ASAP7_75t_SL g231 ( .A1(n_232), .A2(n_244), .B1(n_262), .B2(n_267), .Y(n_231) );
AND2x4_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
NAND4xp25_ASAP7_75t_L g392 ( .A(n_234), .B(n_393), .C(n_394), .D(n_395), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_234), .B(n_293), .Y(n_423) );
INVx4_ASAP7_75t_SL g276 ( .A(n_235), .Y(n_276) );
BUFx2_ASAP7_75t_L g339 ( .A(n_235), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_235), .B(n_284), .Y(n_402) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_240), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g364 ( .A(n_246), .B(n_313), .Y(n_364) );
NOR2x1_ASAP7_75t_L g246 ( .A(n_247), .B(n_249), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x4_ASAP7_75t_L g287 ( .A(n_250), .B(n_265), .Y(n_287) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_251), .B(n_266), .Y(n_311) );
OAI21x1_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_253), .B(n_261), .Y(n_251) );
OAI21x1_ASAP7_75t_L g306 ( .A1(n_252), .A2(n_253), .B(n_261), .Y(n_306) );
OAI21x1_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_257), .B(n_260), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_263), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g329 ( .A(n_263), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g368 ( .A(n_264), .B(n_286), .Y(n_368) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g411 ( .A(n_266), .B(n_321), .Y(n_411) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_267), .A2(n_384), .B1(n_386), .B2(n_389), .C(n_391), .Y(n_383) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx2_ASAP7_75t_L g277 ( .A(n_269), .Y(n_277) );
OR2x2_ASAP7_75t_L g377 ( .A(n_269), .B(n_316), .Y(n_377) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_278), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_273), .A2(n_399), .B1(n_403), .B2(n_406), .Y(n_398) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_277), .Y(n_273) );
AND2x4_ASAP7_75t_L g322 ( .A(n_274), .B(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g434 ( .A(n_274), .B(n_352), .Y(n_434) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x4_ASAP7_75t_L g282 ( .A(n_276), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g298 ( .A(n_276), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g357 ( .A(n_276), .B(n_294), .Y(n_357) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_276), .Y(n_374) );
INVx1_ASAP7_75t_L g388 ( .A(n_276), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_276), .B(n_301), .Y(n_431) );
AND2x4_ASAP7_75t_L g338 ( .A(n_277), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g336 ( .A(n_279), .Y(n_336) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_280), .B(n_321), .Y(n_320) );
NAND2x1_ASAP7_75t_L g440 ( .A(n_280), .B(n_342), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_285), .B1(n_288), .B2(n_290), .Y(n_281) );
AND2x2_ASAP7_75t_L g307 ( .A(n_282), .B(n_300), .Y(n_307) );
INVx1_ASAP7_75t_L g348 ( .A(n_282), .Y(n_348) );
AND2x2_ASAP7_75t_L g455 ( .A(n_282), .B(n_316), .Y(n_455) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x4_ASAP7_75t_SL g285 ( .A(n_286), .B(n_287), .Y(n_285) );
AND2x2_ASAP7_75t_L g288 ( .A(n_286), .B(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g428 ( .A(n_286), .Y(n_428) );
AND2x2_ASAP7_75t_L g445 ( .A(n_286), .B(n_305), .Y(n_445) );
AND2x2_ASAP7_75t_L g461 ( .A(n_286), .B(n_411), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_287), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g384 ( .A(n_287), .B(n_385), .Y(n_384) );
OAI22xp33_ASAP7_75t_L g391 ( .A1(n_287), .A2(n_377), .B1(n_392), .B2(n_396), .Y(n_391) );
INVx1_ASAP7_75t_L g347 ( .A(n_289), .Y(n_347) );
AND2x2_ASAP7_75t_L g378 ( .A(n_289), .B(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_289), .B(n_385), .Y(n_407) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g413 ( .A(n_293), .B(n_414), .Y(n_413) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_293), .A2(n_317), .B1(n_422), .B2(n_424), .Y(n_421) );
INVx3_ASAP7_75t_L g316 ( .A(n_294), .Y(n_316) );
AND2x2_ASAP7_75t_L g448 ( .A(n_294), .B(n_301), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_312), .Y(n_295) );
AOI32xp33_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_302), .A3(n_305), .B1(n_307), .B2(n_308), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_300), .Y(n_297) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_299), .Y(n_394) );
INVx1_ASAP7_75t_L g419 ( .A(n_299), .Y(n_419) );
INVx3_ASAP7_75t_L g375 ( .A(n_300), .Y(n_375) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OAI221xp5_ASAP7_75t_L g450 ( .A1(n_303), .A2(n_451), .B1(n_452), .B2(n_453), .C(n_454), .Y(n_450) );
BUFx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g427 ( .A(n_305), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g463 ( .A(n_305), .B(n_424), .Y(n_463) );
BUFx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g321 ( .A(n_306), .Y(n_321) );
NAND2x1p5_ASAP7_75t_L g335 ( .A(n_308), .B(n_336), .Y(n_335) );
AO22x1_ASAP7_75t_L g365 ( .A1(n_308), .A2(n_366), .B1(n_368), .B2(n_369), .Y(n_365) );
NAND2x1p5_ASAP7_75t_L g469 ( .A(n_308), .B(n_336), .Y(n_469) );
AND2x4_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx2_ASAP7_75t_L g385 ( .A(n_309), .Y(n_385) );
INVx1_ASAP7_75t_L g395 ( .A(n_309), .Y(n_395) );
AND2x2_ASAP7_75t_L g315 ( .A(n_310), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVxp67_ASAP7_75t_SL g397 ( .A(n_311), .Y(n_397) );
INVx1_ASAP7_75t_L g437 ( .A(n_311), .Y(n_437) );
A2O1A1Ixp33_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_315), .B(n_317), .C(n_322), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NOR2x1p5_ASAP7_75t_L g424 ( .A(n_314), .B(n_344), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_315), .B(n_374), .Y(n_451) );
AOI31xp33_ASAP7_75t_L g334 ( .A1(n_316), .A2(n_335), .A3(n_337), .B(n_340), .Y(n_334) );
INVx4_ASAP7_75t_L g393 ( .A(n_316), .Y(n_393) );
OR2x2_ASAP7_75t_L g430 ( .A(n_316), .B(n_431), .Y(n_430) );
INVx2_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AND2x4_ASAP7_75t_L g332 ( .A(n_321), .B(n_333), .Y(n_332) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_323), .Y(n_328) );
AND2x2_ASAP7_75t_L g359 ( .A(n_323), .B(n_357), .Y(n_359) );
NOR2xp67_ASAP7_75t_L g325 ( .A(n_326), .B(n_334), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_L g452 ( .A(n_329), .Y(n_452) );
INVx1_ASAP7_75t_L g360 ( .A(n_330), .Y(n_360) );
AND2x4_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx1_ASAP7_75t_L g390 ( .A(n_331), .Y(n_390) );
AND2x2_ASAP7_75t_L g389 ( .A(n_332), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OAI322xp33_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_348), .A3(n_349), .B1(n_353), .B2(n_356), .C1(n_358), .C2(n_360), .Y(n_346) );
INVxp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AOI211x1_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_364), .B(n_365), .C(n_371), .Y(n_361) );
INVx1_ASAP7_75t_L g466 ( .A(n_362), .Y(n_466) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g420 ( .A(n_364), .Y(n_420) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OA21x2_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_376), .B(n_378), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVx2_ASAP7_75t_L g441 ( .A(n_375), .Y(n_441) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp33_ASAP7_75t_L g436 ( .A(n_379), .B(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_381), .B(n_449), .Y(n_380) );
NOR3xp33_ASAP7_75t_L g381 ( .A(n_382), .B(n_416), .C(n_432), .Y(n_381) );
NAND3xp33_ASAP7_75t_L g382 ( .A(n_383), .B(n_398), .C(n_408), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_385), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OAI21xp33_ASAP7_75t_L g444 ( .A1(n_389), .A2(n_445), .B(n_446), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_393), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_393), .B(n_443), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_394), .B(n_468), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_395), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OAI21xp5_ASAP7_75t_L g454 ( .A1(n_405), .A2(n_455), .B(n_456), .Y(n_454) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OAI21xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_412), .B(n_413), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OAI211xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_420), .B(n_421), .C(n_425), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_429), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_SL g435 ( .A(n_427), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_431), .Y(n_453) );
OAI211xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_435), .B(n_438), .C(n_444), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_443), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g464 ( .A(n_443), .Y(n_464) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g460 ( .A(n_448), .Y(n_460) );
NOR3xp33_ASAP7_75t_L g449 ( .A(n_450), .B(n_458), .C(n_465), .Y(n_449) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AOI21xp33_ASAP7_75t_SL g458 ( .A1(n_459), .A2(n_462), .B(n_464), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AOI21xp33_ASAP7_75t_R g465 ( .A1(n_466), .A2(n_467), .B(n_469), .Y(n_465) );
INVx4_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx12f_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
OAI21xp33_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_486), .B(n_815), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g479 ( .A(n_480), .Y(n_479) );
BUFx12f_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AND2x6_ASAP7_75t_SL g481 ( .A(n_482), .B(n_483), .Y(n_481) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_488), .B1(n_808), .B2(n_814), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x4_ASAP7_75t_L g489 ( .A(n_490), .B(n_713), .Y(n_489) );
NOR3xp33_ASAP7_75t_L g490 ( .A(n_491), .B(n_642), .C(n_684), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_616), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_526), .B1(n_591), .B2(n_602), .Y(n_492) );
INVx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_513), .Y(n_494) );
AOI21xp33_ASAP7_75t_L g635 ( .A1(n_495), .A2(n_636), .B(n_638), .Y(n_635) );
AOI21xp33_ASAP7_75t_L g708 ( .A1(n_495), .A2(n_709), .B(n_710), .Y(n_708) );
OR2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_506), .Y(n_495) );
INVx2_ASAP7_75t_L g628 ( .A(n_496), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_496), .B(n_507), .Y(n_658) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g599 ( .A(n_500), .Y(n_599) );
OAI21x1_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_502), .B(n_503), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_501), .A2(n_539), .B(n_540), .Y(n_538) );
INVx1_ASAP7_75t_L g601 ( .A(n_504), .Y(n_601) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_505), .A2(n_563), .B(n_569), .Y(n_562) );
AND2x2_ASAP7_75t_L g698 ( .A(n_506), .B(n_545), .Y(n_698) );
INVx1_ASAP7_75t_L g731 ( .A(n_506), .Y(n_731) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g593 ( .A(n_507), .B(n_546), .Y(n_593) );
AND2x2_ASAP7_75t_L g624 ( .A(n_507), .B(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g633 ( .A(n_507), .Y(n_633) );
OR2x2_ASAP7_75t_L g652 ( .A(n_507), .B(n_515), .Y(n_652) );
AND2x2_ASAP7_75t_L g667 ( .A(n_507), .B(n_515), .Y(n_667) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_514), .B(n_666), .Y(n_709) );
OR2x2_ASAP7_75t_L g797 ( .A(n_514), .B(n_658), .Y(n_797) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g625 ( .A(n_515), .Y(n_625) );
AND2x2_ASAP7_75t_L g634 ( .A(n_515), .B(n_597), .Y(n_634) );
AND2x2_ASAP7_75t_L g637 ( .A(n_515), .B(n_546), .Y(n_637) );
AND2x2_ASAP7_75t_L g656 ( .A(n_515), .B(n_545), .Y(n_656) );
AND2x4_ASAP7_75t_L g675 ( .A(n_515), .B(n_598), .Y(n_675) );
OAI21xp33_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_543), .B(n_580), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g773 ( .A(n_527), .B(n_670), .Y(n_773) );
CKINVDCx14_ASAP7_75t_R g527 ( .A(n_528), .Y(n_527) );
BUFx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_529), .B(n_590), .Y(n_589) );
INVx3_ASAP7_75t_L g606 ( .A(n_529), .Y(n_606) );
OR2x2_ASAP7_75t_L g614 ( .A(n_529), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_529), .B(n_607), .Y(n_639) );
AND2x2_ASAP7_75t_L g664 ( .A(n_529), .B(n_582), .Y(n_664) );
AND2x2_ASAP7_75t_L g682 ( .A(n_529), .B(n_612), .Y(n_682) );
INVx1_ASAP7_75t_L g721 ( .A(n_529), .Y(n_721) );
AND2x2_ASAP7_75t_L g723 ( .A(n_529), .B(n_724), .Y(n_723) );
NAND2x1p5_ASAP7_75t_SL g742 ( .A(n_529), .B(n_663), .Y(n_742) );
AND2x4_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_538), .B(n_541), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
BUFx4f_ASAP7_75t_L g568 ( .A(n_536), .Y(n_568) );
INVx1_ASAP7_75t_L g558 ( .A(n_542), .Y(n_558) );
OAI32xp33_ASAP7_75t_L g626 ( .A1(n_543), .A2(n_618), .A3(n_627), .B1(n_629), .B2(n_631), .Y(n_626) );
OR2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_559), .Y(n_543) );
INVx1_ASAP7_75t_L g666 ( .A(n_544), .Y(n_666) );
AND2x2_ASAP7_75t_L g674 ( .A(n_544), .B(n_675), .Y(n_674) );
BUFx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g673 ( .A(n_545), .B(n_597), .Y(n_673) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
BUFx3_ASAP7_75t_L g623 ( .A(n_546), .Y(n_623) );
AND2x2_ASAP7_75t_L g632 ( .A(n_546), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g738 ( .A(n_546), .Y(n_738) );
NAND2x1p5_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
OAI21x1_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_554), .B(n_557), .Y(n_548) );
INVx2_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g608 ( .A(n_559), .Y(n_608) );
OR2x2_ASAP7_75t_L g618 ( .A(n_559), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g740 ( .A(n_559), .Y(n_740) );
OR2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_573), .Y(n_559) );
AND2x2_ASAP7_75t_L g641 ( .A(n_560), .B(n_574), .Y(n_641) );
INVx2_ASAP7_75t_L g663 ( .A(n_560), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_560), .B(n_582), .Y(n_683) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g590 ( .A(n_561), .Y(n_590) );
OAI21xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_566), .B(n_568), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_573), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g672 ( .A(n_573), .Y(n_672) );
INVx2_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
BUFx2_ASAP7_75t_L g612 ( .A(n_574), .Y(n_612) );
OR2x2_ASAP7_75t_L g678 ( .A(n_574), .B(n_582), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_574), .B(n_582), .Y(n_711) );
INVx2_ASAP7_75t_L g659 ( .A(n_580), .Y(n_659) );
OR2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_589), .Y(n_580) );
OR2x2_ASAP7_75t_L g646 ( .A(n_581), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g724 ( .A(n_581), .Y(n_724) );
INVx1_ASAP7_75t_L g607 ( .A(n_582), .Y(n_607) );
INVx1_ASAP7_75t_L g615 ( .A(n_582), .Y(n_615) );
INVx1_ASAP7_75t_L g630 ( .A(n_582), .Y(n_630) );
OR2x2_ASAP7_75t_L g734 ( .A(n_589), .B(n_711), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_590), .B(n_606), .Y(n_647) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_590), .Y(n_649) );
OR2x2_ASAP7_75t_L g748 ( .A(n_590), .B(n_672), .Y(n_748) );
INVxp67_ASAP7_75t_L g772 ( .A(n_590), .Y(n_772) );
INVx2_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
NAND2x1_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_593), .B(n_634), .Y(n_701) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g650 ( .A(n_595), .B(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g763 ( .A(n_596), .Y(n_763) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g792 ( .A(n_597), .B(n_625), .Y(n_792) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g718 ( .A(n_598), .B(n_625), .Y(n_718) );
AOI21x1_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_600), .B(n_601), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_609), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_608), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_605), .B(n_641), .Y(n_755) );
AND2x4_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
INVx2_ASAP7_75t_L g619 ( .A(n_606), .Y(n_619) );
AND2x2_ASAP7_75t_L g669 ( .A(n_606), .B(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_606), .B(n_663), .Y(n_712) );
OR2x2_ASAP7_75t_L g784 ( .A(n_606), .B(n_671), .Y(n_784) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g704 ( .A(n_610), .B(n_705), .Y(n_704) );
AND2x4_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
INVx2_ASAP7_75t_L g695 ( .A(n_611), .Y(n_695) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g685 ( .A(n_614), .B(n_686), .Y(n_685) );
INVxp67_ASAP7_75t_SL g696 ( .A(n_614), .Y(n_696) );
OR2x2_ASAP7_75t_L g747 ( .A(n_614), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g802 ( .A(n_614), .Y(n_802) );
AOI211xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_620), .B(n_626), .C(n_635), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g691 ( .A(n_619), .B(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_619), .B(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g764 ( .A(n_619), .B(n_641), .Y(n_764) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_624), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_622), .B(n_667), .Y(n_689) );
NAND2x1p5_ASAP7_75t_L g706 ( .A(n_622), .B(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g774 ( .A(n_622), .B(n_775), .Y(n_774) );
INVx3_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
BUFx2_ASAP7_75t_L g717 ( .A(n_623), .Y(n_717) );
AND2x2_ASAP7_75t_L g745 ( .A(n_624), .B(n_673), .Y(n_745) );
INVx2_ASAP7_75t_L g768 ( .A(n_624), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_624), .B(n_666), .Y(n_800) );
AND2x4_ASAP7_75t_SL g754 ( .A(n_627), .B(n_632), .Y(n_754) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g707 ( .A(n_628), .B(n_633), .Y(n_707) );
OR2x2_ASAP7_75t_L g759 ( .A(n_628), .B(n_652), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_629), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_629), .B(n_641), .Y(n_795) );
BUFx3_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g743 ( .A(n_630), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_634), .Y(n_631) );
INVx1_ASAP7_75t_L g726 ( .A(n_632), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_632), .B(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g776 ( .A(n_633), .Y(n_776) );
BUFx2_ASAP7_75t_L g644 ( .A(n_634), .Y(n_644) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g762 ( .A(n_637), .B(n_763), .Y(n_762) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g686 ( .A(n_641), .Y(n_686) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_641), .Y(n_703) );
NAND3xp33_ASAP7_75t_SL g642 ( .A(n_643), .B(n_653), .C(n_668), .Y(n_642) );
AOI22xp33_ASAP7_75t_SL g643 ( .A1(n_644), .A2(n_645), .B1(n_648), .B2(n_650), .Y(n_643) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AOI222xp33_ASAP7_75t_L g756 ( .A1(n_650), .A2(n_676), .B1(n_757), .B2(n_760), .C1(n_762), .C2(n_764), .Y(n_756) );
AND2x2_ASAP7_75t_L g788 ( .A(n_651), .B(n_737), .Y(n_788) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
OR2x2_ASAP7_75t_L g736 ( .A(n_652), .B(n_737), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_659), .B1(n_660), .B2(n_665), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
INVx2_ASAP7_75t_SL g732 ( .A(n_656), .Y(n_732) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_664), .Y(n_660) );
AND2x2_ASAP7_75t_L g719 ( .A(n_661), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
OR2x2_ASAP7_75t_L g677 ( .A(n_662), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OR2x2_ASAP7_75t_L g671 ( .A(n_663), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g786 ( .A(n_664), .Y(n_786) );
AND2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_667), .B(n_763), .Y(n_782) );
INVx1_ASAP7_75t_L g799 ( .A(n_667), .Y(n_799) );
AOI222xp33_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_673), .B1(n_674), .B2(n_676), .C1(n_679), .C2(n_680), .Y(n_668) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_675), .Y(n_679) );
AND2x2_ASAP7_75t_L g697 ( .A(n_675), .B(n_698), .Y(n_697) );
INVx3_ASAP7_75t_L g728 ( .A(n_675), .Y(n_728) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g692 ( .A(n_678), .Y(n_692) );
OR2x2_ASAP7_75t_L g761 ( .A(n_678), .B(n_742), .Y(n_761) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
OAI211xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_687), .B(n_690), .C(n_699), .Y(n_684) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
OAI21xp33_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_693), .B(n_697), .Y(n_690) );
AOI221xp5_ASAP7_75t_L g777 ( .A1(n_691), .A2(n_729), .B1(n_778), .B2(n_781), .C(n_783), .Y(n_777) );
AND2x4_ASAP7_75t_L g720 ( .A(n_692), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
INVx1_ASAP7_75t_L g751 ( .A(n_698), .Y(n_751) );
AOI211x1_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_702), .B(n_704), .C(n_708), .Y(n_699) );
INVxp67_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g769 ( .A(n_707), .Y(n_769) );
NAND3xp33_ASAP7_75t_L g757 ( .A(n_710), .B(n_758), .C(n_759), .Y(n_757) );
OR2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
INVx1_ASAP7_75t_L g793 ( .A(n_711), .Y(n_793) );
NOR2x1_ASAP7_75t_L g713 ( .A(n_714), .B(n_765), .Y(n_713) );
NAND4xp25_ASAP7_75t_L g714 ( .A(n_715), .B(n_722), .C(n_744), .D(n_756), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_716), .B(n_719), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
AND2x2_ASAP7_75t_L g775 ( .A(n_718), .B(n_776), .Y(n_775) );
AOI221x1_ASAP7_75t_L g744 ( .A1(n_720), .A2(n_745), .B1(n_746), .B2(n_749), .C(n_752), .Y(n_744) );
AND2x2_ASAP7_75t_L g770 ( .A(n_720), .B(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g780 ( .A(n_721), .Y(n_780) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_725), .B1(n_729), .B2(n_733), .C(n_735), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_727), .B(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_732), .A2(n_736), .B1(n_739), .B2(n_741), .Y(n_735) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g752 ( .A1(n_736), .A2(n_753), .B(n_755), .Y(n_752) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g758 ( .A(n_738), .Y(n_758) );
OR2x2_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .Y(n_741) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVxp67_ASAP7_75t_L g779 ( .A(n_748), .Y(n_779) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
OAI22xp33_ASAP7_75t_L g798 ( .A1(n_761), .A2(n_799), .B1(n_800), .B2(n_801), .Y(n_798) );
NAND3xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_777), .C(n_789), .Y(n_765) );
AOI22xp5_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_770), .B1(n_773), .B2(n_774), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
INVxp67_ASAP7_75t_SL g771 ( .A(n_772), .Y(n_771) );
OR2x2_ASAP7_75t_L g785 ( .A(n_772), .B(n_786), .Y(n_785) );
NAND2x1_ASAP7_75t_L g801 ( .A(n_772), .B(n_802), .Y(n_801) );
AND2x2_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
INVx2_ASAP7_75t_SL g781 ( .A(n_782), .Y(n_781) );
AOI21xp5_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_785), .B(n_787), .Y(n_783) );
INVx1_ASAP7_75t_SL g787 ( .A(n_788), .Y(n_787) );
AOI221xp5_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_793), .B1(n_794), .B2(n_796), .C(n_798), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx3_ASAP7_75t_R g796 ( .A(n_797), .Y(n_796) );
INVx4_ASAP7_75t_L g807 ( .A(n_803), .Y(n_807) );
BUFx12f_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
CKINVDCx5p33_ASAP7_75t_R g804 ( .A(n_805), .Y(n_804) );
AND2x2_ASAP7_75t_L g821 ( .A(n_805), .B(n_822), .Y(n_821) );
INVx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
BUFx2_ASAP7_75t_L g831 ( .A(n_806), .Y(n_831) );
CKINVDCx5p33_ASAP7_75t_R g814 ( .A(n_808), .Y(n_814) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx2_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
BUFx10_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_824), .Y(n_823) );
CKINVDCx20_ASAP7_75t_R g824 ( .A(n_825), .Y(n_824) );
CKINVDCx11_ASAP7_75t_R g825 ( .A(n_826), .Y(n_825) );
CKINVDCx10_ASAP7_75t_R g840 ( .A(n_826), .Y(n_840) );
OR2x6_ASAP7_75t_L g826 ( .A(n_827), .B(n_834), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
NOR2x1p5_ASAP7_75t_L g828 ( .A(n_829), .B(n_830), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_831), .B(n_832), .Y(n_830) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
NOR2xp33_ASAP7_75t_L g835 ( .A(n_836), .B(n_837), .Y(n_835) );
INVxp33_ASAP7_75t_SL g837 ( .A(n_838), .Y(n_837) );
CKINVDCx8_ASAP7_75t_R g839 ( .A(n_840), .Y(n_839) );
endmodule