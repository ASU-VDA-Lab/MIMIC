module fake_jpeg_15263_n_307 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_307);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_307;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_41),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_29),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_18),
.B1(n_26),
.B2(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_21),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_46),
.A2(n_56),
.B(n_60),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_21),
.Y(n_49)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_18),
.B1(n_26),
.B2(n_28),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_50),
.A2(n_40),
.B1(n_39),
.B2(n_35),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_18),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_54),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_28),
.B1(n_26),
.B2(n_16),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_52),
.A2(n_31),
.B1(n_40),
.B2(n_35),
.Y(n_74)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_41),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_L g56 ( 
.A1(n_33),
.A2(n_31),
.B(n_23),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_38),
.A2(n_31),
.B1(n_23),
.B2(n_22),
.Y(n_60)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_44),
.B(n_41),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_65),
.B(n_70),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_66),
.B(n_71),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_79),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_37),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_37),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_81),
.B(n_0),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_49),
.B(n_35),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_73),
.B(n_76),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_74),
.A2(n_55),
.B1(n_59),
.B2(n_43),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_37),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_48),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_45),
.A2(n_40),
.B1(n_39),
.B2(n_35),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_80),
.A2(n_55),
.B1(n_43),
.B2(n_42),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_55),
.A2(n_23),
.B1(n_22),
.B2(n_24),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_34),
.C(n_37),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_40),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_47),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_85),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_45),
.B(n_37),
.Y(n_86)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_47),
.B(n_39),
.Y(n_87)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_89),
.A2(n_90),
.B(n_32),
.Y(n_136)
);

OA21x2_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_64),
.B(n_75),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_91),
.B(n_82),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_78),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_100),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_87),
.Y(n_94)
);

INVx3_ASAP7_75t_SL g134 ( 
.A(n_94),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_75),
.A2(n_53),
.B1(n_40),
.B2(n_59),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_113),
.B1(n_114),
.B2(n_68),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_98),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_99),
.A2(n_70),
.B1(n_68),
.B2(n_73),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_16),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_27),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_108),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_66),
.B(n_27),
.Y(n_108)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_71),
.A2(n_43),
.B1(n_25),
.B2(n_19),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_118),
.B(n_138),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_95),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_119),
.B(n_128),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_104),
.B(n_64),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_106),
.Y(n_153)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_130),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_90),
.A2(n_74),
.B1(n_84),
.B2(n_79),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_101),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_90),
.A2(n_65),
.B1(n_68),
.B2(n_80),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_62),
.Y(n_132)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_62),
.Y(n_133)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_136),
.A2(n_137),
.B(n_141),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_97),
.A2(n_92),
.B(n_91),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_109),
.A2(n_112),
.B1(n_110),
.B2(n_99),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_93),
.B(n_61),
.Y(n_139)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_98),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_110),
.A2(n_61),
.B1(n_42),
.B2(n_34),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_129),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_143),
.B(n_151),
.Y(n_191)
);

AOI32xp33_ASAP7_75t_L g144 ( 
.A1(n_136),
.A2(n_103),
.A3(n_89),
.B1(n_104),
.B2(n_94),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_144),
.A2(n_149),
.B(n_119),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_111),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_145),
.A2(n_140),
.B(n_17),
.Y(n_186)
);

AOI22x1_ASAP7_75t_SL g149 ( 
.A1(n_137),
.A2(n_111),
.B1(n_113),
.B2(n_114),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_129),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_131),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_153),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_120),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_156),
.C(n_161),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_106),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_101),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_122),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_167),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_174),
.C(n_161),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_129),
.Y(n_165)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_142),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_168),
.Y(n_178)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_116),
.Y(n_169)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_124),
.Y(n_170)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_125),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_172),
.A2(n_24),
.B1(n_25),
.B2(n_20),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_117),
.B(n_42),
.Y(n_173)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_117),
.B(n_57),
.C(n_34),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_170),
.Y(n_175)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_134),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_183),
.C(n_202),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_180),
.A2(n_184),
.B(n_185),
.Y(n_203)
);

AO22x2_ASAP7_75t_L g181 ( 
.A1(n_149),
.A2(n_134),
.B1(n_121),
.B2(n_141),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_181),
.A2(n_182),
.B1(n_192),
.B2(n_196),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_155),
.A2(n_134),
.B1(n_128),
.B2(n_121),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_171),
.A2(n_115),
.B(n_135),
.Y(n_184)
);

A2O1A1O1Ixp25_ASAP7_75t_L g185 ( 
.A1(n_164),
.A2(n_115),
.B(n_123),
.C(n_30),
.D(n_17),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_186),
.A2(n_181),
.B(n_195),
.Y(n_222)
);

AOI22x1_ASAP7_75t_L g188 ( 
.A1(n_145),
.A2(n_155),
.B1(n_156),
.B2(n_171),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_188),
.A2(n_158),
.B1(n_157),
.B2(n_147),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_148),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_193),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_22),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_146),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_150),
.A2(n_61),
.B1(n_25),
.B2(n_20),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_160),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_145),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_19),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_150),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_199)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_162),
.C(n_159),
.Y(n_202)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_205),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_191),
.Y(n_208)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_209),
.A2(n_221),
.B1(n_225),
.B2(n_181),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_178),
.Y(n_210)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_173),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_212),
.C(n_217),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_166),
.C(n_158),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_176),
.Y(n_213)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_197),
.Y(n_216)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_177),
.B(n_30),
.C(n_25),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_177),
.B(n_30),
.C(n_20),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_182),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_20),
.Y(n_219)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_175),
.Y(n_220)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_222),
.A2(n_19),
.B(n_4),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_187),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_223),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_188),
.Y(n_229)
);

INVx3_ASAP7_75t_SL g225 ( 
.A(n_181),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_229),
.C(n_240),
.Y(n_253)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_222),
.A2(n_185),
.B1(n_186),
.B2(n_192),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_231),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_196),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_238),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_203),
.A2(n_199),
.B(n_190),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_243),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_203),
.B(n_198),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_19),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_214),
.A2(n_219),
.B1(n_212),
.B2(n_216),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_245),
.Y(n_246)
);

BUFx12f_ASAP7_75t_SL g249 ( 
.A(n_238),
.Y(n_249)
);

OAI22x1_ASAP7_75t_L g271 ( 
.A1(n_249),
.A2(n_247),
.B1(n_229),
.B2(n_246),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_206),
.Y(n_252)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_252),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_205),
.Y(n_254)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_254),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_207),
.C(n_218),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_258),
.C(n_236),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_226),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_256),
.B(n_260),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_234),
.B(n_230),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_257),
.B(n_3),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_241),
.A2(n_225),
.B1(n_214),
.B2(n_220),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_204),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_232),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_209),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_243),
.Y(n_261)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_261),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_268),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_227),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_265),
.A2(n_270),
.B(n_262),
.Y(n_283)
);

AOI21x1_ASAP7_75t_SL g266 ( 
.A1(n_251),
.A2(n_231),
.B(n_215),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_266),
.A2(n_273),
.B1(n_6),
.B2(n_9),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_269),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_246),
.B(n_236),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_253),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_247),
.A2(n_215),
.B(n_217),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_272),
.A2(n_253),
.B(n_255),
.Y(n_275)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

MAJx2_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_11),
.C(n_12),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_4),
.C(n_5),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_277),
.C(n_282),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_6),
.C(n_8),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_283),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_265),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_280)
);

INVxp33_ASAP7_75t_L g289 ( 
.A(n_280),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_10),
.C(n_11),
.Y(n_282)
);

OAI21x1_ASAP7_75t_L g295 ( 
.A1(n_286),
.A2(n_293),
.B(n_13),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_281),
.Y(n_287)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_287),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_278),
.B(n_12),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_292),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_277),
.B(n_13),
.Y(n_292)
);

AOI21x1_ASAP7_75t_L g293 ( 
.A1(n_274),
.A2(n_282),
.B(n_276),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_287),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_298),
.Y(n_302)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_295),
.Y(n_300)
);

NOR4xp25_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_13),
.C(n_14),
.D(n_15),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_14),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_299),
.A2(n_288),
.B(n_289),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_301),
.B(n_297),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_302),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_304),
.A2(n_300),
.B(n_296),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_305),
.A2(n_14),
.B(n_15),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_15),
.Y(n_307)
);


endmodule