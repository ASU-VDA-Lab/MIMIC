module real_aes_7559_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_551;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_288;
wire n_147;
wire n_404;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_741;
wire n_314;
wire n_252;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g492 ( .A1(n_0), .A2(n_153), .B(n_493), .C(n_496), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_1), .B(n_488), .Y(n_497) );
INVx1_ASAP7_75t_L g442 ( .A(n_2), .Y(n_442) );
INVx1_ASAP7_75t_L g151 ( .A(n_3), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_4), .B(n_154), .Y(n_561) );
OAI22xp5_ASAP7_75t_SL g106 ( .A1(n_5), .A2(n_107), .B1(n_110), .B2(n_111), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_5), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_6), .A2(n_456), .B(n_532), .Y(n_531) );
AO21x2_ASAP7_75t_L g510 ( .A1(n_7), .A2(n_161), .B(n_511), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g207 ( .A1(n_8), .A2(n_38), .B1(n_141), .B2(n_189), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_9), .B(n_161), .Y(n_169) );
AND2x6_ASAP7_75t_L g156 ( .A(n_10), .B(n_157), .Y(n_156) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_11), .A2(n_156), .B(n_461), .C(n_505), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g107 ( .A1(n_12), .A2(n_42), .B1(n_108), .B2(n_109), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_12), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_13), .B(n_39), .Y(n_443) );
INVx1_ASAP7_75t_L g135 ( .A(n_14), .Y(n_135) );
INVx1_ASAP7_75t_L g132 ( .A(n_15), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_16), .B(n_137), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_17), .B(n_154), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_18), .B(n_128), .Y(n_235) );
AO32x2_ASAP7_75t_L g205 ( .A1(n_19), .A2(n_127), .A3(n_161), .B1(n_180), .B2(n_206), .Y(n_205) );
AOI222xp33_ASAP7_75t_SL g105 ( .A1(n_20), .A2(n_106), .B1(n_112), .B2(n_734), .C1(n_735), .C2(n_737), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_21), .B(n_141), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_22), .B(n_128), .Y(n_158) );
AOI22xp33_ASAP7_75t_L g208 ( .A1(n_23), .A2(n_57), .B1(n_141), .B2(n_189), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g765 ( .A(n_24), .Y(n_765) );
AOI22xp33_ASAP7_75t_SL g191 ( .A1(n_25), .A2(n_83), .B1(n_137), .B2(n_141), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_26), .B(n_141), .Y(n_221) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_27), .A2(n_180), .B(n_461), .C(n_479), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_28), .A2(n_180), .B(n_461), .C(n_514), .Y(n_513) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_29), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_30), .B(n_182), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_31), .A2(n_456), .B(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_32), .B(n_182), .Y(n_223) );
INVx2_ASAP7_75t_L g139 ( .A(n_33), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g458 ( .A1(n_34), .A2(n_459), .B(n_463), .C(n_469), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_35), .B(n_141), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_36), .B(n_182), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_37), .B(n_200), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_40), .B(n_477), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_41), .Y(n_509) );
INVx1_ASAP7_75t_L g109 ( .A(n_42), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_43), .B(n_154), .Y(n_526) );
OAI22xp5_ASAP7_75t_SL g755 ( .A1(n_44), .A2(n_756), .B1(n_758), .B2(n_759), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_44), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_45), .B(n_456), .Y(n_512) );
OAI22xp5_ASAP7_75t_SL g114 ( .A1(n_46), .A2(n_115), .B1(n_116), .B2(n_437), .Y(n_114) );
INVx1_ASAP7_75t_L g437 ( .A(n_46), .Y(n_437) );
OAI22xp5_ASAP7_75t_SL g756 ( .A1(n_46), .A2(n_48), .B1(n_437), .B2(n_757), .Y(n_756) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_47), .A2(n_459), .B(n_469), .C(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_48), .Y(n_757) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_49), .B(n_141), .Y(n_164) );
INVx1_ASAP7_75t_L g494 ( .A(n_50), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_51), .A2(n_91), .B1(n_189), .B2(n_190), .Y(n_188) );
INVx1_ASAP7_75t_L g525 ( .A(n_52), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_53), .B(n_141), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_54), .B(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_55), .B(n_456), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_56), .B(n_149), .Y(n_168) );
AOI22xp33_ASAP7_75t_SL g233 ( .A1(n_58), .A2(n_62), .B1(n_137), .B2(n_141), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_59), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_60), .B(n_141), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_61), .B(n_141), .Y(n_197) );
INVx1_ASAP7_75t_L g157 ( .A(n_63), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_64), .B(n_456), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_65), .B(n_488), .Y(n_537) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_66), .A2(n_143), .B(n_149), .C(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_67), .B(n_141), .Y(n_152) );
INVx1_ASAP7_75t_L g131 ( .A(n_68), .Y(n_131) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_69), .A2(n_104), .B1(n_741), .B2(n_750), .C1(n_766), .C2(n_772), .Y(n_103) );
OAI22xp33_ASAP7_75t_SL g752 ( .A1(n_69), .A2(n_753), .B1(n_760), .B2(n_761), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_69), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_70), .Y(n_746) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_71), .B(n_154), .Y(n_467) );
AO32x2_ASAP7_75t_L g186 ( .A1(n_72), .A2(n_161), .A3(n_180), .B1(n_187), .B2(n_192), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_73), .B(n_155), .Y(n_506) );
INVx1_ASAP7_75t_L g176 ( .A(n_74), .Y(n_176) );
INVx1_ASAP7_75t_L g218 ( .A(n_75), .Y(n_218) );
CKINVDCx16_ASAP7_75t_R g491 ( .A(n_76), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_77), .B(n_466), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g558 ( .A1(n_78), .A2(n_461), .B(n_469), .C(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_79), .B(n_137), .Y(n_219) );
CKINVDCx16_ASAP7_75t_R g533 ( .A(n_80), .Y(n_533) );
INVx1_ASAP7_75t_L g745 ( .A(n_81), .Y(n_745) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_82), .B(n_465), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_84), .B(n_189), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_85), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_86), .B(n_137), .Y(n_222) );
INVx2_ASAP7_75t_L g129 ( .A(n_87), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_88), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_89), .B(n_179), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_90), .B(n_137), .Y(n_165) );
OR2x2_ASAP7_75t_L g440 ( .A(n_92), .B(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g447 ( .A(n_92), .Y(n_447) );
OR2x2_ASAP7_75t_L g749 ( .A(n_92), .B(n_740), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_93), .A2(n_102), .B1(n_137), .B2(n_138), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_94), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g464 ( .A(n_95), .Y(n_464) );
INVxp67_ASAP7_75t_L g536 ( .A(n_96), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_97), .B(n_137), .Y(n_174) );
INVx1_ASAP7_75t_L g502 ( .A(n_98), .Y(n_502) );
INVx1_ASAP7_75t_L g560 ( .A(n_99), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_100), .B(n_745), .Y(n_744) );
AND2x2_ASAP7_75t_L g527 ( .A(n_101), .B(n_182), .Y(n_527) );
INVxp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g734 ( .A(n_106), .Y(n_734) );
CKINVDCx14_ASAP7_75t_R g110 ( .A(n_107), .Y(n_110) );
OAI22x1_ASAP7_75t_SL g112 ( .A1(n_113), .A2(n_438), .B1(n_444), .B2(n_448), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
OAI22xp5_ASAP7_75t_SL g735 ( .A1(n_114), .A2(n_438), .B1(n_446), .B2(n_736), .Y(n_735) );
OAI22xp5_ASAP7_75t_SL g753 ( .A1(n_115), .A2(n_116), .B1(n_754), .B2(n_755), .Y(n_753) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_SL g116 ( .A(n_117), .B(n_403), .Y(n_116) );
NOR3xp33_ASAP7_75t_L g117 ( .A(n_118), .B(n_307), .C(n_391), .Y(n_117) );
NAND4xp25_ASAP7_75t_L g118 ( .A(n_119), .B(n_250), .C(n_272), .D(n_288), .Y(n_118) );
AOI221xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_183), .B1(n_209), .B2(n_228), .C(n_236), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_159), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_122), .B(n_228), .Y(n_262) );
NAND4xp25_ASAP7_75t_L g302 ( .A(n_122), .B(n_290), .C(n_303), .D(n_305), .Y(n_302) );
INVxp67_ASAP7_75t_L g419 ( .A(n_122), .Y(n_419) );
INVx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g301 ( .A(n_123), .B(n_239), .Y(n_301) );
AND2x2_ASAP7_75t_L g325 ( .A(n_123), .B(n_159), .Y(n_325) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g292 ( .A(n_124), .B(n_227), .Y(n_292) );
AND2x2_ASAP7_75t_L g332 ( .A(n_124), .B(n_313), .Y(n_332) );
AND2x2_ASAP7_75t_L g349 ( .A(n_124), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_124), .B(n_160), .Y(n_373) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x2_ASAP7_75t_L g226 ( .A(n_125), .B(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g244 ( .A(n_125), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g256 ( .A(n_125), .B(n_160), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_125), .B(n_170), .Y(n_278) );
OA21x2_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_133), .B(n_158), .Y(n_125) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_126), .A2(n_171), .B(n_181), .Y(n_170) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_127), .B(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_128), .Y(n_161) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
AND2x2_ASAP7_75t_SL g182 ( .A(n_129), .B(n_130), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
OAI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_147), .B(n_156), .Y(n_133) );
O2A1O1Ixp33_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_136), .B(n_140), .C(n_143), .Y(n_134) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_136), .A2(n_506), .B(n_507), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_136), .A2(n_515), .B(n_516), .Y(n_514) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g142 ( .A(n_139), .Y(n_142) );
INVx1_ASAP7_75t_L g150 ( .A(n_139), .Y(n_150) );
INVx3_ASAP7_75t_L g217 ( .A(n_141), .Y(n_217) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_141), .Y(n_562) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g189 ( .A(n_142), .Y(n_189) );
BUFx3_ASAP7_75t_L g190 ( .A(n_142), .Y(n_190) );
AND2x6_ASAP7_75t_L g461 ( .A(n_142), .B(n_462), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_L g559 ( .A1(n_143), .A2(n_560), .B(n_561), .C(n_562), .Y(n_559) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_144), .A2(n_221), .B(n_222), .Y(n_220) );
INVx4_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g466 ( .A(n_145), .Y(n_466) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx3_ASAP7_75t_L g155 ( .A(n_146), .Y(n_155) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_146), .Y(n_179) );
INVx1_ASAP7_75t_L g200 ( .A(n_146), .Y(n_200) );
AND2x2_ASAP7_75t_L g457 ( .A(n_146), .B(n_150), .Y(n_457) );
INVx1_ASAP7_75t_L g462 ( .A(n_146), .Y(n_462) );
O2A1O1Ixp33_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_151), .B(n_152), .C(n_153), .Y(n_147) );
O2A1O1Ixp5_ASAP7_75t_L g175 ( .A1(n_148), .A2(n_176), .B(n_177), .C(n_178), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_148), .A2(n_480), .B(n_481), .Y(n_479) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_153), .A2(n_167), .B(n_168), .Y(n_166) );
OAI22xp5_ASAP7_75t_L g206 ( .A1(n_153), .A2(n_179), .B1(n_207), .B2(n_208), .Y(n_206) );
OAI22xp5_ASAP7_75t_L g231 ( .A1(n_153), .A2(n_179), .B1(n_232), .B2(n_233), .Y(n_231) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_154), .A2(n_164), .B(n_165), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_154), .A2(n_173), .B(n_174), .Y(n_172) );
O2A1O1Ixp5_ASAP7_75t_SL g216 ( .A1(n_154), .A2(n_217), .B(n_218), .C(n_219), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_154), .B(n_536), .Y(n_535) );
INVx5_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
OAI22xp5_ASAP7_75t_SL g187 ( .A1(n_155), .A2(n_179), .B1(n_188), .B2(n_191), .Y(n_187) );
OAI21xp5_ASAP7_75t_L g162 ( .A1(n_156), .A2(n_163), .B(n_166), .Y(n_162) );
BUFx3_ASAP7_75t_L g180 ( .A(n_156), .Y(n_180) );
OAI21xp5_ASAP7_75t_L g195 ( .A1(n_156), .A2(n_196), .B(n_201), .Y(n_195) );
OAI21xp5_ASAP7_75t_L g215 ( .A1(n_156), .A2(n_216), .B(n_220), .Y(n_215) );
AND2x4_ASAP7_75t_L g456 ( .A(n_156), .B(n_457), .Y(n_456) );
INVx4_ASAP7_75t_SL g470 ( .A(n_156), .Y(n_470) );
NAND2x1p5_ASAP7_75t_L g503 ( .A(n_156), .B(n_457), .Y(n_503) );
AND2x2_ASAP7_75t_L g259 ( .A(n_159), .B(n_260), .Y(n_259) );
AOI221xp5_ASAP7_75t_L g308 ( .A1(n_159), .A2(n_309), .B1(n_312), .B2(n_314), .C(n_318), .Y(n_308) );
AND2x2_ASAP7_75t_L g367 ( .A(n_159), .B(n_332), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_159), .B(n_349), .Y(n_401) );
AND2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_170), .Y(n_159) );
INVx3_ASAP7_75t_L g227 ( .A(n_160), .Y(n_227) );
AND2x2_ASAP7_75t_L g276 ( .A(n_160), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g330 ( .A(n_160), .B(n_245), .Y(n_330) );
AND2x2_ASAP7_75t_L g388 ( .A(n_160), .B(n_389), .Y(n_388) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_162), .B(n_169), .Y(n_160) );
INVx4_ASAP7_75t_L g230 ( .A(n_161), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_161), .A2(n_512), .B(n_513), .Y(n_511) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_161), .Y(n_530) );
AND2x2_ASAP7_75t_L g228 ( .A(n_170), .B(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g245 ( .A(n_170), .Y(n_245) );
INVx1_ASAP7_75t_L g300 ( .A(n_170), .Y(n_300) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_170), .Y(n_306) );
AND2x2_ASAP7_75t_L g351 ( .A(n_170), .B(n_227), .Y(n_351) );
OR2x2_ASAP7_75t_L g390 ( .A(n_170), .B(n_229), .Y(n_390) );
OAI21xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_175), .B(n_180), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_178), .A2(n_202), .B(n_203), .Y(n_201) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx4_ASAP7_75t_L g495 ( .A(n_179), .Y(n_495) );
NAND3xp33_ASAP7_75t_L g249 ( .A(n_180), .B(n_230), .C(n_231), .Y(n_249) );
INVx2_ASAP7_75t_L g192 ( .A(n_182), .Y(n_192) );
OA21x2_ASAP7_75t_L g194 ( .A1(n_182), .A2(n_195), .B(n_204), .Y(n_194) );
OA21x2_ASAP7_75t_L g214 ( .A1(n_182), .A2(n_215), .B(n_223), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_182), .A2(n_455), .B(n_458), .Y(n_454) );
INVx1_ASAP7_75t_L g485 ( .A(n_182), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_182), .A2(n_522), .B(n_523), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_183), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g183 ( .A(n_184), .B(n_193), .Y(n_183) );
AND2x2_ASAP7_75t_L g386 ( .A(n_184), .B(n_383), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_184), .B(n_368), .Y(n_418) );
BUFx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g317 ( .A(n_185), .B(n_241), .Y(n_317) );
AND2x2_ASAP7_75t_L g366 ( .A(n_185), .B(n_212), .Y(n_366) );
INVx1_ASAP7_75t_L g412 ( .A(n_185), .Y(n_412) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_186), .Y(n_225) );
AND2x2_ASAP7_75t_L g267 ( .A(n_186), .B(n_241), .Y(n_267) );
INVx1_ASAP7_75t_L g284 ( .A(n_186), .Y(n_284) );
AND2x2_ASAP7_75t_L g290 ( .A(n_186), .B(n_205), .Y(n_290) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_190), .Y(n_468) );
INVx2_ASAP7_75t_L g496 ( .A(n_190), .Y(n_496) );
INVx1_ASAP7_75t_L g482 ( .A(n_192), .Y(n_482) );
AND2x2_ASAP7_75t_L g358 ( .A(n_193), .B(n_266), .Y(n_358) );
INVx2_ASAP7_75t_L g423 ( .A(n_193), .Y(n_423) );
AND2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_205), .Y(n_193) );
AND2x2_ASAP7_75t_L g240 ( .A(n_194), .B(n_241), .Y(n_240) );
OR2x2_ASAP7_75t_L g253 ( .A(n_194), .B(n_213), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_194), .B(n_212), .Y(n_281) );
INVx1_ASAP7_75t_L g287 ( .A(n_194), .Y(n_287) );
INVx1_ASAP7_75t_L g304 ( .A(n_194), .Y(n_304) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_194), .Y(n_316) );
INVx2_ASAP7_75t_L g384 ( .A(n_194), .Y(n_384) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_199), .Y(n_196) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g241 ( .A(n_205), .Y(n_241) );
BUFx2_ASAP7_75t_L g338 ( .A(n_205), .Y(n_338) );
AND2x2_ASAP7_75t_L g383 ( .A(n_205), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_211), .B(n_224), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_211), .B(n_320), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g406 ( .A1(n_211), .A2(n_382), .B(n_396), .Y(n_406) );
AND2x2_ASAP7_75t_L g431 ( .A(n_211), .B(n_317), .Y(n_431) );
BUFx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g353 ( .A(n_213), .Y(n_353) );
AND2x2_ASAP7_75t_L g382 ( .A(n_213), .B(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_214), .Y(n_266) );
INVx2_ASAP7_75t_L g285 ( .A(n_214), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_214), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_226), .Y(n_224) );
INVx2_ASAP7_75t_L g239 ( .A(n_225), .Y(n_239) );
OR2x2_ASAP7_75t_L g252 ( .A(n_225), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g320 ( .A(n_225), .B(n_316), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_225), .B(n_416), .Y(n_415) );
OR2x2_ASAP7_75t_L g421 ( .A(n_225), .B(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_225), .B(n_358), .Y(n_433) );
AND2x2_ASAP7_75t_L g312 ( .A(n_226), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g335 ( .A(n_226), .B(n_228), .Y(n_335) );
INVx2_ASAP7_75t_L g247 ( .A(n_227), .Y(n_247) );
AND2x2_ASAP7_75t_L g275 ( .A(n_227), .B(n_248), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_227), .B(n_300), .Y(n_356) );
AND2x2_ASAP7_75t_L g270 ( .A(n_228), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g417 ( .A(n_228), .Y(n_417) );
AND2x2_ASAP7_75t_L g429 ( .A(n_228), .B(n_292), .Y(n_429) );
AND2x2_ASAP7_75t_L g255 ( .A(n_229), .B(n_245), .Y(n_255) );
INVx1_ASAP7_75t_L g350 ( .A(n_229), .Y(n_350) );
AO21x1_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_234), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_230), .B(n_472), .Y(n_471) );
INVx3_ASAP7_75t_L g488 ( .A(n_230), .Y(n_488) );
AO21x2_ASAP7_75t_L g500 ( .A1(n_230), .A2(n_501), .B(n_508), .Y(n_500) );
AO21x2_ASAP7_75t_L g556 ( .A1(n_230), .A2(n_557), .B(n_564), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_230), .B(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x4_ASAP7_75t_L g248 ( .A(n_235), .B(n_249), .Y(n_248) );
INVxp67_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_242), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_239), .B(n_286), .Y(n_295) );
OR2x2_ASAP7_75t_L g427 ( .A(n_239), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g344 ( .A(n_240), .B(n_285), .Y(n_344) );
AND2x2_ASAP7_75t_L g352 ( .A(n_240), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g411 ( .A(n_240), .B(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g435 ( .A(n_240), .B(n_282), .Y(n_435) );
NOR2xp67_ASAP7_75t_L g393 ( .A(n_241), .B(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g422 ( .A(n_241), .B(n_285), .Y(n_422) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2x1p5_ASAP7_75t_L g243 ( .A(n_244), .B(n_246), .Y(n_243) );
AND2x2_ASAP7_75t_L g274 ( .A(n_244), .B(n_275), .Y(n_274) );
INVxp67_ASAP7_75t_L g436 ( .A(n_244), .Y(n_436) );
NOR2x1_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
INVx1_ASAP7_75t_L g271 ( .A(n_247), .Y(n_271) );
AND2x2_ASAP7_75t_L g322 ( .A(n_247), .B(n_255), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_247), .B(n_390), .Y(n_416) );
INVx2_ASAP7_75t_L g261 ( .A(n_248), .Y(n_261) );
INVx3_ASAP7_75t_L g313 ( .A(n_248), .Y(n_313) );
OR2x2_ASAP7_75t_L g341 ( .A(n_248), .B(n_342), .Y(n_341) );
AOI311xp33_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_254), .A3(n_256), .B(n_257), .C(n_268), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_L g288 ( .A1(n_251), .A2(n_289), .B(n_291), .C(n_293), .Y(n_288) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx2_ASAP7_75t_SL g273 ( .A(n_253), .Y(n_273) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g291 ( .A(n_255), .B(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_255), .B(n_271), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_255), .B(n_256), .Y(n_424) );
AND2x2_ASAP7_75t_L g346 ( .A(n_256), .B(n_260), .Y(n_346) );
AOI21xp33_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_262), .B(n_263), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g404 ( .A(n_260), .B(n_292), .Y(n_404) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_261), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g298 ( .A(n_261), .Y(n_298) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_267), .Y(n_264) );
AND2x2_ASAP7_75t_L g289 ( .A(n_265), .B(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g334 ( .A(n_267), .Y(n_334) );
AND2x4_ASAP7_75t_L g396 ( .A(n_267), .B(n_365), .Y(n_396) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AOI222xp33_ASAP7_75t_L g347 ( .A1(n_270), .A2(n_336), .B1(n_348), .B2(n_352), .C1(n_354), .C2(n_358), .Y(n_347) );
A2O1A1Ixp33_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_274), .B(n_276), .C(n_279), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_273), .B(n_317), .Y(n_340) );
INVx1_ASAP7_75t_L g362 ( .A(n_275), .Y(n_362) );
INVx1_ASAP7_75t_L g296 ( .A(n_277), .Y(n_296) );
OR2x2_ASAP7_75t_L g361 ( .A(n_278), .B(n_362), .Y(n_361) );
OAI21xp33_ASAP7_75t_SL g279 ( .A1(n_280), .A2(n_282), .B(n_286), .Y(n_279) );
NAND3xp33_ASAP7_75t_L g297 ( .A(n_280), .B(n_298), .C(n_299), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g395 ( .A1(n_280), .A2(n_317), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_284), .Y(n_337) );
AND2x2_ASAP7_75t_SL g303 ( .A(n_285), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g394 ( .A(n_285), .Y(n_394) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_285), .Y(n_410) );
INVx2_ASAP7_75t_L g368 ( .A(n_286), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_290), .B(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g342 ( .A(n_292), .Y(n_342) );
OAI221xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_296), .B1(n_297), .B2(n_301), .C(n_302), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_SL g375 ( .A(n_296), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_SL g430 ( .A(n_296), .Y(n_430) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g311 ( .A(n_303), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_303), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g369 ( .A(n_303), .B(n_317), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_303), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g402 ( .A(n_303), .B(n_337), .Y(n_402) );
BUFx3_ASAP7_75t_L g365 ( .A(n_304), .Y(n_365) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND5xp2_ASAP7_75t_L g307 ( .A(n_308), .B(n_326), .C(n_347), .D(n_359), .E(n_374), .Y(n_307) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AOI32xp33_ASAP7_75t_L g399 ( .A1(n_311), .A2(n_338), .A3(n_354), .B1(n_400), .B2(n_402), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_313), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_SL g323 ( .A(n_317), .Y(n_323) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_321), .B1(n_323), .B2(n_324), .Y(n_318) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
AOI221xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_333), .B1(n_335), .B2(n_336), .C(n_339), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_331), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g398 ( .A(n_330), .B(n_349), .Y(n_398) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AOI221xp5_ASAP7_75t_L g413 ( .A1(n_335), .A2(n_396), .B1(n_414), .B2(n_419), .C(n_420), .Y(n_413) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx2_ASAP7_75t_L g379 ( .A(n_338), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_341), .B1(n_343), .B2(n_345), .Y(n_339) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_351), .Y(n_348) );
INVx1_ASAP7_75t_L g357 ( .A(n_349), .Y(n_357) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
AOI222xp33_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_363), .B1(n_367), .B2(n_368), .C1(n_369), .C2(n_370), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_366), .Y(n_363) );
INVxp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OAI22xp33_ASAP7_75t_L g414 ( .A1(n_368), .A2(n_415), .B1(n_417), .B2(n_418), .Y(n_414) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
AOI21xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_377), .B(n_380), .Y(n_374) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AOI21xp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_385), .B(n_387), .Y(n_380) );
INVx2_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g428 ( .A(n_383), .Y(n_428) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
A2O1A1Ixp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_395), .B(n_397), .C(n_399), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AOI211xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B(n_407), .C(n_432), .Y(n_403) );
CKINVDCx16_ASAP7_75t_R g408 ( .A(n_404), .Y(n_408) );
INVxp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OAI211xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_409), .B(n_413), .C(n_425), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
AOI21xp33_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_423), .B(n_424), .Y(n_420) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_429), .B1(n_430), .B2(n_431), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AOI21xp33_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_434), .B(n_436), .Y(n_432) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OR2x2_ASAP7_75t_L g446 ( .A(n_441), .B(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g740 ( .A(n_441), .Y(n_740) );
AND2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NOR2x2_ASAP7_75t_L g739 ( .A(n_447), .B(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g736 ( .A(n_448), .Y(n_736) );
OR3x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_648), .C(n_691), .Y(n_448) );
NAND5xp2_ASAP7_75t_L g449 ( .A(n_450), .B(n_575), .C(n_605), .D(n_622), .E(n_637), .Y(n_449) );
AOI221xp5_ASAP7_75t_SL g450 ( .A1(n_451), .A2(n_498), .B1(n_538), .B2(n_544), .C(n_548), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_473), .Y(n_451) );
OR2x2_ASAP7_75t_L g553 ( .A(n_452), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g592 ( .A(n_452), .B(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g610 ( .A(n_452), .B(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_452), .B(n_546), .Y(n_627) );
OR2x2_ASAP7_75t_L g639 ( .A(n_452), .B(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_452), .B(n_598), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_452), .B(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_452), .B(n_576), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_452), .B(n_584), .Y(n_690) );
AND2x2_ASAP7_75t_L g722 ( .A(n_452), .B(n_486), .Y(n_722) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_452), .Y(n_730) );
INVx5_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_453), .B(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g550 ( .A(n_453), .B(n_528), .Y(n_550) );
BUFx2_ASAP7_75t_L g572 ( .A(n_453), .Y(n_572) );
AND2x2_ASAP7_75t_L g601 ( .A(n_453), .B(n_474), .Y(n_601) );
AND2x2_ASAP7_75t_L g656 ( .A(n_453), .B(n_554), .Y(n_656) );
OR2x6_ASAP7_75t_L g453 ( .A(n_454), .B(n_471), .Y(n_453) );
BUFx2_ASAP7_75t_L g477 ( .A(n_456), .Y(n_477) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
O2A1O1Ixp33_ASAP7_75t_SL g490 ( .A1(n_460), .A2(n_470), .B(n_491), .C(n_492), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_L g532 ( .A1(n_460), .A2(n_470), .B(n_533), .C(n_534), .Y(n_532) );
INVx5_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
O2A1O1Ixp33_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B(n_467), .C(n_468), .Y(n_463) );
O2A1O1Ixp33_ASAP7_75t_L g524 ( .A1(n_465), .A2(n_468), .B(n_525), .C(n_526), .Y(n_524) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_473), .B(n_610), .Y(n_619) );
OAI32xp33_ASAP7_75t_L g633 ( .A1(n_473), .A2(n_569), .A3(n_634), .B1(n_635), .B2(n_636), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_473), .B(n_635), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_473), .B(n_553), .Y(n_676) );
INVx1_ASAP7_75t_SL g705 ( .A(n_473), .Y(n_705) );
NAND4xp25_ASAP7_75t_L g714 ( .A(n_473), .B(n_500), .C(n_656), .D(n_715), .Y(n_714) );
AND2x4_ASAP7_75t_L g473 ( .A(n_474), .B(n_486), .Y(n_473) );
INVx5_ASAP7_75t_L g547 ( .A(n_474), .Y(n_547) );
AND2x2_ASAP7_75t_L g576 ( .A(n_474), .B(n_487), .Y(n_576) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_474), .Y(n_655) );
AND2x2_ASAP7_75t_L g725 ( .A(n_474), .B(n_672), .Y(n_725) );
OR2x6_ASAP7_75t_L g474 ( .A(n_475), .B(n_483), .Y(n_474) );
AOI21xp5_ASAP7_75t_SL g475 ( .A1(n_476), .A2(n_478), .B(n_482), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
AND2x4_ASAP7_75t_L g598 ( .A(n_486), .B(n_547), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_486), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g632 ( .A(n_486), .B(n_554), .Y(n_632) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g546 ( .A(n_487), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g584 ( .A(n_487), .B(n_556), .Y(n_584) );
AND2x2_ASAP7_75t_L g593 ( .A(n_487), .B(n_555), .Y(n_593) );
OA21x2_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_489), .B(n_497), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
AOI222xp33_ASAP7_75t_L g661 ( .A1(n_498), .A2(n_662), .B1(n_664), .B2(n_666), .C1(n_669), .C2(n_670), .Y(n_661) );
AND2x4_ASAP7_75t_L g498 ( .A(n_499), .B(n_517), .Y(n_498) );
AND2x2_ASAP7_75t_L g594 ( .A(n_499), .B(n_595), .Y(n_594) );
NAND3xp33_ASAP7_75t_L g711 ( .A(n_499), .B(n_572), .C(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_510), .Y(n_499) );
INVx5_ASAP7_75t_SL g543 ( .A(n_500), .Y(n_543) );
OAI322xp33_ASAP7_75t_L g548 ( .A1(n_500), .A2(n_549), .A3(n_551), .B1(n_552), .B2(n_566), .C1(n_569), .C2(n_571), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_500), .B(n_541), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_500), .B(n_529), .Y(n_720) );
OAI21xp5_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_503), .B(n_504), .Y(n_501) );
INVx2_ASAP7_75t_L g541 ( .A(n_510), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_510), .B(n_519), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_517), .B(n_579), .Y(n_634) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
OR2x2_ASAP7_75t_L g613 ( .A(n_518), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_528), .Y(n_518) );
OR2x2_ASAP7_75t_L g542 ( .A(n_519), .B(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_519), .B(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g581 ( .A(n_519), .B(n_529), .Y(n_581) );
AND2x2_ASAP7_75t_L g604 ( .A(n_519), .B(n_541), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_519), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g620 ( .A(n_519), .B(n_579), .Y(n_620) );
AND2x2_ASAP7_75t_L g628 ( .A(n_519), .B(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_519), .B(n_588), .Y(n_678) );
INVx5_ASAP7_75t_SL g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g568 ( .A(n_520), .B(n_543), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_520), .B(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g595 ( .A(n_520), .B(n_529), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_520), .B(n_642), .Y(n_683) );
OR2x2_ASAP7_75t_L g699 ( .A(n_520), .B(n_643), .Y(n_699) );
AND2x2_ASAP7_75t_SL g706 ( .A(n_520), .B(n_660), .Y(n_706) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_520), .Y(n_713) );
OR2x6_ASAP7_75t_L g520 ( .A(n_521), .B(n_527), .Y(n_520) );
AND2x2_ASAP7_75t_L g567 ( .A(n_528), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g617 ( .A(n_528), .B(n_541), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_528), .B(n_543), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_528), .B(n_579), .Y(n_701) );
INVx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_529), .B(n_543), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_529), .B(n_541), .Y(n_589) );
OR2x2_ASAP7_75t_L g643 ( .A(n_529), .B(n_541), .Y(n_643) );
AND2x2_ASAP7_75t_L g660 ( .A(n_529), .B(n_540), .Y(n_660) );
INVxp67_ASAP7_75t_L g682 ( .A(n_529), .Y(n_682) );
AND2x2_ASAP7_75t_L g709 ( .A(n_529), .B(n_579), .Y(n_709) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_529), .Y(n_716) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B(n_537), .Y(n_529) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_542), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_540), .B(n_590), .Y(n_663) );
INVx1_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g579 ( .A(n_541), .B(n_543), .Y(n_579) );
OR2x2_ASAP7_75t_L g646 ( .A(n_541), .B(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g590 ( .A(n_542), .Y(n_590) );
OR2x2_ASAP7_75t_L g651 ( .A(n_542), .B(n_643), .Y(n_651) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g551 ( .A(n_546), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_546), .B(n_610), .Y(n_609) );
OR2x2_ASAP7_75t_L g552 ( .A(n_547), .B(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_547), .B(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_547), .B(n_554), .Y(n_586) );
INVx2_ASAP7_75t_L g631 ( .A(n_547), .Y(n_631) );
AND2x2_ASAP7_75t_L g644 ( .A(n_547), .B(n_584), .Y(n_644) );
AND2x2_ASAP7_75t_L g669 ( .A(n_547), .B(n_593), .Y(n_669) );
INVx1_ASAP7_75t_L g621 ( .A(n_552), .Y(n_621) );
INVx2_ASAP7_75t_SL g608 ( .A(n_553), .Y(n_608) );
INVx1_ASAP7_75t_L g611 ( .A(n_554), .Y(n_611) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_555), .Y(n_574) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
BUFx2_ASAP7_75t_L g672 ( .A(n_556), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_563), .Y(n_557) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g641 ( .A(n_568), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g647 ( .A(n_568), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_568), .A2(n_650), .B1(n_652), .B2(n_657), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_568), .B(n_660), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_569), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_SL g603 ( .A(n_570), .Y(n_603) );
OR2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
OR2x2_ASAP7_75t_L g585 ( .A(n_572), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_572), .B(n_576), .Y(n_636) );
AND2x2_ASAP7_75t_L g659 ( .A(n_572), .B(n_660), .Y(n_659) );
BUFx2_ASAP7_75t_L g635 ( .A(n_574), .Y(n_635) );
AOI211xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_577), .B(n_582), .C(n_596), .Y(n_575) );
INVx1_ASAP7_75t_L g599 ( .A(n_576), .Y(n_599) );
OAI221xp5_ASAP7_75t_SL g707 ( .A1(n_576), .A2(n_708), .B1(n_710), .B2(n_711), .C(n_714), .Y(n_707) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
INVx1_ASAP7_75t_L g726 ( .A(n_579), .Y(n_726) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g675 ( .A(n_581), .B(n_614), .Y(n_675) );
A2O1A1Ixp33_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_585), .B(n_587), .C(n_591), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
INVx1_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
OAI32xp33_ASAP7_75t_L g700 ( .A1(n_589), .A2(n_590), .A3(n_653), .B1(n_690), .B2(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_594), .Y(n_591) );
AND2x2_ASAP7_75t_L g732 ( .A(n_592), .B(n_631), .Y(n_732) );
AND2x2_ASAP7_75t_L g679 ( .A(n_593), .B(n_631), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_593), .B(n_601), .Y(n_697) );
AOI31xp33_ASAP7_75t_SL g596 ( .A1(n_597), .A2(n_599), .A3(n_600), .B(n_602), .Y(n_596) );
INVxp67_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_598), .B(n_610), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_598), .B(n_608), .Y(n_695) );
AOI221xp5_ASAP7_75t_L g717 ( .A1(n_598), .A2(n_628), .B1(n_718), .B2(n_721), .C(n_723), .Y(n_717) );
CKINVDCx16_ASAP7_75t_R g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
AND2x2_ASAP7_75t_L g623 ( .A(n_603), .B(n_624), .Y(n_623) );
AOI222xp33_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_612), .B1(n_615), .B2(n_618), .C1(n_620), .C2(n_621), .Y(n_605) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_607), .B(n_609), .Y(n_606) );
INVx1_ASAP7_75t_L g688 ( .A(n_607), .Y(n_688) );
INVx1_ASAP7_75t_L g710 ( .A(n_610), .Y(n_710) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_613), .A2(n_724), .B1(n_726), .B2(n_727), .Y(n_723) );
INVx1_ASAP7_75t_L g629 ( .A(n_614), .Y(n_629) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_626), .B1(n_628), .B2(n_630), .C(n_633), .Y(n_622) );
INVx1_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
OR2x2_ASAP7_75t_L g667 ( .A(n_625), .B(n_668), .Y(n_667) );
OR2x2_ASAP7_75t_L g719 ( .A(n_625), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g694 ( .A(n_630), .Y(n_694) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
INVx1_ASAP7_75t_L g658 ( .A(n_631), .Y(n_658) );
INVx1_ASAP7_75t_L g640 ( .A(n_632), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_635), .B(n_722), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_641), .B1(n_644), .B2(n_645), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_SL g731 ( .A(n_644), .Y(n_731) );
INVxp33_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_646), .B(n_690), .Y(n_689) );
OAI32xp33_ASAP7_75t_L g680 ( .A1(n_647), .A2(n_681), .A3(n_682), .B1(n_683), .B2(n_684), .Y(n_680) );
NAND4xp25_ASAP7_75t_L g648 ( .A(n_649), .B(n_661), .C(n_673), .D(n_685), .Y(n_648) );
INVx1_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
NAND2xp33_ASAP7_75t_SL g652 ( .A(n_653), .B(n_654), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_656), .B(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
CKINVDCx16_ASAP7_75t_R g666 ( .A(n_667), .Y(n_666) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_670), .A2(n_686), .B1(n_703), .B2(n_706), .C(n_707), .Y(n_702) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g721 ( .A(n_672), .B(n_722), .Y(n_721) );
AOI221xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_676), .B1(n_677), .B2(n_679), .C(n_680), .Y(n_673) );
INVx1_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_682), .B(n_713), .Y(n_712) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_688), .B(n_689), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND4xp25_ASAP7_75t_L g691 ( .A(n_692), .B(n_702), .C(n_717), .D(n_728), .Y(n_691) );
O2A1O1Ixp33_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_696), .B(n_698), .C(n_700), .Y(n_692) );
NAND2xp5_ASAP7_75t_SL g693 ( .A(n_694), .B(n_695), .Y(n_693) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVxp67_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g733 ( .A(n_720), .Y(n_733) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
OAI21xp5_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_732), .B(n_733), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
NAND2xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_747), .Y(n_742) );
NOR2xp33_ASAP7_75t_SL g743 ( .A(n_744), .B(n_746), .Y(n_743) );
INVx1_ASAP7_75t_SL g771 ( .A(n_744), .Y(n_771) );
INVx1_ASAP7_75t_L g770 ( .A(n_746), .Y(n_770) );
OA21x2_ASAP7_75t_L g773 ( .A1(n_746), .A2(n_771), .B(n_774), .Y(n_773) );
INVx1_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
HB1xp67_ASAP7_75t_L g762 ( .A(n_749), .Y(n_762) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_749), .Y(n_764) );
BUFx2_ASAP7_75t_L g774 ( .A(n_749), .Y(n_774) );
INVxp67_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
AOI21xp5_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_762), .B(n_763), .Y(n_751) );
INVx1_ASAP7_75t_L g761 ( .A(n_753), .Y(n_761) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_756), .Y(n_759) );
NOR2xp33_ASAP7_75t_SL g763 ( .A(n_764), .B(n_765), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g766 ( .A(n_767), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_768), .Y(n_767) );
AND2x2_ASAP7_75t_L g768 ( .A(n_769), .B(n_771), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_773), .Y(n_772) );
endmodule