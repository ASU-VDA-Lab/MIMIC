module real_jpeg_25746_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_347, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_347;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_1),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_55)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_60),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_60),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_1),
.A2(n_41),
.B1(n_43),
.B2(n_60),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_2),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_2),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_2),
.A2(n_41),
.B1(n_43),
.B2(n_70),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_70),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_70),
.Y(n_278)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_5),
.A2(n_41),
.B1(n_43),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_5),
.A2(n_50),
.B1(n_57),
.B2(n_66),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_50),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_50),
.Y(n_117)
);

INVx8_ASAP7_75t_SL g64 ( 
.A(n_6),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_7),
.A2(n_36),
.B1(n_41),
.B2(n_43),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_7),
.A2(n_36),
.B1(n_58),
.B2(n_59),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_8),
.A2(n_41),
.B1(n_43),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_8),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_8),
.A2(n_58),
.B1(n_59),
.B2(n_127),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_127),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_127),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_9),
.A2(n_41),
.B1(n_43),
.B2(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_9),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_129),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_129),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_9),
.A2(n_58),
.B1(n_59),
.B2(n_129),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_10),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_10),
.B(n_68),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_10),
.B(n_28),
.C(n_32),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_132),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_10),
.B(n_44),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_10),
.A2(n_106),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_12),
.A2(n_71),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_12),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_12),
.A2(n_41),
.B1(n_43),
.B2(n_136),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_136),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_136),
.Y(n_208)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_15),
.Y(n_107)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_15),
.Y(n_150)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_15),
.Y(n_201)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_15),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_96),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_94),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_83),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_19),
.B(n_83),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_74),
.C(n_77),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_20),
.A2(n_74),
.B1(n_331),
.B2(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_20),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_53),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_37),
.B2(n_38),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_22),
.B(n_74),
.C(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_22),
.A2(n_23),
.B1(n_78),
.B2(n_79),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_23),
.B(n_37),
.C(n_53),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_31),
.B(n_34),
.Y(n_23)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_24),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_24),
.A2(n_34),
.B(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_24),
.A2(n_31),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_24),
.A2(n_31),
.B1(n_182),
.B2(n_189),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_24),
.A2(n_248),
.B(n_249),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_24),
.A2(n_31),
.B1(n_115),
.B2(n_278),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_24),
.A2(n_123),
.B(n_278),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_26),
.A2(n_27),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

NAND3xp33_ASAP7_75t_L g227 ( 
.A(n_26),
.B(n_41),
.C(n_47),
.Y(n_227)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_27),
.B(n_178),
.Y(n_177)
);

A2O1A1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_27),
.A2(n_46),
.B(n_226),
.C(n_227),
.Y(n_225)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_31),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_31),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_31),
.B(n_132),
.Y(n_217)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_32),
.B(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_33),
.B(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_35),
.B(n_124),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_48),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_39),
.A2(n_81),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_44),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_40),
.A2(n_44),
.B(n_51),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_40),
.Y(n_271)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_43),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_41),
.A2(n_63),
.B(n_131),
.C(n_152),
.Y(n_151)
);

HAxp5_ASAP7_75t_SL g226 ( 
.A(n_41),
.B(n_132),
.CON(n_226),
.SN(n_226)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND3xp33_ASAP7_75t_L g152 ( 
.A(n_43),
.B(n_57),
.C(n_64),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_44),
.B(n_49),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_44),
.A2(n_51),
.B1(n_126),
.B2(n_128),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_44),
.A2(n_51),
.B1(n_162),
.B2(n_226),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_44),
.A2(n_51),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_45),
.A2(n_81),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_45),
.A2(n_48),
.B(n_301),
.Y(n_300)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_51),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_51),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_61),
.B1(n_68),
.B2(n_69),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_62),
.B(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

HAxp5_ASAP7_75t_SL g131 ( 
.A(n_57),
.B(n_132),
.CON(n_131),
.SN(n_131)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_59),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_65)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_59),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_61),
.A2(n_69),
.B(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_61),
.A2(n_68),
.B1(n_131),
.B2(n_133),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_61),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_61),
.A2(n_68),
.B1(n_143),
.B2(n_268),
.Y(n_267)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_62),
.A2(n_134),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_68),
.B(n_76),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_68),
.B(n_299),
.Y(n_298)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_74),
.A2(n_331),
.B1(n_332),
.B2(n_333),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_74),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_77),
.B(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B(n_82),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_80),
.Y(n_324)
);

OAI21xp33_ASAP7_75t_L g270 ( 
.A1(n_81),
.A2(n_82),
.B(n_271),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_92),
.B2(n_93),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_90),
.B2(n_91),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_86),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_87),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_89),
.A2(n_141),
.B(n_317),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI321xp33_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_328),
.A3(n_339),
.B1(n_344),
.B2(n_345),
.C(n_347),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_306),
.B(n_327),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_283),
.B(n_305),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_170),
.B(n_259),
.C(n_282),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_154),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_101),
.B(n_154),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_137),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_119),
.B2(n_120),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_103),
.B(n_120),
.C(n_137),
.Y(n_260)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_114),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_105),
.B(n_114),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_108),
.B(n_109),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_106),
.A2(n_108),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_106),
.B(n_113),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_106),
.A2(n_191),
.B(n_192),
.Y(n_190)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_106),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_106),
.A2(n_150),
.B1(n_199),
.B2(n_208),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_106),
.A2(n_107),
.B(n_290),
.Y(n_289)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_107),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_110),
.A2(n_193),
.B(n_197),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_113),
.Y(n_110)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_111),
.Y(n_168)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_116),
.B(n_249),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_117),
.B(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_118),
.A2(n_124),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.C(n_130),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_121),
.A2(n_122),
.B1(n_125),
.B2(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_126),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_128),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_130),
.B(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_132),
.B(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_146),
.B2(n_153),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_144),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_140),
.B(n_144),
.C(n_153),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_141),
.A2(n_297),
.B(n_298),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_146),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_151),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_149),
.A2(n_168),
.B(n_169),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.C(n_159),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_155),
.B(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_158),
.B(n_159),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.C(n_166),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_160),
.B(n_243),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_243)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_169),
.B(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_258),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_253),
.B(n_257),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_238),
.B(n_252),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_222),
.B(n_237),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_194),
.B(n_221),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_183),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_176),
.B(n_183),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_177),
.A2(n_179),
.B1(n_180),
.B2(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_177),
.Y(n_204)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_190),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_185),
.B(n_188),
.C(n_190),
.Y(n_236)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_189),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_191),
.Y(n_202)
);

INVxp33_ASAP7_75t_L g275 ( 
.A(n_192),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_193),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_205),
.B(n_220),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_203),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_203),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_200),
.B2(n_202),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_216),
.B(n_219),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_212),
.Y(n_206)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_217),
.B(n_218),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_236),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_236),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_231),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_232),
.C(n_235),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_224)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_225),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_230),
.Y(n_246)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_228),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_235),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_234),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_239),
.B(n_240),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_244),
.B2(n_245),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_247),
.C(n_250),
.Y(n_256)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_250),
.B2(n_251),
.Y(n_245)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_246),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_247),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_256),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_261),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_281),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_272),
.B1(n_279),
.B2(n_280),
.Y(n_262)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_263),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_264),
.B(n_267),
.C(n_269),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_269),
.B2(n_270),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_268),
.Y(n_297)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_272),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_279),
.C(n_281),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_276),
.B2(n_277),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_273),
.B(n_277),
.Y(n_302)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_284),
.B(n_285),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_304),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_293),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_293),
.C(n_304),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_291),
.B2(n_292),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_288),
.A2(n_289),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_288),
.A2(n_312),
.B(n_316),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_291),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_291),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_302),
.B2(n_303),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_300),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_296),
.B(n_300),
.C(n_303),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_299),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_301),
.Y(n_323)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_302),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_307),
.B(n_308),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_326),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_310),
.A2(n_311),
.B1(n_319),
.B2(n_320),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_311),
.B(n_319),
.C(n_326),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_313),
.B1(n_314),
.B2(n_318),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_314),
.Y(n_318)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_321),
.A2(n_322),
.B(n_325),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_322),
.Y(n_325)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_325),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_325),
.A2(n_330),
.B1(n_334),
.B2(n_343),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_336),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_329),
.B(n_336),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_334),
.C(n_335),
.Y(n_329)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_330),
.Y(n_343)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_332),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_335),
.B(n_342),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_340),
.B(n_341),
.Y(n_344)
);


endmodule