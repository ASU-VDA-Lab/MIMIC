module fake_jpeg_28343_n_8 (n_3, n_2, n_1, n_0, n_4, n_8);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_8;

wire n_6;
wire n_5;
wire n_7;

XOR2xp5_ASAP7_75t_L g5 ( 
.A(n_1),
.B(n_0),
.Y(n_5)
);

OA22x2_ASAP7_75t_L g6 ( 
.A1(n_2),
.A2(n_4),
.B1(n_3),
.B2(n_1),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

AOI31xp33_ASAP7_75t_L g8 ( 
.A1(n_6),
.A2(n_5),
.A3(n_7),
.B(n_0),
.Y(n_8)
);


endmodule