module fake_netlist_6_3130_n_163 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_25, n_163);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_25;

output n_163;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_144;
wire n_127;
wire n_125;
wire n_153;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_130;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_108;
wire n_94;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_139;
wire n_41;
wire n_134;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_35;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_24),
.Y(n_34)
);

INVxp67_ASAP7_75t_SL g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_25),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_28),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_23),
.B(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_46),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_32),
.A2(n_0),
.B1(n_4),
.B2(n_6),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_0),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_47),
.B(n_27),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_46),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_33),
.B(n_6),
.Y(n_61)
);

AOI21x1_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_7),
.B(n_8),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_8),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_38),
.B(n_9),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

OR2x6_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_15),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_71)
);

AND2x4_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_19),
.Y(n_72)
);

AND2x4_ASAP7_75t_L g73 ( 
.A(n_37),
.B(n_26),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_43),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_69),
.A2(n_35),
.B(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_41),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_36),
.B(n_52),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_49),
.B(n_17),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_20),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_73),
.B(n_72),
.Y(n_82)
);

NOR3xp33_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_11),
.C(n_12),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

OAI321xp33_ASAP7_75t_L g86 ( 
.A1(n_57),
.A2(n_13),
.A3(n_14),
.B1(n_22),
.B2(n_61),
.C(n_62),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

AOI221x1_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_57),
.B1(n_61),
.B2(n_73),
.C(n_66),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

OR2x6_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_67),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_74),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_73),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g95 ( 
.A1(n_84),
.A2(n_56),
.B(n_71),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_70),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

AOI222xp33_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_56),
.B1(n_71),
.B2(n_65),
.C1(n_63),
.C2(n_53),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_72),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_95),
.B(n_58),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_96),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_92),
.Y(n_109)
);

NAND4xp25_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_53),
.C(n_99),
.D(n_83),
.Y(n_110)
);

NAND3xp33_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_97),
.C(n_77),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_95),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_88),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_112),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_105),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_102),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_104),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_117),
.A2(n_110),
.B1(n_116),
.B2(n_58),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_105),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_101),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_113),
.Y(n_125)
);

NAND2x1_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_106),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_58),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g128 ( 
.A(n_121),
.B(n_90),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_75),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

NAND2xp33_ASAP7_75t_R g131 ( 
.A(n_119),
.B(n_90),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_119),
.Y(n_133)
);

NOR2xp67_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_120),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_SL g135 ( 
.A1(n_128),
.A2(n_121),
.B(n_90),
.Y(n_135)
);

NOR2x1p5_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_124),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_130),
.Y(n_137)
);

O2A1O1Ixp5_ASAP7_75t_L g138 ( 
.A1(n_126),
.A2(n_62),
.B(n_79),
.C(n_125),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_125),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_137),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_136),
.A2(n_131),
.B1(n_90),
.B2(n_66),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_68),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_68),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

OAI21x1_ASAP7_75t_L g148 ( 
.A1(n_146),
.A2(n_138),
.B(n_142),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_144),
.Y(n_149)
);

NOR2x1p5_ASAP7_75t_L g150 ( 
.A(n_147),
.B(n_80),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

NOR2x1_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_90),
.Y(n_152)
);

AND2x4_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_143),
.Y(n_153)
);

XNOR2x1_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_67),
.Y(n_154)
);

OA21x2_ASAP7_75t_L g155 ( 
.A1(n_148),
.A2(n_106),
.B(n_87),
.Y(n_155)
);

NAND5xp2_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_67),
.C(n_107),
.D(n_59),
.E(n_94),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_157),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_149),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_156),
.A2(n_152),
.B1(n_154),
.B2(n_150),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_156),
.A2(n_154),
.B(n_148),
.Y(n_161)
);

NAND3xp33_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_153),
.C(n_155),
.Y(n_162)
);

AOI221xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_160),
.B1(n_159),
.B2(n_153),
.C(n_158),
.Y(n_163)
);


endmodule