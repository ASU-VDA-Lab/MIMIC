module real_aes_12446_n_1 (n_0, n_1);
input n_0;
output n_1;
wire n_4;
wire n_3;
wire n_5;
wire n_2;
BUFx10_ASAP7_75t_L g5 ( .A(n_0), .Y(n_5) );
CKINVDCx5p33_ASAP7_75t_R g1 ( .A(n_2), .Y(n_1) );
BUFx2_ASAP7_75t_R g2 ( .A(n_3), .Y(n_2) );
CKINVDCx5p33_ASAP7_75t_R g3 ( .A(n_4), .Y(n_3) );
CKINVDCx11_ASAP7_75t_R g4 ( .A(n_5), .Y(n_4) );
endmodule