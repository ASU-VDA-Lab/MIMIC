module fake_netlist_6_1566_n_1864 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1864);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1864;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g184 ( 
.A(n_1),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_89),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_110),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_46),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_43),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_32),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_146),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_164),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_31),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_176),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_118),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_22),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_124),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_67),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_152),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_135),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_126),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_87),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_10),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_73),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_7),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_70),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_20),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_61),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_159),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_81),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_168),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_55),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_170),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_116),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_105),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_144),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_154),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_82),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_74),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_52),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_59),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_15),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_162),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_68),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_92),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_183),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_59),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_20),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_145),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_141),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_157),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_38),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_13),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_129),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_166),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_160),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_71),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_111),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_122),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_177),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_4),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_49),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_24),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_19),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_104),
.Y(n_245)
);

BUFx10_ASAP7_75t_L g246 ( 
.A(n_90),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_10),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_180),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_75),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_8),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_158),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_43),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_66),
.Y(n_253)
);

BUFx8_ASAP7_75t_SL g254 ( 
.A(n_17),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_27),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_101),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_123),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_49),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_36),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_134),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_83),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_17),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_142),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_163),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_61),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_21),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_78),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_148),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_18),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_25),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_32),
.Y(n_271)
);

INVxp33_ASAP7_75t_SL g272 ( 
.A(n_76),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_107),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_24),
.Y(n_274)
);

BUFx5_ASAP7_75t_L g275 ( 
.A(n_112),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_3),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_69),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_52),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_6),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_36),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_33),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_33),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_0),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_45),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_156),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_45),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_139),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_21),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_30),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_143),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_79),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_102),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_128),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_115),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_85),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_140),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_50),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_108),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_26),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_98),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_48),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_11),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_153),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_16),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_178),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_147),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_65),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_22),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_29),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_96),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_18),
.Y(n_311)
);

INVx2_ASAP7_75t_SL g312 ( 
.A(n_13),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_29),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_1),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_125),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_94),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_138),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_48),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_181),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_19),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_136),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_4),
.Y(n_322)
);

BUFx5_ASAP7_75t_L g323 ( 
.A(n_171),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_99),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_91),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_12),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_165),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_64),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_26),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_131),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_174),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_7),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_150),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_121),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_39),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_12),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_23),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_117),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_28),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_120),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_50),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_127),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_151),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_30),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_100),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_137),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_97),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_0),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_41),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_35),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_62),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_2),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_14),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_16),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_133),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_35),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_44),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_23),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_93),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_167),
.Y(n_360)
);

BUFx5_ASAP7_75t_L g361 ( 
.A(n_5),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_14),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_72),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_86),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_11),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_84),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_215),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_361),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_361),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_361),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_254),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_216),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_301),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_195),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_361),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_361),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_239),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_332),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_249),
.B(n_2),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_361),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_318),
.B(n_3),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_316),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_296),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_330),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_342),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_220),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_361),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_361),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_221),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_221),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_222),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_187),
.B(n_5),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_217),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_310),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_187),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_309),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_246),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_309),
.Y(n_398)
);

INVxp33_ASAP7_75t_L g399 ( 
.A(n_192),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_365),
.Y(n_400)
);

INVxp67_ASAP7_75t_SL g401 ( 
.A(n_268),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_365),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_227),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_218),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_287),
.B(n_6),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_228),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_221),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_229),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_243),
.B(n_8),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_305),
.B(n_9),
.Y(n_410)
);

INVxp33_ASAP7_75t_SL g411 ( 
.A(n_188),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_294),
.B(n_9),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_294),
.B(n_15),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_221),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_221),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_184),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_189),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_232),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_252),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_266),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_233),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_276),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_241),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_242),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_244),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_279),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_286),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_230),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_231),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_297),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_235),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_313),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_322),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_275),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_275),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_288),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_337),
.Y(n_437)
);

INVxp67_ASAP7_75t_SL g438 ( 
.A(n_202),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_288),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_247),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_299),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_236),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_272),
.B(n_25),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_255),
.Y(n_444)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_202),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_238),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_245),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_253),
.Y(n_448)
);

INVxp33_ASAP7_75t_SL g449 ( 
.A(n_188),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_299),
.Y(n_450)
);

BUFx10_ASAP7_75t_L g451 ( 
.A(n_243),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_256),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_335),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_275),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_335),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_259),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_339),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_261),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_372),
.Y(n_459)
);

AND3x1_ASAP7_75t_L g460 ( 
.A(n_443),
.B(n_312),
.C(n_269),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_404),
.Y(n_461)
);

AND2x6_ASAP7_75t_L g462 ( 
.A(n_409),
.B(n_296),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_377),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_408),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_383),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_428),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_389),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_382),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_429),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_383),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_389),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_R g472 ( 
.A(n_431),
.B(n_442),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_379),
.A2(n_250),
.B1(n_348),
.B2(n_311),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_446),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_383),
.Y(n_475)
);

BUFx8_ASAP7_75t_L g476 ( 
.A(n_381),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_384),
.Y(n_477)
);

BUFx10_ASAP7_75t_L g478 ( 
.A(n_371),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_383),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_438),
.B(n_293),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_447),
.Y(n_481)
);

AND2x6_ASAP7_75t_L g482 ( 
.A(n_409),
.B(n_296),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_390),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_390),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_407),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_448),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_385),
.Y(n_487)
);

OA21x2_ASAP7_75t_L g488 ( 
.A1(n_368),
.A2(n_199),
.B(n_193),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_452),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_401),
.B(n_272),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_458),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_373),
.B(n_246),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_414),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_415),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_445),
.B(n_392),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_392),
.B(n_269),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_371),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_368),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_369),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_388),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_394),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_388),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_374),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_367),
.B(n_293),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_369),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_376),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_386),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_383),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_376),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_370),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_386),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_380),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_380),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_375),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_393),
.B(n_193),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_387),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_374),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_387),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_391),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_434),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_436),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_436),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_395),
.B(n_396),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_398),
.B(n_400),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_439),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_434),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_439),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_391),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_403),
.Y(n_529)
);

AND2x6_ASAP7_75t_L g530 ( 
.A(n_381),
.B(n_296),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_441),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_402),
.B(n_312),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_435),
.B(n_199),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_378),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_403),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_441),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_450),
.Y(n_537)
);

OAI22xp33_ASAP7_75t_SL g538 ( 
.A1(n_515),
.A2(n_412),
.B1(n_413),
.B2(n_397),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_495),
.A2(n_410),
.B1(n_405),
.B2(n_399),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_495),
.B(n_373),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_524),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_496),
.B(n_406),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_524),
.Y(n_543)
);

OR2x6_ASAP7_75t_L g544 ( 
.A(n_504),
.B(n_416),
.Y(n_544)
);

INVxp67_ASAP7_75t_SL g545 ( 
.A(n_520),
.Y(n_545)
);

AND2x6_ASAP7_75t_L g546 ( 
.A(n_496),
.B(n_201),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_490),
.B(n_411),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_476),
.B(n_406),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_465),
.Y(n_549)
);

AO22x2_ASAP7_75t_L g550 ( 
.A1(n_460),
.A2(n_201),
.B1(n_356),
.B2(n_358),
.Y(n_550)
);

NAND2xp33_ASAP7_75t_SL g551 ( 
.A(n_492),
.B(n_258),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_465),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_532),
.B(n_450),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_465),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_520),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_500),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_L g557 ( 
.A1(n_530),
.A2(n_449),
.B1(n_362),
.B2(n_419),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_530),
.A2(n_482),
.B1(n_462),
.B2(n_533),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_498),
.B(n_421),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_476),
.B(n_421),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_520),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_498),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_480),
.B(n_423),
.Y(n_563)
);

OR2x2_ASAP7_75t_L g564 ( 
.A(n_473),
.B(n_378),
.Y(n_564)
);

OR2x6_ASAP7_75t_L g565 ( 
.A(n_523),
.B(n_314),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_530),
.A2(n_457),
.B1(n_427),
.B2(n_430),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_499),
.B(n_423),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_499),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_505),
.B(n_424),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_507),
.B(n_424),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_500),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_505),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_500),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_SL g574 ( 
.A1(n_476),
.A2(n_246),
.B1(n_307),
.B2(n_203),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_476),
.B(n_425),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_506),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_511),
.B(n_425),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_532),
.B(n_521),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_521),
.B(n_453),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_519),
.B(n_440),
.Y(n_580)
);

NAND3xp33_ASAP7_75t_L g581 ( 
.A(n_473),
.B(n_444),
.C(n_440),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_506),
.Y(n_582)
);

BUFx4f_ASAP7_75t_L g583 ( 
.A(n_530),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_465),
.Y(n_584)
);

NOR2x1p5_ASAP7_75t_L g585 ( 
.A(n_497),
.B(n_444),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_472),
.Y(n_586)
);

INVx4_ASAP7_75t_L g587 ( 
.A(n_520),
.Y(n_587)
);

INVx4_ASAP7_75t_SL g588 ( 
.A(n_462),
.Y(n_588)
);

AND2x6_ASAP7_75t_L g589 ( 
.A(n_533),
.B(n_296),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_509),
.Y(n_590)
);

BUFx10_ASAP7_75t_L g591 ( 
.A(n_528),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_460),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_465),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_512),
.Y(n_594)
);

AND2x6_ASAP7_75t_L g595 ( 
.A(n_533),
.B(n_300),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_513),
.Y(n_596)
);

INVxp33_ASAP7_75t_L g597 ( 
.A(n_503),
.Y(n_597)
);

OR2x2_ASAP7_75t_L g598 ( 
.A(n_517),
.B(n_456),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_513),
.B(n_456),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_483),
.Y(n_600)
);

INVxp67_ASAP7_75t_SL g601 ( 
.A(n_470),
.Y(n_601)
);

BUFx8_ASAP7_75t_SL g602 ( 
.A(n_459),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_518),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_529),
.B(n_417),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_535),
.B(n_451),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_SL g606 ( 
.A1(n_534),
.A2(n_307),
.B1(n_336),
.B2(n_341),
.Y(n_606)
);

INVx4_ASAP7_75t_L g607 ( 
.A(n_533),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_522),
.B(n_455),
.Y(n_608)
);

AO21x2_ASAP7_75t_L g609 ( 
.A1(n_518),
.A2(n_194),
.B(n_186),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_522),
.B(n_455),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_SL g611 ( 
.A(n_461),
.B(n_307),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_462),
.B(n_190),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_525),
.B(n_453),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_478),
.B(n_451),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_525),
.B(n_451),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_483),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_510),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_502),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_530),
.A2(n_482),
.B1(n_462),
.B2(n_488),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_510),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_479),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_516),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_462),
.B(n_251),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_462),
.B(n_263),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_462),
.B(n_264),
.Y(n_625)
);

BUFx10_ASAP7_75t_L g626 ( 
.A(n_464),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_482),
.B(n_267),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_502),
.Y(n_628)
);

AND2x6_ASAP7_75t_L g629 ( 
.A(n_516),
.B(n_300),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_530),
.A2(n_432),
.B1(n_437),
.B2(n_420),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_527),
.B(n_418),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_479),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_478),
.B(n_185),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_478),
.B(n_185),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_482),
.B(n_273),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_479),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_514),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_514),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_493),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_527),
.B(n_422),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_478),
.B(n_191),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_493),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_494),
.Y(n_643)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_494),
.B(n_426),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_482),
.B(n_277),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_466),
.B(n_191),
.Y(n_646)
);

BUFx6f_ASAP7_75t_SL g647 ( 
.A(n_530),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_469),
.B(n_197),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_479),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_467),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_526),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_531),
.B(n_197),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_485),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_526),
.Y(n_654)
);

OAI22xp5_ASAP7_75t_L g655 ( 
.A1(n_537),
.A2(n_326),
.B1(n_262),
.B2(n_265),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_531),
.B(n_433),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_485),
.Y(n_657)
);

AND3x2_ASAP7_75t_L g658 ( 
.A(n_536),
.B(n_204),
.C(n_196),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_482),
.B(n_285),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_482),
.B(n_290),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_467),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_470),
.B(n_291),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_471),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_471),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_536),
.B(n_435),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_484),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_537),
.B(n_198),
.Y(n_667)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_474),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_484),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_479),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_488),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_481),
.B(n_198),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_470),
.Y(n_673)
);

INVx4_ASAP7_75t_L g674 ( 
.A(n_508),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_470),
.B(n_200),
.Y(n_675)
);

BUFx4f_ASAP7_75t_L g676 ( 
.A(n_488),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_475),
.Y(n_677)
);

AND2x2_ASAP7_75t_SL g678 ( 
.A(n_488),
.B(n_300),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_475),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_475),
.Y(n_680)
);

OR2x6_ASAP7_75t_L g681 ( 
.A(n_486),
.B(n_219),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_508),
.B(n_292),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_508),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_508),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_489),
.B(n_200),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_491),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_501),
.B(n_206),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_563),
.B(n_206),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_568),
.B(n_223),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_542),
.B(n_547),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_568),
.B(n_224),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_592),
.A2(n_559),
.B1(n_569),
.B2(n_567),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_582),
.B(n_225),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_578),
.B(n_454),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_582),
.B(n_226),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_578),
.B(n_454),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_664),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_599),
.B(n_463),
.Y(n_698)
);

A2O1A1Ixp33_ASAP7_75t_L g699 ( 
.A1(n_562),
.A2(n_317),
.B(n_295),
.C(n_260),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_671),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_664),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_540),
.B(n_209),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_541),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_603),
.B(n_234),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_603),
.B(n_237),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_615),
.B(n_209),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_615),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_538),
.B(n_210),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_604),
.B(n_611),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_546),
.A2(n_345),
.B1(n_298),
.B2(n_257),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_592),
.A2(n_328),
.B1(n_321),
.B2(n_324),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_541),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_685),
.B(n_468),
.Y(n_713)
);

OAI22xp33_ASAP7_75t_L g714 ( 
.A1(n_565),
.A2(n_350),
.B1(n_352),
.B2(n_240),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_661),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_543),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_572),
.B(n_576),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_604),
.B(n_605),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_590),
.B(n_248),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_543),
.B(n_210),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_661),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_594),
.B(n_303),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_574),
.B(n_211),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_553),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_596),
.B(n_306),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_564),
.B(n_203),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_669),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_620),
.B(n_315),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_539),
.B(n_211),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_620),
.B(n_319),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_671),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_669),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_607),
.B(n_213),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_L g734 ( 
.A(n_619),
.B(n_275),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_581),
.B(n_477),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_637),
.B(n_325),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_637),
.B(n_327),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_638),
.B(n_343),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_638),
.B(n_346),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_618),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_665),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_607),
.B(n_213),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_607),
.B(n_214),
.Y(n_743)
);

OAI21xp5_ASAP7_75t_L g744 ( 
.A1(n_676),
.A2(n_333),
.B(n_366),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_618),
.Y(n_745)
);

AND2x2_ASAP7_75t_SL g746 ( 
.A(n_557),
.B(n_300),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_628),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_665),
.Y(n_748)
);

A2O1A1Ixp33_ASAP7_75t_L g749 ( 
.A1(n_676),
.A2(n_331),
.B(n_364),
.C(n_214),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_678),
.B(n_300),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_678),
.B(n_363),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_556),
.Y(n_752)
);

AND2x2_ASAP7_75t_SL g753 ( 
.A(n_558),
.B(n_363),
.Y(n_753)
);

INVxp67_ASAP7_75t_SL g754 ( 
.A(n_676),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_553),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_564),
.B(n_205),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_556),
.Y(n_757)
);

OAI22xp33_ASAP7_75t_L g758 ( 
.A1(n_565),
.A2(n_205),
.B1(n_207),
.B2(n_208),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_644),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_570),
.B(n_487),
.Y(n_760)
);

OAI22x1_ASAP7_75t_SL g761 ( 
.A1(n_586),
.A2(n_207),
.B1(n_208),
.B2(n_212),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_598),
.B(n_334),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_565),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_631),
.B(n_275),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_653),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_544),
.A2(n_364),
.B1(n_347),
.B2(n_360),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_653),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_544),
.A2(n_551),
.B1(n_546),
.B2(n_550),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_546),
.A2(n_323),
.B1(n_275),
.B2(n_363),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_644),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_650),
.B(n_363),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_577),
.B(n_334),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_546),
.A2(n_323),
.B1(n_275),
.B2(n_363),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_663),
.B(n_338),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_666),
.B(n_338),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_601),
.B(n_340),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_580),
.B(n_340),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_631),
.B(n_275),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_571),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_657),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_639),
.B(n_347),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_642),
.B(n_355),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_643),
.B(n_355),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_SL g784 ( 
.A(n_586),
.B(n_591),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_657),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_571),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_675),
.B(n_359),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_545),
.A2(n_360),
.B(n_359),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_680),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_651),
.Y(n_790)
);

O2A1O1Ixp5_ASAP7_75t_L g791 ( 
.A1(n_583),
.A2(n_323),
.B(n_270),
.C(n_271),
.Y(n_791)
);

AND2x6_ASAP7_75t_SL g792 ( 
.A(n_687),
.B(n_212),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_651),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_546),
.A2(n_323),
.B1(n_354),
.B2(n_353),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_654),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_SL g796 ( 
.A(n_591),
.B(n_336),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_617),
.B(n_323),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_646),
.B(n_274),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_652),
.B(n_323),
.Y(n_799)
);

BUFx3_ASAP7_75t_L g800 ( 
.A(n_602),
.Y(n_800)
);

OAI221xp5_ASAP7_75t_L g801 ( 
.A1(n_606),
.A2(n_308),
.B1(n_280),
.B2(n_281),
.C(n_282),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_648),
.B(n_672),
.Y(n_802)
);

OAI22x1_ASAP7_75t_R g803 ( 
.A1(n_602),
.A2(n_357),
.B1(n_354),
.B2(n_353),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_609),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_544),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_573),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_598),
.B(n_320),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_573),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_667),
.B(n_278),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_626),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_600),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_SL g812 ( 
.A(n_591),
.B(n_626),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_600),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_583),
.A2(n_329),
.B(n_284),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_654),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_626),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_616),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_622),
.B(n_283),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_622),
.B(n_289),
.Y(n_819)
);

AOI22xp5_ASAP7_75t_L g820 ( 
.A1(n_544),
.A2(n_304),
.B1(n_302),
.B2(n_349),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_640),
.B(n_357),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_616),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_579),
.Y(n_823)
);

AND2x6_ASAP7_75t_SL g824 ( 
.A(n_681),
.B(n_351),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_609),
.A2(n_550),
.B1(n_551),
.B2(n_623),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_680),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_579),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_597),
.B(n_351),
.Y(n_828)
);

AND2x2_ASAP7_75t_SL g829 ( 
.A(n_583),
.B(n_77),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_609),
.A2(n_344),
.B1(n_341),
.B2(n_349),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_550),
.A2(n_344),
.B1(n_182),
.B2(n_179),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_608),
.Y(n_832)
);

INVx4_ASAP7_75t_L g833 ( 
.A(n_588),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_662),
.B(n_175),
.Y(n_834)
);

O2A1O1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_612),
.A2(n_27),
.B(n_28),
.C(n_31),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_608),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_555),
.B(n_172),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_SL g838 ( 
.A(n_668),
.B(n_34),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_610),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_610),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_614),
.B(n_34),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_555),
.B(n_169),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_683),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_613),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_597),
.B(n_633),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_613),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_640),
.B(n_161),
.Y(n_847)
);

INVxp67_ASAP7_75t_L g848 ( 
.A(n_655),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_634),
.B(n_37),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_555),
.B(n_155),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_641),
.B(n_37),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_656),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_656),
.B(n_149),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_550),
.B(n_132),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_561),
.B(n_130),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_694),
.B(n_565),
.Y(n_856)
);

INVxp67_ASAP7_75t_SL g857 ( 
.A(n_731),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_694),
.B(n_682),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_696),
.B(n_673),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_707),
.B(n_686),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_696),
.B(n_677),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_700),
.A2(n_587),
.B(n_624),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_836),
.B(n_679),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_754),
.A2(n_625),
.B(n_627),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_744),
.A2(n_635),
.B(n_660),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_750),
.A2(n_659),
.B(n_645),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_690),
.B(n_686),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_751),
.A2(n_833),
.B(n_731),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_836),
.B(n_549),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_740),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_692),
.B(n_548),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_718),
.B(n_575),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_839),
.B(n_844),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_707),
.B(n_560),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_848),
.B(n_681),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_790),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_740),
.Y(n_877)
);

BUFx4_ASAP7_75t_SL g878 ( 
.A(n_800),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_712),
.B(n_588),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_802),
.A2(n_585),
.B1(n_681),
.B2(n_647),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_759),
.B(n_681),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_839),
.B(n_549),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_753),
.A2(n_630),
.B1(n_566),
.B2(n_647),
.Y(n_883)
);

O2A1O1Ixp5_ASAP7_75t_L g884 ( 
.A1(n_791),
.A2(n_683),
.B(n_549),
.C(n_554),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_790),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_853),
.A2(n_647),
.B1(n_595),
.B2(n_589),
.Y(n_886)
);

O2A1O1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_724),
.A2(n_554),
.B(n_584),
.C(n_649),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_731),
.B(n_588),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_844),
.B(n_554),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_731),
.Y(n_890)
);

BUFx2_ASAP7_75t_L g891 ( 
.A(n_763),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_753),
.B(n_584),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_745),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_741),
.B(n_584),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_851),
.A2(n_632),
.B(n_649),
.C(n_621),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_712),
.B(n_716),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_746),
.A2(n_632),
.B1(n_649),
.B2(n_674),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_789),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_847),
.B(n_588),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_816),
.Y(n_900)
);

OAI21xp5_ASAP7_75t_L g901 ( 
.A1(n_804),
.A2(n_734),
.B(n_741),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_734),
.A2(n_674),
.B(n_684),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_759),
.B(n_632),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_748),
.A2(n_684),
.B(n_670),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_717),
.A2(n_684),
.B(n_670),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_789),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_847),
.B(n_684),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_789),
.A2(n_670),
.B(n_552),
.Y(n_908)
);

BUFx4f_ASAP7_75t_L g909 ( 
.A(n_854),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_804),
.A2(n_589),
.B(n_595),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_826),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_746),
.A2(n_670),
.B1(n_593),
.B2(n_636),
.Y(n_912)
);

AOI21x1_ASAP7_75t_L g913 ( 
.A1(n_799),
.A2(n_552),
.B(n_636),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_715),
.B(n_552),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_715),
.B(n_552),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_853),
.A2(n_552),
.B(n_636),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_721),
.B(n_636),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_724),
.A2(n_658),
.B(n_595),
.C(n_589),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_721),
.B(n_636),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_834),
.A2(n_621),
.B(n_593),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_770),
.B(n_621),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_755),
.B(n_621),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_798),
.A2(n_621),
.B(n_593),
.C(n_595),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_749),
.A2(n_595),
.B(n_589),
.Y(n_924)
);

OAI21x1_ASAP7_75t_L g925 ( 
.A1(n_843),
.A2(n_595),
.B(n_589),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_770),
.B(n_38),
.Y(n_926)
);

INVxp67_ASAP7_75t_L g927 ( 
.A(n_828),
.Y(n_927)
);

NOR2x1_ASAP7_75t_L g928 ( 
.A(n_810),
.B(n_593),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_755),
.B(n_593),
.Y(n_929)
);

INVx4_ASAP7_75t_L g930 ( 
.A(n_703),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_793),
.Y(n_931)
);

NAND3xp33_ASAP7_75t_L g932 ( 
.A(n_777),
.B(n_39),
.C(n_40),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_703),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_823),
.B(n_629),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_823),
.B(n_629),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_827),
.B(n_629),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_847),
.B(n_629),
.Y(n_937)
);

AOI22xp5_ASAP7_75t_L g938 ( 
.A1(n_768),
.A2(n_629),
.B1(n_119),
.B2(n_114),
.Y(n_938)
);

INVx3_ASAP7_75t_SL g939 ( 
.A(n_816),
.Y(n_939)
);

A2O1A1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_807),
.A2(n_40),
.B(n_41),
.C(n_42),
.Y(n_940)
);

O2A1O1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_729),
.A2(n_42),
.B(n_44),
.C(n_46),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_825),
.A2(n_103),
.B1(n_113),
.B2(n_109),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_727),
.A2(n_629),
.B(n_106),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_827),
.B(n_832),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_843),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_810),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_837),
.A2(n_95),
.B(n_88),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_832),
.B(n_47),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_842),
.A2(n_80),
.B(n_63),
.Y(n_949)
);

OR2x6_ASAP7_75t_SL g950 ( 
.A(n_726),
.B(n_47),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_850),
.A2(n_51),
.B(n_53),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_855),
.A2(n_51),
.B(n_53),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_698),
.B(n_54),
.Y(n_953)
);

INVx3_ASAP7_75t_L g954 ( 
.A(n_843),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_697),
.A2(n_54),
.B(n_55),
.Y(n_955)
);

OAI22xp5_ASAP7_75t_L g956 ( 
.A1(n_840),
.A2(n_62),
.B1(n_57),
.B2(n_58),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_840),
.B(n_56),
.Y(n_957)
);

NAND3xp33_ASAP7_75t_L g958 ( 
.A(n_688),
.B(n_830),
.C(n_702),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_726),
.B(n_756),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_756),
.B(n_56),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_697),
.A2(n_57),
.B(n_58),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_709),
.B(n_60),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_701),
.A2(n_60),
.B(n_776),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_846),
.B(n_852),
.Y(n_964)
);

O2A1O1Ixp5_ASAP7_75t_L g965 ( 
.A1(n_787),
.A2(n_809),
.B(n_691),
.C(n_693),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_701),
.A2(n_743),
.B(n_742),
.Y(n_966)
);

BUFx4f_ASAP7_75t_L g967 ( 
.A(n_854),
.Y(n_967)
);

NOR2x1_ASAP7_75t_L g968 ( 
.A(n_735),
.B(n_845),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_846),
.B(n_852),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_733),
.A2(n_732),
.B(n_727),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_829),
.A2(n_710),
.B1(n_805),
.B2(n_732),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_764),
.A2(n_778),
.B(n_779),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_763),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_764),
.B(n_778),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_728),
.A2(n_739),
.B(n_736),
.Y(n_975)
);

AND2x2_ASAP7_75t_SL g976 ( 
.A(n_829),
.B(n_831),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_708),
.A2(n_706),
.B1(n_738),
.B2(n_737),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_821),
.B(n_841),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_730),
.A2(n_813),
.B(n_822),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_795),
.B(n_815),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_765),
.B(n_767),
.Y(n_981)
);

BUFx2_ASAP7_75t_L g982 ( 
.A(n_821),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_801),
.B(n_713),
.Y(n_983)
);

AOI22xp5_ASAP7_75t_L g984 ( 
.A1(n_818),
.A2(n_819),
.B1(n_849),
.B2(n_720),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_811),
.A2(n_813),
.B(n_822),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_719),
.A2(n_722),
.B1(n_725),
.B2(n_774),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_811),
.A2(n_817),
.B(n_780),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_817),
.A2(n_780),
.B(n_767),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_SL g989 ( 
.A1(n_723),
.A2(n_699),
.B(n_797),
.C(n_771),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_814),
.A2(n_689),
.B(n_695),
.C(n_704),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_705),
.A2(n_794),
.B(n_711),
.C(n_766),
.Y(n_991)
);

HB1xp67_ASAP7_75t_L g992 ( 
.A(n_765),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_785),
.B(n_747),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_785),
.A2(n_747),
.B(n_786),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_SL g995 ( 
.A(n_812),
.B(n_784),
.Y(n_995)
);

NOR2x1_ASAP7_75t_R g996 ( 
.A(n_800),
.B(n_762),
.Y(n_996)
);

NAND3xp33_ASAP7_75t_L g997 ( 
.A(n_820),
.B(n_760),
.C(n_783),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_752),
.A2(n_786),
.B(n_757),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_796),
.B(n_806),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_752),
.A2(n_757),
.B(n_806),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_835),
.A2(n_775),
.B(n_781),
.C(n_782),
.Y(n_1001)
);

AOI21x1_ASAP7_75t_L g1002 ( 
.A1(n_779),
.A2(n_808),
.B(n_788),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_808),
.A2(n_773),
.B(n_769),
.Y(n_1003)
);

OAI321xp33_ASAP7_75t_L g1004 ( 
.A1(n_714),
.A2(n_758),
.A3(n_838),
.B1(n_803),
.B2(n_792),
.C(n_824),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_761),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_746),
.A2(n_753),
.B1(n_734),
.B2(n_829),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_690),
.B(n_547),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_694),
.B(n_696),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_851),
.A2(n_547),
.B(n_802),
.C(n_798),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_790),
.Y(n_1010)
);

AO22x1_ASAP7_75t_L g1011 ( 
.A1(n_851),
.A2(n_547),
.B1(n_777),
.B2(n_772),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_750),
.A2(n_751),
.B(n_676),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_694),
.B(n_696),
.Y(n_1013)
);

BUFx12f_ASAP7_75t_L g1014 ( 
.A(n_824),
.Y(n_1014)
);

OR2x2_ASAP7_75t_L g1015 ( 
.A(n_726),
.B(n_756),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_694),
.B(n_696),
.Y(n_1016)
);

O2A1O1Ixp5_ASAP7_75t_L g1017 ( 
.A1(n_791),
.A2(n_688),
.B(n_744),
.C(n_799),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_700),
.A2(n_676),
.B(n_607),
.Y(n_1018)
);

CKINVDCx8_ASAP7_75t_R g1019 ( 
.A(n_792),
.Y(n_1019)
);

NOR3xp33_ASAP7_75t_L g1020 ( 
.A(n_718),
.B(n_547),
.C(n_687),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_731),
.B(n_700),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_763),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_694),
.B(n_696),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_753),
.A2(n_746),
.B1(n_692),
.B2(n_848),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_694),
.B(n_696),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_790),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_790),
.Y(n_1027)
);

NAND3xp33_ASAP7_75t_L g1028 ( 
.A(n_772),
.B(n_547),
.C(n_777),
.Y(n_1028)
);

OAI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_1006),
.A2(n_967),
.B1(n_909),
.B2(n_1009),
.Y(n_1029)
);

INVxp67_ASAP7_75t_L g1030 ( 
.A(n_1015),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_1002),
.A2(n_920),
.B(n_862),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_R g1032 ( 
.A(n_900),
.B(n_995),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_974),
.A2(n_972),
.B(n_1008),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_1012),
.A2(n_1003),
.B(n_1024),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_1017),
.A2(n_901),
.B(n_1013),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_890),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_1016),
.A2(n_1025),
.B(n_1023),
.Y(n_1037)
);

NOR2x1_ASAP7_75t_L g1038 ( 
.A(n_997),
.B(n_930),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_858),
.A2(n_865),
.B(n_975),
.Y(n_1039)
);

O2A1O1Ixp5_ASAP7_75t_L g1040 ( 
.A1(n_1011),
.A2(n_1028),
.B(n_983),
.C(n_965),
.Y(n_1040)
);

AO31x2_ASAP7_75t_L g1041 ( 
.A1(n_923),
.A2(n_895),
.A3(n_971),
.B(n_990),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_891),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_SL g1043 ( 
.A1(n_857),
.A2(n_883),
.B(n_890),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_1007),
.B(n_1006),
.Y(n_1044)
);

NAND3xp33_ASAP7_75t_SL g1045 ( 
.A(n_983),
.B(n_1020),
.C(n_953),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_871),
.A2(n_967),
.B1(n_909),
.B2(n_1007),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_1018),
.A2(n_884),
.B(n_913),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_873),
.B(n_1027),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_870),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_877),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_927),
.B(n_867),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_907),
.A2(n_864),
.B(n_868),
.Y(n_1052)
);

OAI21x1_ASAP7_75t_L g1053 ( 
.A1(n_979),
.A2(n_916),
.B(n_988),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_992),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_930),
.B(n_933),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_867),
.B(n_875),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_991),
.A2(n_866),
.B(n_998),
.Y(n_1057)
);

AO31x2_ASAP7_75t_L g1058 ( 
.A1(n_912),
.A2(n_897),
.A3(n_970),
.B(n_942),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_876),
.Y(n_1059)
);

OAI21x1_ASAP7_75t_L g1060 ( 
.A1(n_1000),
.A2(n_985),
.B(n_994),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_987),
.A2(n_908),
.B(n_925),
.Y(n_1061)
);

OAI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_892),
.A2(n_958),
.B(n_856),
.Y(n_1062)
);

BUFx8_ASAP7_75t_L g1063 ( 
.A(n_1022),
.Y(n_1063)
);

OA21x2_ASAP7_75t_L g1064 ( 
.A1(n_910),
.A2(n_980),
.B(n_943),
.Y(n_1064)
);

AOI221xp5_ASAP7_75t_L g1065 ( 
.A1(n_960),
.A2(n_953),
.B1(n_871),
.B2(n_962),
.C(n_956),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_SL g1066 ( 
.A1(n_941),
.A2(n_963),
.B(n_966),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_959),
.B(n_982),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_976),
.A2(n_944),
.B1(n_969),
.B2(n_964),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_907),
.A2(n_899),
.B(n_857),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1026),
.B(n_885),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_899),
.A2(n_1021),
.B(n_902),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_893),
.Y(n_1072)
);

NOR2x1_ASAP7_75t_SL g1073 ( 
.A(n_890),
.B(n_888),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_959),
.B(n_978),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_973),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_904),
.A2(n_905),
.B(n_887),
.Y(n_1076)
);

AND2x4_ASAP7_75t_L g1077 ( 
.A(n_933),
.B(n_978),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_914),
.A2(n_919),
.B(n_915),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_875),
.B(n_872),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_917),
.A2(n_993),
.B(n_981),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_960),
.B(n_881),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_946),
.B(n_968),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_1021),
.A2(n_859),
.B(n_861),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_937),
.A2(n_888),
.B(n_898),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_924),
.A2(n_889),
.B(n_882),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_878),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_973),
.Y(n_1087)
);

AO31x2_ASAP7_75t_L g1088 ( 
.A1(n_940),
.A2(n_962),
.A3(n_948),
.B(n_957),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_869),
.A2(n_945),
.B(n_954),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_898),
.A2(n_906),
.B(n_922),
.Y(n_1090)
);

NAND3xp33_ASAP7_75t_SL g1091 ( 
.A(n_872),
.B(n_880),
.C(n_874),
.Y(n_1091)
);

NAND3xp33_ASAP7_75t_SL g1092 ( 
.A(n_874),
.B(n_984),
.C(n_977),
.Y(n_1092)
);

INVxp67_ASAP7_75t_SL g1093 ( 
.A(n_890),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_989),
.A2(n_1001),
.B(n_999),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_906),
.A2(n_929),
.B(n_896),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_945),
.A2(n_954),
.B(n_894),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_931),
.B(n_1010),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_934),
.A2(n_936),
.B(n_935),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_911),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_879),
.A2(n_863),
.B(n_921),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_986),
.B(n_976),
.Y(n_1101)
);

NAND2x1_ASAP7_75t_L g1102 ( 
.A(n_928),
.B(n_921),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_903),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_926),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_918),
.A2(n_932),
.B(n_903),
.C(n_951),
.Y(n_1105)
);

AO21x1_ASAP7_75t_L g1106 ( 
.A1(n_952),
.A2(n_949),
.B(n_947),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_996),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_860),
.B(n_938),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_886),
.A2(n_961),
.B(n_955),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1004),
.A2(n_1005),
.B(n_950),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_939),
.A2(n_878),
.B(n_1019),
.Y(n_1111)
);

AO31x2_ASAP7_75t_L g1112 ( 
.A1(n_939),
.A2(n_1014),
.A3(n_923),
.B(n_1024),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_959),
.B(n_982),
.Y(n_1113)
);

AND2x6_ASAP7_75t_L g1114 ( 
.A(n_890),
.B(n_854),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_992),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_974),
.B(n_1008),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_1002),
.A2(n_920),
.B(n_862),
.Y(n_1117)
);

O2A1O1Ixp5_ASAP7_75t_L g1118 ( 
.A1(n_1011),
.A2(n_1028),
.B(n_1009),
.C(n_983),
.Y(n_1118)
);

INVx8_ASAP7_75t_L g1119 ( 
.A(n_890),
.Y(n_1119)
);

NOR2x1_ASAP7_75t_SL g1120 ( 
.A(n_890),
.B(n_731),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_992),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_1028),
.B(n_1009),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_1009),
.A2(n_1028),
.B(n_983),
.C(n_1007),
.Y(n_1123)
);

OR2x6_ASAP7_75t_L g1124 ( 
.A(n_946),
.B(n_810),
.Y(n_1124)
);

NOR2xp67_ASAP7_75t_L g1125 ( 
.A(n_900),
.B(n_668),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_1028),
.B(n_1007),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_974),
.B(n_1008),
.Y(n_1127)
);

NOR2x1_ASAP7_75t_L g1128 ( 
.A(n_997),
.B(n_810),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_974),
.B(n_1008),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_1002),
.A2(n_920),
.B(n_862),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_974),
.B(n_1008),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_974),
.B(n_1008),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_1009),
.A2(n_1028),
.B(n_983),
.C(n_1007),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1002),
.A2(n_920),
.B(n_862),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_1002),
.A2(n_920),
.B(n_862),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_974),
.B(n_1008),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1012),
.A2(n_974),
.B(n_1003),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_974),
.A2(n_972),
.B(n_1008),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_959),
.B(n_982),
.Y(n_1139)
);

BUFx2_ASAP7_75t_SL g1140 ( 
.A(n_946),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1012),
.A2(n_974),
.B(n_1003),
.Y(n_1141)
);

BUFx12f_ASAP7_75t_L g1142 ( 
.A(n_900),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_973),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1002),
.A2(n_920),
.B(n_862),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_930),
.B(n_703),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1002),
.A2(n_920),
.B(n_862),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_974),
.A2(n_972),
.B(n_1008),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_890),
.Y(n_1148)
);

OAI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1012),
.A2(n_974),
.B(n_1003),
.Y(n_1149)
);

INVx5_ASAP7_75t_L g1150 ( 
.A(n_890),
.Y(n_1150)
);

INVxp67_ASAP7_75t_L g1151 ( 
.A(n_1015),
.Y(n_1151)
);

INVx3_ASAP7_75t_SL g1152 ( 
.A(n_900),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1006),
.A2(n_967),
.B1(n_909),
.B2(n_1009),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1002),
.A2(n_920),
.B(n_862),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1012),
.A2(n_974),
.B(n_1003),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_930),
.B(n_703),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1002),
.A2(n_920),
.B(n_862),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_974),
.B(n_1008),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_1002),
.A2(n_920),
.B(n_862),
.Y(n_1159)
);

OR2x2_ASAP7_75t_L g1160 ( 
.A(n_1015),
.B(n_726),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_974),
.B(n_1008),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1002),
.A2(n_920),
.B(n_862),
.Y(n_1162)
);

AOI21x1_ASAP7_75t_L g1163 ( 
.A1(n_866),
.A2(n_980),
.B(n_865),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_959),
.B(n_982),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1002),
.A2(n_920),
.B(n_862),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_973),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_959),
.B(n_982),
.Y(n_1167)
);

OA21x2_ASAP7_75t_L g1168 ( 
.A1(n_1012),
.A2(n_901),
.B(n_972),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1009),
.A2(n_1028),
.B(n_983),
.C(n_1007),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_992),
.Y(n_1170)
);

AO31x2_ASAP7_75t_L g1171 ( 
.A1(n_923),
.A2(n_1024),
.A3(n_895),
.B(n_865),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_974),
.A2(n_972),
.B(n_1008),
.Y(n_1172)
);

AND2x2_ASAP7_75t_SL g1173 ( 
.A(n_976),
.B(n_909),
.Y(n_1173)
);

BUFx2_ASAP7_75t_L g1174 ( 
.A(n_891),
.Y(n_1174)
);

AO31x2_ASAP7_75t_L g1175 ( 
.A1(n_923),
.A2(n_1024),
.A3(n_895),
.B(n_865),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1012),
.A2(n_974),
.B(n_1003),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_974),
.A2(n_972),
.B(n_1008),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1009),
.A2(n_1028),
.B(n_983),
.C(n_1007),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_1032),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1074),
.B(n_1067),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_1079),
.B(n_1126),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1059),
.Y(n_1182)
);

AO21x1_ASAP7_75t_L g1183 ( 
.A1(n_1029),
.A2(n_1153),
.B(n_1122),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_1063),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1049),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1056),
.B(n_1116),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1145),
.B(n_1156),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_1042),
.Y(n_1188)
);

NAND2x1p5_ASAP7_75t_L g1189 ( 
.A(n_1150),
.B(n_1036),
.Y(n_1189)
);

OR2x2_ASAP7_75t_L g1190 ( 
.A(n_1160),
.B(n_1030),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1039),
.A2(n_1057),
.B(n_1052),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1050),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1145),
.B(n_1156),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1116),
.B(n_1127),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1072),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_1051),
.B(n_1045),
.Y(n_1196)
);

INVx2_ASAP7_75t_SL g1197 ( 
.A(n_1063),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1113),
.B(n_1139),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_1077),
.B(n_1055),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_1087),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1091),
.B(n_1164),
.Y(n_1201)
);

INVx1_ASAP7_75t_SL g1202 ( 
.A(n_1174),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_SL g1203 ( 
.A1(n_1057),
.A2(n_1034),
.B(n_1035),
.C(n_1094),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1034),
.A2(n_1141),
.B(n_1137),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1137),
.A2(n_1149),
.B(n_1141),
.Y(n_1205)
);

INVx2_ASAP7_75t_SL g1206 ( 
.A(n_1124),
.Y(n_1206)
);

OR2x2_ASAP7_75t_L g1207 ( 
.A(n_1151),
.B(n_1167),
.Y(n_1207)
);

AO21x2_ASAP7_75t_L g1208 ( 
.A1(n_1092),
.A2(n_1035),
.B(n_1163),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1081),
.B(n_1104),
.Y(n_1209)
);

AOI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1065),
.A2(n_1046),
.B1(n_1101),
.B2(n_1125),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1142),
.Y(n_1211)
);

AOI21xp33_ASAP7_75t_SL g1212 ( 
.A1(n_1152),
.A2(n_1110),
.B(n_1082),
.Y(n_1212)
);

AO21x1_ASAP7_75t_L g1213 ( 
.A1(n_1029),
.A2(n_1153),
.B(n_1101),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1127),
.B(n_1129),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1054),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_1099),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1149),
.A2(n_1176),
.B(n_1155),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_1124),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1129),
.B(n_1131),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1131),
.B(n_1132),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_1036),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1077),
.B(n_1110),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1155),
.A2(n_1176),
.B(n_1033),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_1099),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1055),
.B(n_1082),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1132),
.B(n_1136),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1115),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_1075),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1121),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1033),
.A2(n_1138),
.B(n_1177),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1170),
.Y(n_1231)
);

A2O1A1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1118),
.A2(n_1065),
.B(n_1169),
.C(n_1123),
.Y(n_1232)
);

BUFx2_ASAP7_75t_L g1233 ( 
.A(n_1143),
.Y(n_1233)
);

AND2x4_ASAP7_75t_L g1234 ( 
.A(n_1124),
.B(n_1038),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1133),
.B(n_1178),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1138),
.A2(n_1177),
.B(n_1172),
.Y(n_1236)
);

O2A1O1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1040),
.A2(n_1068),
.B(n_1105),
.C(n_1044),
.Y(n_1237)
);

NOR2xp67_ASAP7_75t_L g1238 ( 
.A(n_1166),
.B(n_1086),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1136),
.B(n_1158),
.Y(n_1239)
);

CKINVDCx20_ASAP7_75t_R g1240 ( 
.A(n_1107),
.Y(n_1240)
);

AOI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1173),
.A2(n_1128),
.B1(n_1068),
.B2(n_1044),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1070),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1043),
.A2(n_1172),
.B(n_1147),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1158),
.B(n_1161),
.Y(n_1244)
);

INVx2_ASAP7_75t_SL g1245 ( 
.A(n_1119),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_1036),
.Y(n_1246)
);

OAI221xp5_ASAP7_75t_L g1247 ( 
.A1(n_1062),
.A2(n_1161),
.B1(n_1037),
.B2(n_1108),
.C(n_1147),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1070),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1037),
.B(n_1048),
.Y(n_1249)
);

O2A1O1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1108),
.A2(n_1062),
.B(n_1066),
.C(n_1097),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1048),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1099),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1114),
.A2(n_1103),
.B1(n_1106),
.B2(n_1064),
.Y(n_1253)
);

O2A1O1Ixp5_ASAP7_75t_L g1254 ( 
.A1(n_1102),
.A2(n_1071),
.B(n_1100),
.C(n_1098),
.Y(n_1254)
);

INVx2_ASAP7_75t_SL g1255 ( 
.A(n_1119),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1083),
.A2(n_1168),
.B(n_1120),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1119),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1168),
.A2(n_1150),
.B1(n_1064),
.B2(n_1069),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1140),
.B(n_1112),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_1112),
.B(n_1150),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1114),
.B(n_1088),
.Y(n_1261)
);

INVx3_ASAP7_75t_SL g1262 ( 
.A(n_1114),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1112),
.B(n_1150),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1114),
.B(n_1093),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1148),
.B(n_1073),
.Y(n_1265)
);

OR2x6_ASAP7_75t_L g1266 ( 
.A(n_1111),
.B(n_1084),
.Y(n_1266)
);

INVx1_ASAP7_75t_SL g1267 ( 
.A(n_1111),
.Y(n_1267)
);

INVx4_ASAP7_75t_L g1268 ( 
.A(n_1095),
.Y(n_1268)
);

BUFx2_ASAP7_75t_L g1269 ( 
.A(n_1088),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1080),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_1109),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1041),
.B(n_1175),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1098),
.B(n_1090),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_1078),
.B(n_1085),
.Y(n_1274)
);

AO22x1_ASAP7_75t_L g1275 ( 
.A1(n_1041),
.A2(n_1175),
.B1(n_1171),
.B2(n_1058),
.Y(n_1275)
);

NOR2x1_ASAP7_75t_SL g1276 ( 
.A(n_1041),
.B(n_1175),
.Y(n_1276)
);

A2O1A1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1076),
.A2(n_1053),
.B(n_1096),
.C(n_1060),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1089),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1058),
.B(n_1171),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1031),
.A2(n_1135),
.B(n_1165),
.Y(n_1280)
);

INVx1_ASAP7_75t_SL g1281 ( 
.A(n_1047),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_1061),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1117),
.A2(n_1146),
.B(n_1130),
.Y(n_1283)
);

INVxp67_ASAP7_75t_L g1284 ( 
.A(n_1134),
.Y(n_1284)
);

BUFx10_ASAP7_75t_L g1285 ( 
.A(n_1058),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1144),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1154),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1157),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1159),
.Y(n_1289)
);

INVx5_ASAP7_75t_L g1290 ( 
.A(n_1162),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1059),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1036),
.Y(n_1292)
);

OR2x2_ASAP7_75t_SL g1293 ( 
.A(n_1045),
.B(n_1028),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_L g1294 ( 
.A(n_1036),
.Y(n_1294)
);

O2A1O1Ixp5_ASAP7_75t_L g1295 ( 
.A1(n_1106),
.A2(n_1011),
.B(n_1009),
.C(n_1028),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1039),
.A2(n_974),
.B(n_865),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1039),
.A2(n_974),
.B(n_865),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1059),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1074),
.B(n_1067),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1145),
.B(n_1156),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1039),
.A2(n_974),
.B(n_1057),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1056),
.B(n_1116),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1145),
.B(n_1156),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1044),
.A2(n_1006),
.B1(n_909),
.B2(n_967),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1056),
.B(n_1116),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1046),
.B(n_1020),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1087),
.Y(n_1307)
);

INVx5_ASAP7_75t_L g1308 ( 
.A(n_1119),
.Y(n_1308)
);

OR2x2_ASAP7_75t_L g1309 ( 
.A(n_1160),
.B(n_1015),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1045),
.A2(n_983),
.B1(n_1028),
.B2(n_1065),
.Y(n_1310)
);

INVx3_ASAP7_75t_SL g1311 ( 
.A(n_1086),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1045),
.A2(n_983),
.B1(n_1028),
.B2(n_1065),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1039),
.A2(n_974),
.B(n_865),
.Y(n_1313)
);

BUFx6f_ASAP7_75t_L g1314 ( 
.A(n_1036),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1059),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1145),
.B(n_1156),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1039),
.A2(n_974),
.B(n_1057),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1056),
.B(n_1116),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1059),
.Y(n_1319)
);

INVx4_ASAP7_75t_L g1320 ( 
.A(n_1119),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1059),
.Y(n_1321)
);

AOI21xp33_ASAP7_75t_SL g1322 ( 
.A1(n_1126),
.A2(n_983),
.B(n_464),
.Y(n_1322)
);

OA21x2_ASAP7_75t_L g1323 ( 
.A1(n_1034),
.A2(n_1035),
.B(n_1057),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1056),
.B(n_1116),
.Y(n_1324)
);

INVx3_ASAP7_75t_SL g1325 ( 
.A(n_1086),
.Y(n_1325)
);

BUFx2_ASAP7_75t_SL g1326 ( 
.A(n_1125),
.Y(n_1326)
);

NOR2x1_ASAP7_75t_SL g1327 ( 
.A(n_1150),
.B(n_890),
.Y(n_1327)
);

BUFx2_ASAP7_75t_R g1328 ( 
.A(n_1311),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_L g1329 ( 
.A(n_1307),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1235),
.B(n_1310),
.Y(n_1330)
);

BUFx12f_ASAP7_75t_L g1331 ( 
.A(n_1179),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_SL g1332 ( 
.A1(n_1181),
.A2(n_1196),
.B1(n_1304),
.B2(n_1201),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1291),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1312),
.B(n_1186),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1242),
.Y(n_1335)
);

CKINVDCx11_ASAP7_75t_R g1336 ( 
.A(n_1325),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_1271),
.Y(n_1337)
);

NAND2x1p5_ASAP7_75t_L g1338 ( 
.A(n_1308),
.B(n_1267),
.Y(n_1338)
);

AOI222xp33_ASAP7_75t_L g1339 ( 
.A1(n_1232),
.A2(n_1306),
.B1(n_1209),
.B2(n_1180),
.C1(n_1299),
.C2(n_1198),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1186),
.B(n_1302),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1315),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1302),
.B(n_1305),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1183),
.A2(n_1213),
.B1(n_1210),
.B2(n_1222),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1280),
.A2(n_1283),
.B(n_1256),
.Y(n_1344)
);

BUFx3_ASAP7_75t_L g1345 ( 
.A(n_1188),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1304),
.A2(n_1267),
.B1(n_1305),
.B2(n_1324),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1318),
.B(n_1324),
.Y(n_1347)
);

INVx2_ASAP7_75t_SL g1348 ( 
.A(n_1308),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1318),
.A2(n_1309),
.B1(n_1241),
.B2(n_1204),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1194),
.B(n_1214),
.Y(n_1350)
);

INVx3_ASAP7_75t_L g1351 ( 
.A(n_1271),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_SL g1352 ( 
.A(n_1211),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1319),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1182),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1194),
.A2(n_1244),
.B1(n_1214),
.B2(n_1220),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1298),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1204),
.A2(n_1244),
.B1(n_1226),
.B2(n_1220),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1295),
.A2(n_1250),
.B(n_1322),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1219),
.B(n_1226),
.Y(n_1359)
);

INVx3_ASAP7_75t_L g1360 ( 
.A(n_1271),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1321),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1219),
.A2(n_1239),
.B1(n_1269),
.B2(n_1234),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1215),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1260),
.Y(n_1364)
);

BUFx6f_ASAP7_75t_L g1365 ( 
.A(n_1262),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_1308),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1231),
.Y(n_1367)
);

NAND2x1p5_ASAP7_75t_L g1368 ( 
.A(n_1320),
.B(n_1248),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_1240),
.Y(n_1369)
);

BUFx12f_ASAP7_75t_L g1370 ( 
.A(n_1184),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1239),
.A2(n_1266),
.B1(n_1190),
.B2(n_1247),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1225),
.B(n_1199),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1227),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1229),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1185),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1293),
.A2(n_1251),
.B1(n_1202),
.B2(n_1207),
.Y(n_1376)
);

CKINVDCx20_ASAP7_75t_R g1377 ( 
.A(n_1197),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1192),
.Y(n_1378)
);

OA21x2_ASAP7_75t_L g1379 ( 
.A1(n_1243),
.A2(n_1236),
.B(n_1230),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1266),
.A2(n_1247),
.B1(n_1272),
.B2(n_1217),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1195),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1260),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1266),
.A2(n_1205),
.B1(n_1323),
.B2(n_1259),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1276),
.B(n_1249),
.Y(n_1384)
);

AO21x1_ASAP7_75t_L g1385 ( 
.A1(n_1237),
.A2(n_1205),
.B(n_1249),
.Y(n_1385)
);

BUFx6f_ASAP7_75t_SL g1386 ( 
.A(n_1257),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_1326),
.Y(n_1387)
);

INVx3_ASAP7_75t_L g1388 ( 
.A(n_1263),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_SL g1389 ( 
.A1(n_1323),
.A2(n_1225),
.B1(n_1206),
.B2(n_1218),
.Y(n_1389)
);

OAI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1212),
.A2(n_1202),
.B1(n_1200),
.B2(n_1238),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1199),
.B(n_1187),
.Y(n_1391)
);

NAND2x1p5_ASAP7_75t_L g1392 ( 
.A(n_1320),
.B(n_1263),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_SL g1393 ( 
.A1(n_1261),
.A2(n_1200),
.B1(n_1233),
.B2(n_1228),
.Y(n_1393)
);

OAI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1261),
.A2(n_1287),
.B1(n_1273),
.B2(n_1268),
.Y(n_1394)
);

BUFx2_ASAP7_75t_L g1395 ( 
.A(n_1279),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1275),
.B(n_1203),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_SL g1397 ( 
.A1(n_1223),
.A2(n_1264),
.B1(n_1316),
.B2(n_1193),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1252),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1187),
.A2(n_1300),
.B1(n_1303),
.B2(n_1193),
.Y(n_1399)
);

INVx4_ASAP7_75t_L g1400 ( 
.A(n_1257),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_SL g1401 ( 
.A(n_1257),
.Y(n_1401)
);

AOI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1301),
.A2(n_1317),
.B(n_1296),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1300),
.Y(n_1403)
);

BUFx2_ASAP7_75t_L g1404 ( 
.A(n_1265),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1303),
.A2(n_1316),
.B1(n_1285),
.B2(n_1253),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1216),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1285),
.A2(n_1208),
.B1(n_1265),
.B2(n_1289),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1189),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1208),
.A2(n_1288),
.B1(n_1191),
.B2(n_1224),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1224),
.A2(n_1258),
.B1(n_1270),
.B2(n_1278),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1297),
.A2(n_1313),
.B(n_1277),
.Y(n_1411)
);

OA21x2_ASAP7_75t_L g1412 ( 
.A1(n_1254),
.A2(n_1286),
.B(n_1284),
.Y(n_1412)
);

NAND2x1p5_ASAP7_75t_L g1413 ( 
.A(n_1221),
.B(n_1314),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1258),
.A2(n_1245),
.B1(n_1255),
.B2(n_1281),
.Y(n_1414)
);

BUFx6f_ASAP7_75t_L g1415 ( 
.A(n_1246),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1246),
.Y(n_1416)
);

AO21x2_ASAP7_75t_L g1417 ( 
.A1(n_1290),
.A2(n_1327),
.B(n_1282),
.Y(n_1417)
);

AOI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1290),
.A2(n_1282),
.B(n_1189),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_SL g1419 ( 
.A1(n_1290),
.A2(n_1282),
.B(n_1246),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1292),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_SL g1421 ( 
.A1(n_1294),
.A2(n_1181),
.B1(n_611),
.B2(n_995),
.Y(n_1421)
);

OA21x2_ASAP7_75t_L g1422 ( 
.A1(n_1290),
.A2(n_1243),
.B(n_1236),
.Y(n_1422)
);

INVx8_ASAP7_75t_L g1423 ( 
.A(n_1308),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1291),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1181),
.A2(n_983),
.B1(n_1028),
.B2(n_1065),
.Y(n_1425)
);

AOI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1280),
.A2(n_1283),
.B(n_1274),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1291),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1181),
.A2(n_983),
.B1(n_1028),
.B2(n_1065),
.Y(n_1428)
);

INVx8_ASAP7_75t_L g1429 ( 
.A(n_1308),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1291),
.Y(n_1430)
);

OAI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1181),
.A2(n_1028),
.B1(n_838),
.B2(n_611),
.Y(n_1431)
);

INVxp33_ASAP7_75t_L g1432 ( 
.A(n_1309),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1225),
.B(n_1234),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1181),
.A2(n_983),
.B1(n_1028),
.B2(n_1065),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1291),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1291),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_SL g1437 ( 
.A1(n_1181),
.A2(n_611),
.B1(n_995),
.B2(n_983),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1291),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_1307),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1291),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1181),
.A2(n_983),
.B1(n_1028),
.B2(n_1065),
.Y(n_1441)
);

AOI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1280),
.A2(n_1283),
.B(n_1274),
.Y(n_1442)
);

BUFx2_ASAP7_75t_L g1443 ( 
.A(n_1260),
.Y(n_1443)
);

BUFx4_ASAP7_75t_SL g1444 ( 
.A(n_1240),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1181),
.A2(n_983),
.B1(n_1028),
.B2(n_1065),
.Y(n_1445)
);

OR2x6_ASAP7_75t_L g1446 ( 
.A(n_1266),
.B(n_1183),
.Y(n_1446)
);

CKINVDCx20_ASAP7_75t_R g1447 ( 
.A(n_1240),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1291),
.Y(n_1448)
);

AO21x1_ASAP7_75t_L g1449 ( 
.A1(n_1237),
.A2(n_1094),
.B(n_1122),
.Y(n_1449)
);

OAI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1295),
.A2(n_1028),
.B(n_1009),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1291),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_SL g1452 ( 
.A1(n_1181),
.A2(n_611),
.B1(n_995),
.B2(n_983),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1181),
.B(n_1186),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_1444),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1426),
.A2(n_1442),
.B(n_1344),
.Y(n_1455)
);

NOR2xp33_ASAP7_75t_L g1456 ( 
.A(n_1432),
.B(n_1453),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1350),
.B(n_1359),
.Y(n_1457)
);

INVxp67_ASAP7_75t_L g1458 ( 
.A(n_1329),
.Y(n_1458)
);

INVx1_ASAP7_75t_SL g1459 ( 
.A(n_1345),
.Y(n_1459)
);

AO21x2_ASAP7_75t_L g1460 ( 
.A1(n_1411),
.A2(n_1402),
.B(n_1358),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1395),
.B(n_1396),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1361),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1354),
.Y(n_1463)
);

INVxp67_ASAP7_75t_SL g1464 ( 
.A(n_1338),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1395),
.B(n_1396),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1426),
.A2(n_1442),
.B(n_1344),
.Y(n_1466)
);

INVx2_ASAP7_75t_SL g1467 ( 
.A(n_1338),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1439),
.Y(n_1468)
);

BUFx6f_ASAP7_75t_L g1469 ( 
.A(n_1365),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1350),
.B(n_1359),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1340),
.B(n_1342),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1437),
.A2(n_1452),
.B1(n_1445),
.B2(n_1434),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1446),
.B(n_1384),
.Y(n_1473)
);

AND2x4_ASAP7_75t_L g1474 ( 
.A(n_1382),
.B(n_1388),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1330),
.B(n_1384),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1446),
.B(n_1383),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1330),
.B(n_1446),
.Y(n_1477)
);

BUFx2_ASAP7_75t_L g1478 ( 
.A(n_1364),
.Y(n_1478)
);

CKINVDCx8_ASAP7_75t_R g1479 ( 
.A(n_1365),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_SL g1480 ( 
.A(n_1328),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1335),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1356),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1443),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1446),
.B(n_1334),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1385),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1380),
.B(n_1349),
.Y(n_1486)
);

CKINVDCx16_ASAP7_75t_R g1487 ( 
.A(n_1369),
.Y(n_1487)
);

AO21x2_ASAP7_75t_L g1488 ( 
.A1(n_1394),
.A2(n_1449),
.B(n_1450),
.Y(n_1488)
);

INVx3_ASAP7_75t_L g1489 ( 
.A(n_1418),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1334),
.B(n_1343),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1385),
.B(n_1371),
.Y(n_1491)
);

BUFx8_ASAP7_75t_SL g1492 ( 
.A(n_1369),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1412),
.Y(n_1493)
);

BUFx3_ASAP7_75t_L g1494 ( 
.A(n_1345),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_L g1495 ( 
.A(n_1365),
.Y(n_1495)
);

OR2x6_ASAP7_75t_L g1496 ( 
.A(n_1443),
.B(n_1423),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1332),
.B(n_1382),
.Y(n_1497)
);

OR2x6_ASAP7_75t_L g1498 ( 
.A(n_1423),
.B(n_1429),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1412),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1346),
.B(n_1376),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1347),
.B(n_1425),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1422),
.A2(n_1379),
.B(n_1419),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_1336),
.Y(n_1503)
);

OA21x2_ASAP7_75t_L g1504 ( 
.A1(n_1410),
.A2(n_1409),
.B(n_1414),
.Y(n_1504)
);

AO21x2_ASAP7_75t_L g1505 ( 
.A1(n_1419),
.A2(n_1417),
.B(n_1431),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1422),
.A2(n_1379),
.B(n_1351),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1363),
.Y(n_1507)
);

BUFx12f_ASAP7_75t_L g1508 ( 
.A(n_1336),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1428),
.B(n_1441),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1367),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1355),
.B(n_1432),
.Y(n_1511)
);

OAI21x1_ASAP7_75t_L g1512 ( 
.A1(n_1422),
.A2(n_1379),
.B(n_1360),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1333),
.Y(n_1513)
);

OA21x2_ASAP7_75t_L g1514 ( 
.A1(n_1407),
.A2(n_1357),
.B(n_1362),
.Y(n_1514)
);

AO21x2_ASAP7_75t_L g1515 ( 
.A1(n_1417),
.A2(n_1390),
.B(n_1398),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1341),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1353),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1424),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1427),
.Y(n_1519)
);

AOI21xp33_ASAP7_75t_L g1520 ( 
.A1(n_1339),
.A2(n_1421),
.B(n_1397),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_SL g1521 ( 
.A1(n_1405),
.A2(n_1451),
.B(n_1436),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1393),
.B(n_1404),
.Y(n_1522)
);

BUFx2_ASAP7_75t_L g1523 ( 
.A(n_1337),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1430),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1435),
.Y(n_1525)
);

INVx1_ASAP7_75t_SL g1526 ( 
.A(n_1447),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1373),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1438),
.B(n_1448),
.Y(n_1528)
);

CKINVDCx20_ASAP7_75t_R g1529 ( 
.A(n_1447),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1337),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1433),
.B(n_1351),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1374),
.B(n_1381),
.Y(n_1532)
);

BUFx2_ASAP7_75t_L g1533 ( 
.A(n_1368),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1484),
.B(n_1389),
.Y(n_1534)
);

INVxp67_ASAP7_75t_SL g1535 ( 
.A(n_1485),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_SL g1536 ( 
.A(n_1472),
.B(n_1368),
.Y(n_1536)
);

INVx3_ASAP7_75t_L g1537 ( 
.A(n_1506),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1457),
.B(n_1440),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1461),
.B(n_1378),
.Y(n_1539)
);

INVx1_ASAP7_75t_SL g1540 ( 
.A(n_1461),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1484),
.B(n_1375),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1465),
.Y(n_1542)
);

BUFx3_ASAP7_75t_L g1543 ( 
.A(n_1479),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1477),
.B(n_1433),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1477),
.B(n_1406),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1465),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1485),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1493),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1512),
.B(n_1366),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1499),
.Y(n_1550)
);

AOI221xp5_ASAP7_75t_L g1551 ( 
.A1(n_1520),
.A2(n_1509),
.B1(n_1501),
.B2(n_1490),
.C(n_1500),
.Y(n_1551)
);

INVx2_ASAP7_75t_R g1552 ( 
.A(n_1530),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1479),
.Y(n_1553)
);

BUFx3_ASAP7_75t_L g1554 ( 
.A(n_1474),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1515),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1511),
.B(n_1403),
.Y(n_1556)
);

AOI221xp5_ASAP7_75t_L g1557 ( 
.A1(n_1490),
.A2(n_1387),
.B1(n_1399),
.B2(n_1391),
.C(n_1372),
.Y(n_1557)
);

BUFx3_ASAP7_75t_L g1558 ( 
.A(n_1474),
.Y(n_1558)
);

INVxp67_ASAP7_75t_L g1559 ( 
.A(n_1515),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1475),
.B(n_1460),
.Y(n_1560)
);

OAI321xp33_ASAP7_75t_L g1561 ( 
.A1(n_1500),
.A2(n_1392),
.A3(n_1348),
.B1(n_1366),
.B2(n_1416),
.C(n_1413),
.Y(n_1561)
);

AOI21xp33_ASAP7_75t_L g1562 ( 
.A1(n_1488),
.A2(n_1429),
.B(n_1348),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1475),
.B(n_1416),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1460),
.B(n_1392),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1488),
.B(n_1408),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1488),
.B(n_1415),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1473),
.B(n_1415),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1473),
.B(n_1502),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1476),
.B(n_1415),
.Y(n_1569)
);

NAND4xp25_ASAP7_75t_L g1570 ( 
.A(n_1551),
.B(n_1456),
.C(n_1471),
.D(n_1458),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_SL g1571 ( 
.A1(n_1534),
.A2(n_1486),
.B1(n_1497),
.B2(n_1491),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1541),
.B(n_1468),
.Y(n_1572)
);

NAND3xp33_ASAP7_75t_L g1573 ( 
.A(n_1551),
.B(n_1491),
.C(n_1497),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1541),
.B(n_1470),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1541),
.B(n_1527),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1540),
.B(n_1463),
.Y(n_1576)
);

AOI221xp5_ASAP7_75t_L g1577 ( 
.A1(n_1536),
.A2(n_1521),
.B1(n_1513),
.B2(n_1482),
.C(n_1507),
.Y(n_1577)
);

OAI221xp5_ASAP7_75t_L g1578 ( 
.A1(n_1536),
.A2(n_1486),
.B1(n_1526),
.B2(n_1459),
.C(n_1494),
.Y(n_1578)
);

OAI21xp33_ASAP7_75t_L g1579 ( 
.A1(n_1556),
.A2(n_1476),
.B(n_1522),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1557),
.A2(n_1556),
.B1(n_1534),
.B2(n_1514),
.Y(n_1580)
);

NAND3xp33_ASAP7_75t_L g1581 ( 
.A(n_1557),
.B(n_1532),
.C(n_1510),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_SL g1582 ( 
.A(n_1561),
.B(n_1487),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1560),
.B(n_1515),
.Y(n_1583)
);

OA21x2_ASAP7_75t_L g1584 ( 
.A1(n_1559),
.A2(n_1466),
.B(n_1455),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_L g1585 ( 
.A(n_1538),
.B(n_1492),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1548),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1542),
.B(n_1481),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1534),
.A2(n_1514),
.B1(n_1508),
.B2(n_1531),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1560),
.B(n_1567),
.Y(n_1589)
);

NAND3xp33_ASAP7_75t_L g1590 ( 
.A(n_1565),
.B(n_1522),
.C(n_1514),
.Y(n_1590)
);

OAI221xp5_ASAP7_75t_SL g1591 ( 
.A1(n_1559),
.A2(n_1464),
.B1(n_1496),
.B2(n_1494),
.C(n_1533),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1560),
.B(n_1505),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1546),
.B(n_1516),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1534),
.A2(n_1514),
.B1(n_1569),
.B2(n_1508),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1560),
.B(n_1505),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1569),
.A2(n_1531),
.B1(n_1521),
.B2(n_1505),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1543),
.A2(n_1480),
.B1(n_1529),
.B2(n_1387),
.Y(n_1597)
);

OAI221xp5_ASAP7_75t_SL g1598 ( 
.A1(n_1555),
.A2(n_1496),
.B1(n_1533),
.B2(n_1483),
.C(n_1478),
.Y(n_1598)
);

OAI21xp33_ASAP7_75t_L g1599 ( 
.A1(n_1565),
.A2(n_1528),
.B(n_1503),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1538),
.B(n_1517),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1567),
.B(n_1489),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1563),
.B(n_1518),
.Y(n_1602)
);

NAND3xp33_ASAP7_75t_L g1603 ( 
.A(n_1555),
.B(n_1524),
.C(n_1518),
.Y(n_1603)
);

NAND3xp33_ASAP7_75t_L g1604 ( 
.A(n_1565),
.B(n_1519),
.C(n_1524),
.Y(n_1604)
);

NAND2xp33_ASAP7_75t_SL g1605 ( 
.A(n_1539),
.B(n_1503),
.Y(n_1605)
);

NOR3xp33_ASAP7_75t_SL g1606 ( 
.A(n_1561),
.B(n_1454),
.C(n_1530),
.Y(n_1606)
);

AOI21xp5_ASAP7_75t_SL g1607 ( 
.A1(n_1543),
.A2(n_1496),
.B(n_1498),
.Y(n_1607)
);

NAND3xp33_ASAP7_75t_L g1608 ( 
.A(n_1562),
.B(n_1525),
.C(n_1504),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1568),
.B(n_1523),
.Y(n_1609)
);

NAND3xp33_ASAP7_75t_L g1610 ( 
.A(n_1562),
.B(n_1467),
.C(n_1462),
.Y(n_1610)
);

OAI21xp33_ASAP7_75t_SL g1611 ( 
.A1(n_1566),
.A2(n_1467),
.B(n_1535),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1568),
.B(n_1523),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1568),
.B(n_1545),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1613),
.B(n_1589),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1583),
.B(n_1547),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1570),
.B(n_1539),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1613),
.B(n_1552),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1589),
.B(n_1552),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1592),
.B(n_1552),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1586),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1595),
.B(n_1552),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1586),
.Y(n_1622)
);

AOI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1573),
.A2(n_1504),
.B1(n_1529),
.B2(n_1545),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1601),
.B(n_1537),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1595),
.B(n_1552),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1593),
.B(n_1576),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1584),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1584),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1590),
.B(n_1548),
.Y(n_1629)
);

AOI22xp33_ASAP7_75t_SL g1630 ( 
.A1(n_1581),
.A2(n_1553),
.B1(n_1543),
.B2(n_1504),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1584),
.Y(n_1631)
);

NOR2xp33_ASAP7_75t_L g1632 ( 
.A(n_1578),
.B(n_1544),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1584),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1609),
.B(n_1566),
.Y(n_1634)
);

AND2x2_ASAP7_75t_SL g1635 ( 
.A(n_1580),
.B(n_1564),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1612),
.B(n_1566),
.Y(n_1636)
);

INVxp67_ASAP7_75t_L g1637 ( 
.A(n_1610),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1604),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1604),
.Y(n_1639)
);

BUFx2_ASAP7_75t_L g1640 ( 
.A(n_1611),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1603),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1608),
.B(n_1537),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1603),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1611),
.B(n_1550),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1600),
.B(n_1535),
.Y(n_1645)
);

INVx3_ASAP7_75t_L g1646 ( 
.A(n_1624),
.Y(n_1646)
);

OAI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1630),
.A2(n_1571),
.B1(n_1582),
.B2(n_1606),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1637),
.B(n_1579),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1644),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1622),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1622),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1622),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1620),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1644),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1614),
.B(n_1554),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1637),
.B(n_1579),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1616),
.B(n_1574),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1620),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1614),
.B(n_1554),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1614),
.B(n_1554),
.Y(n_1660)
);

INVxp67_ASAP7_75t_SL g1661 ( 
.A(n_1640),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1644),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1620),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1644),
.B(n_1549),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1638),
.B(n_1572),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1614),
.B(n_1554),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1620),
.Y(n_1667)
);

INVx3_ASAP7_75t_L g1668 ( 
.A(n_1624),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1640),
.B(n_1558),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1640),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1638),
.B(n_1602),
.Y(n_1671)
);

OAI21xp33_ASAP7_75t_L g1672 ( 
.A1(n_1623),
.A2(n_1594),
.B(n_1599),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1617),
.B(n_1549),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1616),
.B(n_1575),
.Y(n_1674)
);

NOR2x1_ASAP7_75t_L g1675 ( 
.A(n_1643),
.B(n_1607),
.Y(n_1675)
);

NAND2xp33_ASAP7_75t_SL g1676 ( 
.A(n_1643),
.B(n_1454),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1615),
.B(n_1587),
.Y(n_1677)
);

INVx2_ASAP7_75t_SL g1678 ( 
.A(n_1669),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1669),
.B(n_1617),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1650),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1650),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1649),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1671),
.B(n_1638),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1651),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1661),
.B(n_1617),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1651),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1648),
.B(n_1632),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1670),
.B(n_1618),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1675),
.B(n_1618),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1649),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1648),
.B(n_1632),
.Y(n_1691)
);

OAI22xp33_ASAP7_75t_R g1692 ( 
.A1(n_1647),
.A2(n_1643),
.B1(n_1641),
.B2(n_1629),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1675),
.B(n_1618),
.Y(n_1693)
);

AOI211xp5_ASAP7_75t_L g1694 ( 
.A1(n_1647),
.A2(n_1597),
.B(n_1623),
.C(n_1591),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1671),
.B(n_1639),
.Y(n_1695)
);

OAI21xp33_ASAP7_75t_SL g1696 ( 
.A1(n_1656),
.A2(n_1623),
.B(n_1635),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1655),
.B(n_1634),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1649),
.B(n_1639),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1652),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1652),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1654),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1654),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_L g1703 ( 
.A(n_1657),
.B(n_1585),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1656),
.B(n_1630),
.Y(n_1704)
);

INVx2_ASAP7_75t_SL g1705 ( 
.A(n_1646),
.Y(n_1705)
);

INVx2_ASAP7_75t_SL g1706 ( 
.A(n_1646),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1667),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1667),
.Y(n_1708)
);

INVx2_ASAP7_75t_SL g1709 ( 
.A(n_1646),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1655),
.B(n_1634),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1667),
.Y(n_1711)
);

AO22x1_ASAP7_75t_L g1712 ( 
.A1(n_1676),
.A2(n_1643),
.B1(n_1641),
.B2(n_1639),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1653),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1659),
.B(n_1636),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1674),
.B(n_1665),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1654),
.B(n_1642),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1665),
.B(n_1626),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1677),
.B(n_1626),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1677),
.B(n_1645),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1659),
.B(n_1636),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1687),
.B(n_1672),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1691),
.B(n_1672),
.Y(n_1722)
);

AO21x2_ASAP7_75t_L g1723 ( 
.A1(n_1692),
.A2(n_1641),
.B(n_1662),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1716),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1716),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1680),
.Y(n_1726)
);

INVxp33_ASAP7_75t_L g1727 ( 
.A(n_1703),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1689),
.B(n_1662),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1715),
.B(n_1660),
.Y(n_1729)
);

INVxp67_ASAP7_75t_L g1730 ( 
.A(n_1678),
.Y(n_1730)
);

NAND4xp25_ASAP7_75t_L g1731 ( 
.A(n_1694),
.B(n_1588),
.C(n_1599),
.D(n_1577),
.Y(n_1731)
);

INVxp67_ASAP7_75t_SL g1732 ( 
.A(n_1712),
.Y(n_1732)
);

CKINVDCx16_ASAP7_75t_R g1733 ( 
.A(n_1689),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1692),
.A2(n_1696),
.B1(n_1635),
.B2(n_1704),
.Y(n_1734)
);

AOI22xp33_ASAP7_75t_L g1735 ( 
.A1(n_1696),
.A2(n_1635),
.B1(n_1605),
.B2(n_1608),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1683),
.B(n_1662),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1693),
.B(n_1664),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1717),
.B(n_1660),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1680),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1683),
.B(n_1629),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1681),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1712),
.B(n_1666),
.Y(n_1742)
);

INVxp33_ASAP7_75t_SL g1743 ( 
.A(n_1693),
.Y(n_1743)
);

NOR2xp33_ASAP7_75t_L g1744 ( 
.A(n_1718),
.B(n_1331),
.Y(n_1744)
);

INVx1_ASAP7_75t_SL g1745 ( 
.A(n_1678),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1719),
.B(n_1331),
.Y(n_1746)
);

INVx1_ASAP7_75t_SL g1747 ( 
.A(n_1685),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1681),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1697),
.B(n_1664),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1684),
.Y(n_1750)
);

INVx2_ASAP7_75t_SL g1751 ( 
.A(n_1705),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1694),
.B(n_1666),
.Y(n_1752)
);

INVx3_ASAP7_75t_L g1753 ( 
.A(n_1716),
.Y(n_1753)
);

INVx1_ASAP7_75t_SL g1754 ( 
.A(n_1685),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1684),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1695),
.B(n_1629),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1726),
.Y(n_1757)
);

INVxp67_ASAP7_75t_L g1758 ( 
.A(n_1732),
.Y(n_1758)
);

AOI322xp5_ASAP7_75t_L g1759 ( 
.A1(n_1734),
.A2(n_1721),
.A3(n_1722),
.B1(n_1735),
.B2(n_1752),
.C1(n_1733),
.C2(n_1754),
.Y(n_1759)
);

OAI32xp33_ASAP7_75t_L g1760 ( 
.A1(n_1733),
.A2(n_1695),
.A3(n_1698),
.B1(n_1688),
.B2(n_1679),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1723),
.Y(n_1761)
);

OAI322xp33_ASAP7_75t_L g1762 ( 
.A1(n_1747),
.A2(n_1698),
.A3(n_1690),
.B1(n_1682),
.B2(n_1701),
.C1(n_1702),
.C2(n_1686),
.Y(n_1762)
);

O2A1O1Ixp33_ASAP7_75t_L g1763 ( 
.A1(n_1723),
.A2(n_1642),
.B(n_1688),
.C(n_1705),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1737),
.B(n_1724),
.Y(n_1764)
);

AOI211xp5_ASAP7_75t_L g1765 ( 
.A1(n_1731),
.A2(n_1598),
.B(n_1642),
.C(n_1607),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1726),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1739),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1739),
.Y(n_1768)
);

AOI21xp33_ASAP7_75t_SL g1769 ( 
.A1(n_1727),
.A2(n_1635),
.B(n_1706),
.Y(n_1769)
);

BUFx3_ASAP7_75t_L g1770 ( 
.A(n_1743),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1737),
.B(n_1679),
.Y(n_1771)
);

AOI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1743),
.A2(n_1605),
.B1(n_1642),
.B2(n_1716),
.Y(n_1772)
);

AOI32xp33_ASAP7_75t_L g1773 ( 
.A1(n_1742),
.A2(n_1642),
.A3(n_1619),
.B1(n_1621),
.B2(n_1625),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1745),
.B(n_1697),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1753),
.Y(n_1775)
);

INVxp67_ASAP7_75t_L g1776 ( 
.A(n_1746),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1729),
.B(n_1710),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1723),
.A2(n_1581),
.B1(n_1642),
.B2(n_1596),
.Y(n_1778)
);

AOI21xp5_ASAP7_75t_L g1779 ( 
.A1(n_1744),
.A2(n_1709),
.B(n_1706),
.Y(n_1779)
);

AOI22xp33_ASAP7_75t_L g1780 ( 
.A1(n_1730),
.A2(n_1690),
.B1(n_1701),
.B2(n_1682),
.Y(n_1780)
);

OAI221xp5_ASAP7_75t_L g1781 ( 
.A1(n_1738),
.A2(n_1709),
.B1(n_1686),
.B2(n_1700),
.C(n_1699),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1741),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1736),
.B(n_1710),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1757),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1766),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1767),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1758),
.B(n_1728),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1770),
.B(n_1728),
.Y(n_1788)
);

INVx3_ASAP7_75t_L g1789 ( 
.A(n_1770),
.Y(n_1789)
);

INVxp33_ASAP7_75t_L g1790 ( 
.A(n_1761),
.Y(n_1790)
);

INVxp67_ASAP7_75t_L g1791 ( 
.A(n_1774),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1768),
.Y(n_1792)
);

AND2x4_ASAP7_75t_L g1793 ( 
.A(n_1764),
.B(n_1751),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1759),
.B(n_1724),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1764),
.B(n_1725),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1771),
.B(n_1753),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1761),
.B(n_1783),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1782),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1771),
.B(n_1753),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_SL g1800 ( 
.A(n_1776),
.B(n_1725),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1775),
.Y(n_1801)
);

INVx2_ASAP7_75t_SL g1802 ( 
.A(n_1775),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1769),
.B(n_1749),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1762),
.Y(n_1804)
);

INVxp67_ASAP7_75t_SL g1805 ( 
.A(n_1789),
.Y(n_1805)
);

OAI221xp5_ASAP7_75t_L g1806 ( 
.A1(n_1794),
.A2(n_1778),
.B1(n_1765),
.B2(n_1779),
.C(n_1772),
.Y(n_1806)
);

AOI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1800),
.A2(n_1763),
.B(n_1760),
.Y(n_1807)
);

OAI31xp33_ASAP7_75t_L g1808 ( 
.A1(n_1804),
.A2(n_1778),
.A3(n_1781),
.B(n_1780),
.Y(n_1808)
);

NOR3x1_ASAP7_75t_L g1809 ( 
.A(n_1788),
.B(n_1751),
.C(n_1777),
.Y(n_1809)
);

OAI221xp5_ASAP7_75t_L g1810 ( 
.A1(n_1791),
.A2(n_1773),
.B1(n_1780),
.B2(n_1756),
.C(n_1740),
.Y(n_1810)
);

AOI221xp5_ASAP7_75t_L g1811 ( 
.A1(n_1790),
.A2(n_1748),
.B1(n_1755),
.B2(n_1750),
.C(n_1741),
.Y(n_1811)
);

OAI221xp5_ASAP7_75t_L g1812 ( 
.A1(n_1789),
.A2(n_1756),
.B1(n_1740),
.B2(n_1736),
.C(n_1750),
.Y(n_1812)
);

AOI21xp33_ASAP7_75t_SL g1813 ( 
.A1(n_1789),
.A2(n_1755),
.B(n_1748),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1803),
.B(n_1749),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1802),
.Y(n_1815)
);

OAI221xp5_ASAP7_75t_SL g1816 ( 
.A1(n_1803),
.A2(n_1702),
.B1(n_1699),
.B2(n_1700),
.C(n_1711),
.Y(n_1816)
);

NOR4xp25_ASAP7_75t_SL g1817 ( 
.A(n_1801),
.B(n_1707),
.C(n_1708),
.D(n_1711),
.Y(n_1817)
);

AOI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1790),
.A2(n_1377),
.B(n_1702),
.Y(n_1818)
);

NOR2x1_ASAP7_75t_L g1819 ( 
.A(n_1815),
.B(n_1797),
.Y(n_1819)
);

NOR2x1_ASAP7_75t_L g1820 ( 
.A(n_1818),
.B(n_1797),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1805),
.B(n_1787),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1807),
.B(n_1793),
.Y(n_1822)
);

NAND4xp75_ASAP7_75t_L g1823 ( 
.A(n_1809),
.B(n_1802),
.C(n_1799),
.D(n_1796),
.Y(n_1823)
);

AOI211xp5_ASAP7_75t_L g1824 ( 
.A1(n_1808),
.A2(n_1795),
.B(n_1793),
.C(n_1784),
.Y(n_1824)
);

NAND3xp33_ASAP7_75t_L g1825 ( 
.A(n_1818),
.B(n_1786),
.C(n_1785),
.Y(n_1825)
);

OAI211xp5_ASAP7_75t_SL g1826 ( 
.A1(n_1806),
.A2(n_1798),
.B(n_1792),
.C(n_1793),
.Y(n_1826)
);

NAND3xp33_ASAP7_75t_L g1827 ( 
.A(n_1811),
.B(n_1813),
.C(n_1812),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1814),
.Y(n_1828)
);

AND2x4_ASAP7_75t_L g1829 ( 
.A(n_1816),
.B(n_1796),
.Y(n_1829)
);

AOI22xp33_ASAP7_75t_L g1830 ( 
.A1(n_1810),
.A2(n_1799),
.B1(n_1707),
.B2(n_1708),
.Y(n_1830)
);

AOI211x1_ASAP7_75t_L g1831 ( 
.A1(n_1827),
.A2(n_1817),
.B(n_1713),
.C(n_1714),
.Y(n_1831)
);

AOI211xp5_ASAP7_75t_L g1832 ( 
.A1(n_1826),
.A2(n_1352),
.B(n_1713),
.C(n_1562),
.Y(n_1832)
);

NOR2xp33_ASAP7_75t_L g1833 ( 
.A(n_1821),
.B(n_1370),
.Y(n_1833)
);

NOR2xp67_ASAP7_75t_L g1834 ( 
.A(n_1825),
.B(n_1370),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1820),
.B(n_1720),
.Y(n_1835)
);

AOI21xp33_ASAP7_75t_SL g1836 ( 
.A1(n_1822),
.A2(n_1377),
.B(n_1664),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_SL g1837 ( 
.A(n_1836),
.B(n_1829),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1835),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1831),
.Y(n_1839)
);

AOI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1833),
.A2(n_1828),
.B1(n_1823),
.B2(n_1829),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1834),
.Y(n_1841)
);

NOR2xp67_ASAP7_75t_L g1842 ( 
.A(n_1832),
.B(n_1830),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1835),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1839),
.B(n_1819),
.Y(n_1844)
);

AOI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1837),
.A2(n_1824),
.B(n_1658),
.Y(n_1845)
);

AND2x4_ASAP7_75t_L g1846 ( 
.A(n_1841),
.B(n_1714),
.Y(n_1846)
);

OAI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1840),
.A2(n_1646),
.B1(n_1668),
.B2(n_1664),
.Y(n_1847)
);

NOR2x1_ASAP7_75t_L g1848 ( 
.A(n_1838),
.B(n_1668),
.Y(n_1848)
);

AOI221xp5_ASAP7_75t_L g1849 ( 
.A1(n_1843),
.A2(n_1633),
.B1(n_1631),
.B2(n_1628),
.C(n_1627),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1846),
.Y(n_1850)
);

NOR2x1_ASAP7_75t_L g1851 ( 
.A(n_1844),
.B(n_1842),
.Y(n_1851)
);

INVx2_ASAP7_75t_SL g1852 ( 
.A(n_1848),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1850),
.A2(n_1851),
.B1(n_1847),
.B2(n_1845),
.Y(n_1853)
);

NAND3xp33_ASAP7_75t_SL g1854 ( 
.A(n_1853),
.B(n_1852),
.C(n_1849),
.Y(n_1854)
);

OAI21xp5_ASAP7_75t_L g1855 ( 
.A1(n_1854),
.A2(n_1668),
.B(n_1720),
.Y(n_1855)
);

AOI22xp33_ASAP7_75t_L g1856 ( 
.A1(n_1854),
.A2(n_1668),
.B1(n_1386),
.B2(n_1401),
.Y(n_1856)
);

OAI21xp5_ASAP7_75t_L g1857 ( 
.A1(n_1856),
.A2(n_1658),
.B(n_1653),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1855),
.B(n_1663),
.Y(n_1858)
);

BUFx2_ASAP7_75t_L g1859 ( 
.A(n_1858),
.Y(n_1859)
);

CKINVDCx20_ASAP7_75t_R g1860 ( 
.A(n_1857),
.Y(n_1860)
);

OAI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1860),
.A2(n_1859),
.B(n_1663),
.Y(n_1861)
);

XNOR2xp5_ASAP7_75t_L g1862 ( 
.A(n_1861),
.B(n_1413),
.Y(n_1862)
);

AOI221xp5_ASAP7_75t_L g1863 ( 
.A1(n_1862),
.A2(n_1386),
.B1(n_1401),
.B2(n_1400),
.C(n_1673),
.Y(n_1863)
);

AOI211xp5_ASAP7_75t_L g1864 ( 
.A1(n_1863),
.A2(n_1495),
.B(n_1469),
.C(n_1420),
.Y(n_1864)
);


endmodule