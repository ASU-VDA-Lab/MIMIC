module fake_jpeg_1774_n_36 (n_3, n_2, n_1, n_0, n_4, n_36);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g5 ( 
.A(n_0),
.Y(n_5)
);

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_4),
.Y(n_6)
);

INVx3_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_6),
.B(n_0),
.Y(n_10)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_10),
.B(n_12),
.Y(n_15)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx4_ASAP7_75t_SL g17 ( 
.A(n_11),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_SL g12 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_12)
);

CKINVDCx9p33_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_5),
.A2(n_8),
.B1(n_9),
.B2(n_3),
.Y(n_14)
);

AOI22xp33_ASAP7_75t_L g18 ( 
.A1(n_14),
.A2(n_8),
.B1(n_9),
.B2(n_3),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_18),
.A2(n_12),
.B(n_13),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_SL g19 ( 
.A(n_15),
.B(n_10),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_20),
.C(n_22),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_10),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_21),
.A2(n_16),
.B1(n_17),
.B2(n_12),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_14),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_14),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_17),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_11),
.B1(n_2),
.B2(n_3),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_26),
.C(n_23),
.Y(n_31)
);

NOR2x1_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_25),
.Y(n_30)
);

OAI211xp5_ASAP7_75t_SL g33 ( 
.A1(n_30),
.A2(n_11),
.B(n_1),
.C(n_4),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_28),
.B(n_27),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_34),
.A2(n_33),
.B(n_11),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_4),
.Y(n_36)
);


endmodule