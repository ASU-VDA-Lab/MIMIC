module fake_netlist_6_1362_n_1913 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1913);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1913;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_811;
wire n_683;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1851;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g169 ( 
.A(n_32),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_89),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_66),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_80),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_5),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_144),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_88),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_61),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_77),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_46),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_27),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_152),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_97),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_130),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_135),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_37),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_114),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_91),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_53),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_14),
.Y(n_188)
);

BUFx10_ASAP7_75t_L g189 ( 
.A(n_17),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_11),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_21),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_155),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_25),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_39),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_154),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_64),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_44),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_28),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_16),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_120),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_56),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_22),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_139),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_5),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_60),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_22),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_41),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_151),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_105),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_47),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_158),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_146),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_142),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_50),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_7),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_46),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_168),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_93),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_108),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_24),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_17),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_13),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_29),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_4),
.Y(n_224)
);

INVxp67_ASAP7_75t_SL g225 ( 
.A(n_24),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_52),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_131),
.Y(n_227)
);

BUFx5_ASAP7_75t_L g228 ( 
.A(n_25),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_0),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_69),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_54),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_117),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_163),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_143),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_68),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_72),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_126),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_116),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_54),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_102),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_78),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_71),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_99),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_41),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_40),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_160),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_59),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_82),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_100),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_148),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_4),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_39),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_34),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_49),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_70),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_122),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_112),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_14),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_134),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_118),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_7),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_36),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_140),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_51),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_38),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_0),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_21),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_12),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_149),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_121),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_161),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_18),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_34),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_38),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_94),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_166),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_119),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_40),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_50),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_167),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_12),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_153),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_76),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_81),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_36),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_60),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_67),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_150),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_29),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_132),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_57),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_125),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_28),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_74),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_3),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_79),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_58),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_32),
.Y(n_298)
);

BUFx5_ASAP7_75t_L g299 ( 
.A(n_104),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_44),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_86),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_98),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_6),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_123),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_8),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_53),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_159),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_136),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_52),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_156),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_51),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_129),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_45),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_133),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_87),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_57),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_128),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_45),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_111),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_47),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_11),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_113),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_13),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_19),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_138),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_145),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_3),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_6),
.Y(n_328)
);

BUFx2_ASAP7_75t_SL g329 ( 
.A(n_95),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_157),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_58),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_83),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_65),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_1),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_141),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_96),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_228),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_228),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_228),
.B(n_1),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_293),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_176),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_180),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_208),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_245),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_241),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_335),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_234),
.Y(n_347)
);

BUFx6f_ASAP7_75t_SL g348 ( 
.A(n_280),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_228),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_210),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_189),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_214),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_242),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_196),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_215),
.Y(n_355)
);

INVxp33_ASAP7_75t_L g356 ( 
.A(n_169),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_212),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_228),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_228),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_228),
.Y(n_360)
);

INVxp33_ASAP7_75t_L g361 ( 
.A(n_188),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_288),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_263),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_228),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_209),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_216),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_211),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_194),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_194),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_286),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_277),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_222),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_219),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_187),
.Y(n_374)
);

BUFx2_ASAP7_75t_L g375 ( 
.A(n_286),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_227),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_231),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_283),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_187),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_L g380 ( 
.A(n_226),
.B(n_2),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_189),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_230),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_266),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_252),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_309),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_254),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_189),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_299),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_266),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_258),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_261),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_309),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_232),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_262),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_280),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_198),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_201),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_299),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_264),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_267),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_268),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g402 ( 
.A(n_170),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_202),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g404 ( 
.A(n_171),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_205),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_280),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_308),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_221),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_213),
.B(n_2),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_224),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_184),
.B(n_8),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_229),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_233),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_239),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_247),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_213),
.B(n_9),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_251),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_319),
.B(n_9),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_358),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_358),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_359),
.Y(n_421)
);

AND2x6_ASAP7_75t_L g422 ( 
.A(n_337),
.B(n_246),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_359),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_402),
.B(n_319),
.Y(n_424)
);

AND2x6_ASAP7_75t_L g425 ( 
.A(n_337),
.B(n_246),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_344),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_349),
.Y(n_427)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_407),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_364),
.B(n_304),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_350),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_338),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_404),
.B(n_304),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_338),
.B(n_308),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_360),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_360),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_407),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_365),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_407),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_407),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_407),
.Y(n_440)
);

NAND2xp33_ASAP7_75t_L g441 ( 
.A(n_409),
.B(n_226),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_339),
.B(n_308),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g443 ( 
.A(n_350),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_388),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_388),
.B(n_308),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_398),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_398),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_374),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_374),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_379),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_379),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_383),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_416),
.B(n_308),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g454 ( 
.A(n_375),
.B(n_392),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_383),
.Y(n_455)
);

BUFx12f_ASAP7_75t_L g456 ( 
.A(n_352),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_389),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_389),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_396),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_418),
.B(n_172),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_396),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_405),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_380),
.B(n_307),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_405),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_368),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_397),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_412),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_415),
.B(n_175),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_375),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_417),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_392),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_369),
.Y(n_472)
);

AND2x2_ASAP7_75t_SL g473 ( 
.A(n_395),
.B(n_185),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_370),
.B(n_186),
.Y(n_474)
);

AND2x4_ASAP7_75t_SL g475 ( 
.A(n_367),
.B(n_307),
.Y(n_475)
);

BUFx12f_ASAP7_75t_L g476 ( 
.A(n_352),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_385),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_356),
.B(n_200),
.Y(n_478)
);

OA21x2_ASAP7_75t_L g479 ( 
.A1(n_403),
.A2(n_265),
.B(n_253),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_408),
.B(n_217),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_410),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_414),
.B(n_243),
.Y(n_482)
);

BUFx8_ASAP7_75t_L g483 ( 
.A(n_348),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_345),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_355),
.Y(n_485)
);

INVx6_ASAP7_75t_L g486 ( 
.A(n_406),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_346),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_363),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_371),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_378),
.B(n_248),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_361),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_351),
.B(n_255),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_419),
.Y(n_493)
);

INVx8_ASAP7_75t_L g494 ( 
.A(n_485),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_435),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_419),
.Y(n_496)
);

BUFx10_ASAP7_75t_L g497 ( 
.A(n_486),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_435),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_473),
.A2(n_362),
.B1(n_373),
.B2(n_413),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_487),
.B(n_355),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_445),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_440),
.Y(n_502)
);

INVx8_ASAP7_75t_L g503 ( 
.A(n_485),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_487),
.B(n_366),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_435),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_488),
.B(n_376),
.Y(n_506)
);

INVx5_ASAP7_75t_L g507 ( 
.A(n_422),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_465),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_419),
.Y(n_509)
);

NOR2x1p5_ASAP7_75t_L g510 ( 
.A(n_491),
.B(n_366),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_419),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_L g512 ( 
.A1(n_460),
.A2(n_334),
.B1(n_306),
.B2(n_300),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_465),
.Y(n_513)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_426),
.B(n_340),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_465),
.Y(n_515)
);

INVxp67_ASAP7_75t_SL g516 ( 
.A(n_439),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_487),
.B(n_372),
.Y(n_517)
);

AND3x2_ASAP7_75t_L g518 ( 
.A(n_426),
.B(n_443),
.C(n_430),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_488),
.B(n_489),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_420),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_491),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_440),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_487),
.B(n_453),
.Y(n_523)
);

NOR2x1p5_ASAP7_75t_L g524 ( 
.A(n_491),
.B(n_372),
.Y(n_524)
);

AND2x6_ASAP7_75t_L g525 ( 
.A(n_442),
.B(n_284),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_420),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_453),
.B(n_377),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_440),
.Y(n_528)
);

INVx4_ASAP7_75t_L g529 ( 
.A(n_445),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_453),
.B(n_377),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_453),
.B(n_384),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_465),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_460),
.A2(n_432),
.B1(n_424),
.B2(n_442),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_466),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_420),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_473),
.A2(n_382),
.B1(n_393),
.B2(n_357),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_488),
.B(n_384),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_489),
.B(n_460),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_466),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_440),
.Y(n_540)
);

NAND2xp33_ASAP7_75t_L g541 ( 
.A(n_422),
.B(n_299),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_424),
.B(n_386),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_440),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_469),
.Y(n_544)
);

AND2x6_ASAP7_75t_L g545 ( 
.A(n_442),
.B(n_294),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_453),
.B(n_386),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_420),
.Y(n_547)
);

AND3x2_ASAP7_75t_L g548 ( 
.A(n_430),
.B(n_225),
.C(n_381),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_430),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g550 ( 
.A(n_443),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_440),
.Y(n_551)
);

BUFx2_ASAP7_75t_L g552 ( 
.A(n_443),
.Y(n_552)
);

AOI21x1_ASAP7_75t_L g553 ( 
.A1(n_429),
.A2(n_314),
.B(n_296),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_424),
.B(n_390),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_466),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_421),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_467),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_440),
.Y(n_558)
);

AND2x6_ASAP7_75t_L g559 ( 
.A(n_442),
.B(n_315),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_453),
.B(n_390),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_467),
.Y(n_561)
);

AND3x2_ASAP7_75t_L g562 ( 
.A(n_469),
.B(n_326),
.C(n_325),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_473),
.B(n_391),
.Y(n_563)
);

CKINVDCx14_ASAP7_75t_R g564 ( 
.A(n_486),
.Y(n_564)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_445),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_454),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_440),
.Y(n_567)
);

AO21x1_ASAP7_75t_L g568 ( 
.A1(n_490),
.A2(n_295),
.B(n_279),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_489),
.B(n_391),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_473),
.B(n_411),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_440),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_467),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_472),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_437),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_421),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_424),
.B(n_394),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_432),
.B(n_394),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_473),
.A2(n_354),
.B1(n_401),
.B2(n_400),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_432),
.B(n_399),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_454),
.B(n_387),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_421),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_427),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_428),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_421),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_427),
.Y(n_585)
);

BUFx10_ASAP7_75t_L g586 ( 
.A(n_486),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_454),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_444),
.Y(n_588)
);

AO22x2_ASAP7_75t_L g589 ( 
.A1(n_442),
.A2(n_334),
.B1(n_303),
.B2(n_206),
.Y(n_589)
);

AOI21x1_ASAP7_75t_L g590 ( 
.A1(n_429),
.A2(n_332),
.B(n_330),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_444),
.Y(n_591)
);

AND2x6_ASAP7_75t_L g592 ( 
.A(n_442),
.B(n_333),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_444),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_432),
.B(n_399),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_433),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_484),
.B(n_400),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_474),
.B(n_218),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_472),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_444),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_474),
.B(n_235),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_484),
.B(n_401),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_474),
.B(n_307),
.Y(n_602)
);

AND2x2_ASAP7_75t_SL g603 ( 
.A(n_475),
.B(n_329),
.Y(n_603)
);

BUFx10_ASAP7_75t_L g604 ( 
.A(n_486),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_446),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_427),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_446),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_446),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_454),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_446),
.Y(n_610)
);

OAI21xp33_ASAP7_75t_SL g611 ( 
.A1(n_463),
.A2(n_193),
.B(n_299),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_484),
.B(n_236),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_447),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_474),
.B(n_480),
.Y(n_614)
);

NAND2xp33_ASAP7_75t_L g615 ( 
.A(n_422),
.B(n_299),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_427),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_447),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_474),
.B(n_237),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_SL g619 ( 
.A(n_456),
.B(n_341),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_L g620 ( 
.A1(n_485),
.A2(n_278),
.B1(n_272),
.B2(n_273),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_428),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_485),
.B(n_348),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_433),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_433),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_479),
.A2(n_348),
.B1(n_299),
.B2(n_191),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_472),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_433),
.Y(n_627)
);

AND2x6_ASAP7_75t_L g628 ( 
.A(n_485),
.B(n_299),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_479),
.B(n_238),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_447),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_433),
.Y(n_631)
);

INVxp33_ASAP7_75t_L g632 ( 
.A(n_478),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_479),
.B(n_240),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_433),
.Y(n_634)
);

AND2x6_ASAP7_75t_L g635 ( 
.A(n_485),
.B(n_474),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_479),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_431),
.Y(n_637)
);

NAND2xp33_ASAP7_75t_L g638 ( 
.A(n_422),
.B(n_299),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_431),
.Y(n_639)
);

NOR2x1p5_ASAP7_75t_L g640 ( 
.A(n_456),
.B(n_173),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_428),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_431),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_431),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_533),
.B(n_479),
.Y(n_644)
);

NOR3xp33_ASAP7_75t_L g645 ( 
.A(n_499),
.B(n_463),
.C(n_437),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_595),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_538),
.B(n_479),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_632),
.B(n_475),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_632),
.B(n_475),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_517),
.B(n_479),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_SL g651 ( 
.A(n_603),
.B(n_456),
.Y(n_651)
);

AND2x2_ASAP7_75t_SL g652 ( 
.A(n_625),
.B(n_475),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_510),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_595),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_623),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_566),
.B(n_490),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_501),
.B(n_445),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_517),
.B(n_481),
.Y(n_658)
);

INVxp33_ASAP7_75t_L g659 ( 
.A(n_514),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_501),
.B(n_445),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_501),
.B(n_445),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_544),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_493),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_493),
.Y(n_664)
);

BUFx4f_ASAP7_75t_L g665 ( 
.A(n_603),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_523),
.B(n_478),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_624),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_523),
.B(n_478),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_627),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_519),
.B(n_478),
.Y(n_670)
);

OAI22xp33_ASAP7_75t_L g671 ( 
.A1(n_542),
.A2(n_490),
.B1(n_486),
.B2(n_482),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_631),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_504),
.B(n_486),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_514),
.Y(n_674)
);

NAND2xp33_ASAP7_75t_L g675 ( 
.A(n_635),
.B(n_422),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_508),
.B(n_513),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_515),
.B(n_472),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_529),
.B(n_472),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_634),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_534),
.Y(n_680)
);

INVxp67_ASAP7_75t_SL g681 ( 
.A(n_583),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_495),
.B(n_498),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_505),
.B(n_472),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_524),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_529),
.B(n_565),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_568),
.A2(n_480),
.B1(n_441),
.B2(n_492),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_496),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_532),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_563),
.A2(n_486),
.B1(n_456),
.B2(n_476),
.Y(n_689)
);

INVxp67_ASAP7_75t_SL g690 ( 
.A(n_583),
.Y(n_690)
);

INVxp33_ASAP7_75t_L g691 ( 
.A(n_537),
.Y(n_691)
);

NOR3xp33_ASAP7_75t_L g692 ( 
.A(n_536),
.B(n_563),
.C(n_506),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_579),
.B(n_481),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_496),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_529),
.B(n_472),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_597),
.B(n_472),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_597),
.B(n_472),
.Y(n_697)
);

NOR2xp67_ASAP7_75t_L g698 ( 
.A(n_622),
.B(n_476),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_565),
.B(n_471),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_527),
.A2(n_476),
.B1(n_492),
.B2(n_353),
.Y(n_700)
);

AND2x6_ASAP7_75t_L g701 ( 
.A(n_602),
.B(n_492),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_597),
.B(n_434),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_509),
.Y(n_703)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_549),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_539),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_555),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_574),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_569),
.B(n_342),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_557),
.B(n_434),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_596),
.B(n_343),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_527),
.A2(n_476),
.B1(n_492),
.B2(n_347),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_561),
.Y(n_712)
);

INVx8_ASAP7_75t_L g713 ( 
.A(n_635),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_565),
.B(n_471),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_614),
.B(n_471),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_614),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_614),
.B(n_471),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_572),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_509),
.Y(n_719)
);

NOR3xp33_ASAP7_75t_L g720 ( 
.A(n_580),
.B(n_482),
.C(n_441),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_601),
.B(n_492),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_554),
.B(n_434),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_568),
.A2(n_480),
.B1(n_492),
.B2(n_425),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_636),
.B(n_471),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_500),
.B(n_481),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_636),
.B(n_471),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_566),
.B(n_482),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_521),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_500),
.B(n_480),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_576),
.B(n_434),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_577),
.B(n_471),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_594),
.B(n_471),
.Y(n_732)
);

INVxp67_ASAP7_75t_L g733 ( 
.A(n_550),
.Y(n_733)
);

INVxp67_ASAP7_75t_L g734 ( 
.A(n_552),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_579),
.B(n_480),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_629),
.B(n_471),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_587),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_532),
.B(n_480),
.Y(n_738)
);

INVx8_ASAP7_75t_L g739 ( 
.A(n_635),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_580),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_587),
.B(n_477),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_633),
.B(n_429),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_602),
.B(n_464),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_611),
.B(n_497),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_522),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_516),
.B(n_464),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_497),
.B(n_483),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_609),
.Y(n_748)
);

INVxp67_ASAP7_75t_L g749 ( 
.A(n_620),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_612),
.B(n_464),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_609),
.B(n_477),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_628),
.B(n_464),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_511),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_497),
.B(n_483),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_511),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_628),
.B(n_464),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_520),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_586),
.B(n_483),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_562),
.Y(n_759)
);

AO22x2_ASAP7_75t_L g760 ( 
.A1(n_530),
.A2(n_411),
.B1(n_468),
.B2(n_477),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_578),
.B(n_477),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_586),
.B(n_604),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_628),
.B(n_464),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_530),
.B(n_468),
.Y(n_764)
);

OAI22xp33_ASAP7_75t_L g765 ( 
.A1(n_531),
.A2(n_468),
.B1(n_320),
.B2(n_199),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_520),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_628),
.B(n_464),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_583),
.A2(n_428),
.B(n_447),
.Y(n_768)
);

NOR3xp33_ASAP7_75t_L g769 ( 
.A(n_531),
.B(n_285),
.C(n_274),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_526),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_586),
.B(n_604),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_628),
.B(n_464),
.Y(n_772)
);

INVx1_ASAP7_75t_SL g773 ( 
.A(n_574),
.Y(n_773)
);

NOR3xp33_ASAP7_75t_L g774 ( 
.A(n_546),
.B(n_281),
.C(n_297),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_526),
.Y(n_775)
);

AND2x6_ASAP7_75t_SL g776 ( 
.A(n_570),
.B(n_197),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_546),
.B(n_560),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_604),
.B(n_483),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_512),
.B(n_470),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_535),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_525),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_535),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_628),
.B(n_494),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_494),
.B(n_464),
.Y(n_784)
);

NAND2xp33_ASAP7_75t_L g785 ( 
.A(n_635),
.B(n_422),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_494),
.B(n_423),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_494),
.B(n_503),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_503),
.B(n_423),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_547),
.Y(n_789)
);

INVxp67_ASAP7_75t_SL g790 ( 
.A(n_621),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_503),
.B(n_423),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_560),
.B(n_470),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_547),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_503),
.B(n_458),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_518),
.B(n_640),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_548),
.B(n_174),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_621),
.B(n_458),
.Y(n_797)
);

A2O1A1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_541),
.A2(n_449),
.B(n_450),
.C(n_455),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_556),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_600),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_621),
.B(n_483),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_556),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_600),
.A2(n_276),
.B1(n_249),
.B2(n_250),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_522),
.Y(n_804)
);

BUFx6f_ASAP7_75t_SL g805 ( 
.A(n_600),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_641),
.B(n_458),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_575),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_575),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_581),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_570),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_525),
.A2(n_422),
.B1(n_425),
.B2(n_470),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_641),
.B(n_458),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_641),
.B(n_458),
.Y(n_813)
);

NAND2x1_ASAP7_75t_L g814 ( 
.A(n_635),
.B(n_428),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_618),
.B(n_483),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_670),
.B(n_635),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_721),
.B(n_618),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_L g818 ( 
.A1(n_647),
.A2(n_639),
.B(n_637),
.Y(n_818)
);

O2A1O1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_650),
.A2(n_638),
.B(n_541),
.C(n_615),
.Y(n_819)
);

NAND3xp33_ASAP7_75t_L g820 ( 
.A(n_692),
.B(n_619),
.C(n_618),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_777),
.B(n_589),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_729),
.A2(n_764),
.B1(n_691),
.B2(n_644),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_663),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_693),
.B(n_589),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_783),
.A2(n_787),
.B(n_771),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_725),
.B(n_589),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_681),
.B(n_589),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_707),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_690),
.B(n_790),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_762),
.A2(n_502),
.B(n_522),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_741),
.B(n_525),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_742),
.A2(n_643),
.B(n_642),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_655),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_663),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_L g835 ( 
.A1(n_691),
.A2(n_564),
.B1(n_207),
.B2(n_244),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_664),
.Y(n_836)
);

OAI22xp5_ASAP7_75t_L g837 ( 
.A1(n_749),
.A2(n_666),
.B1(n_668),
.B2(n_652),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_662),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_751),
.B(n_658),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_652),
.A2(n_564),
.B1(n_220),
.B2(n_223),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_667),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_762),
.A2(n_502),
.B(n_522),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_735),
.B(n_525),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_722),
.B(n_525),
.Y(n_844)
);

A2O1A1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_673),
.A2(n_638),
.B(n_615),
.C(n_606),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_730),
.B(n_525),
.Y(n_846)
);

O2A1O1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_727),
.A2(n_582),
.B(n_616),
.C(n_585),
.Y(n_847)
);

NOR3xp33_ASAP7_75t_L g848 ( 
.A(n_708),
.B(n_765),
.C(n_710),
.Y(n_848)
);

O2A1O1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_671),
.A2(n_470),
.B(n_617),
.C(n_613),
.Y(n_849)
);

A2O1A1Ixp33_ASAP7_75t_L g850 ( 
.A1(n_792),
.A2(n_543),
.B(n_551),
.C(n_567),
.Y(n_850)
);

INVx6_ASAP7_75t_L g851 ( 
.A(n_688),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_664),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_771),
.A2(n_788),
.B(n_786),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_669),
.Y(n_854)
);

AOI21xp33_ASAP7_75t_L g855 ( 
.A1(n_659),
.A2(n_178),
.B(n_173),
.Y(n_855)
);

AOI21xp33_ASAP7_75t_L g856 ( 
.A1(n_659),
.A2(n_649),
.B(n_648),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_791),
.A2(n_502),
.B(n_522),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_687),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_656),
.B(n_680),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_687),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_694),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_800),
.B(n_449),
.Y(n_862)
);

OAI21xp33_ASAP7_75t_L g863 ( 
.A1(n_728),
.A2(n_179),
.B(n_178),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_716),
.A2(n_292),
.B1(n_177),
.B2(n_181),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_705),
.B(n_545),
.Y(n_865)
);

OAI21xp33_ASAP7_75t_L g866 ( 
.A1(n_748),
.A2(n_190),
.B(n_179),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_706),
.B(n_545),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_712),
.B(n_545),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_672),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_718),
.B(n_702),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_685),
.A2(n_502),
.B(n_528),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_779),
.B(n_545),
.Y(n_872)
);

AOI21x1_ASAP7_75t_L g873 ( 
.A1(n_724),
.A2(n_590),
.B(n_553),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_740),
.B(n_543),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_731),
.B(n_545),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_685),
.A2(n_697),
.B(n_696),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_679),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_657),
.A2(n_540),
.B(n_528),
.Y(n_878)
);

A2O1A1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_720),
.A2(n_543),
.B(n_551),
.C(n_567),
.Y(n_879)
);

O2A1O1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_798),
.A2(n_630),
.B(n_617),
.C(n_613),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_732),
.B(n_545),
.Y(n_881)
);

INVx3_ASAP7_75t_SL g882 ( 
.A(n_707),
.Y(n_882)
);

BUFx2_ASAP7_75t_L g883 ( 
.A(n_704),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_737),
.B(n_559),
.Y(n_884)
);

BUFx12f_ASAP7_75t_L g885 ( 
.A(n_776),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_694),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_716),
.B(n_528),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_759),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_703),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_703),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_682),
.B(n_559),
.Y(n_891)
);

INVx1_ASAP7_75t_SL g892 ( 
.A(n_773),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_657),
.A2(n_540),
.B(n_528),
.Y(n_893)
);

CKINVDCx20_ASAP7_75t_R g894 ( 
.A(n_810),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_716),
.B(n_528),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_719),
.Y(n_896)
);

NOR2x2_ASAP7_75t_L g897 ( 
.A(n_760),
.B(n_190),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_660),
.A2(n_540),
.B(n_558),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_761),
.B(n_559),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_745),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_686),
.B(n_738),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_646),
.B(n_559),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_674),
.B(n_551),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_733),
.B(n_567),
.Y(n_904)
);

O2A1O1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_798),
.A2(n_630),
.B(n_610),
.C(n_608),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_654),
.B(n_559),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_676),
.Y(n_907)
);

NOR2xp67_ASAP7_75t_R g908 ( 
.A(n_781),
.B(n_507),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_660),
.A2(n_540),
.B(n_558),
.Y(n_909)
);

AOI33xp33_ASAP7_75t_L g910 ( 
.A1(n_653),
.A2(n_449),
.A3(n_450),
.B1(n_452),
.B2(n_455),
.B3(n_457),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_701),
.B(n_559),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_661),
.A2(n_742),
.B(n_752),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_734),
.B(n_571),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_701),
.B(n_592),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_661),
.A2(n_540),
.B(n_558),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_701),
.B(n_592),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_651),
.B(n_700),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_745),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_701),
.B(n_592),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_701),
.B(n_592),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_711),
.B(n_571),
.Y(n_921)
);

A2O1A1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_665),
.A2(n_571),
.B(n_610),
.C(n_608),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_688),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_756),
.A2(n_558),
.B(n_428),
.Y(n_924)
);

O2A1O1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_815),
.A2(n_581),
.B(n_607),
.C(n_605),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_665),
.B(n_558),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_684),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_688),
.B(n_592),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_689),
.A2(n_290),
.B1(n_177),
.B2(n_181),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_688),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_763),
.A2(n_626),
.B(n_573),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_723),
.B(n_592),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_743),
.B(n_584),
.Y(n_933)
);

OAI21xp33_ASAP7_75t_L g934 ( 
.A1(n_760),
.A2(n_316),
.B(n_289),
.Y(n_934)
);

A2O1A1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_774),
.A2(n_458),
.B(n_313),
.C(n_328),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_767),
.A2(n_626),
.B(n_573),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_719),
.B(n_584),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_724),
.A2(n_588),
.B(n_607),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_713),
.B(n_573),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_713),
.A2(n_287),
.B1(n_182),
.B2(n_183),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_755),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_796),
.B(n_191),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_755),
.B(n_588),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_770),
.B(n_591),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_770),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_805),
.B(n_204),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_713),
.B(n_573),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_775),
.B(n_591),
.Y(n_948)
);

BUFx8_ASAP7_75t_L g949 ( 
.A(n_795),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_769),
.A2(n_259),
.B1(n_256),
.B2(n_260),
.Y(n_950)
);

O2A1O1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_815),
.A2(n_605),
.B(n_599),
.C(n_593),
.Y(n_951)
);

NAND3xp33_ASAP7_75t_SL g952 ( 
.A(n_645),
.B(n_313),
.C(n_204),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_745),
.Y(n_953)
);

OAI321xp33_ASAP7_75t_L g954 ( 
.A1(n_803),
.A2(n_801),
.A3(n_746),
.B1(n_760),
.B2(n_744),
.C(n_709),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_750),
.A2(n_593),
.B(n_599),
.C(n_257),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_805),
.B(n_289),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_775),
.B(n_459),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_804),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_772),
.A2(n_626),
.B(n_598),
.Y(n_959)
);

OR2x2_ASAP7_75t_L g960 ( 
.A(n_810),
.B(n_291),
.Y(n_960)
);

BUFx4f_ASAP7_75t_L g961 ( 
.A(n_745),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_789),
.B(n_459),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_726),
.A2(n_626),
.B(n_598),
.Y(n_963)
);

OAI21xp5_ASAP7_75t_L g964 ( 
.A1(n_726),
.A2(n_425),
.B(n_422),
.Y(n_964)
);

NAND3xp33_ASAP7_75t_L g965 ( 
.A(n_715),
.B(n_203),
.C(n_182),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_784),
.A2(n_794),
.B(n_736),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_698),
.A2(n_203),
.B(n_174),
.C(n_183),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_713),
.A2(n_290),
.B1(n_336),
.B2(n_322),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_736),
.A2(n_806),
.B(n_797),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_812),
.A2(n_626),
.B(n_598),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_805),
.B(n_291),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_813),
.A2(n_598),
.B(n_573),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_715),
.B(n_459),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_717),
.A2(n_598),
.B(n_507),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_717),
.A2(n_507),
.B(n_439),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_781),
.B(n_459),
.Y(n_976)
);

OAI321xp33_ASAP7_75t_L g977 ( 
.A1(n_801),
.A2(n_450),
.A3(n_452),
.B1(n_455),
.B2(n_457),
.C(n_462),
.Y(n_977)
);

AOI22xp33_ASAP7_75t_L g978 ( 
.A1(n_675),
.A2(n_425),
.B1(n_422),
.B2(n_318),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_804),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_789),
.B(n_461),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_768),
.A2(n_422),
.B(n_425),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_753),
.B(n_297),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_744),
.A2(n_675),
.B(n_785),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_785),
.A2(n_678),
.B(n_695),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_809),
.Y(n_985)
);

CKINVDCx10_ASAP7_75t_R g986 ( 
.A(n_747),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_809),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_804),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_757),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_739),
.A2(n_192),
.B1(n_195),
.B2(n_257),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_766),
.B(n_780),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_695),
.A2(n_507),
.B(n_439),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_782),
.B(n_461),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_699),
.A2(n_439),
.B(n_438),
.Y(n_994)
);

OAI21xp33_ASAP7_75t_L g995 ( 
.A1(n_811),
.A2(n_298),
.B(n_305),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_793),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_799),
.B(n_298),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_802),
.B(n_807),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_808),
.B(n_461),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_739),
.B(n_461),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_739),
.B(n_683),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_677),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_739),
.A2(n_814),
.B(n_714),
.C(n_699),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_714),
.A2(n_439),
.B(n_438),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_747),
.B(n_192),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_754),
.B(n_462),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_778),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_900),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_883),
.Y(n_1009)
);

BUFx2_ASAP7_75t_L g1010 ( 
.A(n_838),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_900),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_823),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_848),
.B(n_754),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_848),
.B(n_778),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_838),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_817),
.A2(n_758),
.B(n_438),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_901),
.A2(n_758),
.B(n_438),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_834),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_900),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_839),
.B(n_462),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_836),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_917),
.A2(n_282),
.B1(n_269),
.B2(n_270),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_942),
.B(n_824),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_942),
.B(n_452),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_816),
.A2(n_881),
.B(n_875),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_876),
.A2(n_436),
.B(n_462),
.Y(n_1026)
);

INVxp67_ASAP7_75t_L g1027 ( 
.A(n_859),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_907),
.B(n_457),
.Y(n_1028)
);

AOI221xp5_ASAP7_75t_L g1029 ( 
.A1(n_917),
.A2(n_305),
.B1(n_311),
.B2(n_316),
.C(n_318),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_844),
.A2(n_436),
.B(n_451),
.Y(n_1030)
);

OAI22x1_ASAP7_75t_L g1031 ( 
.A1(n_882),
.A2(n_331),
.B1(n_328),
.B2(n_327),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_856),
.B(n_195),
.Y(n_1032)
);

CKINVDCx8_ASAP7_75t_R g1033 ( 
.A(n_986),
.Y(n_1033)
);

INVx6_ASAP7_75t_L g1034 ( 
.A(n_949),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_833),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_841),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_821),
.A2(n_451),
.B(n_448),
.C(n_436),
.Y(n_1037)
);

OAI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_837),
.A2(n_425),
.B(n_422),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_870),
.B(n_287),
.Y(n_1039)
);

OAI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_912),
.A2(n_425),
.B(n_422),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_846),
.A2(n_436),
.B(n_451),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_932),
.A2(n_317),
.B1(n_292),
.B2(n_336),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_852),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_835),
.B(n_311),
.Y(n_1044)
);

INVx2_ASAP7_75t_SL g1045 ( 
.A(n_888),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_855),
.B(n_321),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_SL g1047 ( 
.A(n_894),
.B(n_312),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_820),
.A2(n_271),
.B1(n_275),
.B2(n_302),
.Y(n_1048)
);

CKINVDCx14_ASAP7_75t_R g1049 ( 
.A(n_828),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_960),
.B(n_321),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_900),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_892),
.B(n_331),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_858),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_918),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_854),
.B(n_322),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_966),
.A2(n_451),
.B(n_448),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_983),
.A2(n_448),
.B(n_317),
.Y(n_1057)
);

OAI221xp5_ASAP7_75t_L g1058 ( 
.A1(n_934),
.A2(n_323),
.B1(n_327),
.B2(n_324),
.C(n_312),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_869),
.B(n_310),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_819),
.A2(n_448),
.B(n_310),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_877),
.B(n_302),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_853),
.A2(n_301),
.B(n_425),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_840),
.B(n_301),
.Y(n_1063)
);

INVx3_ASAP7_75t_L g1064 ( 
.A(n_918),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_982),
.B(n_323),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_918),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_952),
.B(n_324),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_941),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_945),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_985),
.Y(n_1070)
);

NAND2x1_ASAP7_75t_SL g1071 ( 
.A(n_882),
.B(n_10),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_982),
.B(n_10),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_822),
.B(n_15),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_997),
.B(n_946),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_997),
.B(n_15),
.Y(n_1075)
);

BUFx3_ASAP7_75t_L g1076 ( 
.A(n_927),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_904),
.B(n_425),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_923),
.Y(n_1078)
);

CKINVDCx14_ASAP7_75t_R g1079 ( 
.A(n_885),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_984),
.A2(n_425),
.B(n_73),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_904),
.B(n_16),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_913),
.B(n_425),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_913),
.B(n_425),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_860),
.Y(n_1084)
);

BUFx4f_ASAP7_75t_L g1085 ( 
.A(n_851),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_845),
.A2(n_63),
.B(n_164),
.Y(n_1086)
);

CKINVDCx11_ASAP7_75t_R g1087 ( 
.A(n_949),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_891),
.A2(n_62),
.B(n_162),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_946),
.B(n_18),
.Y(n_1089)
);

BUFx4f_ASAP7_75t_L g1090 ( 
.A(n_851),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_961),
.B(n_75),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_899),
.A2(n_165),
.B1(n_147),
.B2(n_137),
.Y(n_1092)
);

AOI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_921),
.A2(n_127),
.B1(n_124),
.B2(n_115),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_861),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_921),
.A2(n_110),
.B1(n_109),
.B2(n_107),
.Y(n_1095)
);

NOR2xp67_ASAP7_75t_L g1096 ( 
.A(n_965),
.B(n_106),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_956),
.B(n_19),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_956),
.B(n_20),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_874),
.B(n_20),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_825),
.A2(n_101),
.B(n_92),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_874),
.B(n_23),
.Y(n_1101)
);

AO32x1_ASAP7_75t_L g1102 ( 
.A1(n_929),
.A2(n_23),
.A3(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_886),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_903),
.B(n_26),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_889),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_918),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_971),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_818),
.A2(n_103),
.B(n_90),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_890),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_SL g1110 ( 
.A1(n_826),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_896),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_987),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_953),
.Y(n_1113)
);

BUFx3_ASAP7_75t_L g1114 ( 
.A(n_851),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_923),
.Y(n_1115)
);

HB1xp67_ASAP7_75t_L g1116 ( 
.A(n_930),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_953),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_996),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_903),
.B(n_31),
.Y(n_1119)
);

AOI222xp33_ASAP7_75t_L g1120 ( 
.A1(n_863),
.A2(n_33),
.B1(n_35),
.B2(n_37),
.C1(n_42),
.C2(n_43),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_961),
.B(n_85),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_SL g1122 ( 
.A1(n_971),
.A2(n_35),
.B1(n_42),
.B2(n_43),
.Y(n_1122)
);

CKINVDCx8_ASAP7_75t_R g1123 ( 
.A(n_953),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_989),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_969),
.A2(n_84),
.B(n_49),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_862),
.B(n_48),
.Y(n_1126)
);

O2A1O1Ixp5_ASAP7_75t_L g1127 ( 
.A1(n_955),
.A2(n_48),
.B(n_55),
.C(n_56),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_998),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_977),
.A2(n_55),
.B(n_59),
.Y(n_1129)
);

NOR2xp67_ASAP7_75t_SL g1130 ( 
.A(n_953),
.B(n_954),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_935),
.A2(n_827),
.B(n_1005),
.C(n_847),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1000),
.A2(n_933),
.B(n_831),
.Y(n_1132)
);

NOR2xp67_ASAP7_75t_SL g1133 ( 
.A(n_1007),
.B(n_930),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_862),
.B(n_950),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_843),
.A2(n_872),
.B(n_1003),
.Y(n_1135)
);

AO32x1_ASAP7_75t_L g1136 ( 
.A1(n_1002),
.A2(n_864),
.A3(n_990),
.B1(n_968),
.B2(n_940),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_958),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_989),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_973),
.A2(n_995),
.B1(n_1005),
.B2(n_976),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_958),
.B(n_979),
.Y(n_1140)
);

NOR2xp67_ASAP7_75t_L g1141 ( 
.A(n_866),
.B(n_884),
.Y(n_1141)
);

AND2x4_ASAP7_75t_L g1142 ( 
.A(n_979),
.B(n_988),
.Y(n_1142)
);

BUFx3_ASAP7_75t_L g1143 ( 
.A(n_988),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_829),
.A2(n_1006),
.B(n_931),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_910),
.B(n_991),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_926),
.A2(n_867),
.B1(n_868),
.B2(n_865),
.Y(n_1146)
);

OR2x2_ASAP7_75t_L g1147 ( 
.A(n_935),
.B(n_926),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_887),
.B(n_895),
.Y(n_1148)
);

AND3x1_ASAP7_75t_SL g1149 ( 
.A(n_897),
.B(n_978),
.C(n_967),
.Y(n_1149)
);

AO32x1_ASAP7_75t_L g1150 ( 
.A1(n_873),
.A2(n_849),
.A3(n_879),
.B1(n_832),
.B2(n_922),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_936),
.A2(n_959),
.B(n_1001),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_928),
.B(n_902),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_R g1153 ( 
.A(n_991),
.B(n_906),
.Y(n_1153)
);

NOR2x1_ASAP7_75t_R g1154 ( 
.A(n_887),
.B(n_895),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_964),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_850),
.A2(n_916),
.B1(n_911),
.B2(n_920),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_993),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_937),
.B(n_944),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_1001),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_857),
.A2(n_970),
.B(n_972),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_914),
.B(n_919),
.Y(n_1161)
);

INVx4_ASAP7_75t_L g1162 ( 
.A(n_908),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_978),
.B(n_909),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_938),
.B(n_999),
.Y(n_1164)
);

OAI22x1_ASAP7_75t_L g1165 ( 
.A1(n_939),
.A2(n_947),
.B1(n_948),
.B2(n_943),
.Y(n_1165)
);

OAI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_939),
.A2(n_947),
.B1(n_915),
.B2(n_878),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_957),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_1074),
.B(n_898),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_1076),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1128),
.B(n_962),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1073),
.A2(n_1098),
.B(n_1089),
.C(n_1081),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1035),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1135),
.A2(n_905),
.B(n_880),
.Y(n_1173)
);

BUFx10_ASAP7_75t_L g1174 ( 
.A(n_1052),
.Y(n_1174)
);

AO31x2_ASAP7_75t_L g1175 ( 
.A1(n_1165),
.A2(n_830),
.A3(n_842),
.B(n_893),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1036),
.Y(n_1176)
);

OA21x2_ASAP7_75t_L g1177 ( 
.A1(n_1135),
.A2(n_980),
.B(n_1004),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1073),
.A2(n_951),
.B(n_925),
.C(n_994),
.Y(n_1178)
);

NAND3xp33_ASAP7_75t_SL g1179 ( 
.A(n_1107),
.B(n_981),
.C(n_975),
.Y(n_1179)
);

INVx1_ASAP7_75t_SL g1180 ( 
.A(n_1009),
.Y(n_1180)
);

AO31x2_ASAP7_75t_L g1181 ( 
.A1(n_1017),
.A2(n_963),
.A3(n_871),
.B(n_924),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1144),
.A2(n_974),
.B(n_992),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1118),
.Y(n_1183)
);

A2O1A1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1080),
.A2(n_1131),
.B(n_1072),
.C(n_1075),
.Y(n_1184)
);

BUFx10_ASAP7_75t_L g1185 ( 
.A(n_1034),
.Y(n_1185)
);

INVx4_ASAP7_75t_L g1186 ( 
.A(n_1085),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1068),
.Y(n_1187)
);

OAI22x1_ASAP7_75t_L g1188 ( 
.A1(n_1159),
.A2(n_1097),
.B1(n_1067),
.B2(n_1023),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1024),
.B(n_1027),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1069),
.Y(n_1190)
);

CKINVDCx11_ASAP7_75t_R g1191 ( 
.A(n_1087),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_1123),
.Y(n_1192)
);

INVx5_ASAP7_75t_L g1193 ( 
.A(n_1011),
.Y(n_1193)
);

O2A1O1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1013),
.A2(n_1014),
.B(n_1032),
.C(n_1120),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_1010),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_1015),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1030),
.A2(n_1041),
.B(n_1160),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1027),
.B(n_1028),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1041),
.A2(n_1056),
.B(n_1144),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1050),
.B(n_1015),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1132),
.A2(n_1025),
.B(n_1156),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1070),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1131),
.A2(n_1108),
.B(n_1141),
.C(n_1065),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_1039),
.B(n_1047),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_1034),
.Y(n_1205)
);

NAND2xp33_ASAP7_75t_L g1206 ( 
.A(n_1153),
.B(n_1145),
.Y(n_1206)
);

OA21x2_ASAP7_75t_L g1207 ( 
.A1(n_1016),
.A2(n_1125),
.B(n_1060),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1112),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1012),
.Y(n_1209)
);

AOI211x1_ASAP7_75t_L g1210 ( 
.A1(n_1129),
.A2(n_1058),
.B(n_1130),
.C(n_1104),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1157),
.B(n_1020),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_1140),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1044),
.B(n_1046),
.Y(n_1213)
);

AO21x1_ASAP7_75t_L g1214 ( 
.A1(n_1108),
.A2(n_1125),
.B(n_1086),
.Y(n_1214)
);

AOI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1134),
.A2(n_1029),
.B1(n_1063),
.B2(n_1022),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1152),
.A2(n_1161),
.B(n_1146),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1163),
.A2(n_1150),
.B(n_1158),
.Y(n_1217)
);

AO31x2_ASAP7_75t_L g1218 ( 
.A1(n_1086),
.A2(n_1062),
.A3(n_1060),
.B(n_1057),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1018),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_1140),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1021),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1078),
.B(n_1055),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1115),
.B(n_1116),
.Y(n_1223)
);

A2O1A1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1147),
.A2(n_1148),
.B(n_1119),
.C(n_1099),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1034),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1059),
.B(n_1061),
.Y(n_1226)
);

AOI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1029),
.A2(n_1149),
.B1(n_1049),
.B2(n_1122),
.Y(n_1227)
);

AO31x2_ASAP7_75t_L g1228 ( 
.A1(n_1062),
.A2(n_1057),
.A3(n_1100),
.B(n_1088),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1150),
.A2(n_1164),
.B(n_1100),
.Y(n_1229)
);

AO32x2_ASAP7_75t_L g1230 ( 
.A1(n_1042),
.A2(n_1092),
.A3(n_1095),
.B1(n_1136),
.B2(n_1102),
.Y(n_1230)
);

AOI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1133),
.A2(n_1101),
.B(n_1088),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1150),
.A2(n_1083),
.B(n_1082),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1038),
.A2(n_1040),
.B(n_1037),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1043),
.Y(n_1234)
);

AOI21xp33_ASAP7_75t_L g1235 ( 
.A1(n_1037),
.A2(n_1139),
.B(n_1154),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1077),
.A2(n_1139),
.B(n_1155),
.Y(n_1236)
);

BUFx10_ASAP7_75t_L g1237 ( 
.A(n_1045),
.Y(n_1237)
);

OR2x6_ASAP7_75t_L g1238 ( 
.A(n_1011),
.B(n_1113),
.Y(n_1238)
);

AOI31xp67_ASAP7_75t_L g1239 ( 
.A1(n_1136),
.A2(n_1093),
.A3(n_1121),
.B(n_1091),
.Y(n_1239)
);

OAI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1127),
.A2(n_1129),
.B(n_1096),
.Y(n_1240)
);

INVx6_ASAP7_75t_L g1241 ( 
.A(n_1114),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1053),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1085),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1084),
.Y(n_1244)
);

O2A1O1Ixp5_ASAP7_75t_L g1245 ( 
.A1(n_1127),
.A2(n_1162),
.B(n_1138),
.C(n_1124),
.Y(n_1245)
);

AO21x1_ASAP7_75t_L g1246 ( 
.A1(n_1162),
.A2(n_1136),
.B(n_1142),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1094),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1103),
.A2(n_1105),
.B(n_1111),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_1090),
.B(n_1126),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1167),
.A2(n_1142),
.B(n_1137),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1137),
.A2(n_1109),
.B(n_1106),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1008),
.A2(n_1066),
.B(n_1064),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1115),
.B(n_1116),
.Y(n_1253)
);

O2A1O1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1143),
.A2(n_1008),
.B(n_1064),
.C(n_1066),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1110),
.A2(n_1048),
.B1(n_1167),
.B2(n_1031),
.Y(n_1255)
);

O2A1O1Ixp5_ASAP7_75t_SL g1256 ( 
.A1(n_1102),
.A2(n_1106),
.B(n_1110),
.C(n_1149),
.Y(n_1256)
);

AOI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1167),
.A2(n_1102),
.B(n_1019),
.Y(n_1257)
);

OA21x2_ASAP7_75t_L g1258 ( 
.A1(n_1071),
.A2(n_1011),
.B(n_1019),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1019),
.B(n_1051),
.Y(n_1259)
);

AO31x2_ASAP7_75t_L g1260 ( 
.A1(n_1051),
.A2(n_1054),
.A3(n_1113),
.B(n_1117),
.Y(n_1260)
);

NAND2x1p5_ASAP7_75t_L g1261 ( 
.A(n_1090),
.B(n_1051),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1054),
.Y(n_1262)
);

INVxp67_ASAP7_75t_SL g1263 ( 
.A(n_1054),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1113),
.Y(n_1264)
);

BUFx4f_ASAP7_75t_SL g1265 ( 
.A(n_1117),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1033),
.B(n_1117),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1079),
.B(n_1128),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_1074),
.B(n_691),
.Y(n_1268)
);

AOI31xp67_ASAP7_75t_L g1269 ( 
.A1(n_1013),
.A2(n_1014),
.A3(n_1005),
.B(n_801),
.Y(n_1269)
);

CKINVDCx16_ASAP7_75t_R g1270 ( 
.A(n_1047),
.Y(n_1270)
);

NAND3xp33_ASAP7_75t_L g1271 ( 
.A(n_1089),
.B(n_848),
.C(n_692),
.Y(n_1271)
);

O2A1O1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1073),
.A2(n_848),
.B(n_692),
.C(n_1089),
.Y(n_1272)
);

A2O1A1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1073),
.A2(n_848),
.B(n_777),
.C(n_692),
.Y(n_1273)
);

AO31x2_ASAP7_75t_L g1274 ( 
.A1(n_1165),
.A2(n_1017),
.A3(n_1166),
.B(n_1160),
.Y(n_1274)
);

O2A1O1Ixp5_ASAP7_75t_L g1275 ( 
.A1(n_1013),
.A2(n_1014),
.B(n_917),
.C(n_1005),
.Y(n_1275)
);

AOI21x1_ASAP7_75t_SL g1276 ( 
.A1(n_1072),
.A2(n_1075),
.B(n_1099),
.Y(n_1276)
);

AOI221xp5_ASAP7_75t_L g1277 ( 
.A1(n_1029),
.A2(n_848),
.B1(n_1098),
.B2(n_1089),
.C(n_538),
.Y(n_1277)
);

INVx2_ASAP7_75t_SL g1278 ( 
.A(n_1076),
.Y(n_1278)
);

AOI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1130),
.A2(n_1014),
.B(n_1013),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1035),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1035),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1151),
.A2(n_1026),
.B(n_1030),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1135),
.A2(n_1025),
.B(n_1132),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1074),
.B(n_1023),
.Y(n_1284)
);

INVxp67_ASAP7_75t_L g1285 ( 
.A(n_1015),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1009),
.B(n_960),
.Y(n_1286)
);

NAND3xp33_ASAP7_75t_SL g1287 ( 
.A(n_1089),
.B(n_848),
.C(n_692),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1151),
.A2(n_1026),
.B(n_1030),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_SL g1289 ( 
.A1(n_1107),
.A2(n_570),
.B1(n_708),
.B2(n_411),
.Y(n_1289)
);

O2A1O1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1073),
.A2(n_848),
.B(n_692),
.C(n_1089),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1128),
.B(n_839),
.Y(n_1291)
);

BUFx12f_ASAP7_75t_L g1292 ( 
.A(n_1087),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1151),
.A2(n_1026),
.B(n_1030),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1151),
.A2(n_1026),
.B(n_1030),
.Y(n_1294)
);

O2A1O1Ixp33_ASAP7_75t_SL g1295 ( 
.A1(n_1013),
.A2(n_1014),
.B(n_1003),
.C(n_926),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1140),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1128),
.B(n_839),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1128),
.B(n_839),
.Y(n_1298)
);

O2A1O1Ixp33_ASAP7_75t_SL g1299 ( 
.A1(n_1013),
.A2(n_1014),
.B(n_1003),
.C(n_926),
.Y(n_1299)
);

AOI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1130),
.A2(n_1014),
.B(n_1013),
.Y(n_1300)
);

O2A1O1Ixp5_ASAP7_75t_L g1301 ( 
.A1(n_1013),
.A2(n_1014),
.B(n_917),
.C(n_1005),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1035),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1114),
.B(n_1078),
.Y(n_1303)
);

O2A1O1Ixp33_ASAP7_75t_L g1304 ( 
.A1(n_1073),
.A2(n_848),
.B(n_692),
.C(n_1089),
.Y(n_1304)
);

NOR2xp67_ASAP7_75t_L g1305 ( 
.A(n_1027),
.B(n_653),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1035),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1128),
.B(n_839),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1128),
.B(n_839),
.Y(n_1308)
);

AOI221x1_ASAP7_75t_L g1309 ( 
.A1(n_1073),
.A2(n_848),
.B1(n_692),
.B2(n_1108),
.C(n_1125),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1128),
.A2(n_777),
.B1(n_533),
.B2(n_652),
.Y(n_1310)
);

BUFx10_ASAP7_75t_L g1311 ( 
.A(n_1052),
.Y(n_1311)
);

OA21x2_ASAP7_75t_L g1312 ( 
.A1(n_1135),
.A2(n_1025),
.B(n_1017),
.Y(n_1312)
);

AND2x4_ASAP7_75t_L g1313 ( 
.A(n_1114),
.B(n_1078),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1151),
.A2(n_1026),
.B(n_1030),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1144),
.A2(n_783),
.B(n_817),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_SL g1316 ( 
.A(n_1074),
.B(n_1107),
.Y(n_1316)
);

O2A1O1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1073),
.A2(n_848),
.B(n_692),
.C(n_1089),
.Y(n_1317)
);

NAND3xp33_ASAP7_75t_L g1318 ( 
.A(n_1089),
.B(n_848),
.C(n_692),
.Y(n_1318)
);

OR2x2_ASAP7_75t_L g1319 ( 
.A(n_1009),
.B(n_960),
.Y(n_1319)
);

AO31x2_ASAP7_75t_L g1320 ( 
.A1(n_1165),
.A2(n_1017),
.A3(n_1166),
.B(n_1160),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1140),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1144),
.A2(n_783),
.B(n_817),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1135),
.A2(n_1025),
.B(n_1132),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1074),
.B(n_1023),
.Y(n_1324)
);

A2O1A1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1073),
.A2(n_848),
.B(n_777),
.C(n_692),
.Y(n_1325)
);

BUFx2_ASAP7_75t_L g1326 ( 
.A(n_1223),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1277),
.A2(n_1287),
.B1(n_1271),
.B2(n_1318),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1252),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1277),
.A2(n_1215),
.B1(n_1213),
.B2(n_1188),
.Y(n_1329)
);

BUFx3_ASAP7_75t_L g1330 ( 
.A(n_1241),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_SL g1331 ( 
.A1(n_1289),
.A2(n_1204),
.B1(n_1270),
.B2(n_1311),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1226),
.A2(n_1268),
.B1(n_1227),
.B2(n_1255),
.Y(n_1332)
);

INVx3_ASAP7_75t_L g1333 ( 
.A(n_1279),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1176),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1171),
.A2(n_1200),
.B1(n_1189),
.B2(n_1184),
.Y(n_1335)
);

OAI21xp5_ASAP7_75t_SL g1336 ( 
.A1(n_1171),
.A2(n_1290),
.B(n_1272),
.Y(n_1336)
);

HB1xp67_ASAP7_75t_SL g1337 ( 
.A(n_1169),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1183),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_L g1339 ( 
.A(n_1193),
.Y(n_1339)
);

BUFx8_ASAP7_75t_L g1340 ( 
.A(n_1292),
.Y(n_1340)
);

CKINVDCx11_ASAP7_75t_R g1341 ( 
.A(n_1191),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_1193),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1180),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1253),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1306),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1189),
.A2(n_1325),
.B1(n_1273),
.B2(n_1198),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1172),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1206),
.A2(n_1324),
.B1(n_1284),
.B2(n_1316),
.Y(n_1348)
);

BUFx2_ASAP7_75t_L g1349 ( 
.A(n_1196),
.Y(n_1349)
);

BUFx12f_ASAP7_75t_L g1350 ( 
.A(n_1185),
.Y(n_1350)
);

OAI22xp33_ASAP7_75t_SL g1351 ( 
.A1(n_1198),
.A2(n_1240),
.B1(n_1298),
.B2(n_1308),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1185),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1222),
.A2(n_1179),
.B1(n_1310),
.B2(n_1311),
.Y(n_1353)
);

CKINVDCx11_ASAP7_75t_R g1354 ( 
.A(n_1192),
.Y(n_1354)
);

INVx3_ASAP7_75t_L g1355 ( 
.A(n_1300),
.Y(n_1355)
);

INVx1_ASAP7_75t_SL g1356 ( 
.A(n_1286),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1310),
.A2(n_1174),
.B1(n_1235),
.B2(n_1214),
.Y(n_1357)
);

CKINVDCx11_ASAP7_75t_R g1358 ( 
.A(n_1192),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1174),
.A2(n_1235),
.B1(n_1240),
.B2(n_1236),
.Y(n_1359)
);

INVx1_ASAP7_75t_SL g1360 ( 
.A(n_1319),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1280),
.Y(n_1361)
);

BUFx6f_ASAP7_75t_L g1362 ( 
.A(n_1193),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1236),
.A2(n_1168),
.B1(n_1267),
.B2(n_1249),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1267),
.A2(n_1195),
.B1(n_1297),
.B2(n_1308),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1291),
.B(n_1297),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1272),
.A2(n_1304),
.B1(n_1290),
.B2(n_1317),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1281),
.Y(n_1367)
);

AO22x1_ASAP7_75t_L g1368 ( 
.A1(n_1186),
.A2(n_1266),
.B1(n_1291),
.B2(n_1298),
.Y(n_1368)
);

BUFx10_ASAP7_75t_L g1369 ( 
.A(n_1243),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1302),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1307),
.A2(n_1305),
.B1(n_1211),
.B2(n_1220),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1304),
.A2(n_1317),
.B1(n_1307),
.B2(n_1203),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1211),
.B(n_1170),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1187),
.Y(n_1374)
);

OAI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1309),
.A2(n_1186),
.B1(n_1192),
.B2(n_1225),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1224),
.B(n_1190),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1212),
.A2(n_1321),
.B1(n_1296),
.B2(n_1220),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_SL g1378 ( 
.A1(n_1205),
.A2(n_1243),
.B1(n_1283),
.B2(n_1323),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1170),
.B(n_1285),
.Y(n_1379)
);

OAI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1243),
.A2(n_1212),
.B1(n_1321),
.B2(n_1296),
.Y(n_1380)
);

CKINVDCx20_ASAP7_75t_R g1381 ( 
.A(n_1265),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_SL g1382 ( 
.A1(n_1283),
.A2(n_1323),
.B1(n_1194),
.B2(n_1173),
.Y(n_1382)
);

INVx3_ASAP7_75t_L g1383 ( 
.A(n_1216),
.Y(n_1383)
);

AOI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1303),
.A2(n_1313),
.B1(n_1278),
.B2(n_1241),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1202),
.Y(n_1385)
);

INVx1_ASAP7_75t_SL g1386 ( 
.A(n_1303),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1246),
.A2(n_1313),
.B1(n_1244),
.B2(n_1234),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1208),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1209),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1219),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1194),
.B(n_1221),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1242),
.A2(n_1247),
.B1(n_1250),
.B2(n_1258),
.Y(n_1392)
);

CKINVDCx11_ASAP7_75t_R g1393 ( 
.A(n_1237),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_SL g1394 ( 
.A1(n_1173),
.A2(n_1258),
.B1(n_1201),
.B2(n_1207),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1250),
.A2(n_1248),
.B1(n_1207),
.B2(n_1312),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_1261),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_1237),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1251),
.Y(n_1398)
);

INVxp67_ASAP7_75t_SL g1399 ( 
.A(n_1259),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1264),
.A2(n_1233),
.B1(n_1322),
.B2(n_1315),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1259),
.Y(n_1401)
);

BUFx2_ASAP7_75t_SL g1402 ( 
.A(n_1193),
.Y(n_1402)
);

BUFx10_ASAP7_75t_L g1403 ( 
.A(n_1238),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_SL g1404 ( 
.A(n_1275),
.B(n_1301),
.Y(n_1404)
);

CKINVDCx6p67_ASAP7_75t_R g1405 ( 
.A(n_1238),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1210),
.A2(n_1261),
.B1(n_1178),
.B2(n_1263),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1322),
.A2(n_1315),
.B1(n_1262),
.B2(n_1229),
.Y(n_1407)
);

BUFx12f_ASAP7_75t_L g1408 ( 
.A(n_1238),
.Y(n_1408)
);

INVx6_ASAP7_75t_L g1409 ( 
.A(n_1260),
.Y(n_1409)
);

INVx1_ASAP7_75t_SL g1410 ( 
.A(n_1177),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_SL g1411 ( 
.A1(n_1256),
.A2(n_1229),
.B1(n_1239),
.B2(n_1276),
.Y(n_1411)
);

CKINVDCx11_ASAP7_75t_R g1412 ( 
.A(n_1260),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_SL g1413 ( 
.A1(n_1231),
.A2(n_1217),
.B(n_1254),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1245),
.Y(n_1414)
);

INVx1_ASAP7_75t_SL g1415 ( 
.A(n_1177),
.Y(n_1415)
);

BUFx4f_ASAP7_75t_SL g1416 ( 
.A(n_1254),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1274),
.B(n_1320),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_SL g1418 ( 
.A1(n_1217),
.A2(n_1295),
.B1(n_1299),
.B2(n_1230),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1320),
.Y(n_1419)
);

BUFx2_ASAP7_75t_L g1420 ( 
.A(n_1320),
.Y(n_1420)
);

CKINVDCx20_ASAP7_75t_R g1421 ( 
.A(n_1232),
.Y(n_1421)
);

OAI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1257),
.A2(n_1232),
.B1(n_1182),
.B2(n_1230),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1269),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1182),
.A2(n_1197),
.B1(n_1199),
.B2(n_1282),
.Y(n_1424)
);

BUFx2_ASAP7_75t_SL g1425 ( 
.A(n_1175),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_1175),
.Y(n_1426)
);

BUFx2_ASAP7_75t_L g1427 ( 
.A(n_1218),
.Y(n_1427)
);

CKINVDCx6p67_ASAP7_75t_R g1428 ( 
.A(n_1218),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1288),
.A2(n_1314),
.B1(n_1294),
.B2(n_1293),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1181),
.Y(n_1430)
);

AOI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1230),
.A2(n_1218),
.B1(n_1228),
.B2(n_1181),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_SL g1432 ( 
.A1(n_1228),
.A2(n_708),
.B1(n_619),
.B2(n_1289),
.Y(n_1432)
);

AOI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1228),
.A2(n_848),
.B1(n_708),
.B2(n_1277),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1181),
.Y(n_1434)
);

BUFx2_ASAP7_75t_L g1435 ( 
.A(n_1223),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1176),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1277),
.A2(n_848),
.B1(n_1287),
.B2(n_692),
.Y(n_1437)
);

INVx1_ASAP7_75t_SL g1438 ( 
.A(n_1180),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1277),
.A2(n_848),
.B1(n_1287),
.B2(n_692),
.Y(n_1439)
);

OAI21xp33_ASAP7_75t_L g1440 ( 
.A1(n_1277),
.A2(n_848),
.B(n_708),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1176),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1277),
.A2(n_848),
.B1(n_1287),
.B2(n_692),
.Y(n_1442)
);

BUFx4f_ASAP7_75t_SL g1443 ( 
.A(n_1292),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1176),
.Y(n_1444)
);

CKINVDCx20_ASAP7_75t_R g1445 ( 
.A(n_1191),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1176),
.Y(n_1446)
);

OAI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1227),
.A2(n_1215),
.B1(n_619),
.B2(n_651),
.Y(n_1447)
);

BUFx6f_ASAP7_75t_L g1448 ( 
.A(n_1193),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1176),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1277),
.A2(n_848),
.B1(n_1287),
.B2(n_692),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1176),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1277),
.A2(n_848),
.B1(n_1287),
.B2(n_692),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1176),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1180),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1176),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1176),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1171),
.A2(n_708),
.B1(n_1277),
.B2(n_1215),
.Y(n_1457)
);

CKINVDCx20_ASAP7_75t_R g1458 ( 
.A(n_1191),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1176),
.Y(n_1459)
);

OAI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1227),
.A2(n_1215),
.B1(n_619),
.B2(n_651),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1176),
.Y(n_1461)
);

CKINVDCx20_ASAP7_75t_R g1462 ( 
.A(n_1191),
.Y(n_1462)
);

BUFx10_ASAP7_75t_L g1463 ( 
.A(n_1266),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1180),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1429),
.A2(n_1424),
.B(n_1383),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1366),
.B(n_1372),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1412),
.Y(n_1467)
);

AOI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1457),
.A2(n_1440),
.B1(n_1327),
.B2(n_1336),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1326),
.B(n_1344),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1326),
.B(n_1344),
.Y(n_1470)
);

OAI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1437),
.A2(n_1442),
.B(n_1439),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1349),
.Y(n_1472)
);

INVx2_ASAP7_75t_SL g1473 ( 
.A(n_1403),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1430),
.Y(n_1474)
);

NAND2x1p5_ASAP7_75t_L g1475 ( 
.A(n_1404),
.B(n_1376),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1349),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1434),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1365),
.B(n_1373),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1419),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1346),
.B(n_1364),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1328),
.B(n_1383),
.Y(n_1481)
);

INVx3_ASAP7_75t_L g1482 ( 
.A(n_1409),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1435),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1435),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1356),
.B(n_1360),
.Y(n_1485)
);

INVx2_ASAP7_75t_SL g1486 ( 
.A(n_1403),
.Y(n_1486)
);

INVxp33_ASAP7_75t_SL g1487 ( 
.A(n_1354),
.Y(n_1487)
);

INVx3_ASAP7_75t_L g1488 ( 
.A(n_1409),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_SL g1489 ( 
.A1(n_1391),
.A2(n_1406),
.B(n_1363),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1343),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1412),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1433),
.B(n_1382),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1431),
.B(n_1427),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1427),
.B(n_1420),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1423),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1420),
.Y(n_1496)
);

CKINVDCx20_ASAP7_75t_R g1497 ( 
.A(n_1445),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1426),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1426),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1454),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1414),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1376),
.B(n_1401),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1418),
.B(n_1374),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1398),
.Y(n_1504)
);

INVx1_ASAP7_75t_SL g1505 ( 
.A(n_1438),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1398),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1408),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1398),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1417),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1417),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1417),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1428),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_SL g1513 ( 
.A1(n_1335),
.A2(n_1416),
.B1(n_1421),
.B2(n_1447),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1374),
.B(n_1385),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1385),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1388),
.B(n_1357),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1425),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1410),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1428),
.Y(n_1519)
);

BUFx12f_ASAP7_75t_L g1520 ( 
.A(n_1341),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1415),
.Y(n_1521)
);

AOI221xp5_ASAP7_75t_L g1522 ( 
.A1(n_1450),
.A2(n_1452),
.B1(n_1460),
.B2(n_1329),
.C(n_1332),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1333),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1464),
.Y(n_1524)
);

OAI222xp33_ASAP7_75t_L g1525 ( 
.A1(n_1432),
.A2(n_1359),
.B1(n_1353),
.B2(n_1331),
.C1(n_1348),
.C2(n_1371),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_SL g1526 ( 
.A1(n_1445),
.A2(n_1462),
.B1(n_1458),
.B2(n_1381),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1333),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1355),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1421),
.B(n_1334),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1386),
.B(n_1463),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1379),
.B(n_1399),
.Y(n_1531)
);

OA21x2_ASAP7_75t_L g1532 ( 
.A1(n_1413),
.A2(n_1404),
.B(n_1407),
.Y(n_1532)
);

OA21x2_ASAP7_75t_L g1533 ( 
.A1(n_1395),
.A2(n_1400),
.B(n_1387),
.Y(n_1533)
);

OAI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1355),
.A2(n_1392),
.B(n_1370),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1347),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1453),
.Y(n_1536)
);

INVx2_ASAP7_75t_SL g1537 ( 
.A(n_1403),
.Y(n_1537)
);

BUFx4f_ASAP7_75t_L g1538 ( 
.A(n_1339),
.Y(n_1538)
);

INVx8_ASAP7_75t_L g1539 ( 
.A(n_1339),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1456),
.B(n_1367),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1361),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1351),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1422),
.Y(n_1543)
);

OAI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1378),
.A2(n_1375),
.B(n_1394),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1389),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1390),
.Y(n_1546)
);

BUFx3_ASAP7_75t_L g1547 ( 
.A(n_1408),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1338),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1345),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1436),
.Y(n_1550)
);

INVx11_ASAP7_75t_L g1551 ( 
.A(n_1340),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1441),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1444),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1446),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1449),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1451),
.Y(n_1556)
);

AO21x2_ASAP7_75t_L g1557 ( 
.A1(n_1380),
.A2(n_1461),
.B(n_1459),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1455),
.Y(n_1558)
);

NOR2x1p5_ASAP7_75t_L g1559 ( 
.A(n_1405),
.B(n_1396),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1497),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1529),
.B(n_1411),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1535),
.Y(n_1562)
);

OAI21x1_ASAP7_75t_SL g1563 ( 
.A1(n_1489),
.A2(n_1377),
.B(n_1368),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1468),
.A2(n_1337),
.B1(n_1384),
.B2(n_1397),
.Y(n_1564)
);

AOI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1468),
.A2(n_1462),
.B1(n_1458),
.B2(n_1463),
.Y(n_1565)
);

INVx4_ASAP7_75t_L g1566 ( 
.A(n_1539),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1529),
.B(n_1463),
.Y(n_1567)
);

AO21x2_ASAP7_75t_L g1568 ( 
.A1(n_1489),
.A2(n_1402),
.B(n_1405),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1469),
.B(n_1358),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1469),
.B(n_1358),
.Y(n_1570)
);

AOI21xp5_ASAP7_75t_L g1571 ( 
.A1(n_1471),
.A2(n_1448),
.B(n_1339),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1470),
.B(n_1354),
.Y(n_1572)
);

AO32x2_ASAP7_75t_L g1573 ( 
.A1(n_1473),
.A2(n_1393),
.A3(n_1397),
.B1(n_1369),
.B2(n_1341),
.Y(n_1573)
);

OR2x6_ASAP7_75t_L g1574 ( 
.A(n_1475),
.B(n_1350),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1470),
.B(n_1543),
.Y(n_1575)
);

AOI221xp5_ASAP7_75t_L g1576 ( 
.A1(n_1522),
.A2(n_1352),
.B1(n_1330),
.B2(n_1381),
.C(n_1342),
.Y(n_1576)
);

AO21x2_ASAP7_75t_L g1577 ( 
.A1(n_1544),
.A2(n_1448),
.B(n_1339),
.Y(n_1577)
);

AOI221xp5_ASAP7_75t_L g1578 ( 
.A1(n_1492),
.A2(n_1352),
.B1(n_1330),
.B2(n_1342),
.C(n_1362),
.Y(n_1578)
);

INVxp67_ASAP7_75t_L g1579 ( 
.A(n_1485),
.Y(n_1579)
);

A2O1A1Ixp33_ASAP7_75t_L g1580 ( 
.A1(n_1492),
.A2(n_1466),
.B(n_1513),
.C(n_1480),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1483),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1466),
.B(n_1393),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1546),
.Y(n_1583)
);

A2O1A1Ixp33_ASAP7_75t_L g1584 ( 
.A1(n_1478),
.A2(n_1342),
.B(n_1362),
.C(n_1369),
.Y(n_1584)
);

A2O1A1Ixp33_ASAP7_75t_L g1585 ( 
.A1(n_1542),
.A2(n_1342),
.B(n_1362),
.C(n_1369),
.Y(n_1585)
);

A2O1A1Ixp33_ASAP7_75t_L g1586 ( 
.A1(n_1542),
.A2(n_1350),
.B(n_1340),
.C(n_1443),
.Y(n_1586)
);

AND2x4_ASAP7_75t_L g1587 ( 
.A(n_1509),
.B(n_1510),
.Y(n_1587)
);

A2O1A1Ixp33_ASAP7_75t_L g1588 ( 
.A1(n_1516),
.A2(n_1340),
.B(n_1503),
.C(n_1467),
.Y(n_1588)
);

AO32x2_ASAP7_75t_L g1589 ( 
.A1(n_1473),
.A2(n_1486),
.A3(n_1537),
.B1(n_1475),
.B2(n_1494),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1484),
.B(n_1490),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1502),
.B(n_1503),
.Y(n_1591)
);

OAI21x1_ASAP7_75t_L g1592 ( 
.A1(n_1465),
.A2(n_1534),
.B(n_1495),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1472),
.B(n_1476),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1514),
.B(n_1500),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1514),
.B(n_1524),
.Y(n_1595)
);

A2O1A1Ixp33_ASAP7_75t_SL g1596 ( 
.A1(n_1530),
.A2(n_1519),
.B(n_1512),
.C(n_1501),
.Y(n_1596)
);

AO21x2_ASAP7_75t_L g1597 ( 
.A1(n_1517),
.A2(n_1495),
.B(n_1501),
.Y(n_1597)
);

AO32x2_ASAP7_75t_L g1598 ( 
.A1(n_1486),
.A2(n_1537),
.A3(n_1475),
.B1(n_1494),
.B2(n_1493),
.Y(n_1598)
);

OA21x2_ASAP7_75t_L g1599 ( 
.A1(n_1534),
.A2(n_1477),
.B(n_1474),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1531),
.B(n_1493),
.Y(n_1600)
);

O2A1O1Ixp33_ASAP7_75t_SL g1601 ( 
.A1(n_1525),
.A2(n_1519),
.B(n_1487),
.C(n_1496),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1516),
.B(n_1540),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1467),
.A2(n_1491),
.B1(n_1520),
.B2(n_1547),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1540),
.B(n_1467),
.Y(n_1604)
);

INVx3_ASAP7_75t_L g1605 ( 
.A(n_1481),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1511),
.B(n_1541),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1541),
.B(n_1527),
.Y(n_1607)
);

OAI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1532),
.A2(n_1538),
.B(n_1505),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1515),
.Y(n_1609)
);

O2A1O1Ixp33_ASAP7_75t_SL g1610 ( 
.A1(n_1496),
.A2(n_1498),
.B(n_1499),
.C(n_1556),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1540),
.B(n_1536),
.Y(n_1611)
);

AND2x4_ASAP7_75t_L g1612 ( 
.A(n_1482),
.B(n_1488),
.Y(n_1612)
);

OAI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1532),
.A2(n_1538),
.B(n_1533),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1518),
.B(n_1521),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1523),
.B(n_1528),
.Y(n_1615)
);

AOI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1491),
.A2(n_1520),
.B1(n_1507),
.B2(n_1547),
.Y(n_1616)
);

BUFx6f_ASAP7_75t_L g1617 ( 
.A(n_1507),
.Y(n_1617)
);

A2O1A1Ixp33_ASAP7_75t_L g1618 ( 
.A1(n_1491),
.A2(n_1538),
.B(n_1559),
.C(n_1512),
.Y(n_1618)
);

AOI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1532),
.A2(n_1538),
.B(n_1533),
.Y(n_1619)
);

A2O1A1Ixp33_ASAP7_75t_L g1620 ( 
.A1(n_1559),
.A2(n_1512),
.B(n_1507),
.C(n_1547),
.Y(n_1620)
);

O2A1O1Ixp33_ASAP7_75t_L g1621 ( 
.A1(n_1532),
.A2(n_1558),
.B(n_1549),
.C(n_1556),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1551),
.A2(n_1526),
.B1(n_1555),
.B2(n_1554),
.Y(n_1622)
);

AO21x1_ASAP7_75t_L g1623 ( 
.A1(n_1548),
.A2(n_1558),
.B(n_1555),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1523),
.B(n_1528),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1598),
.B(n_1506),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1583),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1600),
.B(n_1498),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1583),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1598),
.B(n_1508),
.Y(n_1629)
);

INVxp67_ASAP7_75t_SL g1630 ( 
.A(n_1623),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1597),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1614),
.B(n_1599),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1598),
.B(n_1506),
.Y(n_1633)
);

INVxp67_ASAP7_75t_L g1634 ( 
.A(n_1581),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1615),
.Y(n_1635)
);

INVxp67_ASAP7_75t_L g1636 ( 
.A(n_1607),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1609),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1605),
.B(n_1508),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1615),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1576),
.A2(n_1533),
.B1(n_1557),
.B2(n_1553),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1562),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1609),
.Y(n_1642)
);

AOI222xp33_ASAP7_75t_L g1643 ( 
.A1(n_1580),
.A2(n_1564),
.B1(n_1579),
.B2(n_1582),
.C1(n_1622),
.C2(n_1578),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1624),
.Y(n_1644)
);

INVxp67_ASAP7_75t_L g1645 ( 
.A(n_1590),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1589),
.B(n_1504),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1575),
.B(n_1545),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1611),
.B(n_1606),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1606),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1592),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1575),
.B(n_1479),
.Y(n_1651)
);

BUFx3_ASAP7_75t_L g1652 ( 
.A(n_1574),
.Y(n_1652)
);

AOI221xp5_ASAP7_75t_L g1653 ( 
.A1(n_1630),
.A2(n_1601),
.B1(n_1580),
.B2(n_1621),
.C(n_1582),
.Y(n_1653)
);

OAI33xp33_ASAP7_75t_L g1654 ( 
.A1(n_1645),
.A2(n_1553),
.A3(n_1554),
.B1(n_1552),
.B2(n_1550),
.B3(n_1549),
.Y(n_1654)
);

OAI21xp5_ASAP7_75t_SL g1655 ( 
.A1(n_1643),
.A2(n_1565),
.B(n_1640),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1635),
.B(n_1589),
.Y(n_1656)
);

INVx3_ASAP7_75t_L g1657 ( 
.A(n_1635),
.Y(n_1657)
);

BUFx6f_ASAP7_75t_L g1658 ( 
.A(n_1652),
.Y(n_1658)
);

AND2x4_ASAP7_75t_L g1659 ( 
.A(n_1652),
.B(n_1587),
.Y(n_1659)
);

NAND4xp25_ASAP7_75t_L g1660 ( 
.A(n_1643),
.B(n_1603),
.C(n_1601),
.D(n_1616),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1645),
.B(n_1593),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1640),
.A2(n_1563),
.B1(n_1577),
.B2(n_1561),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1637),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1635),
.B(n_1589),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1637),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1635),
.B(n_1591),
.Y(n_1666)
);

INVx4_ASAP7_75t_L g1667 ( 
.A(n_1652),
.Y(n_1667)
);

AOI222xp33_ASAP7_75t_L g1668 ( 
.A1(n_1630),
.A2(n_1613),
.B1(n_1561),
.B2(n_1608),
.C1(n_1588),
.C2(n_1591),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1637),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1652),
.A2(n_1577),
.B1(n_1567),
.B2(n_1604),
.Y(n_1670)
);

NAND3xp33_ASAP7_75t_L g1671 ( 
.A(n_1634),
.B(n_1571),
.C(n_1588),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1642),
.Y(n_1672)
);

NOR3xp33_ASAP7_75t_SL g1673 ( 
.A(n_1647),
.B(n_1586),
.C(n_1620),
.Y(n_1673)
);

NAND3xp33_ASAP7_75t_L g1674 ( 
.A(n_1634),
.B(n_1619),
.C(n_1596),
.Y(n_1674)
);

AOI221xp5_ASAP7_75t_L g1675 ( 
.A1(n_1647),
.A2(n_1586),
.B1(n_1602),
.B2(n_1610),
.C(n_1596),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1648),
.B(n_1594),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1642),
.Y(n_1677)
);

AOI221xp5_ASAP7_75t_L g1678 ( 
.A1(n_1651),
.A2(n_1610),
.B1(n_1595),
.B2(n_1550),
.C(n_1552),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1639),
.B(n_1587),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1642),
.Y(n_1680)
);

INVx2_ASAP7_75t_SL g1681 ( 
.A(n_1649),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1626),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1639),
.B(n_1644),
.Y(n_1683)
);

INVx3_ASAP7_75t_L g1684 ( 
.A(n_1644),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1628),
.Y(n_1685)
);

BUFx2_ASAP7_75t_L g1686 ( 
.A(n_1638),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1628),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1644),
.B(n_1587),
.Y(n_1688)
);

NOR3xp33_ASAP7_75t_L g1689 ( 
.A(n_1650),
.B(n_1620),
.C(n_1618),
.Y(n_1689)
);

BUFx3_ASAP7_75t_L g1690 ( 
.A(n_1627),
.Y(n_1690)
);

OAI22xp5_ASAP7_75t_SL g1691 ( 
.A1(n_1641),
.A2(n_1560),
.B1(n_1574),
.B2(n_1617),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1657),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1656),
.B(n_1625),
.Y(n_1693)
);

INVx3_ASAP7_75t_L g1694 ( 
.A(n_1657),
.Y(n_1694)
);

BUFx2_ASAP7_75t_L g1695 ( 
.A(n_1667),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1663),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1656),
.B(n_1625),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1664),
.B(n_1625),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1664),
.B(n_1629),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1686),
.B(n_1629),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1678),
.B(n_1636),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1681),
.B(n_1632),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1663),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1681),
.B(n_1632),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1665),
.B(n_1636),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1657),
.B(n_1632),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1665),
.Y(n_1707)
);

INVx1_ASAP7_75t_SL g1708 ( 
.A(n_1690),
.Y(n_1708)
);

AND2x4_ASAP7_75t_L g1709 ( 
.A(n_1667),
.B(n_1646),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1686),
.B(n_1629),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1669),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1669),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1684),
.B(n_1633),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1672),
.Y(n_1714)
);

HB1xp67_ASAP7_75t_L g1715 ( 
.A(n_1672),
.Y(n_1715)
);

INVx1_ASAP7_75t_SL g1716 ( 
.A(n_1690),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1684),
.B(n_1631),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1684),
.B(n_1633),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1677),
.B(n_1680),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1660),
.B(n_1560),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1661),
.B(n_1551),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1677),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1683),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1680),
.Y(n_1724)
);

INVx2_ASAP7_75t_SL g1725 ( 
.A(n_1658),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1682),
.Y(n_1726)
);

AOI22xp33_ASAP7_75t_L g1727 ( 
.A1(n_1653),
.A2(n_1574),
.B1(n_1568),
.B2(n_1612),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1682),
.B(n_1685),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1683),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1666),
.B(n_1633),
.Y(n_1730)
);

AND2x4_ASAP7_75t_L g1731 ( 
.A(n_1667),
.B(n_1646),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1715),
.Y(n_1732)
);

INVx3_ASAP7_75t_L g1733 ( 
.A(n_1709),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1701),
.B(n_1655),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1701),
.B(n_1675),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1708),
.B(n_1666),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1715),
.Y(n_1737)
);

INVxp67_ASAP7_75t_SL g1738 ( 
.A(n_1695),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1702),
.Y(n_1739)
);

INVx1_ASAP7_75t_SL g1740 ( 
.A(n_1708),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1702),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1709),
.B(n_1658),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1696),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1696),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1703),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1702),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1716),
.B(n_1674),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1716),
.B(n_1668),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1703),
.Y(n_1749)
);

INVxp67_ASAP7_75t_L g1750 ( 
.A(n_1720),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1704),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1704),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1707),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1709),
.B(n_1731),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1709),
.B(n_1658),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1727),
.B(n_1679),
.Y(n_1756)
);

NAND2x1p5_ASAP7_75t_L g1757 ( 
.A(n_1695),
.B(n_1658),
.Y(n_1757)
);

AND2x4_ASAP7_75t_L g1758 ( 
.A(n_1709),
.B(n_1689),
.Y(n_1758)
);

AOI32xp33_ASAP7_75t_SL g1759 ( 
.A1(n_1721),
.A2(n_1673),
.A3(n_1573),
.B1(n_1687),
.B2(n_1685),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1725),
.B(n_1679),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1707),
.Y(n_1761)
);

AND2x4_ASAP7_75t_SL g1762 ( 
.A(n_1731),
.B(n_1658),
.Y(n_1762)
);

NOR2x1_ASAP7_75t_L g1763 ( 
.A(n_1731),
.B(n_1671),
.Y(n_1763)
);

NAND2x1_ASAP7_75t_L g1764 ( 
.A(n_1731),
.B(n_1659),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_SL g1765 ( 
.A(n_1725),
.B(n_1691),
.Y(n_1765)
);

AOI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1725),
.A2(n_1662),
.B1(n_1574),
.B2(n_1659),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1711),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1704),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1706),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1711),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1712),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1705),
.B(n_1688),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1712),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1714),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_SL g1775 ( 
.A(n_1763),
.B(n_1670),
.Y(n_1775)
);

NAND5xp2_ASAP7_75t_L g1776 ( 
.A(n_1734),
.B(n_1618),
.C(n_1569),
.D(n_1570),
.E(n_1572),
.Y(n_1776)
);

INVx4_ASAP7_75t_L g1777 ( 
.A(n_1757),
.Y(n_1777)
);

INVx1_ASAP7_75t_SL g1778 ( 
.A(n_1740),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1735),
.B(n_1705),
.Y(n_1779)
);

BUFx2_ASAP7_75t_SL g1780 ( 
.A(n_1738),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1732),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1763),
.B(n_1731),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1772),
.B(n_1723),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1748),
.B(n_1723),
.Y(n_1784)
);

AOI22xp5_ASAP7_75t_SL g1785 ( 
.A1(n_1750),
.A2(n_1617),
.B1(n_1659),
.B2(n_1573),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1743),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_SL g1787 ( 
.A(n_1747),
.B(n_1659),
.Y(n_1787)
);

HB1xp67_ASAP7_75t_L g1788 ( 
.A(n_1732),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1743),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1765),
.B(n_1676),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1736),
.B(n_1723),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1757),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1744),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1739),
.B(n_1729),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1762),
.B(n_1693),
.Y(n_1795)
);

INVxp67_ASAP7_75t_SL g1796 ( 
.A(n_1757),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1739),
.B(n_1729),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1758),
.B(n_1729),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1737),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1758),
.B(n_1688),
.Y(n_1800)
);

NOR2x1p5_ASAP7_75t_SL g1801 ( 
.A(n_1741),
.B(n_1717),
.Y(n_1801)
);

OAI211xp5_ASAP7_75t_SL g1802 ( 
.A1(n_1766),
.A2(n_1717),
.B(n_1714),
.C(n_1722),
.Y(n_1802)
);

INVxp67_ASAP7_75t_L g1803 ( 
.A(n_1742),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1758),
.B(n_1730),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1758),
.B(n_1730),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1762),
.B(n_1693),
.Y(n_1806)
);

NOR2x1_ASAP7_75t_L g1807 ( 
.A(n_1737),
.B(n_1722),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1756),
.B(n_1730),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1744),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1746),
.B(n_1706),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_L g1811 ( 
.A(n_1778),
.B(n_1742),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1786),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1790),
.B(n_1779),
.Y(n_1813)
);

XNOR2x2_ASAP7_75t_L g1814 ( 
.A(n_1775),
.B(n_1759),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1781),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1786),
.Y(n_1816)
);

HB1xp67_ASAP7_75t_L g1817 ( 
.A(n_1780),
.Y(n_1817)
);

INVxp67_ASAP7_75t_SL g1818 ( 
.A(n_1782),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1803),
.B(n_1760),
.Y(n_1819)
);

INVxp67_ASAP7_75t_L g1820 ( 
.A(n_1780),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1784),
.B(n_1788),
.Y(n_1821)
);

INVx1_ASAP7_75t_SL g1822 ( 
.A(n_1782),
.Y(n_1822)
);

OAI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1785),
.A2(n_1764),
.B1(n_1759),
.B2(n_1762),
.Y(n_1823)
);

OAI21xp5_ASAP7_75t_L g1824 ( 
.A1(n_1802),
.A2(n_1755),
.B(n_1764),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1795),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1789),
.Y(n_1826)
);

AOI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1776),
.A2(n_1787),
.B(n_1796),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1799),
.B(n_1755),
.Y(n_1828)
);

OAI21xp5_ASAP7_75t_L g1829 ( 
.A1(n_1807),
.A2(n_1754),
.B(n_1749),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1795),
.B(n_1746),
.Y(n_1830)
);

AOI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1806),
.A2(n_1754),
.B1(n_1733),
.B2(n_1654),
.Y(n_1831)
);

AOI22xp5_ASAP7_75t_L g1832 ( 
.A1(n_1806),
.A2(n_1733),
.B1(n_1768),
.B2(n_1771),
.Y(n_1832)
);

AOI222xp33_ASAP7_75t_L g1833 ( 
.A1(n_1801),
.A2(n_1768),
.B1(n_1733),
.B2(n_1752),
.C1(n_1751),
.C2(n_1741),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1777),
.B(n_1733),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1798),
.B(n_1741),
.Y(n_1835)
);

NAND3xp33_ASAP7_75t_L g1836 ( 
.A(n_1777),
.B(n_1751),
.C(n_1752),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1820),
.B(n_1804),
.Y(n_1837)
);

BUFx2_ASAP7_75t_L g1838 ( 
.A(n_1817),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1815),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1815),
.Y(n_1840)
);

OAI32xp33_ASAP7_75t_L g1841 ( 
.A1(n_1814),
.A2(n_1777),
.A3(n_1805),
.B1(n_1792),
.B2(n_1808),
.Y(n_1841)
);

AOI32xp33_ASAP7_75t_L g1842 ( 
.A1(n_1823),
.A2(n_1807),
.A3(n_1792),
.B1(n_1800),
.B2(n_1791),
.Y(n_1842)
);

OR2x2_ASAP7_75t_L g1843 ( 
.A(n_1821),
.B(n_1830),
.Y(n_1843)
);

NAND3xp33_ASAP7_75t_L g1844 ( 
.A(n_1833),
.B(n_1793),
.C(n_1789),
.Y(n_1844)
);

HB1xp67_ASAP7_75t_L g1845 ( 
.A(n_1814),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1825),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1825),
.B(n_1783),
.Y(n_1847)
);

OAI22x1_ASAP7_75t_L g1848 ( 
.A1(n_1818),
.A2(n_1793),
.B1(n_1809),
.B2(n_1751),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1811),
.B(n_1809),
.Y(n_1849)
);

A2O1A1Ixp33_ASAP7_75t_L g1850 ( 
.A1(n_1827),
.A2(n_1813),
.B(n_1829),
.C(n_1836),
.Y(n_1850)
);

NOR2xp33_ASAP7_75t_L g1851 ( 
.A(n_1811),
.B(n_1783),
.Y(n_1851)
);

INVxp67_ASAP7_75t_L g1852 ( 
.A(n_1828),
.Y(n_1852)
);

INVxp67_ASAP7_75t_L g1853 ( 
.A(n_1822),
.Y(n_1853)
);

INVx2_ASAP7_75t_SL g1854 ( 
.A(n_1834),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1812),
.Y(n_1855)
);

INVx1_ASAP7_75t_SL g1856 ( 
.A(n_1834),
.Y(n_1856)
);

O2A1O1Ixp33_ASAP7_75t_L g1857 ( 
.A1(n_1845),
.A2(n_1824),
.B(n_1816),
.C(n_1826),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1838),
.B(n_1819),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1846),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1856),
.B(n_1854),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1846),
.Y(n_1861)
);

HB1xp67_ASAP7_75t_L g1862 ( 
.A(n_1845),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1847),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1839),
.Y(n_1864)
);

O2A1O1Ixp5_ASAP7_75t_L g1865 ( 
.A1(n_1841),
.A2(n_1835),
.B(n_1794),
.C(n_1797),
.Y(n_1865)
);

AOI222xp33_ASAP7_75t_L g1866 ( 
.A1(n_1850),
.A2(n_1801),
.B1(n_1752),
.B2(n_1769),
.C1(n_1773),
.C2(n_1745),
.Y(n_1866)
);

AOI222xp33_ASAP7_75t_L g1867 ( 
.A1(n_1850),
.A2(n_1769),
.B1(n_1745),
.B2(n_1749),
.C1(n_1753),
.C2(n_1761),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1848),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1859),
.Y(n_1869)
);

NOR2xp33_ASAP7_75t_L g1870 ( 
.A(n_1858),
.B(n_1852),
.Y(n_1870)
);

OAI211xp5_ASAP7_75t_SL g1871 ( 
.A1(n_1866),
.A2(n_1842),
.B(n_1853),
.C(n_1837),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1861),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1862),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1863),
.B(n_1851),
.Y(n_1874)
);

NOR3xp33_ASAP7_75t_L g1875 ( 
.A(n_1860),
.B(n_1840),
.C(n_1851),
.Y(n_1875)
);

AOI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1857),
.A2(n_1844),
.B(n_1849),
.Y(n_1876)
);

NAND3xp33_ASAP7_75t_SL g1877 ( 
.A(n_1867),
.B(n_1843),
.C(n_1832),
.Y(n_1877)
);

AOI22xp5_ASAP7_75t_L g1878 ( 
.A1(n_1862),
.A2(n_1831),
.B1(n_1855),
.B2(n_1794),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1868),
.Y(n_1879)
);

AOI221xp5_ASAP7_75t_L g1880 ( 
.A1(n_1876),
.A2(n_1868),
.B1(n_1865),
.B2(n_1864),
.C(n_1797),
.Y(n_1880)
);

OAI211xp5_ASAP7_75t_SL g1881 ( 
.A1(n_1874),
.A2(n_1810),
.B(n_1769),
.C(n_1773),
.Y(n_1881)
);

AOI221x1_ASAP7_75t_L g1882 ( 
.A1(n_1879),
.A2(n_1767),
.B1(n_1774),
.B2(n_1771),
.C(n_1770),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1873),
.Y(n_1883)
);

AOI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1871),
.A2(n_1810),
.B1(n_1774),
.B2(n_1770),
.Y(n_1884)
);

AOI22xp33_ASAP7_75t_L g1885 ( 
.A1(n_1877),
.A2(n_1767),
.B1(n_1761),
.B2(n_1753),
.Y(n_1885)
);

OAI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1878),
.A2(n_1717),
.B1(n_1694),
.B2(n_1700),
.Y(n_1886)
);

AOI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1880),
.A2(n_1870),
.B1(n_1875),
.B2(n_1872),
.Y(n_1887)
);

AOI211xp5_ASAP7_75t_L g1888 ( 
.A1(n_1881),
.A2(n_1869),
.B(n_1617),
.C(n_1584),
.Y(n_1888)
);

AOI22xp5_ASAP7_75t_L g1889 ( 
.A1(n_1886),
.A2(n_1617),
.B1(n_1700),
.B2(n_1710),
.Y(n_1889)
);

O2A1O1Ixp33_ASAP7_75t_L g1890 ( 
.A1(n_1883),
.A2(n_1584),
.B(n_1585),
.C(n_1706),
.Y(n_1890)
);

AOI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1885),
.A2(n_1884),
.B1(n_1710),
.B2(n_1700),
.Y(n_1891)
);

OAI221xp5_ASAP7_75t_SL g1892 ( 
.A1(n_1882),
.A2(n_1585),
.B1(n_1573),
.B2(n_1710),
.C(n_1693),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1887),
.Y(n_1893)
);

NOR2x1_ASAP7_75t_L g1894 ( 
.A(n_1890),
.B(n_1694),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1891),
.Y(n_1895)
);

BUFx3_ASAP7_75t_L g1896 ( 
.A(n_1889),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1888),
.Y(n_1897)
);

NOR3xp33_ASAP7_75t_L g1898 ( 
.A(n_1893),
.B(n_1892),
.C(n_1566),
.Y(n_1898)
);

AOI322xp5_ASAP7_75t_L g1899 ( 
.A1(n_1893),
.A2(n_1895),
.A3(n_1897),
.B1(n_1896),
.B2(n_1894),
.C1(n_1699),
.C2(n_1698),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1895),
.Y(n_1900)
);

HB1xp67_ASAP7_75t_L g1901 ( 
.A(n_1900),
.Y(n_1901)
);

OAI22xp5_ASAP7_75t_SL g1902 ( 
.A1(n_1901),
.A2(n_1899),
.B1(n_1898),
.B2(n_1573),
.Y(n_1902)
);

AOI22x1_ASAP7_75t_L g1903 ( 
.A1(n_1902),
.A2(n_1726),
.B1(n_1724),
.B2(n_1692),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1902),
.B(n_1694),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1904),
.Y(n_1905)
);

OAI22xp5_ASAP7_75t_L g1906 ( 
.A1(n_1903),
.A2(n_1692),
.B1(n_1694),
.B2(n_1697),
.Y(n_1906)
);

INVxp33_ASAP7_75t_SL g1907 ( 
.A(n_1905),
.Y(n_1907)
);

OAI21x1_ASAP7_75t_L g1908 ( 
.A1(n_1906),
.A2(n_1692),
.B(n_1699),
.Y(n_1908)
);

AOI22xp5_ASAP7_75t_L g1909 ( 
.A1(n_1907),
.A2(n_1699),
.B1(n_1697),
.B2(n_1698),
.Y(n_1909)
);

AOI222xp33_ASAP7_75t_L g1910 ( 
.A1(n_1909),
.A2(n_1908),
.B1(n_1726),
.B2(n_1724),
.C1(n_1728),
.C2(n_1719),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1910),
.Y(n_1911)
);

AOI221xp5_ASAP7_75t_L g1912 ( 
.A1(n_1911),
.A2(n_1719),
.B1(n_1728),
.B2(n_1698),
.C(n_1697),
.Y(n_1912)
);

AOI211xp5_ASAP7_75t_L g1913 ( 
.A1(n_1912),
.A2(n_1713),
.B(n_1718),
.C(n_1687),
.Y(n_1913)
);


endmodule