module fake_jpeg_18921_n_324 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_44),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_16),
.Y(n_44)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_44),
.A2(n_26),
.B1(n_22),
.B2(n_29),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_53),
.B1(n_44),
.B2(n_43),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_22),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_59),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_19),
.B1(n_32),
.B2(n_24),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_52),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_26),
.B1(n_29),
.B2(n_20),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_18),
.Y(n_94)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_19),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_30),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_41),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_51),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_88),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_59),
.B(n_28),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_66),
.B(n_69),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_50),
.A2(n_36),
.B(n_27),
.C(n_38),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_67),
.A2(n_92),
.B(n_40),
.C(n_55),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_36),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_68),
.Y(n_123)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_72),
.A2(n_43),
.B1(n_40),
.B2(n_42),
.Y(n_97)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_76),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_52),
.A2(n_26),
.B1(n_29),
.B2(n_27),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_47),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_77),
.A2(n_55),
.B1(n_40),
.B2(n_49),
.Y(n_108)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_79),
.Y(n_101)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_83),
.Y(n_113)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_45),
.A2(n_29),
.B1(n_20),
.B2(n_27),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

BUFx8_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_85),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_45),
.A2(n_20),
.B1(n_44),
.B2(n_28),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_47),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_24),
.B1(n_32),
.B2(n_25),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_17),
.B1(n_25),
.B2(n_34),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_63),
.Y(n_107)
);

FAx1_ASAP7_75t_SL g92 ( 
.A(n_57),
.B(n_43),
.CI(n_42),
.CON(n_92),
.SN(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_97),
.A2(n_105),
.B1(n_34),
.B2(n_70),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_61),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_98),
.A2(n_124),
.B(n_41),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_107),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_63),
.C(n_42),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_106),
.B(n_109),
.C(n_16),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_68),
.B(n_92),
.C(n_75),
.Y(n_109)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_65),
.A2(n_40),
.B1(n_49),
.B2(n_17),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_67),
.B(n_41),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_114),
.B(n_68),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_127),
.B(n_137),
.Y(n_180)
);

AO22x1_ASAP7_75t_SL g129 ( 
.A1(n_100),
.A2(n_77),
.B1(n_64),
.B2(n_71),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_136),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_131),
.A2(n_143),
.B1(n_116),
.B2(n_102),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_80),
.B1(n_64),
.B2(n_96),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_132),
.A2(n_153),
.B1(n_97),
.B2(n_111),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_116),
.A2(n_110),
.B1(n_125),
.B2(n_123),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_134),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_95),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_114),
.B(n_34),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_93),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_151),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_140),
.A2(n_148),
.B(n_102),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_87),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_141),
.B(n_146),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_109),
.A2(n_82),
.B1(n_78),
.B2(n_70),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_112),
.A2(n_85),
.B1(n_30),
.B2(n_21),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_106),
.B(n_85),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_155),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_119),
.B(n_21),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_113),
.B(n_21),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_147),
.B(n_149),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_31),
.B(n_18),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_33),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_18),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_107),
.B(n_60),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_152),
.B(n_102),
.Y(n_169)
);

OA21x2_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_31),
.B(n_60),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_104),
.Y(n_154)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_104),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_117),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_157),
.A2(n_0),
.B(n_1),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_158),
.A2(n_161),
.B1(n_172),
.B2(n_178),
.Y(n_193)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_128),
.A2(n_131),
.B1(n_133),
.B2(n_152),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_101),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_163),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_133),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_165),
.A2(n_164),
.B(n_169),
.Y(n_209)
);

NAND3xp33_ASAP7_75t_SL g166 ( 
.A(n_128),
.B(n_98),
.C(n_105),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_166),
.B(n_171),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_169),
.B(n_190),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_115),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_170),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_126),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_117),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_173),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_111),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_150),
.A2(n_98),
.B(n_97),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_175),
.A2(n_179),
.B(n_150),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_148),
.A2(n_97),
.B1(n_103),
.B2(n_99),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_155),
.A2(n_103),
.B1(n_99),
.B2(n_31),
.Y(n_179)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_130),
.Y(n_184)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_130),
.B(n_33),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_185),
.Y(n_218)
);

INVx13_ASAP7_75t_L g186 ( 
.A(n_136),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_145),
.B(n_16),
.C(n_30),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_153),
.C(n_142),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_138),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_129),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_144),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_192),
.A2(n_203),
.B(n_209),
.Y(n_238)
);

OA21x2_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_129),
.B(n_135),
.Y(n_195)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_195),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_181),
.Y(n_196)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_196),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_202),
.C(n_214),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_212),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_139),
.C(n_140),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_176),
.A2(n_135),
.B(n_151),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_143),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_198),
.Y(n_225)
);

OAI22x1_ASAP7_75t_SL g208 ( 
.A1(n_159),
.A2(n_153),
.B1(n_132),
.B2(n_31),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_208),
.A2(n_177),
.B1(n_175),
.B2(n_164),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_162),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_215),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_161),
.B(n_33),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_16),
.Y(n_213)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_30),
.C(n_21),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_162),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_172),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_216),
.A2(n_177),
.B1(n_167),
.B2(n_176),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_219),
.A2(n_165),
.B(n_157),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_204),
.Y(n_221)
);

NAND3xp33_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_207),
.C(n_209),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_223),
.A2(n_233),
.B1(n_239),
.B2(n_241),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_199),
.B(n_180),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_224),
.B(n_229),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_234),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_191),
.Y(n_228)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_228),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_200),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_230),
.A2(n_219),
.B1(n_208),
.B2(n_212),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_232),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_179),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_213),
.Y(n_235)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_200),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_SL g252 ( 
.A(n_236),
.B(n_217),
.C(n_218),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_216),
.A2(n_183),
.B1(n_167),
.B2(n_180),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_165),
.C(n_158),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_214),
.C(n_193),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_193),
.A2(n_189),
.B1(n_184),
.B2(n_182),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_207),
.Y(n_242)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_206),
.B(n_181),
.Y(n_243)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_192),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_247),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_191),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_257),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_203),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_248),
.A2(n_232),
.B(n_220),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_255),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_227),
.A2(n_218),
.B(n_194),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_250),
.A2(n_194),
.B(n_197),
.Y(n_274)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_252),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_211),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_195),
.C(n_217),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_259),
.C(n_223),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_195),
.C(n_168),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_220),
.B(n_186),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_261),
.A2(n_222),
.B1(n_196),
.B2(n_8),
.Y(n_276)
);

OAI21x1_ASAP7_75t_L g264 ( 
.A1(n_263),
.A2(n_230),
.B(n_228),
.Y(n_264)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_264),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_265),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_253),
.A2(n_226),
.B1(n_242),
.B2(n_235),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_272),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_276),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_241),
.C(n_226),
.Y(n_272)
);

A2O1A1Ixp33_ASAP7_75t_SL g273 ( 
.A1(n_259),
.A2(n_231),
.B(n_186),
.C(n_237),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_273),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_275),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_258),
.A2(n_231),
.B1(n_168),
.B2(n_190),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_245),
.B(n_7),
.C(n_13),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_255),
.C(n_257),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_251),
.A2(n_7),
.B(n_13),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_261),
.Y(n_287)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_254),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_6),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_281),
.B(n_287),
.Y(n_298)
);

BUFx24_ASAP7_75t_SL g282 ( 
.A(n_271),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_290),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_270),
.A2(n_262),
.B(n_256),
.Y(n_285)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_285),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_268),
.A2(n_272),
.B1(n_277),
.B2(n_244),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_286),
.B(n_5),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_260),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_245),
.C(n_248),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_293),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_269),
.C(n_266),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_300),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_284),
.A2(n_273),
.B(n_266),
.Y(n_299)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_299),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_276),
.C(n_273),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_288),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_301),
.A2(n_303),
.B1(n_290),
.B2(n_289),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_283),
.A2(n_6),
.B(n_11),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_304),
.C(n_287),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_6),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_296),
.B(n_292),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_308),
.C(n_312),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_307),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_5),
.C(n_11),
.Y(n_308)
);

OAI322xp33_ASAP7_75t_L g311 ( 
.A1(n_304),
.A2(n_5),
.A3(n_11),
.B1(n_10),
.B2(n_8),
.C1(n_15),
.C2(n_4),
.Y(n_311)
);

OA21x2_ASAP7_75t_L g316 ( 
.A1(n_311),
.A2(n_303),
.B(n_10),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_297),
.A2(n_8),
.B(n_10),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_294),
.C(n_301),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_316),
.Y(n_318)
);

A2O1A1Ixp33_ASAP7_75t_SL g317 ( 
.A1(n_309),
.A2(n_0),
.B(n_2),
.C(n_3),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_317),
.A2(n_311),
.B1(n_2),
.B2(n_4),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_319),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_314),
.A2(n_0),
.B(n_4),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_318),
.C(n_313),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_322),
.A2(n_317),
.B(n_320),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_4),
.Y(n_324)
);


endmodule