module fake_jpeg_6761_n_318 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_37),
.Y(n_50)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_8),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_0),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_21),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_16),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_44),
.B(n_55),
.Y(n_66)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_21),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_30),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_56),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_25),
.B(n_32),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_57),
.B(n_19),
.C(n_32),
.Y(n_72)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_53),
.Y(n_86)
);

OR2x4_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_27),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_34),
.A2(n_21),
.B1(n_17),
.B2(n_22),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_58),
.A2(n_17),
.B1(n_33),
.B2(n_23),
.Y(n_92)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_34),
.A2(n_31),
.B1(n_17),
.B2(n_32),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_17),
.B1(n_57),
.B2(n_22),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_30),
.Y(n_62)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_63),
.A2(n_92),
.B1(n_73),
.B2(n_84),
.Y(n_95)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_64),
.B(n_70),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_31),
.B1(n_16),
.B2(n_24),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_65),
.A2(n_83),
.B1(n_88),
.B2(n_23),
.Y(n_94)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_71),
.B(n_80),
.Y(n_117)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

AND2x4_ASAP7_75t_SL g73 ( 
.A(n_56),
.B(n_42),
.Y(n_73)
);

MAJx2_ASAP7_75t_L g115 ( 
.A(n_73),
.B(n_27),
.C(n_26),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_42),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_90),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_55),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_77),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_25),
.B(n_24),
.C(n_19),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_79),
.B(n_84),
.Y(n_114)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_54),
.A2(n_31),
.B1(n_17),
.B2(n_25),
.Y(n_81)
);

OAI22x1_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_27),
.B1(n_33),
.B2(n_23),
.Y(n_103)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_87),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_54),
.A2(n_24),
.B1(n_19),
.B2(n_38),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_56),
.B(n_28),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_85),
.Y(n_109)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_47),
.A2(n_39),
.B1(n_38),
.B2(n_18),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_42),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_91),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_94),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_95),
.A2(n_113),
.B1(n_68),
.B2(n_74),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_80),
.A2(n_38),
.B1(n_39),
.B2(n_46),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_97),
.A2(n_104),
.B1(n_112),
.B2(n_68),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_90),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_99),
.Y(n_138)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_92),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_101),
.B(n_111),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_73),
.A2(n_46),
.B1(n_53),
.B2(n_27),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_102),
.A2(n_103),
.B1(n_106),
.B2(n_119),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_72),
.A2(n_39),
.B1(n_46),
.B2(n_29),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_73),
.A2(n_46),
.B1(n_53),
.B2(n_27),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_76),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_53),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_46),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_64),
.A2(n_48),
.B1(n_61),
.B2(n_42),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_67),
.A2(n_61),
.B1(n_48),
.B2(n_29),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_115),
.A2(n_75),
.B(n_86),
.Y(n_127)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_118),
.B(n_28),
.Y(n_148)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_70),
.B1(n_69),
.B2(n_77),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_121),
.A2(n_122),
.B1(n_128),
.B2(n_136),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_95),
.A2(n_69),
.B1(n_78),
.B2(n_87),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_132),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_142),
.B1(n_145),
.B2(n_146),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_100),
.B(n_78),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_125),
.B(n_147),
.Y(n_156)
);

NOR2x1_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_114),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_126),
.A2(n_140),
.B(n_0),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_26),
.Y(n_172)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_130),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_120),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_133),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_75),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_74),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_144),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_135),
.B(n_0),
.C(n_1),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_93),
.A2(n_61),
.B1(n_29),
.B2(n_23),
.Y(n_136)
);

AND2x4_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_27),
.Y(n_140)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_137),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_104),
.A2(n_29),
.B1(n_33),
.B2(n_26),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_45),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_93),
.A2(n_71),
.B1(n_33),
.B2(n_45),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_111),
.A2(n_71),
.B1(n_45),
.B2(n_20),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_100),
.B(n_28),
.Y(n_147)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_94),
.A2(n_26),
.B1(n_20),
.B2(n_28),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_149),
.A2(n_119),
.B1(n_99),
.B2(n_26),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_98),
.B(n_45),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_112),
.Y(n_166)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_151),
.B(n_157),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_139),
.A2(n_109),
.B1(n_114),
.B2(n_105),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_153),
.B(n_159),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_138),
.B(n_118),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_113),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_171),
.C(n_176),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_150),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_161),
.B(n_165),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_125),
.B(n_109),
.Y(n_162)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_162),
.Y(n_207)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_166),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_145),
.Y(n_165)
);

AO21x1_ASAP7_75t_L g201 ( 
.A1(n_167),
.A2(n_139),
.B(n_133),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_128),
.Y(n_168)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_168),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_107),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_169),
.A2(n_179),
.B(n_140),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_107),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_180),
.Y(n_189)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_20),
.Y(n_175)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_177),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_7),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_184),
.C(n_129),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_146),
.Y(n_180)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_126),
.Y(n_181)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_182),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_124),
.Y(n_183)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_183),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_127),
.B(n_0),
.C(n_1),
.Y(n_184)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_154),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_196),
.Y(n_226)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_131),
.Y(n_197)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_203),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_199),
.A2(n_201),
.B1(n_212),
.B2(n_141),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_159),
.B(n_121),
.Y(n_200)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_166),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_206),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_151),
.B(n_155),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_209),
.Y(n_235)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_173),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_155),
.B(n_177),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_210),
.Y(n_232)
);

AOI222xp33_ASAP7_75t_SL g211 ( 
.A1(n_181),
.A2(n_153),
.B1(n_143),
.B2(n_173),
.C1(n_160),
.C2(n_182),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_179),
.Y(n_220)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_152),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_214),
.A2(n_215),
.B1(n_219),
.B2(n_221),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_209),
.A2(n_212),
.B1(n_211),
.B2(n_213),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_192),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_216),
.B(n_223),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_171),
.C(n_176),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_218),
.C(n_224),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_172),
.C(n_122),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_190),
.A2(n_205),
.B1(n_191),
.B2(n_185),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_227),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_190),
.A2(n_169),
.B1(n_142),
.B2(n_149),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_197),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_208),
.C(n_187),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_178),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_191),
.A2(n_169),
.B1(n_136),
.B2(n_184),
.Y(n_229)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

AO21x2_ASAP7_75t_L g231 ( 
.A1(n_195),
.A2(n_156),
.B(n_170),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_231),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_254)
);

OA21x2_ASAP7_75t_L g233 ( 
.A1(n_210),
.A2(n_2),
.B(n_3),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_236),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_189),
.B(n_187),
.C(n_204),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_206),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_195),
.Y(n_236)
);

O2A1O1Ixp33_ASAP7_75t_L g237 ( 
.A1(n_200),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_237)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_202),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_245),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_241),
.B(n_253),
.C(n_234),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_228),
.A2(n_198),
.B(n_193),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_242),
.A2(n_250),
.B(n_235),
.Y(n_263)
);

NAND3xp33_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_196),
.C(n_194),
.Y(n_243)
);

NAND3xp33_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_237),
.C(n_222),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_201),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_188),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_249),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_247),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_188),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_228),
.A2(n_185),
.B(n_207),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_215),
.B(n_203),
.Y(n_253)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_254),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_233),
.Y(n_255)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_255),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_231),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_233),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_248),
.A2(n_235),
.B1(n_230),
.B2(n_232),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_259),
.A2(n_263),
.B1(n_269),
.B2(n_244),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_224),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_251),
.Y(n_282)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_265),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_225),
.Y(n_266)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_266),
.Y(n_279)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_240),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_270),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_256),
.A2(n_231),
.B1(n_221),
.B2(n_229),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_253),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_241),
.C(n_239),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_226),
.Y(n_272)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_272),
.Y(n_285)
);

A2O1A1Ixp33_ASAP7_75t_L g280 ( 
.A1(n_273),
.A2(n_263),
.B(n_259),
.C(n_265),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_260),
.B(n_264),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_284),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_272),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_247),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_278),
.B(n_261),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_280),
.A2(n_286),
.B(n_258),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_251),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_282),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_287),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_266),
.B(n_245),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_239),
.C(n_243),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_258),
.B(n_10),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_288),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_294),
.C(n_298),
.Y(n_305)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_292),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_275),
.B(n_261),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_295),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_283),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_280),
.B(n_10),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_286),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_7),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_4),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_297),
.A2(n_15),
.B(n_6),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_288),
.A2(n_279),
.B1(n_274),
.B2(n_287),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_300),
.A2(n_297),
.B1(n_289),
.B2(n_290),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_5),
.C(n_6),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_305),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_303),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_304),
.B(n_11),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_307),
.A2(n_309),
.B(n_311),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_9),
.Y(n_309)
);

NOR2x1_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_306),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_312),
.A2(n_313),
.B(n_12),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_308),
.A2(n_300),
.B(n_301),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_314),
.Y(n_316)
);

OAI311xp33_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_13),
.A3(n_14),
.B1(n_15),
.C1(n_312),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_13),
.Y(n_318)
);


endmodule