module fake_jpeg_17350_n_314 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_314);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_10),
.B(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_13),
.B(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_35),
.B(n_31),
.Y(n_52)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_37),
.B(n_26),
.Y(n_45)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_42),
.Y(n_61)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_30),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_64),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_0),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_47),
.A2(n_53),
.B(n_46),
.Y(n_73)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_30),
.B1(n_25),
.B2(n_24),
.Y(n_49)
);

AO22x2_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_42),
.B1(n_19),
.B2(n_32),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_52),
.B(n_27),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_26),
.B1(n_34),
.B2(n_21),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_31),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_55),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_38),
.B1(n_43),
.B2(n_40),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_33),
.B1(n_32),
.B2(n_28),
.Y(n_86)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_42),
.Y(n_71)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_33),
.Y(n_64)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_67),
.A2(n_81),
.B1(n_82),
.B2(n_61),
.Y(n_107)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_34),
.B1(n_21),
.B2(n_25),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_70),
.A2(n_73),
.B1(n_97),
.B2(n_28),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_44),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_74),
.Y(n_110)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_87),
.Y(n_103)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_51),
.A2(n_42),
.B1(n_19),
.B2(n_21),
.Y(n_82)
);

CKINVDCx12_ASAP7_75t_R g83 ( 
.A(n_44),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_84),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_47),
.A2(n_34),
.B1(n_22),
.B2(n_33),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_86),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_22),
.Y(n_87)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_88),
.Y(n_130)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_90),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_49),
.B(n_29),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_96),
.Y(n_124)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_62),
.A2(n_25),
.B1(n_24),
.B2(n_27),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_100),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_99),
.Y(n_122)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_101),
.B(n_29),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_47),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_104),
.B(n_106),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_47),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_107),
.A2(n_67),
.B1(n_100),
.B2(n_89),
.Y(n_136)
);

AOI32xp33_ASAP7_75t_L g109 ( 
.A1(n_73),
.A2(n_53),
.A3(n_56),
.B1(n_42),
.B2(n_29),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_123),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_67),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_85),
.Y(n_131)
);

AND2x6_ASAP7_75t_L g117 ( 
.A(n_67),
.B(n_12),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_117),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_50),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_118),
.A2(n_86),
.B(n_28),
.Y(n_145)
);

CKINVDCx12_ASAP7_75t_R g119 ( 
.A(n_66),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_74),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_68),
.B(n_23),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_121),
.B(n_129),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_65),
.B(n_20),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_68),
.B(n_23),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_131),
.B(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_134),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_107),
.A2(n_98),
.B1(n_96),
.B2(n_94),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_135),
.A2(n_159),
.B1(n_124),
.B2(n_118),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_136),
.A2(n_142),
.B1(n_144),
.B2(n_154),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_139),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_110),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_140),
.A2(n_78),
.B1(n_108),
.B2(n_61),
.Y(n_193)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_76),
.B1(n_88),
.B2(n_91),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_126),
.A2(n_76),
.B1(n_91),
.B2(n_69),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_145),
.A2(n_153),
.B(n_78),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_103),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_158),
.Y(n_165)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_104),
.B(n_77),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

NOR2x1_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_82),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_115),
.A2(n_61),
.B1(n_79),
.B2(n_72),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_99),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_156),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_116),
.B(n_23),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_102),
.Y(n_157)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_112),
.B(n_80),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_115),
.A2(n_61),
.B1(n_78),
.B2(n_66),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_84),
.Y(n_160)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_160),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_106),
.B(n_32),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g179 ( 
.A1(n_161),
.A2(n_103),
.B(n_129),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_162),
.A2(n_185),
.B1(n_189),
.B2(n_153),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_111),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_163),
.A2(n_108),
.B1(n_90),
.B2(n_114),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_140),
.A2(n_124),
.B1(n_109),
.B2(n_117),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_168),
.A2(n_171),
.B1(n_132),
.B2(n_160),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_133),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_173),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_118),
.B1(n_121),
.B2(n_105),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_141),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_157),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_174),
.B(n_189),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_123),
.C(n_105),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_182),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_122),
.Y(n_178)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_179),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_122),
.Y(n_180)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_180),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_113),
.C(n_102),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_150),
.C(n_132),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_183),
.B(n_161),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_147),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_190),
.B(n_152),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_127),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_131),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_142),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_192),
.B(n_184),
.Y(n_194)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_194),
.Y(n_236)
);

NOR2x1_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_153),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_170),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_196),
.A2(n_203),
.B(n_205),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_165),
.B(n_148),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_197),
.B(n_212),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_199),
.B(n_202),
.Y(n_233)
);

INVxp33_ASAP7_75t_L g201 ( 
.A(n_164),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_211),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_171),
.Y(n_225)
);

XOR2x2_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_145),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_183),
.A2(n_135),
.B1(n_144),
.B2(n_156),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_207),
.A2(n_220),
.B1(n_167),
.B2(n_174),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_148),
.Y(n_209)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_193),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_172),
.B(n_151),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_213),
.B(n_217),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_137),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_17),
.C(n_8),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_168),
.B(n_20),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_163),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_120),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_187),
.B(n_128),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_219),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_120),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_203),
.A2(n_163),
.B1(n_162),
.B2(n_167),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_222),
.A2(n_231),
.B1(n_234),
.B2(n_240),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_216),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_225),
.B(n_202),
.Y(n_245)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_227),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_228),
.A2(n_214),
.B(n_200),
.Y(n_256)
);

OAI322xp33_ASAP7_75t_L g230 ( 
.A1(n_205),
.A2(n_191),
.A3(n_188),
.B1(n_166),
.B2(n_169),
.C1(n_176),
.C2(n_186),
.Y(n_230)
);

NAND3xp33_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_199),
.C(n_207),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_203),
.A2(n_188),
.B1(n_166),
.B2(n_169),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_186),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_241),
.C(n_8),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_196),
.A2(n_181),
.B1(n_176),
.B2(n_175),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_210),
.A2(n_181),
.B1(n_175),
.B2(n_114),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_235),
.A2(n_238),
.B1(n_198),
.B2(n_224),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_114),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_194),
.Y(n_247)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_215),
.Y(n_239)
);

INVx13_ASAP7_75t_L g249 ( 
.A(n_239),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_211),
.A2(n_20),
.B1(n_1),
.B2(n_3),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_222),
.A2(n_195),
.B1(n_220),
.B2(n_204),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_244),
.A2(n_246),
.B1(n_225),
.B2(n_227),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_233),
.Y(n_273)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_259),
.C(n_260),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_206),
.Y(n_250)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_236),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_239),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_229),
.B(n_208),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_254),
.B(n_255),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_226),
.B(n_201),
.Y(n_255)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_0),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_257),
.A2(n_258),
.B(n_1),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_228),
.A2(n_10),
.B(n_15),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_17),
.C(n_3),
.Y(n_260)
);

MAJx2_ASAP7_75t_L g261 ( 
.A(n_221),
.B(n_17),
.C(n_11),
.Y(n_261)
);

BUFx24_ASAP7_75t_SL g271 ( 
.A(n_261),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_242),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_268),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_265),
.B(n_269),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_253),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_258),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_257),
.A2(n_234),
.B1(n_221),
.B2(n_223),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_272),
.A2(n_257),
.B1(n_261),
.B2(n_244),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_274),
.C(n_248),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_233),
.C(n_241),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_280),
.C(n_274),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_246),
.C(n_245),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_281),
.B(n_288),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_282),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_262),
.B(n_250),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_286),
.Y(n_293)
);

XOR2x2_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_243),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_284),
.A2(n_287),
.B(n_273),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_249),
.Y(n_285)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_285),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_249),
.Y(n_286)
);

OA21x2_ASAP7_75t_SL g287 ( 
.A1(n_276),
.A2(n_243),
.B(n_259),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_240),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_287),
.A2(n_275),
.B(n_263),
.Y(n_291)
);

AOI21xp33_ASAP7_75t_L g301 ( 
.A1(n_291),
.A2(n_271),
.B(n_260),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_277),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_294),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_266),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_284),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_8),
.Y(n_304)
);

MAJx2_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_295),
.C(n_298),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_290),
.C(n_293),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_289),
.A2(n_280),
.B(n_278),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_299),
.A2(n_302),
.B(n_13),
.Y(n_308)
);

AOI322xp5_ASAP7_75t_L g307 ( 
.A1(n_300),
.A2(n_301),
.A3(n_305),
.B1(n_15),
.B2(n_14),
.C1(n_13),
.C2(n_6),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_304),
.B(n_12),
.Y(n_306)
);

NAND4xp25_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_12),
.C(n_15),
.D(n_14),
.Y(n_305)
);

AOI322xp5_ASAP7_75t_L g310 ( 
.A1(n_306),
.A2(n_307),
.A3(n_309),
.B1(n_1),
.B2(n_4),
.C1(n_5),
.C2(n_7),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_308),
.A2(n_300),
.B(n_302),
.Y(n_311)
);

AOI322xp5_ASAP7_75t_L g309 ( 
.A1(n_303),
.A2(n_17),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_1),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_310),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_312),
.A2(n_311),
.B1(n_7),
.B2(n_4),
.Y(n_313)
);

AO21x2_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_4),
.B(n_17),
.Y(n_314)
);


endmodule