module fake_jpeg_17126_n_114 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_114);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_114;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_36),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_0),
.B(n_11),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_25),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_15),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_0),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_1),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_2),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_2),
.Y(n_71)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_61),
.A2(n_47),
.B1(n_45),
.B2(n_56),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_67),
.A2(n_76),
.B1(n_58),
.B2(n_57),
.Y(n_81)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_77),
.Y(n_82)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_47),
.B1(n_53),
.B2(n_55),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_60),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_79),
.Y(n_89)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_76),
.B1(n_73),
.B2(n_3),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_70),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_84),
.Y(n_90)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_87),
.B(n_88),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_43),
.Y(n_88)
);

INVx6_ASAP7_75t_SL g91 ( 
.A(n_85),
.Y(n_91)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_89),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_93),
.A2(n_86),
.B1(n_82),
.B2(n_67),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_97),
.B1(n_94),
.B2(n_90),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_92),
.A2(n_68),
.B1(n_75),
.B2(n_4),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_99),
.A2(n_101),
.B1(n_98),
.B2(n_82),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_93),
.B(n_54),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_100),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_103),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_105),
.A2(n_103),
.B1(n_51),
.B2(n_49),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_41),
.C(n_46),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_16),
.Y(n_108)
);

AOI21x1_ASAP7_75t_SL g109 ( 
.A1(n_108),
.A2(n_19),
.B(n_37),
.Y(n_109)
);

AOI322xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_14),
.A3(n_34),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_110),
.A2(n_22),
.B(n_33),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_20),
.B(n_31),
.Y(n_112)
);

AOI322xp5_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_13),
.A3(n_30),
.B1(n_9),
.B2(n_10),
.C1(n_12),
.C2(n_38),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_23),
.Y(n_114)
);


endmodule