module fake_jpeg_28903_n_251 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_251);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_220;
wire n_137;
wire n_31;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_45;
wire n_61;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_218;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx5_ASAP7_75t_SL g98 ( 
.A(n_38),
.Y(n_98)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_50),
.Y(n_62)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_0),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_35),
.Y(n_80)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_18),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_18),
.B(n_15),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_57),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_15),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_60),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_66),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_48),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_45),
.A2(n_59),
.B1(n_58),
.B2(n_56),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_73),
.A2(n_77),
.B1(n_97),
.B2(n_37),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_44),
.A2(n_31),
.B(n_33),
.C(n_32),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_76),
.A2(n_30),
.B(n_26),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_42),
.A2(n_35),
.B1(n_27),
.B2(n_34),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_25),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_81),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_0),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_43),
.B(n_16),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_38),
.B(n_25),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_83),
.B(n_84),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_39),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_85),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_41),
.B(n_21),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_86),
.B(n_90),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_54),
.A2(n_19),
.B1(n_34),
.B2(n_37),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_89),
.A2(n_37),
.B1(n_26),
.B2(n_2),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_28),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_47),
.B(n_28),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_93),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_46),
.B(n_24),
.Y(n_93)
);

CKINVDCx12_ASAP7_75t_R g94 ( 
.A(n_43),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_53),
.B(n_24),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_96),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_45),
.A2(n_19),
.B1(n_21),
.B2(n_30),
.Y(n_97)
);

CKINVDCx12_ASAP7_75t_R g100 ( 
.A(n_43),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_32),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_116),
.Y(n_133)
);

OR2x2_ASAP7_75t_SL g147 ( 
.A(n_105),
.B(n_99),
.Y(n_147)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_77),
.B1(n_65),
.B2(n_74),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_112),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_82),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_113),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_62),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_87),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_93),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_80),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_118),
.A2(n_121),
.B(n_126),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_1),
.C(n_2),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_5),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_127),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_76),
.A2(n_5),
.B(n_6),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_7),
.Y(n_127)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_104),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_131),
.B(n_136),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_120),
.B(n_72),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_103),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_109),
.B(n_75),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_138),
.A2(n_88),
.B1(n_74),
.B2(n_69),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_141),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_102),
.B(n_122),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_99),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_142),
.B(n_150),
.Y(n_181)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

NOR2xp67_ASAP7_75t_SL g168 ( 
.A(n_147),
.B(n_155),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_125),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_87),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_153),
.Y(n_182)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_98),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_116),
.A2(n_120),
.B1(n_127),
.B2(n_118),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_154),
.A2(n_157),
.B1(n_111),
.B2(n_117),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_105),
.A2(n_88),
.B1(n_65),
.B2(n_71),
.Y(n_157)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_156),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_161),
.Y(n_194)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_158),
.A2(n_126),
.B(n_112),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_165),
.A2(n_166),
.B(n_115),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_123),
.B(n_121),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_167),
.A2(n_172),
.B1(n_178),
.B2(n_61),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_168),
.A2(n_135),
.B(n_145),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_174),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_133),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_171),
.B(n_177),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_149),
.B(n_128),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_173),
.B(n_149),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_103),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_130),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_176),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_132),
.B(n_72),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_154),
.A2(n_71),
.B1(n_69),
.B2(n_91),
.Y(n_178)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_180),
.Y(n_186)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_135),
.Y(n_180)
);

NOR4xp25_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_170),
.C(n_136),
.D(n_131),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_188),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_172),
.Y(n_205)
);

AOI221xp5_ASAP7_75t_L g188 ( 
.A1(n_166),
.A2(n_168),
.B1(n_171),
.B2(n_165),
.C(n_155),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_174),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_199),
.C(n_178),
.Y(n_203)
);

AOI221xp5_ASAP7_75t_L g190 ( 
.A1(n_175),
.A2(n_133),
.B1(n_149),
.B2(n_158),
.C(n_143),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_191),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_163),
.B(n_133),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_193),
.A2(n_195),
.B(n_176),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_150),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_200),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_167),
.B(n_128),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_169),
.B(n_115),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_206),
.Y(n_218)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_197),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_205),
.Y(n_216)
);

MAJx2_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_195),
.C(n_199),
.Y(n_219)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_197),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_177),
.C(n_164),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_211),
.C(n_185),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_180),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_210),
.Y(n_224)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_160),
.C(n_159),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_148),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_213),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_208),
.Y(n_215)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_215),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_201),
.A2(n_193),
.B1(n_192),
.B2(n_159),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_217),
.A2(n_194),
.B1(n_144),
.B2(n_162),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_221),
.C(n_196),
.Y(n_231)
);

NAND3xp33_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_196),
.C(n_194),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_223),
.Y(n_225)
);

BUFx24_ASAP7_75t_SL g223 ( 
.A(n_214),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_218),
.A2(n_204),
.B(n_212),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_226),
.A2(n_229),
.B(n_148),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_224),
.A2(n_205),
.B1(n_212),
.B2(n_160),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_227),
.A2(n_220),
.B1(n_219),
.B2(n_162),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_222),
.A2(n_211),
.B(n_203),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_207),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_231),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_232),
.A2(n_152),
.B1(n_140),
.B2(n_137),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_233),
.B(n_234),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_231),
.B(n_144),
.C(n_137),
.Y(n_234)
);

AOI322xp5_ASAP7_75t_L g241 ( 
.A1(n_235),
.A2(n_179),
.A3(n_161),
.B1(n_113),
.B2(n_70),
.C1(n_85),
.C2(n_61),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_230),
.Y(n_240)
);

A2O1A1Ixp33_ASAP7_75t_L g237 ( 
.A1(n_225),
.A2(n_140),
.B(n_161),
.C(n_179),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_237),
.A2(n_226),
.B(n_228),
.Y(n_239)
);

NOR2x1_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_237),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_240),
.A2(n_241),
.B(n_243),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_113),
.C(n_124),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_246),
.Y(n_247)
);

NOR2x1_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_234),
.Y(n_246)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_236),
.C(n_113),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_98),
.Y(n_249)
);

AOI322xp5_ASAP7_75t_L g250 ( 
.A1(n_249),
.A2(n_247),
.A3(n_63),
.B1(n_12),
.B2(n_14),
.C1(n_10),
.C2(n_9),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_12),
.Y(n_251)
);


endmodule