module fake_jpeg_22947_n_301 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_300;
wire n_211;
wire n_299;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_2),
.B(n_3),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_36),
.B(n_44),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_28),
.B1(n_31),
.B2(n_33),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_35),
.B(n_10),
.Y(n_44)
);

AND2x2_ASAP7_75t_SL g45 ( 
.A(n_38),
.B(n_19),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_55),
.Y(n_85)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_40),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_30),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_58),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_36),
.A2(n_24),
.B1(n_27),
.B2(n_33),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_68),
.B1(n_69),
.B2(n_26),
.Y(n_75)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_24),
.B1(n_31),
.B2(n_27),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_60),
.A2(n_32),
.B1(n_39),
.B2(n_43),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_30),
.Y(n_64)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_43),
.B(n_35),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_65),
.B(n_30),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_38),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_66),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_37),
.A2(n_31),
.B1(n_26),
.B2(n_28),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_37),
.A2(n_26),
.B1(n_33),
.B2(n_27),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_73),
.B(n_93),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_75),
.A2(n_77),
.B1(n_90),
.B2(n_103),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_76),
.B(n_45),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_32),
.B1(n_19),
.B2(n_35),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_79),
.Y(n_110)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_40),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_81),
.B(n_82),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_42),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_86),
.A2(n_39),
.B1(n_61),
.B2(n_68),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_41),
.Y(n_89)
);

NAND2x1_ASAP7_75t_SL g112 ( 
.A(n_89),
.B(n_92),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_57),
.A2(n_41),
.B(n_32),
.C(n_20),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_42),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_85),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_41),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_59),
.B(n_65),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_96),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_48),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_66),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_99),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_101),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_17),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_102),
.B(n_63),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_60),
.A2(n_17),
.B1(n_29),
.B2(n_20),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_61),
.B(n_63),
.Y(n_104)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_45),
.A2(n_37),
.B1(n_42),
.B2(n_22),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_105),
.A2(n_42),
.B1(n_51),
.B2(n_48),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_63),
.A2(n_37),
.B1(n_39),
.B2(n_43),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_106),
.A2(n_69),
.B(n_56),
.Y(n_120)
);

NAND3xp33_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_45),
.C(n_4),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_109),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_132),
.B1(n_133),
.B2(n_96),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_116),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_95),
.B(n_58),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_117),
.A2(n_122),
.B(n_124),
.Y(n_152)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_121),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_120),
.A2(n_70),
.B(n_99),
.Y(n_148)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_81),
.A2(n_29),
.B(n_18),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_131),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_74),
.A2(n_61),
.B1(n_37),
.B2(n_39),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_82),
.B(n_50),
.Y(n_129)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_84),
.B(n_50),
.Y(n_130)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_76),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_74),
.A2(n_101),
.B1(n_90),
.B2(n_100),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_85),
.B(n_53),
.Y(n_134)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_135),
.A2(n_143),
.B1(n_154),
.B2(n_159),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_126),
.A2(n_85),
.B1(n_105),
.B2(n_88),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_136),
.A2(n_144),
.B1(n_122),
.B2(n_128),
.Y(n_181)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_140),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_110),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_139),
.Y(n_185)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_132),
.A2(n_89),
.B1(n_70),
.B2(n_92),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_126),
.A2(n_88),
.B1(n_97),
.B2(n_89),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_117),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_150),
.Y(n_169)
);

MAJx2_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_92),
.C(n_80),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_153),
.C(n_157),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_148),
.A2(n_112),
.B(n_115),
.Y(n_179)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_116),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_155),
.Y(n_184)
);

A2O1A1O1Ixp25_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_102),
.B(n_95),
.C(n_83),
.D(n_80),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_131),
.B1(n_127),
.B2(n_129),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_110),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_158),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_83),
.C(n_102),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_72),
.B1(n_87),
.B2(n_79),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_165),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_120),
.A2(n_72),
.B1(n_87),
.B2(n_78),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_164),
.A2(n_135),
.B1(n_160),
.B2(n_165),
.Y(n_188)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_162),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_166),
.B(n_168),
.Y(n_214)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

AO21x1_ASAP7_75t_L g170 ( 
.A1(n_152),
.A2(n_109),
.B(n_108),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_170),
.A2(n_182),
.B(n_190),
.Y(n_209)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_163),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_172),
.Y(n_197)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_123),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_176),
.Y(n_196)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_175),
.B(n_178),
.Y(n_213)
);

AOI221xp5_ASAP7_75t_L g176 ( 
.A1(n_136),
.A2(n_123),
.B1(n_112),
.B2(n_122),
.C(n_121),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_148),
.Y(n_177)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_179),
.A2(n_183),
.B(n_107),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_157),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_141),
.C(n_53),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_181),
.A2(n_189),
.B1(n_194),
.B2(n_22),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_137),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_142),
.A2(n_147),
.B(n_149),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_188),
.A2(n_195),
.B1(n_146),
.B2(n_156),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_160),
.A2(n_122),
.B1(n_111),
.B2(n_118),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_145),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_153),
.Y(n_191)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_191),
.Y(n_200)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_150),
.A2(n_72),
.B1(n_94),
.B2(n_111),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_149),
.A2(n_115),
.B1(n_107),
.B2(n_42),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_138),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_201),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_138),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_184),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_205),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_203),
.A2(n_168),
.B1(n_187),
.B2(n_175),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_181),
.B(n_158),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_204),
.B(n_211),
.Y(n_221)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

AO21x1_ASAP7_75t_L g224 ( 
.A1(n_206),
.A2(n_193),
.B(n_178),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_186),
.C(n_195),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_208),
.Y(n_232)
);

A2O1A1O1Ixp25_ASAP7_75t_L g211 ( 
.A1(n_179),
.A2(n_18),
.B(n_51),
.C(n_25),
.D(n_22),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_167),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_215),
.Y(n_233)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_172),
.A2(n_51),
.B1(n_22),
.B2(n_18),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_216),
.A2(n_21),
.B1(n_4),
.B2(n_5),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_174),
.B(n_25),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_169),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_185),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_166),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_219),
.A2(n_21),
.B1(n_4),
.B2(n_5),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_220),
.A2(n_205),
.B1(n_197),
.B2(n_213),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_196),
.B(n_174),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_229),
.Y(n_242)
);

OAI322xp33_ASAP7_75t_L g223 ( 
.A1(n_206),
.A2(n_183),
.A3(n_170),
.B1(n_189),
.B2(n_185),
.C1(n_171),
.C2(n_190),
.Y(n_223)
);

NOR2xp67_ASAP7_75t_SL g246 ( 
.A(n_223),
.B(n_211),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_224),
.A2(n_239),
.B(n_7),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_234),
.C(n_237),
.Y(n_243)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_227),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_214),
.Y(n_228)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_228),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_230),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_51),
.C(n_25),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_198),
.A2(n_18),
.B1(n_51),
.B2(n_21),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_235),
.A2(n_236),
.B1(n_238),
.B2(n_203),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_196),
.B(n_21),
.C(n_2),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_213),
.A2(n_11),
.B(n_5),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_229),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_231),
.A2(n_197),
.B1(n_209),
.B2(n_204),
.Y(n_244)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_244),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_226),
.A2(n_209),
.B1(n_224),
.B2(n_200),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_245),
.A2(n_248),
.B1(n_252),
.B2(n_225),
.Y(n_259)
);

OAI31xp33_ASAP7_75t_L g268 ( 
.A1(n_246),
.A2(n_250),
.A3(n_255),
.B(n_248),
.Y(n_268)
);

AOI21x1_ASAP7_75t_L g247 ( 
.A1(n_239),
.A2(n_201),
.B(n_216),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_247),
.A2(n_250),
.B(n_254),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_234),
.A2(n_232),
.B1(n_237),
.B2(n_221),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_221),
.A2(n_199),
.B(n_217),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_233),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_21),
.C(n_9),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_236),
.Y(n_256)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_256),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_225),
.Y(n_258)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_258),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_266),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_8),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_262),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_9),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_247),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_263),
.A2(n_268),
.B1(n_249),
.B2(n_12),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_253),
.B(n_10),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_264),
.B(n_11),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

AOI21x1_ASAP7_75t_L g271 ( 
.A1(n_265),
.A2(n_240),
.B(n_254),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_271),
.A2(n_265),
.B(n_259),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_252),
.Y(n_275)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_275),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_245),
.Y(n_276)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_276),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_279),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_260),
.A2(n_243),
.B1(n_13),
.B2(n_14),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_263),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_262),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_281),
.B(n_285),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_243),
.C(n_261),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_272),
.C(n_274),
.Y(n_290)
);

AOI21x1_ASAP7_75t_L g288 ( 
.A1(n_286),
.A2(n_287),
.B(n_271),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_273),
.A2(n_13),
.B(n_14),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_288),
.A2(n_291),
.B(n_293),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_292),
.C(n_16),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_280),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_282),
.A2(n_285),
.B1(n_276),
.B2(n_277),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_280),
.B(n_278),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_294),
.A2(n_297),
.B1(n_15),
.B2(n_16),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_291),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_296),
.Y(n_299)
);

OAI21x1_ASAP7_75t_L g297 ( 
.A1(n_289),
.A2(n_13),
.B(n_15),
.Y(n_297)
);

MAJx2_ASAP7_75t_L g300 ( 
.A(n_298),
.B(n_295),
.C(n_15),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_299),
.Y(n_301)
);


endmodule