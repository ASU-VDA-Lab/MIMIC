module real_aes_7811_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_357;
wire n_287;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_519;
wire n_92;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_478;
wire n_356;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_527;
wire n_505;
wire n_502;
wire n_434;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_500;
wire n_307;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_0), .Y(n_111) );
AOI22xp33_ASAP7_75t_L g138 ( .A1(n_1), .A2(n_3), .B1(n_139), .B2(n_144), .Y(n_138) );
INVx1_ASAP7_75t_L g317 ( .A(n_2), .Y(n_317) );
AOI21xp33_ASAP7_75t_L g224 ( .A1(n_4), .A2(n_225), .B(n_226), .Y(n_224) );
INVx1_ASAP7_75t_L g182 ( .A(n_5), .Y(n_182) );
AND2x6_ASAP7_75t_L g199 ( .A(n_5), .B(n_180), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_5), .B(n_527), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_6), .A2(n_293), .B(n_294), .Y(n_292) );
INVx1_ASAP7_75t_L g233 ( .A(n_7), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_8), .B(n_285), .Y(n_284) );
AO22x2_ASAP7_75t_L g88 ( .A1(n_9), .A2(n_25), .B1(n_89), .B2(n_90), .Y(n_88) );
INVx1_ASAP7_75t_L g196 ( .A(n_10), .Y(n_196) );
INVx1_ASAP7_75t_L g299 ( .A(n_11), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_12), .B(n_244), .Y(n_271) );
AO22x2_ASAP7_75t_L g92 ( .A1(n_13), .A2(n_26), .B1(n_89), .B2(n_93), .Y(n_92) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_14), .B(n_225), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_15), .B(n_221), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_16), .A2(n_505), .B1(n_506), .B2(n_507), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_16), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g164 ( .A1(n_17), .A2(n_34), .B1(n_165), .B2(n_169), .Y(n_164) );
A2O1A1Ixp33_ASAP7_75t_L g296 ( .A1(n_18), .A2(n_297), .B(n_298), .C(n_300), .Y(n_296) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_19), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_20), .B(n_231), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g158 ( .A1(n_21), .A2(n_33), .B1(n_159), .B2(n_162), .Y(n_158) );
AOI22xp33_ASAP7_75t_L g149 ( .A1(n_22), .A2(n_27), .B1(n_150), .B2(n_154), .Y(n_149) );
INVx1_ASAP7_75t_L g209 ( .A(n_23), .Y(n_209) );
INVx2_ASAP7_75t_L g203 ( .A(n_24), .Y(n_203) );
OAI221xp5_ASAP7_75t_L g517 ( .A1(n_26), .A2(n_41), .B1(n_49), .B2(n_518), .C(n_519), .Y(n_517) );
INVxp67_ASAP7_75t_L g520 ( .A(n_26), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_28), .A2(n_199), .B(n_210), .C(n_255), .Y(n_254) );
OAI22xp5_ASAP7_75t_SL g510 ( .A1(n_29), .A2(n_46), .B1(n_511), .B2(n_512), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_29), .Y(n_511) );
INVx1_ASAP7_75t_L g207 ( .A(n_30), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_31), .B(n_231), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_32), .B(n_122), .Y(n_121) );
CKINVDCx16_ASAP7_75t_R g213 ( .A(n_35), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_36), .B(n_225), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_37), .Y(n_99) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_38), .A2(n_201), .B1(n_204), .B2(n_210), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_38), .A2(n_502), .B1(n_516), .B2(n_522), .Y(n_501) );
CKINVDCx16_ASAP7_75t_R g535 ( .A(n_38), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g264 ( .A(n_39), .Y(n_264) );
CKINVDCx16_ASAP7_75t_R g314 ( .A(n_40), .Y(n_314) );
AO22x2_ASAP7_75t_L g98 ( .A1(n_41), .A2(n_59), .B1(n_89), .B2(n_93), .Y(n_98) );
INVxp67_ASAP7_75t_L g521 ( .A(n_41), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_42), .A2(n_230), .B(n_232), .C(n_235), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g274 ( .A(n_43), .Y(n_274) );
INVx1_ASAP7_75t_L g227 ( .A(n_44), .Y(n_227) );
INVx1_ASAP7_75t_L g180 ( .A(n_45), .Y(n_180) );
INVx1_ASAP7_75t_L g512 ( .A(n_46), .Y(n_512) );
INVx1_ASAP7_75t_L g195 ( .A(n_47), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_48), .Y(n_518) );
AO22x2_ASAP7_75t_L g96 ( .A1(n_49), .A2(n_64), .B1(n_89), .B2(n_90), .Y(n_96) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_50), .Y(n_126) );
A2O1A1Ixp33_ASAP7_75t_SL g243 ( .A1(n_51), .A2(n_235), .B(n_244), .C(n_245), .Y(n_243) );
INVxp67_ASAP7_75t_L g246 ( .A(n_52), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_53), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_54), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g218 ( .A(n_55), .Y(n_218) );
INVx1_ASAP7_75t_L g267 ( .A(n_56), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g268 ( .A1(n_57), .A2(n_199), .B(n_210), .C(n_269), .Y(n_268) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_57), .A2(n_509), .B1(n_510), .B2(n_513), .Y(n_508) );
INVx1_ASAP7_75t_L g513 ( .A(n_57), .Y(n_513) );
INVx1_ASAP7_75t_L g506 ( .A(n_58), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_60), .B(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g193 ( .A(n_61), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_62), .B(n_244), .Y(n_258) );
A2O1A1Ixp33_ASAP7_75t_L g315 ( .A1(n_63), .A2(n_199), .B(n_210), .C(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_65), .B(n_238), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g321 ( .A(n_66), .Y(n_321) );
A2O1A1Ixp33_ASAP7_75t_L g281 ( .A1(n_67), .A2(n_199), .B(n_210), .C(n_282), .Y(n_281) );
CKINVDCx20_ASAP7_75t_R g289 ( .A(n_68), .Y(n_289) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_69), .A2(n_80), .B1(n_173), .B2(n_174), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_69), .Y(n_173) );
INVx1_ASAP7_75t_L g242 ( .A(n_70), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_71), .B(n_257), .Y(n_283) );
CKINVDCx16_ASAP7_75t_R g295 ( .A(n_72), .Y(n_295) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_73), .Y(n_83) );
INVx1_ASAP7_75t_L g89 ( .A(n_74), .Y(n_89) );
INVx1_ASAP7_75t_L g91 ( .A(n_74), .Y(n_91) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_75), .B(n_223), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_76), .A2(n_225), .B(n_241), .Y(n_240) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_175), .B1(n_183), .B2(n_495), .C(n_498), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_79), .Y(n_78) );
INVx1_ASAP7_75t_L g174 ( .A(n_80), .Y(n_174) );
OAI322xp33_ASAP7_75t_L g498 ( .A1(n_80), .A2(n_213), .A3(n_499), .B1(n_500), .B2(n_501), .C1(n_528), .C2(n_532), .Y(n_498) );
AND2x2_ASAP7_75t_L g80 ( .A(n_81), .B(n_136), .Y(n_80) );
INVxp67_ASAP7_75t_L g500 ( .A(n_81), .Y(n_500) );
NOR3xp33_ASAP7_75t_L g81 ( .A(n_82), .B(n_104), .C(n_125), .Y(n_81) );
OAI22xp5_ASAP7_75t_L g82 ( .A1(n_83), .A2(n_84), .B1(n_99), .B2(n_100), .Y(n_82) );
BUFx6f_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
OR2x2_ASAP7_75t_L g85 ( .A(n_86), .B(n_94), .Y(n_85) );
INVx2_ASAP7_75t_L g153 ( .A(n_86), .Y(n_153) );
OR2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_92), .Y(n_86) );
AND2x2_ASAP7_75t_L g103 ( .A(n_87), .B(n_92), .Y(n_103) );
AND2x2_ASAP7_75t_L g143 ( .A(n_87), .B(n_118), .Y(n_143) );
INVx2_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
AND2x2_ASAP7_75t_L g108 ( .A(n_88), .B(n_92), .Y(n_108) );
AND2x2_ASAP7_75t_L g119 ( .A(n_88), .B(n_98), .Y(n_119) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g93 ( .A(n_91), .Y(n_93) );
INVx2_ASAP7_75t_L g118 ( .A(n_92), .Y(n_118) );
INVx1_ASAP7_75t_L g172 ( .A(n_92), .Y(n_172) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
NAND2x1p5_ASAP7_75t_L g102 ( .A(n_95), .B(n_103), .Y(n_102) );
AND2x4_ASAP7_75t_L g163 ( .A(n_95), .B(n_143), .Y(n_163) );
AND2x2_ASAP7_75t_L g95 ( .A(n_96), .B(n_97), .Y(n_95) );
INVx1_ASAP7_75t_L g110 ( .A(n_96), .Y(n_110) );
INVx1_ASAP7_75t_L g117 ( .A(n_96), .Y(n_117) );
INVx1_ASAP7_75t_L g135 ( .A(n_96), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_96), .B(n_98), .Y(n_148) );
AND2x2_ASAP7_75t_L g109 ( .A(n_97), .B(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND2x2_ASAP7_75t_L g142 ( .A(n_98), .B(n_135), .Y(n_142) );
INVx1_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x4_ASAP7_75t_L g156 ( .A(n_103), .B(n_109), .Y(n_156) );
AND2x2_ASAP7_75t_L g168 ( .A(n_103), .B(n_142), .Y(n_168) );
OAI221xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_111), .B1(n_112), .B2(n_120), .C(n_121), .Y(n_104) );
INVx2_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x6_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
INVx1_ASAP7_75t_L g132 ( .A(n_108), .Y(n_132) );
AND2x6_ASAP7_75t_L g152 ( .A(n_109), .B(n_153), .Y(n_152) );
AND2x2_ASAP7_75t_L g161 ( .A(n_109), .B(n_143), .Y(n_161) );
INVx2_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x4_ASAP7_75t_L g115 ( .A(n_116), .B(n_119), .Y(n_115) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
INVx1_ASAP7_75t_L g124 ( .A(n_117), .Y(n_124) );
INVx1_ASAP7_75t_L g128 ( .A(n_118), .Y(n_128) );
AND2x4_ASAP7_75t_L g123 ( .A(n_119), .B(n_124), .Y(n_123) );
NAND2x1p5_ASAP7_75t_L g127 ( .A(n_119), .B(n_128), .Y(n_127) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI22xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_127), .B1(n_129), .B2(n_130), .Y(n_125) );
BUFx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OR2x6_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVxp67_ASAP7_75t_L g499 ( .A(n_136), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_137), .B(n_157), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_149), .Y(n_137) );
BUFx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
AND2x4_ASAP7_75t_L g146 ( .A(n_143), .B(n_147), .Y(n_146) );
BUFx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
BUFx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
OR2x6_ASAP7_75t_L g171 ( .A(n_148), .B(n_172), .Y(n_171) );
INVx4_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx11_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx6_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_158), .B(n_164), .Y(n_157) );
BUFx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
BUFx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx5_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx8_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx6_ASAP7_75t_SL g170 ( .A(n_171), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_176), .Y(n_175) );
OR2x2_ASAP7_75t_SL g176 ( .A(n_177), .B(n_181), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AND3x1_ASAP7_75t_SL g516 ( .A(n_178), .B(n_181), .C(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g524 ( .A(n_178), .B(n_525), .Y(n_524) );
OA21x2_ASAP7_75t_L g530 ( .A1(n_178), .A2(n_215), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_179), .B(n_182), .Y(n_531) );
HB1xp67_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AND3x1_ASAP7_75t_L g184 ( .A(n_185), .B(n_420), .C(n_469), .Y(n_184) );
NOR3xp33_ASAP7_75t_SL g185 ( .A(n_186), .B(n_327), .C(n_365), .Y(n_185) );
OAI222xp33_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_248), .B1(n_302), .B2(n_308), .C1(n_322), .C2(n_325), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_188), .B(n_219), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_188), .B(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_188), .B(n_370), .Y(n_461) );
BUFx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
OR2x2_ASAP7_75t_L g338 ( .A(n_189), .B(n_239), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_189), .B(n_220), .Y(n_346) );
AND2x2_ASAP7_75t_L g381 ( .A(n_189), .B(n_358), .Y(n_381) );
OR2x2_ASAP7_75t_L g405 ( .A(n_189), .B(n_220), .Y(n_405) );
OR2x2_ASAP7_75t_L g413 ( .A(n_189), .B(n_312), .Y(n_413) );
AND2x2_ASAP7_75t_L g416 ( .A(n_189), .B(n_239), .Y(n_416) );
INVx3_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
OR2x2_ASAP7_75t_L g310 ( .A(n_190), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g324 ( .A(n_190), .B(n_239), .Y(n_324) );
AND2x2_ASAP7_75t_L g374 ( .A(n_190), .B(n_312), .Y(n_374) );
AND2x2_ASAP7_75t_L g387 ( .A(n_190), .B(n_220), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_190), .B(n_473), .Y(n_494) );
AO21x2_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_197), .B(n_217), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_191), .B(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g262 ( .A(n_191), .Y(n_262) );
AO21x2_ASAP7_75t_L g312 ( .A1(n_191), .A2(n_313), .B(n_320), .Y(n_312) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_192), .Y(n_223) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .Y(n_192) );
AND2x2_ASAP7_75t_SL g238 ( .A(n_193), .B(n_194), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
OAI22xp33_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_200), .B1(n_213), .B2(n_214), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_198), .A2(n_227), .B(n_228), .C(n_229), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_L g241 ( .A1(n_198), .A2(n_228), .B(n_242), .C(n_243), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_L g294 ( .A1(n_198), .A2(n_228), .B(n_295), .C(n_296), .Y(n_294) );
INVx4_ASAP7_75t_SL g198 ( .A(n_199), .Y(n_198) );
NAND2x1p5_ASAP7_75t_L g214 ( .A(n_199), .B(n_215), .Y(n_214) );
AND2x4_ASAP7_75t_L g225 ( .A(n_199), .B(n_215), .Y(n_225) );
INVx2_ASAP7_75t_L g319 ( .A(n_201), .Y(n_319) );
INVx3_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g211 ( .A(n_203), .Y(n_211) );
INVx1_ASAP7_75t_L g216 ( .A(n_203), .Y(n_216) );
OAI22xp5_ASAP7_75t_SL g204 ( .A1(n_205), .A2(n_207), .B1(n_208), .B2(n_209), .Y(n_204) );
INVx2_ASAP7_75t_L g208 ( .A(n_205), .Y(n_208) );
INVx4_ASAP7_75t_L g297 ( .A(n_205), .Y(n_297) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g212 ( .A(n_206), .Y(n_212) );
AND2x2_ASAP7_75t_L g215 ( .A(n_206), .B(n_216), .Y(n_215) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_206), .Y(n_231) );
INVx3_ASAP7_75t_L g234 ( .A(n_206), .Y(n_234) );
INVx1_ASAP7_75t_L g244 ( .A(n_206), .Y(n_244) );
INVx5_ASAP7_75t_L g228 ( .A(n_210), .Y(n_228) );
AND2x6_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_211), .Y(n_236) );
BUFx3_ASAP7_75t_L g261 ( .A(n_211), .Y(n_261) );
OAI21xp5_ASAP7_75t_L g266 ( .A1(n_214), .A2(n_267), .B(n_268), .Y(n_266) );
OAI21xp5_ASAP7_75t_L g313 ( .A1(n_214), .A2(n_314), .B(n_315), .Y(n_313) );
O2A1O1Ixp33_ASAP7_75t_L g412 ( .A1(n_219), .A2(n_413), .B(n_414), .C(n_417), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_219), .B(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_219), .B(n_357), .Y(n_479) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_239), .Y(n_219) );
AND2x2_ASAP7_75t_SL g323 ( .A(n_220), .B(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g337 ( .A(n_220), .Y(n_337) );
AND2x2_ASAP7_75t_L g364 ( .A(n_220), .B(n_358), .Y(n_364) );
INVx1_ASAP7_75t_SL g372 ( .A(n_220), .Y(n_372) );
AND2x2_ASAP7_75t_L g395 ( .A(n_220), .B(n_396), .Y(n_395) );
BUFx2_ASAP7_75t_L g473 ( .A(n_220), .Y(n_473) );
OA21x2_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_224), .B(n_237), .Y(n_220) );
INVx3_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_SL g263 ( .A(n_222), .B(n_264), .Y(n_263) );
INVx4_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_223), .A2(n_240), .B(n_247), .Y(n_239) );
BUFx2_ASAP7_75t_L g293 ( .A(n_225), .Y(n_293) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx4_ASAP7_75t_L g285 ( .A(n_231), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_234), .B(n_246), .Y(n_245) );
INVx5_ASAP7_75t_L g257 ( .A(n_234), .Y(n_257) );
INVx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_236), .Y(n_286) );
INVx1_ASAP7_75t_L g275 ( .A(n_238), .Y(n_275) );
INVx2_ASAP7_75t_L g279 ( .A(n_238), .Y(n_279) );
OA21x2_ASAP7_75t_L g291 ( .A1(n_238), .A2(n_292), .B(n_301), .Y(n_291) );
BUFx2_ASAP7_75t_L g309 ( .A(n_239), .Y(n_309) );
INVx1_ASAP7_75t_L g371 ( .A(n_239), .Y(n_371) );
INVx3_ASAP7_75t_L g396 ( .A(n_239), .Y(n_396) );
NAND2xp5_ASAP7_75t_SL g329 ( .A(n_248), .B(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_276), .Y(n_248) );
INVx1_ASAP7_75t_L g392 ( .A(n_249), .Y(n_392) );
OAI32xp33_ASAP7_75t_L g398 ( .A1(n_249), .A2(n_337), .A3(n_399), .B1(n_400), .B2(n_401), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_249), .A2(n_403), .B1(n_406), .B2(n_411), .Y(n_402) );
INVx4_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g340 ( .A(n_250), .B(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g418 ( .A(n_250), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g488 ( .A(n_250), .B(n_434), .Y(n_488) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_265), .Y(n_250) );
AND2x2_ASAP7_75t_L g303 ( .A(n_251), .B(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g333 ( .A(n_251), .Y(n_333) );
INVx1_ASAP7_75t_L g352 ( .A(n_251), .Y(n_352) );
OR2x2_ASAP7_75t_L g360 ( .A(n_251), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g367 ( .A(n_251), .B(n_341), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_251), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g388 ( .A(n_251), .B(n_306), .Y(n_388) );
INVx3_ASAP7_75t_L g410 ( .A(n_251), .Y(n_410) );
AND2x2_ASAP7_75t_L g435 ( .A(n_251), .B(n_307), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_251), .B(n_400), .Y(n_483) );
OR2x6_ASAP7_75t_L g251 ( .A(n_252), .B(n_263), .Y(n_251) );
AOI21xp5_ASAP7_75t_SL g252 ( .A1(n_253), .A2(n_254), .B(n_262), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_258), .B(n_259), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_L g316 ( .A1(n_257), .A2(n_317), .B(n_318), .C(n_319), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_259), .A2(n_270), .B(n_271), .Y(n_269) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g300 ( .A(n_261), .Y(n_300) );
INVx1_ASAP7_75t_L g272 ( .A(n_262), .Y(n_272) );
INVx2_ASAP7_75t_L g307 ( .A(n_265), .Y(n_307) );
AND2x2_ASAP7_75t_L g439 ( .A(n_265), .B(n_277), .Y(n_439) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_272), .B(n_273), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_275), .B(n_289), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_275), .B(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g481 ( .A(n_276), .Y(n_481) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_290), .Y(n_276) );
INVx1_ASAP7_75t_L g326 ( .A(n_277), .Y(n_326) );
AND2x2_ASAP7_75t_L g353 ( .A(n_277), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_277), .B(n_307), .Y(n_361) );
AND2x2_ASAP7_75t_L g419 ( .A(n_277), .B(n_342), .Y(n_419) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g305 ( .A(n_278), .Y(n_305) );
AND2x2_ASAP7_75t_L g332 ( .A(n_278), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g341 ( .A(n_278), .B(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_278), .B(n_307), .Y(n_407) );
AO21x2_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_280), .B(n_288), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_287), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_284), .B(n_286), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_290), .B(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g354 ( .A(n_290), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_290), .B(n_307), .Y(n_400) );
AND2x2_ASAP7_75t_L g409 ( .A(n_290), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g434 ( .A(n_290), .Y(n_434) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g306 ( .A(n_291), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g342 ( .A(n_291), .Y(n_342) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_293), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_297), .B(n_299), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_302), .A2(n_312), .B1(n_471), .B2(n_474), .Y(n_470) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
OAI21xp5_ASAP7_75t_SL g493 ( .A1(n_304), .A2(n_415), .B(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_305), .B(n_410), .Y(n_427) );
INVx1_ASAP7_75t_L g452 ( .A(n_305), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_306), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g379 ( .A(n_306), .B(n_332), .Y(n_379) );
INVx2_ASAP7_75t_L g335 ( .A(n_307), .Y(n_335) );
INVx1_ASAP7_75t_L g385 ( .A(n_307), .Y(n_385) );
OAI221xp5_ASAP7_75t_L g476 ( .A1(n_308), .A2(n_460), .B1(n_477), .B2(n_480), .C(n_482), .Y(n_476) );
OR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx1_ASAP7_75t_L g347 ( .A(n_309), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_309), .B(n_358), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_310), .B(n_369), .Y(n_368) );
OR2x2_ASAP7_75t_L g401 ( .A(n_310), .B(n_347), .Y(n_401) );
INVx3_ASAP7_75t_SL g442 ( .A(n_310), .Y(n_442) );
AND2x2_ASAP7_75t_L g386 ( .A(n_311), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g415 ( .A(n_311), .B(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_311), .B(n_324), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_311), .B(n_370), .Y(n_456) );
INVx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx3_ASAP7_75t_L g358 ( .A(n_312), .Y(n_358) );
OAI322xp33_ASAP7_75t_L g453 ( .A1(n_312), .A2(n_384), .A3(n_406), .B1(n_454), .B2(n_456), .C1(n_457), .C2(n_458), .Y(n_453) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AOI21xp33_ASAP7_75t_L g477 ( .A1(n_323), .A2(n_326), .B(n_478), .Y(n_477) );
NOR2xp33_ASAP7_75t_SL g403 ( .A(n_324), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g425 ( .A(n_324), .B(n_337), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_324), .B(n_364), .Y(n_440) );
INVxp67_ASAP7_75t_L g391 ( .A(n_326), .Y(n_391) );
AOI211xp5_ASAP7_75t_L g397 ( .A1(n_326), .A2(n_398), .B(n_402), .C(n_412), .Y(n_397) );
OAI221xp5_ASAP7_75t_SL g327 ( .A1(n_328), .A2(n_336), .B1(n_339), .B2(n_343), .C(n_348), .Y(n_327) );
INVxp67_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_334), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g351 ( .A(n_335), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g468 ( .A(n_335), .Y(n_468) );
OAI221xp5_ASAP7_75t_L g484 ( .A1(n_336), .A2(n_485), .B1(n_490), .B2(n_491), .C(n_493), .Y(n_484) );
OR2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_337), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_SL g384 ( .A(n_337), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_337), .B(n_415), .Y(n_422) );
AND2x2_ASAP7_75t_L g464 ( .A(n_337), .B(n_442), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_338), .B(n_363), .Y(n_362) );
OAI22xp33_ASAP7_75t_L g459 ( .A1(n_338), .A2(n_350), .B1(n_460), .B2(n_461), .Y(n_459) );
OR2x2_ASAP7_75t_L g490 ( .A(n_338), .B(n_358), .Y(n_490) );
CKINVDCx16_ASAP7_75t_R g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g467 ( .A(n_341), .Y(n_467) );
AND2x2_ASAP7_75t_L g492 ( .A(n_341), .B(n_435), .Y(n_492) );
INVxp67_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NOR2xp33_ASAP7_75t_SL g344 ( .A(n_345), .B(n_347), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g356 ( .A(n_346), .B(n_357), .Y(n_356) );
AOI22xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_355), .B1(n_359), .B2(n_362), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
INVx1_ASAP7_75t_L g423 ( .A(n_351), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_351), .B(n_391), .Y(n_458) );
AOI322xp5_ASAP7_75t_L g382 ( .A1(n_353), .A2(n_383), .A3(n_385), .B1(n_386), .B2(n_388), .C1(n_389), .C2(n_393), .Y(n_382) );
INVxp67_ASAP7_75t_L g376 ( .A(n_354), .Y(n_376) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_356), .A2(n_361), .B1(n_378), .B2(n_380), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_357), .B(n_370), .Y(n_457) );
INVx1_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_358), .B(n_396), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_358), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OR2x2_ASAP7_75t_L g454 ( .A(n_360), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
NAND3xp33_ASAP7_75t_SL g365 ( .A(n_366), .B(n_382), .C(n_397), .Y(n_365) );
AOI221xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .B1(n_373), .B2(n_375), .C(n_377), .Y(n_366) );
AND2x2_ASAP7_75t_L g373 ( .A(n_369), .B(n_374), .Y(n_373) );
INVx3_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
AND2x4_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
AND2x2_ASAP7_75t_L g383 ( .A(n_374), .B(n_384), .Y(n_383) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_376), .Y(n_455) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_381), .B(n_395), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_384), .B(n_442), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_385), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_SL g460 ( .A(n_388), .Y(n_460) );
AND2x2_ASAP7_75t_L g475 ( .A(n_388), .B(n_452), .Y(n_475) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AOI211xp5_ASAP7_75t_L g469 ( .A1(n_399), .A2(n_470), .B(n_476), .C(n_484), .Y(n_469) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OR2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g438 ( .A(n_409), .B(n_439), .Y(n_438) );
NAND2x1_ASAP7_75t_SL g480 ( .A(n_410), .B(n_481), .Y(n_480) );
CKINVDCx16_ASAP7_75t_R g450 ( .A(n_413), .Y(n_450) );
INVx1_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g445 ( .A(n_419), .Y(n_445) );
AND2x2_ASAP7_75t_L g449 ( .A(n_419), .B(n_435), .Y(n_449) );
NOR5xp2_ASAP7_75t_L g420 ( .A(n_421), .B(n_436), .C(n_453), .D(n_459), .E(n_462), .Y(n_420) );
OAI221xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_423), .B1(n_424), .B2(n_426), .C(n_428), .Y(n_421) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_425), .B(n_483), .Y(n_482) );
INVxp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_431), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_433), .B(n_435), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g451 ( .A(n_435), .B(n_452), .Y(n_451) );
OAI221xp5_ASAP7_75t_SL g436 ( .A1(n_437), .A2(n_440), .B1(n_441), .B2(n_443), .C(n_446), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_449), .B1(n_450), .B2(n_451), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g489 ( .A(n_449), .Y(n_489) );
AOI211xp5_ASAP7_75t_SL g462 ( .A1(n_463), .A2(n_465), .B(n_467), .C(n_468), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVxp67_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_487), .B(n_489), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
CKINVDCx14_ASAP7_75t_R g491 ( .A(n_492), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_496), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_497), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_503), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_503), .A2(n_524), .B1(n_533), .B2(n_535), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_508), .B1(n_514), .B2(n_515), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_504), .Y(n_514) );
INVx1_ASAP7_75t_L g507 ( .A(n_506), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_508), .Y(n_515) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_516), .Y(n_534) );
INVxp67_ASAP7_75t_L g527 ( .A(n_517), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
CKINVDCx16_ASAP7_75t_R g522 ( .A(n_523), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_526), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_529), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_530), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_534), .Y(n_533) );
endmodule