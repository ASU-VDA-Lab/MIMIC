module fake_jpeg_2163_n_651 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_651);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_651;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_60),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_61),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_62),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_63),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_64),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_23),
.B(n_10),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_65),
.B(n_66),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_23),
.B(n_10),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_67),
.Y(n_214)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_69),
.Y(n_157)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_70),
.Y(n_139)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_71),
.Y(n_217)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_73),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_75),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_29),
.B(n_8),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_76),
.B(n_80),
.Y(n_130)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_77),
.Y(n_180)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_78),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_33),
.B(n_8),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_79),
.B(n_95),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_11),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_81),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_35),
.B(n_11),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_82),
.B(n_102),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_83),
.Y(n_164)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_86),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_87),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_90),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_93),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_94),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_30),
.B(n_11),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_96),
.Y(n_216)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_97),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g185 ( 
.A(n_98),
.Y(n_185)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_99),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVxp67_ASAP7_75t_SL g187 ( 
.A(n_100),
.Y(n_187)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_7),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_104),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_105),
.Y(n_137)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_106),
.Y(n_173)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_21),
.Y(n_108)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_108),
.Y(n_193)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_43),
.Y(n_109)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_109),
.Y(n_181)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_43),
.Y(n_110)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_110),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_28),
.B(n_12),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_111),
.B(n_114),
.Y(n_156)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_46),
.Y(n_112)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_112),
.Y(n_202)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_46),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_113),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_57),
.B(n_41),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_31),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_115),
.B(n_121),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_28),
.B(n_12),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_116),
.B(n_125),
.Y(n_160)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_46),
.Y(n_117)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_117),
.Y(n_184)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_26),
.Y(n_118)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_50),
.Y(n_119)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_119),
.Y(n_188)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_37),
.Y(n_120)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_120),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_30),
.B(n_12),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_45),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_50),
.Y(n_123)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_123),
.Y(n_195)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_50),
.Y(n_124)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_124),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_42),
.B(n_18),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_26),
.Y(n_126)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_45),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g210 ( 
.A(n_127),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_37),
.Y(n_128)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_128),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_79),
.A2(n_25),
.B1(n_53),
.B2(n_37),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g277 ( 
.A1(n_133),
.A2(n_167),
.B1(n_179),
.B2(n_32),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_77),
.A2(n_53),
.B1(n_52),
.B2(n_50),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_136),
.A2(n_154),
.B1(n_163),
.B2(n_192),
.Y(n_242)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_142),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_64),
.A2(n_20),
.B1(n_25),
.B2(n_47),
.Y(n_154)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_100),
.Y(n_159)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_159),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_59),
.B(n_34),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_161),
.B(n_170),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_73),
.A2(n_53),
.B1(n_52),
.B2(n_40),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_67),
.A2(n_25),
.B1(n_19),
.B2(n_52),
.Y(n_167)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_105),
.A2(n_40),
.B(n_34),
.C(n_44),
.Y(n_169)
);

AOI21xp33_ASAP7_75t_L g232 ( 
.A1(n_169),
.A2(n_160),
.B(n_156),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_71),
.B(n_44),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_68),
.B(n_41),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_178),
.B(n_194),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_84),
.A2(n_19),
.B1(n_20),
.B2(n_42),
.Y(n_179)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_90),
.Y(n_182)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_182),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_91),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_186),
.B(n_81),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_106),
.B(n_27),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_190),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_75),
.A2(n_20),
.B1(n_47),
.B2(n_27),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_74),
.B(n_36),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_83),
.B(n_36),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_200),
.Y(n_227)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_96),
.Y(n_199)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_199),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_108),
.B(n_14),
.Y(n_200)
);

AND2x2_ASAP7_75t_SL g203 ( 
.A(n_98),
.B(n_31),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_99),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_87),
.A2(n_31),
.B1(n_45),
.B2(n_19),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_205),
.A2(n_32),
.B1(n_1),
.B2(n_2),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_128),
.B(n_13),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_219),
.Y(n_234)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_92),
.Y(n_211)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_211),
.Y(n_247)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_94),
.Y(n_212)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_212),
.Y(n_259)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_88),
.Y(n_215)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_215),
.Y(n_260)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_89),
.Y(n_218)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_218),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_78),
.B(n_13),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_137),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_220),
.B(n_226),
.Y(n_327)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_155),
.Y(n_221)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_221),
.Y(n_304)
);

O2A1O1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_169),
.A2(n_31),
.B(n_124),
.C(n_123),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_223),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_224),
.B(n_249),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_217),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_228),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_193),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_229),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_166),
.B(n_97),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_230),
.B(n_241),
.Y(n_306)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

INVx4_ASAP7_75t_SL g326 ( 
.A(n_231),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_232),
.A2(n_238),
.B(n_187),
.Y(n_300)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_155),
.Y(n_233)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_233),
.Y(n_328)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_168),
.Y(n_235)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_235),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_137),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_237),
.B(n_252),
.Y(n_309)
);

NAND2xp33_ASAP7_75t_SL g238 ( 
.A(n_190),
.B(n_0),
.Y(n_238)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_168),
.Y(n_239)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_239),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_130),
.B(n_93),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_154),
.A2(n_86),
.B1(n_63),
.B2(n_62),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_243),
.A2(n_279),
.B1(n_172),
.B2(n_174),
.Y(n_344)
);

BUFx12f_ASAP7_75t_L g244 ( 
.A(n_142),
.Y(n_244)
);

INVx11_ASAP7_75t_L g305 ( 
.A(n_244),
.Y(n_305)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_162),
.Y(n_245)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_245),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_175),
.Y(n_246)
);

INVx5_ASAP7_75t_L g308 ( 
.A(n_246),
.Y(n_308)
);

BUFx12_ASAP7_75t_L g248 ( 
.A(n_214),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g302 ( 
.A(n_248),
.Y(n_302)
);

AO22x2_ASAP7_75t_L g249 ( 
.A1(n_203),
.A2(n_31),
.B1(n_60),
.B2(n_61),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_129),
.B(n_13),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_250),
.B(n_258),
.Y(n_333)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_189),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_251),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_217),
.Y(n_252)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_175),
.Y(n_253)
);

INVx8_ASAP7_75t_L g313 ( 
.A(n_253),
.Y(n_313)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_213),
.Y(n_254)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_254),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_255),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_209),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_256),
.Y(n_343)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_213),
.Y(n_257)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_257),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_131),
.B(n_13),
.Y(n_258)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_139),
.Y(n_261)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_261),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_165),
.B(n_6),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_262),
.B(n_292),
.Y(n_321)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_216),
.Y(n_263)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_263),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_140),
.B(n_14),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_264),
.B(n_266),
.Y(n_314)
);

INVx6_ASAP7_75t_L g265 ( 
.A(n_176),
.Y(n_265)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_265),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_146),
.B(n_14),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_158),
.B(n_5),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_267),
.B(n_271),
.Y(n_334)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_193),
.Y(n_268)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_268),
.Y(n_324)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_173),
.Y(n_269)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_269),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_132),
.B(n_15),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_176),
.Y(n_272)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_272),
.Y(n_331)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_209),
.Y(n_273)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_273),
.Y(n_353)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_181),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_274),
.B(n_281),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_132),
.A2(n_32),
.B1(n_4),
.B2(n_16),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_167),
.A2(n_32),
.B1(n_4),
.B2(n_16),
.Y(n_276)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_188),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_278),
.B(n_290),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_192),
.A2(n_32),
.B1(n_1),
.B2(n_2),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_184),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_150),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_282),
.B(n_286),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_147),
.A2(n_4),
.B1(n_17),
.B2(n_18),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_283),
.A2(n_295),
.B1(n_296),
.B2(n_297),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_135),
.A2(n_18),
.B1(n_1),
.B2(n_2),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_284),
.A2(n_179),
.B1(n_148),
.B2(n_138),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_177),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_285),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_134),
.B(n_3),
.Y(n_286)
);

INVx8_ASAP7_75t_L g287 ( 
.A(n_185),
.Y(n_287)
);

BUFx8_ASAP7_75t_L g338 ( 
.A(n_287),
.Y(n_338)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_164),
.Y(n_288)
);

INVx6_ASAP7_75t_SL g322 ( 
.A(n_288),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_216),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_289),
.Y(n_355)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_195),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_153),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_143),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_294),
.Y(n_352)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_201),
.Y(n_295)
);

INVx11_ASAP7_75t_L g296 ( 
.A(n_185),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_171),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_300),
.B(n_244),
.Y(n_398)
);

INVx2_ASAP7_75t_R g301 ( 
.A(n_232),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_301),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_242),
.A2(n_157),
.B1(n_191),
.B2(n_202),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_311),
.A2(n_318),
.B1(n_344),
.B2(n_253),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_293),
.A2(n_249),
.B1(n_223),
.B2(n_224),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_316),
.A2(n_320),
.B1(n_325),
.B2(n_329),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_243),
.A2(n_187),
.B1(n_204),
.B2(n_207),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_249),
.A2(n_151),
.B1(n_143),
.B2(n_135),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_249),
.A2(n_151),
.B1(n_138),
.B2(n_180),
.Y(n_329)
);

OAI22xp33_ASAP7_75t_L g332 ( 
.A1(n_276),
.A2(n_177),
.B1(n_207),
.B2(n_204),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_332),
.A2(n_347),
.B1(n_351),
.B2(n_289),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_234),
.B(n_180),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_339),
.B(n_346),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_238),
.B(n_197),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_222),
.A2(n_208),
.B1(n_172),
.B2(n_141),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_279),
.A2(n_183),
.B1(n_145),
.B2(n_152),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_348),
.A2(n_244),
.B1(n_231),
.B2(n_296),
.Y(n_359)
);

BUFx12_ASAP7_75t_L g349 ( 
.A(n_280),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_349),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_227),
.A2(n_208),
.B1(n_196),
.B2(n_141),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_225),
.B(n_152),
.C(n_174),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_356),
.B(n_257),
.C(n_288),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_L g424 ( 
.A1(n_357),
.A2(n_331),
.B1(n_303),
.B2(n_342),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_345),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_358),
.B(n_377),
.Y(n_433)
);

OAI22xp33_ASAP7_75t_L g435 ( 
.A1(n_359),
.A2(n_363),
.B1(n_395),
.B2(n_305),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_306),
.B(n_291),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_362),
.B(n_381),
.Y(n_440)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_313),
.Y(n_364)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_364),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_307),
.B(n_277),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_365),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_307),
.A2(n_277),
.B1(n_149),
.B2(n_196),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_366),
.A2(n_373),
.B1(n_374),
.B2(n_394),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_322),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_367),
.Y(n_423)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_353),
.Y(n_368)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_368),
.Y(n_406)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_353),
.Y(n_370)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_370),
.Y(n_407)
);

O2A1O1Ixp33_ASAP7_75t_L g371 ( 
.A1(n_319),
.A2(n_240),
.B(n_260),
.C(n_247),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_371),
.B(n_372),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_339),
.B(n_259),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_307),
.A2(n_149),
.B1(n_275),
.B2(n_265),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_319),
.A2(n_344),
.B1(n_323),
.B2(n_316),
.Y(n_374)
);

NAND2xp33_ASAP7_75t_SL g375 ( 
.A(n_346),
.B(n_229),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_375),
.A2(n_398),
.B(n_342),
.Y(n_414)
);

BUFx5_ASAP7_75t_L g376 ( 
.A(n_338),
.Y(n_376)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_376),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_345),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_326),
.Y(n_379)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_379),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_329),
.A2(n_270),
.B1(n_269),
.B2(n_290),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_380),
.A2(n_388),
.B1(n_336),
.B2(n_310),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_345),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_306),
.B(n_239),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_382),
.A2(n_396),
.B(n_338),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_308),
.Y(n_383)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_383),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_350),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_384),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_322),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_385),
.B(n_386),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_354),
.B(n_268),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_337),
.B(n_221),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_387),
.B(n_391),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_320),
.A2(n_246),
.B1(n_285),
.B2(n_272),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_298),
.Y(n_389)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_389),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_314),
.B(n_236),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_390),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_301),
.B(n_333),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_298),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_392),
.B(n_393),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_301),
.B(n_233),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_300),
.A2(n_283),
.B1(n_263),
.B2(n_254),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_L g395 ( 
.A1(n_352),
.A2(n_336),
.B1(n_327),
.B2(n_309),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_352),
.A2(n_251),
.B(n_245),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_397),
.B(n_324),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_334),
.B(n_235),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_399),
.B(n_401),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_308),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_400),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_343),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_343),
.B(n_287),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_402),
.B(n_385),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_398),
.A2(n_338),
.B(n_356),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_404),
.A2(n_414),
.B(n_421),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_410),
.A2(n_411),
.B1(n_412),
.B2(n_418),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_374),
.A2(n_351),
.B1(n_332),
.B2(n_321),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_361),
.A2(n_321),
.B1(n_340),
.B2(n_310),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_413),
.B(n_397),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_417),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_361),
.A2(n_331),
.B1(n_313),
.B2(n_333),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_365),
.A2(n_326),
.B1(n_303),
.B2(n_338),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_424),
.A2(n_426),
.B1(n_428),
.B2(n_430),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g426 ( 
.A1(n_357),
.A2(n_355),
.B1(n_330),
.B2(n_324),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_363),
.A2(n_330),
.B1(n_315),
.B2(n_326),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_L g430 ( 
.A1(n_358),
.A2(n_335),
.B1(n_299),
.B2(n_315),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_367),
.Y(n_431)
);

CKINVDCx14_ASAP7_75t_R g445 ( 
.A(n_431),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_434),
.B(n_436),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_435),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_372),
.B(n_335),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_360),
.B(n_299),
.Y(n_438)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_438),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_366),
.A2(n_312),
.B1(n_341),
.B2(n_328),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_439),
.A2(n_389),
.B1(n_379),
.B2(n_364),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_408),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g508 ( 
.A(n_442),
.Y(n_508)
);

XOR2x2_ASAP7_75t_L g446 ( 
.A(n_415),
.B(n_391),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_446),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_448),
.B(n_465),
.Y(n_503)
);

OR2x6_ASAP7_75t_L g450 ( 
.A(n_416),
.B(n_378),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_450),
.B(n_460),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_409),
.A2(n_365),
.B1(n_394),
.B2(n_373),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_452),
.A2(n_453),
.B1(n_457),
.B2(n_469),
.Y(n_493)
);

CKINVDCx14_ASAP7_75t_R g453 ( 
.A(n_432),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_404),
.A2(n_393),
.B(n_378),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_454),
.A2(n_473),
.B(n_475),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_413),
.B(n_360),
.C(n_387),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_455),
.B(n_456),
.C(n_459),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_415),
.B(n_382),
.C(n_401),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_409),
.A2(n_382),
.B1(n_388),
.B2(n_381),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_408),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_458),
.B(n_470),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_404),
.B(n_386),
.C(n_377),
.Y(n_459)
);

A2O1A1Ixp33_ASAP7_75t_L g460 ( 
.A1(n_403),
.A2(n_371),
.B(n_362),
.C(n_375),
.Y(n_460)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_406),
.Y(n_463)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_463),
.Y(n_486)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_406),
.Y(n_464)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_464),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_433),
.B(n_368),
.C(n_370),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_434),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_466),
.B(n_476),
.Y(n_504)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_407),
.Y(n_467)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_467),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_440),
.B(n_399),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_468),
.B(n_419),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_418),
.A2(n_380),
.B1(n_396),
.B2(n_392),
.Y(n_469)
);

CKINVDCx14_ASAP7_75t_R g470 ( 
.A(n_432),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_407),
.Y(n_471)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_471),
.Y(n_495)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_472),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_412),
.A2(n_367),
.B1(n_402),
.B2(n_369),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_440),
.B(n_371),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_474),
.B(n_429),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_414),
.A2(n_376),
.B(n_305),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_437),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_437),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_477),
.B(n_430),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_463),
.Y(n_479)
);

BUFx12f_ASAP7_75t_L g515 ( 
.A(n_479),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_SL g480 ( 
.A(n_448),
.B(n_433),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_480),
.B(n_505),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_445),
.Y(n_481)
);

NOR3xp33_ASAP7_75t_L g530 ( 
.A(n_481),
.B(n_369),
.C(n_441),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_455),
.B(n_419),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_482),
.B(n_489),
.Y(n_514)
);

XOR2x2_ASAP7_75t_L g540 ( 
.A(n_483),
.B(n_450),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_443),
.A2(n_416),
.B(n_429),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_484),
.A2(n_502),
.B(n_450),
.Y(n_535)
);

NOR2x1p5_ASAP7_75t_L g487 ( 
.A(n_474),
.B(n_403),
.Y(n_487)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_487),
.Y(n_517)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_464),
.Y(n_488)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_488),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_461),
.A2(n_416),
.B1(n_438),
.B2(n_428),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_492),
.A2(n_497),
.B1(n_500),
.B2(n_510),
.Y(n_526)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_465),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_496),
.B(n_369),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_452),
.A2(n_442),
.B1(n_451),
.B2(n_466),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_457),
.A2(n_411),
.B1(n_424),
.B2(n_439),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_499),
.A2(n_506),
.B1(n_477),
.B2(n_476),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_451),
.A2(n_417),
.B1(n_410),
.B2(n_436),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_449),
.A2(n_421),
.B(n_431),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_446),
.B(n_421),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_473),
.A2(n_444),
.B1(n_469),
.B2(n_443),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_507),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_444),
.A2(n_405),
.B1(n_425),
.B2(n_422),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_459),
.B(n_420),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_511),
.B(n_450),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_478),
.B(n_447),
.Y(n_512)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_512),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_485),
.B(n_405),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g544 ( 
.A(n_513),
.B(n_529),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_503),
.B(n_456),
.C(n_454),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_516),
.B(n_519),
.C(n_522),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_493),
.A2(n_447),
.B1(n_462),
.B2(n_449),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_518),
.A2(n_520),
.B1(n_524),
.B2(n_537),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_503),
.B(n_460),
.C(n_420),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_497),
.A2(n_450),
.B1(n_475),
.B2(n_426),
.Y(n_520)
);

INVxp33_ASAP7_75t_L g521 ( 
.A(n_504),
.Y(n_521)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_521),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_485),
.B(n_480),
.C(n_511),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_508),
.B(n_471),
.Y(n_527)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_527),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_504),
.B(n_467),
.Y(n_528)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_528),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_509),
.B(n_427),
.Y(n_529)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_530),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_532),
.B(n_540),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_509),
.B(n_427),
.Y(n_533)
);

CKINVDCx16_ASAP7_75t_R g559 ( 
.A(n_533),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_479),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_534),
.B(n_539),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_L g546 ( 
.A1(n_535),
.A2(n_542),
.B(n_491),
.Y(n_546)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_488),
.Y(n_536)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_536),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_492),
.A2(n_450),
.B1(n_425),
.B2(n_422),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_538),
.B(n_484),
.Y(n_547)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_510),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_483),
.B(n_423),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_541),
.B(n_502),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_491),
.A2(n_441),
.B(n_423),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_546),
.B(n_537),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_547),
.B(n_526),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_526),
.A2(n_506),
.B1(n_499),
.B2(n_498),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_550),
.A2(n_525),
.B1(n_517),
.B2(n_528),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_518),
.A2(n_500),
.B1(n_498),
.B2(n_494),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_551),
.B(n_555),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_519),
.B(n_505),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_554),
.B(n_565),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_524),
.A2(n_494),
.B1(n_487),
.B2(n_507),
.Y(n_555)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_558),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_514),
.B(n_423),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_560),
.B(n_562),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_539),
.A2(n_487),
.B1(n_495),
.B2(n_490),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_522),
.B(n_486),
.C(n_495),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_563),
.B(n_564),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_516),
.B(n_486),
.C(n_501),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_531),
.B(n_312),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_538),
.B(n_341),
.C(n_304),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_567),
.B(n_540),
.C(n_535),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_569),
.B(n_572),
.Y(n_603)
);

XOR2xp5_ASAP7_75t_L g591 ( 
.A(n_570),
.B(n_571),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_563),
.B(n_531),
.C(n_542),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_564),
.B(n_545),
.C(n_554),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_573),
.B(n_576),
.Y(n_605)
);

MAJx2_ASAP7_75t_L g593 ( 
.A(n_575),
.B(n_556),
.C(n_543),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_545),
.B(n_540),
.C(n_520),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_SL g577 ( 
.A(n_548),
.B(n_514),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_577),
.B(n_581),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_567),
.B(n_527),
.C(n_517),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_578),
.B(n_580),
.C(n_582),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_557),
.B(n_536),
.C(n_523),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_566),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_565),
.B(n_523),
.C(n_512),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_551),
.B(n_525),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g595 ( 
.A(n_584),
.B(n_585),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_547),
.B(n_534),
.Y(n_585)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_566),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_587),
.B(n_584),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_561),
.B(n_400),
.C(n_383),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_588),
.B(n_546),
.C(n_561),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g606 ( 
.A(n_590),
.B(n_599),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_573),
.B(n_556),
.C(n_552),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_592),
.B(n_594),
.Y(n_614)
);

XOR2xp5_ASAP7_75t_L g615 ( 
.A(n_593),
.B(n_515),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_583),
.B(n_550),
.C(n_553),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_579),
.B(n_557),
.C(n_559),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_597),
.B(n_602),
.Y(n_610)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_598),
.Y(n_612)
);

XOR2xp5_ASAP7_75t_L g599 ( 
.A(n_572),
.B(n_562),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_SL g600 ( 
.A1(n_575),
.A2(n_549),
.B(n_568),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_L g608 ( 
.A1(n_600),
.A2(n_569),
.B(n_582),
.Y(n_608)
);

OAI21xp5_ASAP7_75t_SL g601 ( 
.A1(n_574),
.A2(n_543),
.B(n_549),
.Y(n_601)
);

OAI21xp5_ASAP7_75t_SL g609 ( 
.A1(n_601),
.A2(n_588),
.B(n_515),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_576),
.B(n_555),
.C(n_544),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_586),
.B(n_400),
.C(n_383),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_604),
.B(n_317),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_594),
.A2(n_571),
.B1(n_585),
.B2(n_578),
.Y(n_607)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_607),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_608),
.B(n_609),
.Y(n_625)
);

OAI21xp5_ASAP7_75t_SL g611 ( 
.A1(n_605),
.A2(n_515),
.B(n_302),
.Y(n_611)
);

OAI21xp5_ASAP7_75t_SL g622 ( 
.A1(n_611),
.A2(n_618),
.B(n_619),
.Y(n_622)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_603),
.B(n_515),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_613),
.B(n_616),
.Y(n_629)
);

XNOR2xp5_ASAP7_75t_L g628 ( 
.A(n_615),
.B(n_617),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_589),
.B(n_304),
.C(n_328),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_SL g618 ( 
.A1(n_600),
.A2(n_302),
.B(n_349),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_591),
.A2(n_317),
.B(n_302),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_613),
.Y(n_620)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_620),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_614),
.B(n_592),
.C(n_599),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_621),
.B(n_626),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_SL g624 ( 
.A1(n_610),
.A2(n_596),
.B(n_593),
.Y(n_624)
);

AO21x1_ASAP7_75t_L g637 ( 
.A1(n_624),
.A2(n_302),
.B(n_349),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_606),
.B(n_591),
.C(n_595),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_606),
.B(n_595),
.C(n_317),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_627),
.B(n_607),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_612),
.B(n_615),
.Y(n_630)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_630),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_620),
.B(n_608),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_631),
.B(n_635),
.Y(n_640)
);

AOI21x1_ASAP7_75t_L g635 ( 
.A1(n_625),
.A2(n_616),
.B(n_619),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_636),
.B(n_637),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_623),
.B(n_185),
.Y(n_638)
);

NOR2xp67_ASAP7_75t_SL g642 ( 
.A(n_638),
.B(n_628),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g639 ( 
.A(n_634),
.B(n_629),
.C(n_630),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_639),
.B(n_643),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g644 ( 
.A(n_642),
.B(n_632),
.C(n_633),
.Y(n_644)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_631),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_SL g646 ( 
.A1(n_644),
.A2(n_640),
.B(n_641),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_646),
.A2(n_645),
.B1(n_622),
.B2(n_349),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_L g648 ( 
.A1(n_647),
.A2(n_144),
.B(n_210),
.Y(n_648)
);

XNOR2xp5_ASAP7_75t_L g649 ( 
.A(n_648),
.B(n_248),
.Y(n_649)
);

XOR2xp5_ASAP7_75t_L g650 ( 
.A(n_649),
.B(n_248),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_SL g651 ( 
.A1(n_650),
.A2(n_0),
.B(n_2),
.Y(n_651)
);


endmodule