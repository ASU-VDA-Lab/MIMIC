module fake_jpeg_25664_n_198 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_198);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_198;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_11),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_12),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_26),
.B(n_27),
.Y(n_45)
);

HAxp5_ASAP7_75t_SL g27 ( 
.A(n_12),
.B(n_6),
.CON(n_27),
.SN(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_6),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_33),
.Y(n_41)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_24),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_24),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_31),
.Y(n_64)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_29),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_18),
.B1(n_21),
.B2(n_14),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_17),
.B1(n_18),
.B2(n_25),
.Y(n_62)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_17),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_47),
.B(n_26),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_32),
.B1(n_29),
.B2(n_31),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_48),
.A2(n_62),
.B1(n_52),
.B2(n_61),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_49),
.B(n_54),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_57),
.Y(n_84)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_16),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_56),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_16),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_14),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_37),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_63),
.A2(n_66),
.B1(n_70),
.B2(n_39),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_33),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_65),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_67),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_15),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_68),
.A2(n_41),
.B(n_20),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_28),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_44),
.C(n_35),
.Y(n_85)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_60),
.A2(n_43),
.B1(n_40),
.B2(n_39),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_72),
.A2(n_78),
.B1(n_79),
.B2(n_65),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_74),
.B(n_25),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_40),
.B(n_0),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_75),
.A2(n_58),
.B(n_54),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_85),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_64),
.A2(n_39),
.B1(n_33),
.B2(n_35),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_52),
.A2(n_35),
.B1(n_44),
.B2(n_36),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_87),
.B1(n_90),
.B2(n_55),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_51),
.A2(n_36),
.B1(n_15),
.B2(n_21),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_44),
.C(n_34),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_34),
.C(n_24),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_51),
.A2(n_20),
.B1(n_25),
.B2(n_22),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_92),
.Y(n_94)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_SL g119 ( 
.A1(n_95),
.A2(n_111),
.B(n_116),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_80),
.A2(n_70),
.B1(n_53),
.B2(n_67),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_98),
.B1(n_100),
.B2(n_78),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_75),
.A2(n_59),
.B(n_49),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_97),
.B(n_74),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_68),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_101),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_66),
.B1(n_63),
.B2(n_57),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_73),
.Y(n_101)
);

NOR2x1_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_34),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_104),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_103),
.B(n_107),
.Y(n_135)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_81),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_106),
.Y(n_122)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_24),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_110),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_56),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_113),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_34),
.C(n_19),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_81),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_114),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_82),
.B(n_19),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_79),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_0),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_124),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_111),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_128),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_85),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_84),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_127),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_113),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_130),
.A2(n_116),
.B(n_104),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_93),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_133),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_93),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_88),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_94),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_111),
.A2(n_65),
.B1(n_92),
.B2(n_77),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_136),
.A2(n_103),
.B1(n_107),
.B2(n_105),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_140),
.Y(n_162)
);

AO21x1_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_105),
.B(n_95),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_96),
.B1(n_102),
.B2(n_116),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_147),
.B1(n_150),
.B2(n_151),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_143),
.B(n_144),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_120),
.Y(n_145)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_145),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_91),
.Y(n_146)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_131),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_121),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_135),
.A2(n_94),
.B(n_91),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_149),
.B(n_129),
.C(n_124),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_154),
.C(n_158),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_129),
.C(n_133),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_145),
.A2(n_128),
.B1(n_117),
.B2(n_132),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_126),
.C(n_127),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_134),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_143),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_162),
.A2(n_147),
.B1(n_139),
.B2(n_151),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_165),
.Y(n_179)
);

INVx11_ASAP7_75t_L g165 ( 
.A(n_159),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_148),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_166),
.A2(n_169),
.B(n_170),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_154),
.C(n_152),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_137),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_150),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_153),
.Y(n_171)
);

NAND4xp25_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_23),
.C(n_2),
.D(n_3),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_157),
.A2(n_138),
.B1(n_140),
.B2(n_137),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_157),
.B1(n_140),
.B2(n_141),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_173),
.A2(n_175),
.B1(n_176),
.B2(n_180),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_177),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_168),
.A2(n_158),
.B1(n_125),
.B2(n_130),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_168),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_176)
);

MAJx2_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_22),
.C(n_23),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_169),
.Y(n_181)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_181),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_179),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_182),
.Y(n_190)
);

A2O1A1O1Ixp25_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_172),
.B(n_167),
.C(n_163),
.D(n_165),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_183),
.A2(n_184),
.B1(n_177),
.B2(n_174),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_175),
.A2(n_8),
.B1(n_4),
.B2(n_5),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_187),
.A2(n_188),
.B(n_183),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_186),
.A2(n_9),
.B1(n_5),
.B2(n_6),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_191),
.A2(n_192),
.B(n_189),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_190),
.A2(n_185),
.B(n_7),
.Y(n_192)
);

NOR3xp33_ASAP7_75t_L g195 ( 
.A(n_193),
.B(n_194),
.C(n_7),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_191),
.A2(n_185),
.B(n_7),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_195),
.A2(n_9),
.B(n_10),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_11),
.C(n_1),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_1),
.Y(n_198)
);


endmodule