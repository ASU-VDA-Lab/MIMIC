module real_jpeg_32334_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_0),
.A2(n_43),
.B1(n_48),
.B2(n_50),
.Y(n_42)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_0),
.Y(n_131)
);

AO22x1_ASAP7_75t_L g207 ( 
.A1(n_0),
.A2(n_50),
.B1(n_208),
.B2(n_211),
.Y(n_207)
);

AOI22x1_ASAP7_75t_L g275 ( 
.A1(n_0),
.A2(n_50),
.B1(n_276),
.B2(n_279),
.Y(n_275)
);

BUFx12f_ASAP7_75t_L g233 ( 
.A(n_1),
.Y(n_233)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_1),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_1),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_2),
.A2(n_15),
.B(n_527),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_2),
.B(n_528),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_4),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_5),
.Y(n_165)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_5),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_5),
.Y(n_243)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_5),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_6),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_86)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_6),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g221 ( 
.A1(n_6),
.A2(n_89),
.B1(n_222),
.B2(n_225),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_6),
.A2(n_89),
.B1(n_287),
.B2(n_290),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_6),
.A2(n_89),
.B1(n_276),
.B2(n_350),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_7),
.Y(n_106)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_7),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_7),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_7),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_9),
.A2(n_54),
.B1(n_59),
.B2(n_64),
.Y(n_53)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_9),
.A2(n_64),
.B1(n_133),
.B2(n_136),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_9),
.A2(n_64),
.B1(n_142),
.B2(n_146),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_9),
.A2(n_64),
.B1(n_241),
.B2(n_244),
.Y(n_240)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_10),
.Y(n_154)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_10),
.Y(n_159)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_11),
.Y(n_528)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_12),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_12),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_13),
.A2(n_79),
.B1(n_80),
.B2(n_83),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_13),
.Y(n_79)
);

OAI22x1_ASAP7_75t_SL g178 ( 
.A1(n_13),
.A2(n_79),
.B1(n_179),
.B2(n_183),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_13),
.A2(n_79),
.B1(n_252),
.B2(n_255),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_13),
.A2(n_79),
.B1(n_314),
.B2(n_316),
.Y(n_313)
);

INVx2_ASAP7_75t_R g340 ( 
.A(n_13),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_13),
.B(n_139),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_13),
.B(n_218),
.Y(n_386)
);

NAND2xp33_ASAP7_75t_SL g416 ( 
.A(n_13),
.B(n_21),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_13),
.B(n_430),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_67),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_66),
.Y(n_16)
);

OR2x2_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_65),
.Y(n_17)
);

NAND2x1_ASAP7_75t_SL g66 ( 
.A(n_18),
.B(n_65),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_18),
.B(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_18),
.B(n_196),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_42),
.B1(n_51),
.B2(n_53),
.Y(n_18)
);

AO21x1_ASAP7_75t_L g65 ( 
.A1(n_19),
.A2(n_51),
.B(n_53),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_19),
.A2(n_52),
.B(n_77),
.Y(n_259)
);

INVxp67_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_20),
.B(n_78),
.Y(n_172)
);

NOR2x1_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_32),
.Y(n_20)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

AO22x2_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_24),
.B1(n_27),
.B2(n_29),
.Y(n_21)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_23),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_23),
.Y(n_446)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_26),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_26),
.Y(n_124)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_27),
.Y(n_136)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_35),
.Y(n_441)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_40),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_42),
.A2(n_51),
.B(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_50),
.A2(n_122),
.B(n_125),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_52),
.A2(n_77),
.B1(n_86),
.B2(n_93),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_52),
.A2(n_86),
.B(n_172),
.Y(n_171)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21x1_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_296),
.B(n_515),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_197),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_195),
.Y(n_69)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_70),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_185),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g524 ( 
.A(n_71),
.B(n_185),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_168),
.C(n_173),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g199 ( 
.A1(n_73),
.A2(n_74),
.B1(n_168),
.B2(n_169),
.Y(n_199)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_94),
.B2(n_95),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_75),
.A2(n_76),
.B1(n_219),
.B2(n_417),
.Y(n_462)
);

OAI22x1_ASAP7_75t_L g491 ( 
.A1(n_75),
.A2(n_76),
.B1(n_271),
.B2(n_492),
.Y(n_491)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

HB1xp67_ASAP7_75t_SL g193 ( 
.A(n_76),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_76),
.B(n_219),
.C(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI211xp5_ASAP7_75t_SL g320 ( 
.A1(n_79),
.A2(n_321),
.B(n_324),
.C(n_327),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_79),
.B(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_79),
.B(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_140),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_96),
.B(n_193),
.C(n_194),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_121),
.B1(n_132),
.B2(n_137),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_97),
.B(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_98),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g219 ( 
.A1(n_98),
.A2(n_138),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

OA22x2_ASAP7_75t_L g271 ( 
.A1(n_98),
.A2(n_138),
.B1(n_220),
.B2(n_221),
.Y(n_271)
);

AOI21x1_ASAP7_75t_L g477 ( 
.A1(n_98),
.A2(n_138),
.B(n_220),
.Y(n_477)
);

NAND2x1p5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_112),
.Y(n_98)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

AOI22x1_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_104),
.B1(n_107),
.B2(n_109),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_103),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_106),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_106),
.Y(n_257)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_111),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_116),
.B1(n_117),
.B2(n_120),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_115),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_119),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_121),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_131),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_129),
.Y(n_338)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_132),
.B(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_136),
.B(n_443),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g137 ( 
.A(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_138),
.A2(n_176),
.B(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_138),
.B(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_168),
.C(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_140),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_140),
.A2(n_174),
.B1(n_175),
.B2(n_194),
.Y(n_203)
);

NAND2x1_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_149),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_141),
.A2(n_207),
.B1(n_213),
.B2(n_218),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_142),
.B(n_340),
.Y(n_339)
);

INVx4_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_145),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_148),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_149),
.B(n_251),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_162),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_150),
.B(n_250),
.Y(n_249)
);

OAI21xp33_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_157),
.B(n_162),
.Y(n_150)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_151),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_156),
.Y(n_289)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_156),
.Y(n_292)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_157),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_159),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_159),
.Y(n_166)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_162),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_162),
.Y(n_218)
);

OA22x2_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_166),
.B2(n_167),
.Y(n_162)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_164),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_164),
.Y(n_280)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_165),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_165),
.Y(n_383)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_169),
.B(n_203),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_170),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_170),
.B(n_271),
.C(n_452),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_171),
.B(n_477),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

XOR2x2_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_178),
.Y(n_220)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_181),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_182),
.Y(n_331)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_192),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_190),
.C(n_192),
.Y(n_196)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_193),
.Y(n_272)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_195),
.Y(n_517)
);

OA21x2_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_200),
.B(n_260),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_198),
.B(n_200),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_198),
.B(n_200),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.C(n_226),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_L g294 ( 
.A1(n_202),
.A2(n_204),
.B1(n_205),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_202),
.Y(n_295)
);

INVxp67_ASAP7_75t_SL g204 ( 
.A(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_205),
.A2(n_206),
.B(n_219),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_219),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_207),
.A2(n_218),
.B(n_249),
.Y(n_248)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AO22x2_ASAP7_75t_L g285 ( 
.A1(n_214),
.A2(n_218),
.B1(n_251),
.B2(n_286),
.Y(n_285)
);

AO22x2_ASAP7_75t_L g305 ( 
.A1(n_214),
.A2(n_218),
.B1(n_251),
.B2(n_286),
.Y(n_305)
);

AOI21x1_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B(n_217),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_215),
.A2(n_372),
.B1(n_377),
.B2(n_381),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_219),
.A2(n_413),
.B1(n_414),
.B2(n_417),
.Y(n_412)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_219),
.Y(n_417)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_226),
.B(n_294),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_247),
.B(n_258),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_227),
.B(n_248),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_227),
.A2(n_228),
.B1(n_247),
.B2(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XNOR2x1_ASAP7_75t_L g265 ( 
.A(n_228),
.B(n_259),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_240),
.Y(n_228)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_229),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_237),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_230),
.A2(n_275),
.B1(n_281),
.B2(n_282),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_230),
.Y(n_347)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_231),
.B(n_313),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g389 ( 
.A(n_232),
.B(n_340),
.Y(n_389)
);

INVx4_ASAP7_75t_SL g232 ( 
.A(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_236),
.Y(n_246)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_236),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_236),
.Y(n_318)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_236),
.Y(n_376)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_238),
.Y(n_284)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVxp33_ASAP7_75t_SL g281 ( 
.A(n_240),
.Y(n_281)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_243),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_247),
.Y(n_495)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_252),
.Y(n_380)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_257),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_293),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_261),
.B(n_293),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_266),
.C(n_268),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_262),
.A2(n_263),
.B1(n_266),
.B2(n_267),
.Y(n_499)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2x1_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_268),
.B(n_499),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_272),
.C(n_273),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_269),
.B(n_409),
.C(n_410),
.Y(n_408)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_271),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_271),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_271),
.A2(n_307),
.B1(n_452),
.B2(n_453),
.Y(n_451)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_271),
.Y(n_492)
);

XNOR2x1_ASAP7_75t_L g490 ( 
.A(n_273),
.B(n_491),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_285),
.Y(n_273)
);

XOR2x2_ASAP7_75t_L g479 ( 
.A(n_274),
.B(n_359),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_275),
.A2(n_365),
.B(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_285),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_285),
.B(n_401),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_285),
.A2(n_359),
.B1(n_419),
.B2(n_420),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_285),
.B(n_420),
.C(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

NAND2x1p5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_507),
.Y(n_297)
);

AOI21x1_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_455),
.B(n_506),
.Y(n_298)
);

AO21x2_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_422),
.B(n_454),
.Y(n_299)
);

AO21x1_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_407),
.B(n_421),
.Y(n_300)
);

OAI21x1_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_360),
.B(n_406),
.Y(n_301)
);

NOR2xp67_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_343),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_303),
.B(n_343),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_308),
.Y(n_303)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_305),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_305),
.A2(n_306),
.B1(n_370),
.B2(n_371),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_305),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_305),
.A2(n_306),
.B1(n_464),
.B2(n_468),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_305),
.B(n_464),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_306),
.B(n_370),
.Y(n_399)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_308),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_341),
.Y(n_308)
);

NAND3xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_320),
.C(n_332),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

OAI21xp33_ASAP7_75t_L g341 ( 
.A1(n_311),
.A2(n_333),
.B(n_342),
.Y(n_341)
);

OAI21xp33_ASAP7_75t_SL g419 ( 
.A1(n_311),
.A2(n_333),
.B(n_342),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_319),
.Y(n_311)
);

OA22x2_ASAP7_75t_L g402 ( 
.A1(n_312),
.A2(n_347),
.B1(n_348),
.B2(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_313),
.B(n_354),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_320),
.Y(n_342)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_330),
.Y(n_434)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_339),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_358),
.C(n_359),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_345),
.B(n_386),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_345),
.B(n_386),
.Y(n_396)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

OAI21xp33_ASAP7_75t_L g427 ( 
.A1(n_346),
.A2(n_428),
.B(n_447),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_346),
.B(n_428),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_348),
.B(n_353),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_349),
.B(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_357),
.Y(n_368)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_357),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_358),
.B(n_402),
.Y(n_401)
);

AOI21x1_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_398),
.B(n_405),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_384),
.B(n_397),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_369),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_363),
.B(n_369),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_363),
.A2(n_364),
.B1(n_415),
.B2(n_416),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_363),
.B(n_415),
.C(n_417),
.Y(n_448)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_364),
.B(n_388),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

BUFx2_ASAP7_75t_R g404 ( 
.A(n_368),
.Y(n_404)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g373 ( 
.A(n_374),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_385),
.A2(n_387),
.B(n_396),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_389),
.B(n_390),
.Y(n_388)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

OR2x2_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_400),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_399),
.B(n_400),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_404),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_411),
.Y(n_407)
);

NOR2xp67_ASAP7_75t_L g421 ( 
.A(n_408),
.B(n_411),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_418),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_412),
.Y(n_424)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_419),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_425),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_423),
.B(n_425),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_426),
.B(n_449),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_448),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_427),
.Y(n_484)
);

AO22x1_ASAP7_75t_L g428 ( 
.A1(n_429),
.A2(n_432),
.B1(n_438),
.B2(n_442),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_431),
.Y(n_430)
);

NAND2xp33_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_435),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx4_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx11_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

BUFx12f_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_447),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_448),
.Y(n_485)
);

MAJx2_ASAP7_75t_L g483 ( 
.A(n_449),
.B(n_484),
.C(n_485),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_450),
.B(n_477),
.C(n_478),
.Y(n_497)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_452),
.Y(n_453)
);

NOR2x1_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_486),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_480),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_457),
.B(n_512),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_471),
.Y(n_457)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_458),
.B(n_471),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_463),
.C(n_469),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_460),
.B(n_482),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_462),
.Y(n_460)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_461),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_463),
.B(n_470),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g468 ( 
.A(n_464),
.Y(n_468)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_474),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_472),
.B(n_502),
.C(n_503),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_479),
.Y(n_474)
);

INVxp33_ASAP7_75t_L g502 ( 
.A(n_475),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_478),
.Y(n_475)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_479),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_483),
.Y(n_480)
);

NOR2x1_ASAP7_75t_L g512 ( 
.A(n_481),
.B(n_483),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_500),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_487),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_498),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_488),
.B(n_498),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_493),
.C(n_496),
.Y(n_488)
);

INVxp33_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_490),
.B(n_494),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVxp33_ASAP7_75t_SL g496 ( 
.A(n_497),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_497),
.B(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_500),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_504),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_501),
.B(n_504),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_509),
.Y(n_507)
);

A2O1A1Ixp33_ASAP7_75t_L g509 ( 
.A1(n_510),
.A2(n_511),
.B(n_513),
.C(n_514),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_516),
.A2(n_519),
.B(n_523),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_518),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_517),
.A2(n_524),
.B(n_525),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_520),
.A2(n_521),
.B(n_522),
.Y(n_519)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);


endmodule