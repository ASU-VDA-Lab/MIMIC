module fake_jpeg_13397_n_445 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_445);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_445;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_16),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_8),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_60),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_28),
.B(n_15),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_61),
.B(n_66),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_33),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_62),
.B(n_87),
.Y(n_118)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_63),
.Y(n_141)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_28),
.B(n_15),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_32),
.B(n_15),
.Y(n_68)
);

NOR2xp67_ASAP7_75t_R g171 ( 
.A(n_68),
.B(n_104),
.Y(n_171)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_32),
.B(n_14),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_70),
.B(n_79),
.Y(n_136)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

BUFx4f_ASAP7_75t_SL g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_73),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_75),
.Y(n_153)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_40),
.Y(n_76)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_76),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_77),
.Y(n_157)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_78),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_41),
.B(n_14),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_80),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_81),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_41),
.B(n_10),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_82),
.B(n_90),
.Y(n_156)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_83),
.Y(n_159)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_84),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_85),
.Y(n_163)
);

BUFx12_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx6_ASAP7_75t_SL g164 ( 
.A(n_86),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_23),
.B(n_10),
.Y(n_87)
);

INVx6_ASAP7_75t_SL g88 ( 
.A(n_24),
.Y(n_88)
);

INVx5_ASAP7_75t_SL g142 ( 
.A(n_88),
.Y(n_142)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_46),
.B(n_10),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_23),
.Y(n_91)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_22),
.Y(n_92)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_92),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_46),
.B(n_2),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_100),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_22),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g174 ( 
.A(n_95),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_98),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_50),
.B(n_2),
.Y(n_100)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_35),
.Y(n_101)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_102),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_50),
.B(n_3),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_105),
.Y(n_131)
);

HAxp5_ASAP7_75t_SL g104 ( 
.A(n_35),
.B(n_3),
.CON(n_104),
.SN(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_56),
.B(n_8),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_106),
.Y(n_151)
);

BUFx10_ASAP7_75t_L g107 ( 
.A(n_35),
.Y(n_107)
);

INVx11_ASAP7_75t_L g155 ( 
.A(n_107),
.Y(n_155)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_40),
.Y(n_109)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_56),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_26),
.Y(n_140)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_27),
.Y(n_111)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_19),
.Y(n_112)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_112),
.Y(n_168)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_27),
.Y(n_113)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_113),
.Y(n_169)
);

AOI21xp33_ASAP7_75t_L g114 ( 
.A1(n_17),
.A2(n_4),
.B(n_5),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_114),
.A2(n_55),
.B(n_52),
.Y(n_124)
);

NAND2xp33_ASAP7_75t_SL g117 ( 
.A(n_87),
.B(n_38),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_117),
.B(n_124),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_59),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_129),
.B(n_140),
.Y(n_238)
);

OR2x2_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_26),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_133),
.B(n_175),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_89),
.A2(n_38),
.B1(n_29),
.B2(n_18),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_143),
.A2(n_176),
.B1(n_178),
.B2(n_51),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_94),
.B(n_29),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_144),
.B(n_160),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_94),
.B(n_55),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_104),
.A2(n_53),
.B1(n_18),
.B2(n_48),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_161),
.A2(n_165),
.B1(n_166),
.B2(n_173),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_76),
.A2(n_53),
.B1(n_18),
.B2(n_54),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_60),
.A2(n_53),
.B1(n_37),
.B2(n_44),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_97),
.B(n_52),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_180),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_64),
.A2(n_44),
.B1(n_42),
.B2(n_37),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_107),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_77),
.A2(n_54),
.B1(n_42),
.B2(n_34),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_80),
.A2(n_21),
.B1(n_47),
.B2(n_43),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_97),
.B(n_21),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_101),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_181),
.Y(n_200)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_122),
.Y(n_182)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_182),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_142),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_184),
.B(n_194),
.Y(n_243)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_185),
.Y(n_248)
);

AND2x4_ASAP7_75t_SL g186 ( 
.A(n_171),
.B(n_78),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_186),
.Y(n_267)
);

O2A1O1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_142),
.A2(n_161),
.B(n_118),
.C(n_178),
.Y(n_187)
);

NAND2xp33_ASAP7_75t_L g268 ( 
.A(n_187),
.B(n_240),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_150),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_188),
.A2(n_191),
.B1(n_213),
.B2(n_215),
.Y(n_271)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_169),
.Y(n_189)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_189),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_146),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_190),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_148),
.A2(n_65),
.B1(n_81),
.B2(n_99),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_192),
.A2(n_163),
.B1(n_132),
.B2(n_120),
.Y(n_261)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_128),
.Y(n_193)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_193),
.Y(n_259)
);

O2A1O1Ixp33_ASAP7_75t_SL g194 ( 
.A1(n_176),
.A2(n_73),
.B(n_109),
.C(n_86),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_141),
.Y(n_195)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_195),
.Y(n_255)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_139),
.Y(n_196)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_196),
.Y(n_269)
);

INVxp33_ASAP7_75t_L g197 ( 
.A(n_155),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_197),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_198),
.Y(n_280)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_152),
.Y(n_199)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_199),
.Y(n_263)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_116),
.Y(n_201)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_201),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_202),
.Y(n_282)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_203),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_164),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_204),
.B(n_217),
.Y(n_247)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_151),
.Y(n_205)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_205),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_131),
.A2(n_106),
.B1(n_102),
.B2(n_96),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_206),
.A2(n_220),
.B1(n_234),
.B2(n_239),
.Y(n_246)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_126),
.Y(n_209)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_209),
.Y(n_276)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_139),
.Y(n_210)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_210),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_155),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_211),
.B(n_224),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_130),
.A2(n_98),
.B1(n_95),
.B2(n_36),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_115),
.A2(n_34),
.B1(n_51),
.B2(n_47),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_127),
.B(n_20),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_216),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_167),
.B(n_20),
.C(n_43),
.Y(n_217)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_116),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_218),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_115),
.A2(n_130),
.B1(n_145),
.B2(n_153),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_219),
.A2(n_145),
.B1(n_162),
.B2(n_172),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_156),
.A2(n_17),
.B1(n_36),
.B2(n_71),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_135),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_221),
.Y(n_284)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_174),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_222),
.B(n_225),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_157),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_223),
.A2(n_226),
.B1(n_231),
.B2(n_236),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_134),
.B(n_6),
.Y(n_224)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_174),
.Y(n_225)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_137),
.Y(n_226)
);

INVx13_ASAP7_75t_L g227 ( 
.A(n_119),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_227),
.Y(n_257)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_159),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_228),
.Y(n_281)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_158),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_229),
.B(n_230),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_136),
.B(n_6),
.Y(n_230)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_137),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_179),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_232),
.B(n_233),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_119),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_165),
.A2(n_7),
.B1(n_8),
.B2(n_166),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_147),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_147),
.Y(n_242)
);

INVx8_ASAP7_75t_L g236 ( 
.A(n_121),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_237),
.A2(n_120),
.B1(n_163),
.B2(n_226),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_173),
.A2(n_7),
.B1(n_121),
.B2(n_125),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_137),
.B(n_149),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_242),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_194),
.A2(n_172),
.B1(n_153),
.B2(n_125),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_244),
.A2(n_258),
.B1(n_231),
.B2(n_200),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_177),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_249),
.B(n_252),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_250),
.A2(n_279),
.B1(n_223),
.B2(n_198),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_186),
.B(n_123),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_186),
.B(n_138),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_254),
.B(n_277),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_234),
.A2(n_162),
.B1(n_132),
.B2(n_174),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_261),
.A2(n_258),
.B1(n_262),
.B2(n_252),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_265),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_207),
.A2(n_120),
.B1(n_163),
.B2(n_187),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_270),
.A2(n_197),
.B1(n_225),
.B2(n_222),
.Y(n_298)
);

AO22x1_ASAP7_75t_L g273 ( 
.A1(n_207),
.A2(n_239),
.B1(n_213),
.B2(n_211),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_273),
.A2(n_261),
.B(n_243),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_183),
.B(n_230),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_188),
.A2(n_191),
.B1(n_215),
.B2(n_219),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_216),
.B(n_238),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_283),
.B(n_251),
.Y(n_315)
);

INVx8_ASAP7_75t_L g287 ( 
.A(n_257),
.Y(n_287)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_287),
.Y(n_331)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_242),
.Y(n_289)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_289),
.Y(n_324)
);

OAI21xp33_ASAP7_75t_SL g341 ( 
.A1(n_290),
.A2(n_312),
.B(n_286),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_272),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_291),
.B(n_292),
.Y(n_337)
);

NAND3xp33_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_214),
.C(n_227),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g346 ( 
.A(n_293),
.Y(n_346)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_259),
.Y(n_294)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_294),
.Y(n_328)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_259),
.Y(n_295)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_295),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_296),
.A2(n_273),
.B1(n_260),
.B2(n_279),
.Y(n_326)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_263),
.Y(n_297)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_297),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_298),
.A2(n_303),
.B(n_310),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_245),
.B(n_208),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_300),
.B(n_302),
.Y(n_347)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_263),
.Y(n_301)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_301),
.Y(n_344)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_274),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_268),
.A2(n_208),
.B(n_214),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_249),
.B(n_217),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_304),
.Y(n_322)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_274),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_305),
.B(n_307),
.Y(n_325)
);

INVx11_ASAP7_75t_L g306 ( 
.A(n_257),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_306),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_246),
.A2(n_190),
.B1(n_201),
.B2(n_218),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_277),
.B(n_196),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_309),
.B(n_271),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_267),
.A2(n_210),
.B1(n_205),
.B2(n_236),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_283),
.B(n_247),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_311),
.A2(n_282),
.B(n_284),
.Y(n_345)
);

BUFx12f_ASAP7_75t_L g313 ( 
.A(n_281),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_313),
.B(n_315),
.Y(n_330)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_241),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_316),
.B(n_318),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_246),
.A2(n_254),
.B1(n_273),
.B2(n_271),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_317),
.B(n_253),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_256),
.B(n_241),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_248),
.B(n_256),
.C(n_266),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_319),
.B(n_320),
.C(n_285),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_248),
.B(n_266),
.C(n_276),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_276),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_321),
.B(n_319),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_323),
.B(n_335),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_326),
.A2(n_327),
.B1(n_334),
.B2(n_341),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_296),
.A2(n_250),
.B1(n_260),
.B2(n_280),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_299),
.B(n_278),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_333),
.B(n_309),
.C(n_299),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_289),
.A2(n_280),
.B1(n_281),
.B2(n_264),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_335),
.B(n_339),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_336),
.B(n_343),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_308),
.B(n_264),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_308),
.B(n_285),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_345),
.B(n_306),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_348),
.A2(n_288),
.B1(n_310),
.B2(n_318),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_322),
.B(n_291),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_349),
.B(n_352),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_348),
.A2(n_303),
.B(n_314),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_350),
.A2(n_355),
.B(n_360),
.Y(n_384)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_328),
.Y(n_351)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_351),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_336),
.B(n_288),
.C(n_315),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_353),
.B(n_364),
.C(n_365),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_356),
.A2(n_363),
.B1(n_366),
.B2(n_370),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_345),
.Y(n_357)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_357),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_322),
.B(n_311),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_358),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_326),
.A2(n_317),
.B1(n_312),
.B2(n_314),
.Y(n_360)
);

BUFx24_ASAP7_75t_SL g361 ( 
.A(n_337),
.Y(n_361)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_361),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_331),
.Y(n_362)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_362),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_324),
.A2(n_290),
.B1(n_293),
.B2(n_316),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_SL g364 ( 
.A(n_337),
.B(n_347),
.C(n_341),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_333),
.B(n_320),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_324),
.A2(n_294),
.B1(n_301),
.B2(n_297),
.Y(n_366)
);

XNOR2x1_ASAP7_75t_L g374 ( 
.A(n_367),
.B(n_332),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_323),
.B(n_347),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_368),
.B(n_343),
.C(n_332),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_323),
.A2(n_295),
.B1(n_321),
.B2(n_287),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_357),
.A2(n_346),
.B1(n_330),
.B2(n_327),
.Y(n_372)
);

XNOR2x1_ASAP7_75t_L g394 ( 
.A(n_372),
.B(n_374),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_363),
.A2(n_346),
.B1(n_330),
.B2(n_339),
.Y(n_373)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_373),
.Y(n_393)
);

AO22x1_ASAP7_75t_SL g376 ( 
.A1(n_369),
.A2(n_338),
.B1(n_325),
.B2(n_331),
.Y(n_376)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_376),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_382),
.B(n_387),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_370),
.A2(n_325),
.B1(n_334),
.B2(n_340),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_383),
.B(n_359),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_360),
.A2(n_338),
.B1(n_340),
.B2(n_342),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_385),
.A2(n_369),
.B1(n_367),
.B2(n_366),
.Y(n_395)
);

OAI21xp33_ASAP7_75t_SL g386 ( 
.A1(n_350),
.A2(n_344),
.B(n_342),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_386),
.A2(n_313),
.B1(n_302),
.B2(n_362),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_354),
.B(n_344),
.C(n_329),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_359),
.A2(n_364),
.B(n_352),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_388),
.A2(n_328),
.B(n_305),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_379),
.B(n_353),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_390),
.B(n_391),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_379),
.B(n_365),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_392),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_395),
.A2(n_396),
.B1(n_402),
.B2(n_372),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_385),
.A2(n_368),
.B1(n_351),
.B2(n_329),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_373),
.B(n_351),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_397),
.B(n_371),
.C(n_382),
.Y(n_412)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_381),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_400),
.B(n_401),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_380),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_381),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_403),
.A2(n_378),
.B(n_384),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_404),
.B(n_383),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g405 ( 
.A(n_394),
.B(n_374),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_405),
.B(n_407),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_394),
.B(n_375),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_408),
.A2(n_403),
.B(n_404),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_410),
.B(n_413),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_412),
.B(n_414),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g413 ( 
.A(n_396),
.B(n_375),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_398),
.A2(n_371),
.B1(n_384),
.B2(n_377),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_415),
.A2(n_414),
.B1(n_398),
.B2(n_393),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_416),
.B(n_423),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_SL g417 ( 
.A1(n_409),
.A2(n_393),
.B1(n_376),
.B2(n_392),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_417),
.A2(n_422),
.B(n_376),
.Y(n_429)
);

AOI21x1_ASAP7_75t_L g425 ( 
.A1(n_419),
.A2(n_420),
.B(n_413),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_412),
.A2(n_399),
.B(n_388),
.Y(n_420)
);

AO21x1_ASAP7_75t_L g422 ( 
.A1(n_411),
.A2(n_395),
.B(n_397),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_406),
.B(n_387),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_425),
.B(n_431),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_418),
.B(n_389),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_426),
.B(n_428),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_424),
.B(n_407),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_429),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_418),
.B(n_389),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_430),
.B(n_405),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_421),
.B(n_424),
.Y(n_431)
);

OR2x2_ASAP7_75t_L g434 ( 
.A(n_427),
.B(n_417),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_434),
.A2(n_422),
.B(n_429),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_435),
.B(n_431),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_437),
.B(n_438),
.Y(n_440)
);

AOI31xp67_ASAP7_75t_L g439 ( 
.A1(n_432),
.A2(n_313),
.A3(n_282),
.B(n_284),
.Y(n_439)
);

A2O1A1O1Ixp25_ASAP7_75t_L g441 ( 
.A1(n_439),
.A2(n_313),
.B(n_286),
.C(n_253),
.D(n_433),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_441),
.B(n_436),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_442),
.B(n_434),
.C(n_440),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_443),
.A2(n_255),
.B1(n_269),
.B2(n_440),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_444),
.B(n_269),
.Y(n_445)
);


endmodule