module fake_netlist_5_731_n_771 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_771);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_771;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_667;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_452;
wire n_397;
wire n_525;
wire n_493;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_155;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_564;
wire n_467;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_443;
wire n_372;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_150;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_152;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_379;
wire n_308;
wire n_428;
wire n_267;
wire n_570;
wire n_457;
wire n_514;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_185;
wire n_183;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_169;
wire n_550;
wire n_522;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_432;
wire n_164;
wire n_553;
wire n_395;
wire n_727;
wire n_311;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_517;
wire n_482;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_477;
wire n_338;
wire n_149;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_151;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_729;
wire n_730;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_710;
wire n_707;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_409;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_766;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_162;
wire n_759;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_140),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_31),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_78),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_65),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_5),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_48),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_62),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_64),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_54),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_0),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_141),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_91),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_67),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_74),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_60),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_3),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_59),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_13),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_46),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_86),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_26),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_124),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_61),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_144),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_137),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_49),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_23),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_47),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_108),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_76),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_2),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_50),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_143),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_53),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_17),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_132),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_101),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_68),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_71),
.Y(n_189)
);

BUFx8_ASAP7_75t_SL g190 ( 
.A(n_125),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_32),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_34),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_7),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_99),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_88),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_85),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_23),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_5),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_89),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_52),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_116),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

AND2x4_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_148),
.Y(n_203)
);

AND2x4_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_24),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_0),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_1),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

AND2x4_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_25),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_151),
.Y(n_211)
);

AND2x4_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_147),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_1),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_153),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

AND2x4_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_146),
.Y(n_217)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_155),
.B(n_2),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_177),
.B(n_3),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_152),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_156),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_157),
.B(n_4),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_161),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

AND2x6_ASAP7_75t_L g228 ( 
.A(n_167),
.B(n_27),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_169),
.B(n_176),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_180),
.B(n_4),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g231 ( 
.A(n_152),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_188),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_168),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_189),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_199),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_150),
.B(n_6),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_168),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_158),
.Y(n_238)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_190),
.Y(n_239)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_160),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_162),
.B(n_6),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_206),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_234),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

OR2x6_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_181),
.Y(n_246)
);

AO22x2_ASAP7_75t_L g247 ( 
.A1(n_203),
.A2(n_204),
.B1(n_210),
.B2(n_212),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_206),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_163),
.Y(n_249)
);

AO22x2_ASAP7_75t_L g250 ( 
.A1(n_203),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_205),
.A2(n_201),
.B1(n_200),
.B2(n_154),
.Y(n_251)
);

OR2x6_ASAP7_75t_L g252 ( 
.A(n_215),
.B(n_181),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_211),
.B(n_154),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_236),
.A2(n_201),
.B1(n_200),
.B2(n_196),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_202),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_216),
.A2(n_149),
.B1(n_192),
.B2(n_191),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_202),
.B(n_164),
.Y(n_258)
);

AO22x2_ASAP7_75t_L g259 ( 
.A1(n_203),
.A2(n_204),
.B1(n_210),
.B2(n_212),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_211),
.B(n_166),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_241),
.A2(n_194),
.B1(n_187),
.B2(n_186),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_170),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_L g263 ( 
.A1(n_227),
.A2(n_149),
.B1(n_183),
.B2(n_178),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_206),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_206),
.Y(n_265)
);

OR2x6_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_8),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_223),
.B(n_171),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_224),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_206),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_213),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_L g271 ( 
.A1(n_233),
.A2(n_237),
.B1(n_221),
.B2(n_214),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_235),
.Y(n_272)
);

INVx8_ASAP7_75t_L g273 ( 
.A(n_239),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_235),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_211),
.B(n_226),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_231),
.A2(n_184),
.B1(n_175),
.B2(n_174),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_239),
.B(n_28),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_219),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_222),
.A2(n_225),
.B1(n_230),
.B2(n_207),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_239),
.B(n_226),
.Y(n_280)
);

AO22x2_ASAP7_75t_L g281 ( 
.A1(n_203),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_281)
);

AO22x2_ASAP7_75t_L g282 ( 
.A1(n_204),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_238),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_232),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_226),
.B(n_222),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_219),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_232),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_238),
.B(n_29),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_239),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_254),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_233),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_268),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_238),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_261),
.B(n_217),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_229),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_274),
.Y(n_297)
);

INVxp33_ASAP7_75t_L g298 ( 
.A(n_258),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

BUFx6f_ASAP7_75t_SL g300 ( 
.A(n_246),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_287),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_275),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_249),
.B(n_240),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_242),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_275),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_244),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_245),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_264),
.Y(n_308)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_253),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_243),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_264),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_264),
.Y(n_312)
);

INVx4_ASAP7_75t_SL g313 ( 
.A(n_277),
.Y(n_313)
);

NAND2x1p5_ASAP7_75t_L g314 ( 
.A(n_280),
.B(n_217),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_253),
.B(n_239),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_285),
.B(n_260),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_269),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_269),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_257),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_262),
.B(n_240),
.Y(n_320)
);

INVxp33_ASAP7_75t_L g321 ( 
.A(n_267),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_243),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_269),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_255),
.B(n_251),
.Y(n_324)
);

INVxp33_ASAP7_75t_L g325 ( 
.A(n_285),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_260),
.B(n_240),
.Y(n_326)
);

OR2x2_ASAP7_75t_SL g327 ( 
.A(n_263),
.B(n_220),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_248),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_248),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_278),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_263),
.B(n_240),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_256),
.B(n_240),
.Y(n_332)
);

XNOR2x2_ASAP7_75t_L g333 ( 
.A(n_250),
.B(n_213),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_278),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_286),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_286),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_265),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_265),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_265),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_265),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_247),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_247),
.Y(n_342)
);

INVxp33_ASAP7_75t_L g343 ( 
.A(n_250),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_247),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_259),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_259),
.B(n_240),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_246),
.B(n_204),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_256),
.B(n_239),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_246),
.B(n_210),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_259),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_283),
.B(n_220),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_R g352 ( 
.A(n_304),
.B(n_288),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_325),
.B(n_250),
.Y(n_353)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_344),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_325),
.B(n_281),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_293),
.B(n_283),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_293),
.B(n_283),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_316),
.B(n_281),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_344),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_296),
.B(n_281),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_296),
.B(n_210),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_310),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_351),
.B(n_212),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_298),
.B(n_271),
.Y(n_364)
);

AND2x4_ASAP7_75t_L g365 ( 
.A(n_302),
.B(n_212),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_341),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_310),
.Y(n_367)
);

INVxp33_ASAP7_75t_L g368 ( 
.A(n_291),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_342),
.B(n_228),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_345),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_305),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_350),
.B(n_228),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_290),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_332),
.B(n_217),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_309),
.B(n_282),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_332),
.B(n_217),
.Y(n_376)
);

AND2x6_ASAP7_75t_L g377 ( 
.A(n_346),
.B(n_282),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_298),
.B(n_271),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_295),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_322),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_309),
.B(n_228),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_292),
.B(n_266),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_294),
.B(n_228),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_295),
.Y(n_384)
);

OAI21xp33_ASAP7_75t_L g385 ( 
.A1(n_331),
.A2(n_282),
.B(n_214),
.Y(n_385)
);

AND2x2_ASAP7_75t_SL g386 ( 
.A(n_331),
.B(n_228),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_322),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_348),
.B(n_209),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_328),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_329),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_297),
.B(n_228),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_321),
.B(n_209),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_315),
.B(n_228),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_311),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_314),
.B(n_232),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_314),
.B(n_232),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_321),
.B(n_266),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_289),
.B(n_299),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_343),
.B(n_266),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_301),
.B(n_326),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_337),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_327),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_324),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_326),
.B(n_232),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_343),
.A2(n_208),
.B1(n_252),
.B2(n_219),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_319),
.B(n_306),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_307),
.B(n_208),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_330),
.Y(n_408)
);

BUFx5_ASAP7_75t_L g409 ( 
.A(n_334),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_335),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_347),
.B(n_252),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_336),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_333),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_308),
.B(n_208),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_312),
.B(n_219),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_317),
.B(n_219),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_318),
.B(n_218),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_338),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_361),
.B(n_313),
.Y(n_419)
);

OR2x2_ASAP7_75t_L g420 ( 
.A(n_402),
.B(n_252),
.Y(n_420)
);

OR2x6_ASAP7_75t_L g421 ( 
.A(n_354),
.B(n_273),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_362),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_359),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_406),
.B(n_300),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_378),
.B(n_349),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_366),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_359),
.B(n_313),
.Y(n_427)
);

NAND2x1p5_ASAP7_75t_L g428 ( 
.A(n_354),
.B(n_323),
.Y(n_428)
);

BUFx12f_ASAP7_75t_L g429 ( 
.A(n_382),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_392),
.B(n_313),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_362),
.Y(n_431)
);

NAND2xp33_ASAP7_75t_L g432 ( 
.A(n_356),
.B(n_339),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_366),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_392),
.B(n_340),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_354),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g436 ( 
.A(n_413),
.B(n_12),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_399),
.Y(n_437)
);

AND2x6_ASAP7_75t_L g438 ( 
.A(n_366),
.B(n_303),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_360),
.B(n_303),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_357),
.B(n_320),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_379),
.B(n_320),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_412),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_412),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_366),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_373),
.B(n_30),
.Y(n_445)
);

AND2x6_ASAP7_75t_L g446 ( 
.A(n_366),
.B(n_300),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_370),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_370),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_367),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_364),
.B(n_384),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_370),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_397),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_373),
.B(n_33),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_371),
.B(n_13),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_370),
.B(n_358),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_367),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_403),
.B(n_14),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_388),
.B(n_218),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_399),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_411),
.B(n_273),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_380),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_352),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_370),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_360),
.B(n_35),
.Y(n_464)
);

BUFx4f_ASAP7_75t_L g465 ( 
.A(n_377),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_358),
.B(n_36),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_353),
.Y(n_467)
);

NAND2x1p5_ASAP7_75t_L g468 ( 
.A(n_394),
.B(n_218),
.Y(n_468)
);

OR2x6_ASAP7_75t_L g469 ( 
.A(n_353),
.B(n_273),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_385),
.B(n_218),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_380),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_387),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_388),
.B(n_365),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_365),
.B(n_218),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_422),
.Y(n_475)
);

BUFx4f_ASAP7_75t_SL g476 ( 
.A(n_429),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_442),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_429),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_433),
.Y(n_479)
);

INVx3_ASAP7_75t_SL g480 ( 
.A(n_462),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_433),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_443),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_455),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_450),
.B(n_355),
.Y(n_484)
);

INVx5_ASAP7_75t_L g485 ( 
.A(n_421),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_467),
.Y(n_486)
);

BUFx12f_ASAP7_75t_L g487 ( 
.A(n_462),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_425),
.B(n_375),
.Y(n_488)
);

INVx8_ASAP7_75t_L g489 ( 
.A(n_446),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_422),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_450),
.B(n_355),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_437),
.Y(n_492)
);

NAND2x1p5_ASAP7_75t_L g493 ( 
.A(n_430),
.B(n_401),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_431),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_431),
.Y(n_495)
);

INVx6_ASAP7_75t_L g496 ( 
.A(n_445),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_449),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_449),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_426),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g500 ( 
.A1(n_439),
.A2(n_385),
.B1(n_386),
.B2(n_377),
.Y(n_500)
);

BUFx4f_ASAP7_75t_SL g501 ( 
.A(n_446),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_446),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_434),
.B(n_386),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_426),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_455),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_456),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_456),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_420),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_425),
.B(n_375),
.Y(n_509)
);

CKINVDCx11_ASAP7_75t_R g510 ( 
.A(n_445),
.Y(n_510)
);

BUFx8_ASAP7_75t_L g511 ( 
.A(n_446),
.Y(n_511)
);

NAND2x1_ASAP7_75t_L g512 ( 
.A(n_426),
.B(n_394),
.Y(n_512)
);

BUFx2_ASAP7_75t_SL g513 ( 
.A(n_446),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_444),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_461),
.Y(n_515)
);

NAND2x1p5_ASAP7_75t_L g516 ( 
.A(n_430),
.B(n_401),
.Y(n_516)
);

CKINVDCx8_ASAP7_75t_R g517 ( 
.A(n_466),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_461),
.Y(n_518)
);

BUFx5_ASAP7_75t_L g519 ( 
.A(n_438),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_471),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_471),
.Y(n_521)
);

CKINVDCx6p67_ASAP7_75t_R g522 ( 
.A(n_480),
.Y(n_522)
);

CKINVDCx11_ASAP7_75t_R g523 ( 
.A(n_480),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_479),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_488),
.A2(n_466),
.B1(n_452),
.B2(n_386),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_517),
.A2(n_465),
.B1(n_455),
.B2(n_435),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_509),
.A2(n_466),
.B1(n_464),
.B2(n_459),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_517),
.A2(n_465),
.B1(n_473),
.B2(n_451),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_503),
.A2(n_439),
.B(n_440),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_492),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_508),
.Y(n_531)
);

INVx4_ASAP7_75t_L g532 ( 
.A(n_489),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_475),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_SL g534 ( 
.A1(n_496),
.A2(n_424),
.B1(n_436),
.B2(n_470),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_477),
.Y(n_535)
);

CKINVDCx11_ASAP7_75t_R g536 ( 
.A(n_487),
.Y(n_536)
);

BUFx2_ASAP7_75t_SL g537 ( 
.A(n_478),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_478),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_487),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_482),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_484),
.A2(n_377),
.B1(n_464),
.B2(n_453),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_491),
.A2(n_445),
.B1(n_453),
.B2(n_454),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_490),
.Y(n_543)
);

OAI22xp33_ASAP7_75t_L g544 ( 
.A1(n_496),
.A2(n_405),
.B1(n_457),
.B2(n_465),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_SL g545 ( 
.A1(n_500),
.A2(n_368),
.B(n_405),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_SL g546 ( 
.A1(n_496),
.A2(n_453),
.B1(n_377),
.B2(n_460),
.Y(n_546)
);

BUFx2_ASAP7_75t_SL g547 ( 
.A(n_479),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_476),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_500),
.A2(n_463),
.B1(n_444),
.B2(n_448),
.Y(n_549)
);

INVx1_ASAP7_75t_SL g550 ( 
.A(n_508),
.Y(n_550)
);

INVx6_ASAP7_75t_L g551 ( 
.A(n_511),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_483),
.A2(n_382),
.B1(n_377),
.B2(n_365),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_489),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_476),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_SL g555 ( 
.A1(n_511),
.A2(n_377),
.B1(n_382),
.B2(n_438),
.Y(n_555)
);

CKINVDCx11_ASAP7_75t_R g556 ( 
.A(n_510),
.Y(n_556)
);

BUFx6f_ASAP7_75t_SL g557 ( 
.A(n_486),
.Y(n_557)
);

INVx4_ASAP7_75t_L g558 ( 
.A(n_489),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_SL g559 ( 
.A1(n_511),
.A2(n_501),
.B1(n_489),
.B2(n_377),
.Y(n_559)
);

BUFx12f_ASAP7_75t_L g560 ( 
.A(n_510),
.Y(n_560)
);

BUFx12f_ASAP7_75t_L g561 ( 
.A(n_479),
.Y(n_561)
);

BUFx10_ASAP7_75t_L g562 ( 
.A(n_479),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_483),
.Y(n_563)
);

OAI22xp33_ASAP7_75t_L g564 ( 
.A1(n_545),
.A2(n_535),
.B1(n_540),
.B2(n_544),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_542),
.A2(n_501),
.B1(n_483),
.B2(n_505),
.Y(n_565)
);

INVx4_ASAP7_75t_L g566 ( 
.A(n_561),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_543),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_534),
.A2(n_441),
.B1(n_483),
.B2(n_505),
.Y(n_568)
);

BUFx8_ASAP7_75t_SL g569 ( 
.A(n_548),
.Y(n_569)
);

OAI21xp33_ASAP7_75t_L g570 ( 
.A1(n_527),
.A2(n_398),
.B(n_407),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_534),
.A2(n_505),
.B1(n_407),
.B2(n_502),
.Y(n_571)
);

INVx4_ASAP7_75t_R g572 ( 
.A(n_554),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_525),
.A2(n_505),
.B1(n_519),
.B2(n_438),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_531),
.B(n_481),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_550),
.A2(n_519),
.B1(n_438),
.B2(n_432),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_529),
.A2(n_519),
.B1(n_438),
.B2(n_432),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_SL g577 ( 
.A1(n_546),
.A2(n_381),
.B(n_493),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_SL g578 ( 
.A1(n_551),
.A2(n_519),
.B1(n_513),
.B2(n_485),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_530),
.B(n_423),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_533),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_538),
.B(n_481),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_SL g582 ( 
.A1(n_551),
.A2(n_519),
.B1(n_485),
.B2(n_493),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_544),
.A2(n_519),
.B1(n_481),
.B2(n_389),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_546),
.A2(n_519),
.B1(n_516),
.B2(n_363),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g585 ( 
.A1(n_541),
.A2(n_516),
.B1(n_448),
.B2(n_447),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_541),
.A2(n_448),
.B1(n_447),
.B2(n_444),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_530),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_552),
.A2(n_447),
.B1(n_428),
.B2(n_485),
.Y(n_588)
);

AOI222xp33_ASAP7_75t_L g589 ( 
.A1(n_560),
.A2(n_521),
.B1(n_494),
.B2(n_518),
.C1(n_515),
.C2(n_497),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_562),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_523),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_557),
.A2(n_481),
.B1(n_390),
.B2(n_408),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_524),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_524),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_524),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_563),
.B(n_507),
.Y(n_596)
);

BUFx8_ASAP7_75t_SL g597 ( 
.A(n_539),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_551),
.A2(n_520),
.B1(n_498),
.B2(n_475),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_562),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_536),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_L g601 ( 
.A1(n_555),
.A2(n_428),
.B1(n_485),
.B2(n_427),
.Y(n_601)
);

OAI21xp5_ASAP7_75t_SL g602 ( 
.A1(n_555),
.A2(n_374),
.B(n_376),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_557),
.A2(n_410),
.B1(n_389),
.B2(n_390),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_547),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_549),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g606 ( 
.A(n_537),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_SL g607 ( 
.A1(n_559),
.A2(n_400),
.B(n_419),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_532),
.B(n_504),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_526),
.B(n_495),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_559),
.A2(n_528),
.B1(n_522),
.B2(n_553),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_564),
.A2(n_556),
.B1(n_410),
.B2(n_408),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_564),
.A2(n_396),
.B1(n_395),
.B2(n_418),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_568),
.A2(n_558),
.B1(n_553),
.B2(n_532),
.Y(n_613)
);

NAND3xp33_ASAP7_75t_L g614 ( 
.A(n_589),
.B(n_414),
.C(n_404),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_568),
.A2(n_558),
.B1(n_499),
.B2(n_512),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_570),
.A2(n_514),
.B1(n_504),
.B2(n_401),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_571),
.A2(n_573),
.B1(n_605),
.B2(n_610),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_567),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_575),
.A2(n_514),
.B1(n_504),
.B2(n_401),
.Y(n_619)
);

NOR3xp33_ASAP7_75t_L g620 ( 
.A(n_565),
.B(n_383),
.C(n_391),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_574),
.A2(n_514),
.B1(n_401),
.B2(n_499),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_580),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_583),
.A2(n_469),
.B1(n_394),
.B2(n_498),
.Y(n_623)
);

AOI21xp33_ASAP7_75t_L g624 ( 
.A1(n_607),
.A2(n_520),
.B(n_506),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_SL g625 ( 
.A1(n_596),
.A2(n_469),
.B1(n_506),
.B2(n_495),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_SL g626 ( 
.A1(n_588),
.A2(n_601),
.B1(n_606),
.B2(n_566),
.Y(n_626)
);

OAI221xp5_ASAP7_75t_L g627 ( 
.A1(n_603),
.A2(n_469),
.B1(n_393),
.B2(n_369),
.C(n_372),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_L g628 ( 
.A1(n_592),
.A2(n_469),
.B1(n_372),
.B2(n_369),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_576),
.A2(n_472),
.B1(n_458),
.B2(n_387),
.Y(n_629)
);

OAI222xp33_ASAP7_75t_L g630 ( 
.A1(n_582),
.A2(n_472),
.B1(n_15),
.B2(n_16),
.C1(n_17),
.C2(n_18),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_SL g631 ( 
.A1(n_600),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_609),
.Y(n_632)
);

OAI221xp5_ASAP7_75t_SL g633 ( 
.A1(n_602),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.C(n_21),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_587),
.A2(n_409),
.B1(n_474),
.B2(n_421),
.Y(n_634)
);

NOR3xp33_ASAP7_75t_L g635 ( 
.A(n_606),
.B(n_416),
.C(n_415),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_SL g636 ( 
.A1(n_591),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_582),
.A2(n_409),
.B1(n_421),
.B2(n_468),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_584),
.A2(n_409),
.B1(n_421),
.B2(n_468),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_566),
.A2(n_604),
.B1(n_578),
.B2(n_599),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_578),
.A2(n_409),
.B1(n_417),
.B2(n_218),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_598),
.A2(n_22),
.B1(n_409),
.B2(n_38),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_SL g642 ( 
.A1(n_585),
.A2(n_22),
.B1(n_409),
.B2(n_39),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_581),
.A2(n_579),
.B1(n_598),
.B2(n_594),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_581),
.A2(n_409),
.B1(n_40),
.B2(n_41),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_595),
.A2(n_409),
.B1(n_42),
.B2(n_43),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_SL g646 ( 
.A1(n_590),
.A2(n_593),
.B1(n_608),
.B2(n_572),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_618),
.B(n_632),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_L g648 ( 
.A1(n_633),
.A2(n_577),
.B1(n_590),
.B2(n_608),
.Y(n_648)
);

NAND3xp33_ASAP7_75t_L g649 ( 
.A(n_611),
.B(n_593),
.C(n_586),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_631),
.A2(n_569),
.B1(n_597),
.B2(n_45),
.Y(n_650)
);

OAI21xp33_ASAP7_75t_L g651 ( 
.A1(n_617),
.A2(n_37),
.B(n_44),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_632),
.B(n_51),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_618),
.B(n_145),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_622),
.B(n_55),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_622),
.B(n_56),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_SL g656 ( 
.A1(n_636),
.A2(n_57),
.B1(n_58),
.B2(n_63),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_642),
.A2(n_612),
.B1(n_641),
.B2(n_614),
.Y(n_657)
);

OAI21xp33_ASAP7_75t_L g658 ( 
.A1(n_626),
.A2(n_66),
.B(n_69),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_625),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_639),
.B(n_75),
.Y(n_660)
);

OAI221xp5_ASAP7_75t_SL g661 ( 
.A1(n_612),
.A2(n_77),
.B1(n_79),
.B2(n_80),
.C(n_81),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_643),
.B(n_82),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_646),
.B(n_83),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_616),
.B(n_84),
.Y(n_664)
);

AOI221xp5_ASAP7_75t_L g665 ( 
.A1(n_630),
.A2(n_87),
.B1(n_90),
.B2(n_92),
.C(n_93),
.Y(n_665)
);

AOI221xp5_ASAP7_75t_L g666 ( 
.A1(n_624),
.A2(n_94),
.B1(n_95),
.B2(n_97),
.C(n_98),
.Y(n_666)
);

OAI22xp5_ASAP7_75t_L g667 ( 
.A1(n_644),
.A2(n_623),
.B1(n_645),
.B2(n_619),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_621),
.B(n_100),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_615),
.Y(n_669)
);

NAND3xp33_ASAP7_75t_L g670 ( 
.A(n_635),
.B(n_102),
.C(n_103),
.Y(n_670)
);

NAND3xp33_ASAP7_75t_L g671 ( 
.A(n_634),
.B(n_104),
.C(n_105),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_613),
.B(n_106),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_628),
.B(n_107),
.Y(n_673)
);

NAND4xp25_ASAP7_75t_SL g674 ( 
.A(n_638),
.B(n_109),
.C(n_110),
.D(n_111),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_SL g675 ( 
.A1(n_667),
.A2(n_627),
.B1(n_637),
.B2(n_640),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_647),
.B(n_620),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_647),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_669),
.B(n_629),
.Y(n_678)
);

OAI211xp5_ASAP7_75t_L g679 ( 
.A1(n_650),
.A2(n_112),
.B(n_113),
.C(n_114),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_653),
.B(n_115),
.Y(n_680)
);

NAND3xp33_ASAP7_75t_L g681 ( 
.A(n_657),
.B(n_665),
.C(n_661),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_654),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_652),
.B(n_117),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_655),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_673),
.B(n_118),
.Y(n_685)
);

NAND4xp75_ASAP7_75t_L g686 ( 
.A(n_672),
.B(n_673),
.C(n_660),
.D(n_663),
.Y(n_686)
);

AO21x2_ASAP7_75t_L g687 ( 
.A1(n_672),
.A2(n_670),
.B(n_662),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_648),
.B(n_119),
.Y(n_688)
);

NOR3xp33_ASAP7_75t_SL g689 ( 
.A(n_674),
.B(n_658),
.C(n_659),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_657),
.B(n_120),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_649),
.Y(n_691)
);

XOR2x2_ASAP7_75t_L g692 ( 
.A(n_686),
.B(n_650),
.Y(n_692)
);

HB1xp67_ASAP7_75t_L g693 ( 
.A(n_677),
.Y(n_693)
);

NAND4xp25_ASAP7_75t_SL g694 ( 
.A(n_681),
.B(n_656),
.C(n_666),
.D(n_671),
.Y(n_694)
);

NOR3xp33_ASAP7_75t_L g695 ( 
.A(n_686),
.B(n_679),
.C(n_691),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_677),
.B(n_668),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_676),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_676),
.Y(n_698)
);

HB1xp67_ASAP7_75t_L g699 ( 
.A(n_684),
.Y(n_699)
);

INVxp67_ASAP7_75t_L g700 ( 
.A(n_691),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_684),
.Y(n_701)
);

INVxp67_ASAP7_75t_L g702 ( 
.A(n_699),
.Y(n_702)
);

INVxp67_ASAP7_75t_L g703 ( 
.A(n_697),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_698),
.B(n_682),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_698),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_701),
.Y(n_706)
);

XOR2x2_ASAP7_75t_L g707 ( 
.A(n_704),
.B(n_692),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_705),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_706),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_705),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_705),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_709),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_709),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_708),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_710),
.Y(n_715)
);

OA22x2_ASAP7_75t_L g716 ( 
.A1(n_714),
.A2(n_700),
.B1(n_698),
.B2(n_702),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_712),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_713),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_716),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_717),
.A2(n_695),
.B1(n_692),
.B2(n_707),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_718),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_717),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_721),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_720),
.B(n_715),
.Y(n_724)
);

NOR4xp25_ASAP7_75t_L g725 ( 
.A(n_722),
.B(n_694),
.C(n_690),
.D(n_688),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_719),
.B(n_711),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_721),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_719),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_719),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_728),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_729),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_728),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_726),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_723),
.Y(n_734)
);

OR2x2_ASAP7_75t_L g735 ( 
.A(n_725),
.B(n_703),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_727),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_724),
.B(n_704),
.Y(n_737)
);

NOR4xp75_ASAP7_75t_L g738 ( 
.A(n_737),
.B(n_690),
.C(n_688),
.D(n_651),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_731),
.A2(n_689),
.B1(n_675),
.B2(n_693),
.Y(n_739)
);

HB1xp67_ASAP7_75t_L g740 ( 
.A(n_730),
.Y(n_740)
);

OA22x2_ASAP7_75t_L g741 ( 
.A1(n_732),
.A2(n_685),
.B1(n_696),
.B2(n_680),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_731),
.Y(n_742)
);

NOR4xp25_ASAP7_75t_L g743 ( 
.A(n_733),
.B(n_685),
.C(n_683),
.D(n_680),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_L g744 ( 
.A1(n_735),
.A2(n_696),
.B1(n_682),
.B2(n_683),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_734),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_740),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_SL g747 ( 
.A1(n_739),
.A2(n_736),
.B1(n_687),
.B2(n_664),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_742),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_741),
.Y(n_749)
);

HB1xp67_ASAP7_75t_L g750 ( 
.A(n_745),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_744),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_738),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_743),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_746),
.Y(n_754)
);

AO22x2_ASAP7_75t_L g755 ( 
.A1(n_749),
.A2(n_678),
.B1(n_687),
.B2(n_123),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_752),
.A2(n_751),
.B1(n_748),
.B2(n_753),
.Y(n_756)
);

INVx3_ASAP7_75t_L g757 ( 
.A(n_750),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_747),
.A2(n_687),
.B1(n_678),
.B2(n_126),
.Y(n_758)
);

OAI211xp5_ASAP7_75t_L g759 ( 
.A1(n_747),
.A2(n_121),
.B(n_122),
.C(n_127),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_757),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_754),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_756),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_755),
.Y(n_763)
);

AO22x2_ASAP7_75t_L g764 ( 
.A1(n_763),
.A2(n_760),
.B1(n_762),
.B2(n_761),
.Y(n_764)
);

OAI22xp5_ASAP7_75t_SL g765 ( 
.A1(n_762),
.A2(n_758),
.B1(n_759),
.B2(n_130),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_764),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_765),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_766),
.A2(n_128),
.B1(n_129),
.B2(n_131),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_768),
.Y(n_769)
);

AOI221xp5_ASAP7_75t_L g770 ( 
.A1(n_769),
.A2(n_767),
.B1(n_134),
.B2(n_135),
.C(n_138),
.Y(n_770)
);

AOI211xp5_ASAP7_75t_L g771 ( 
.A1(n_770),
.A2(n_133),
.B(n_139),
.C(n_142),
.Y(n_771)
);


endmodule