module real_aes_4790_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_560;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_656;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_449;
wire n_363;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_646;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g282 ( .A(n_0), .Y(n_282) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_1), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_1), .B(n_297), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_2), .B(n_417), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_3), .A2(n_28), .B1(n_296), .B2(n_361), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g336 ( .A1(n_4), .A2(n_32), .B1(n_271), .B2(n_337), .Y(n_336) );
AOI22xp5_ASAP7_75t_L g261 ( .A1(n_5), .A2(n_51), .B1(n_245), .B2(n_248), .Y(n_261) );
INVx1_ASAP7_75t_L g277 ( .A(n_6), .Y(n_277) );
INVx1_ASAP7_75t_L g109 ( .A(n_7), .Y(n_109) );
INVxp67_ASAP7_75t_L g125 ( .A(n_7), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_7), .B(n_58), .Y(n_148) );
INVx1_ASAP7_75t_L g187 ( .A(n_8), .Y(n_187) );
INVx1_ASAP7_75t_L g280 ( .A(n_9), .Y(n_280) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_10), .A2(n_55), .B(n_241), .Y(n_240) );
OA21x2_ASAP7_75t_L g256 ( .A1(n_10), .A2(n_55), .B(n_241), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g105 ( .A(n_11), .B(n_93), .Y(n_105) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_12), .A2(n_83), .B1(n_84), .B2(n_651), .Y(n_650) );
CKINVDCx20_ASAP7_75t_R g651 ( .A(n_12), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_13), .A2(n_53), .B1(n_245), .B2(n_248), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g112 ( .A1(n_14), .A2(n_74), .B1(n_113), .B2(n_117), .Y(n_112) );
INVx1_ASAP7_75t_L g270 ( .A(n_15), .Y(n_270) );
BUFx3_ASAP7_75t_L g202 ( .A(n_16), .Y(n_202) );
INVx1_ASAP7_75t_L g142 ( .A(n_17), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_18), .Y(n_196) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_19), .Y(n_93) );
AO22x1_ASAP7_75t_L g410 ( .A1(n_20), .A2(n_61), .B1(n_283), .B2(n_411), .Y(n_410) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_21), .Y(n_300) );
AND2x2_ASAP7_75t_L g314 ( .A(n_22), .B(n_271), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_23), .B(n_283), .Y(n_306) );
AOI22xp5_ASAP7_75t_L g153 ( .A1(n_24), .A2(n_75), .B1(n_154), .B2(n_160), .Y(n_153) );
AOI22x1_ASAP7_75t_L g343 ( .A1(n_25), .A2(n_71), .B1(n_245), .B2(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g97 ( .A(n_26), .Y(n_97) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_26), .B(n_57), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_27), .B(n_346), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g87 ( .A(n_29), .B(n_88), .Y(n_87) );
AOI22xp33_ASAP7_75t_L g127 ( .A1(n_30), .A2(n_37), .B1(n_128), .B2(n_130), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g322 ( .A(n_31), .B(n_323), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_33), .Y(n_82) );
AOI21xp33_ASAP7_75t_L g138 ( .A1(n_34), .A2(n_139), .B(n_141), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_35), .B(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_36), .B(n_275), .Y(n_305) );
INVx1_ASAP7_75t_L g241 ( .A(n_38), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g163 ( .A1(n_39), .A2(n_46), .B1(n_164), .B2(n_169), .Y(n_163) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_40), .Y(n_213) );
AND2x4_ASAP7_75t_L g216 ( .A(n_40), .B(n_211), .Y(n_216) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_41), .Y(n_221) );
INVx2_ASAP7_75t_L g252 ( .A(n_42), .Y(n_252) );
AOI22xp33_ASAP7_75t_SL g178 ( .A1(n_43), .A2(n_72), .B1(n_179), .B2(n_181), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_44), .A2(n_73), .B1(n_172), .B2(n_176), .Y(n_171) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_45), .A2(n_59), .B1(n_296), .B2(n_344), .Y(n_357) );
AND2x2_ASAP7_75t_L g320 ( .A(n_47), .B(n_283), .Y(n_320) );
CKINVDCx14_ASAP7_75t_R g419 ( .A(n_48), .Y(n_419) );
OA22x2_ASAP7_75t_L g91 ( .A1(n_49), .A2(n_58), .B1(n_92), .B2(n_93), .Y(n_91) );
INVx1_ASAP7_75t_L g136 ( .A(n_49), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_50), .B(n_382), .Y(n_381) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_51), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_52), .B(n_373), .Y(n_372) );
NAND2x1p5_ASAP7_75t_L g324 ( .A(n_54), .B(n_254), .Y(n_324) );
CKINVDCx14_ASAP7_75t_R g349 ( .A(n_56), .Y(n_349) );
INVx1_ASAP7_75t_L g111 ( .A(n_57), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_57), .B(n_134), .Y(n_151) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_57), .Y(n_205) );
OAI21xp33_ASAP7_75t_L g137 ( .A1(n_58), .A2(n_62), .B(n_126), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_60), .B(n_297), .Y(n_377) );
INVx1_ASAP7_75t_L g99 ( .A(n_62), .Y(n_99) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_62), .B(n_70), .Y(n_149) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_63), .Y(n_225) );
BUFx5_ASAP7_75t_L g247 ( .A(n_63), .Y(n_247) );
INVx1_ASAP7_75t_L g340 ( .A(n_63), .Y(n_340) );
INVx2_ASAP7_75t_L g285 ( .A(n_64), .Y(n_285) );
NAND2xp33_ASAP7_75t_L g316 ( .A(n_65), .B(n_317), .Y(n_316) );
INVx2_ASAP7_75t_SL g211 ( .A(n_66), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_67), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_68), .B(n_323), .Y(n_376) );
HB1xp67_ASAP7_75t_L g186 ( .A(n_69), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_70), .B(n_104), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_76), .B(n_311), .Y(n_310) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_197), .B1(n_214), .B2(n_226), .C(n_644), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_183), .Y(n_78) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_80), .A2(n_81), .B1(n_83), .B2(n_84), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
XNOR2xp5_ASAP7_75t_L g645 ( .A(n_83), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
INVxp33_ASAP7_75t_SL g84 ( .A(n_85), .Y(n_84) );
NOR2x1_ASAP7_75t_L g85 ( .A(n_86), .B(n_152), .Y(n_85) );
NAND4xp25_ASAP7_75t_L g86 ( .A(n_87), .B(n_112), .C(n_127), .D(n_138), .Y(n_86) );
BUFx8_ASAP7_75t_SL g88 ( .A(n_89), .Y(n_88) );
AND2x4_ASAP7_75t_L g89 ( .A(n_90), .B(n_100), .Y(n_89) );
AND2x4_ASAP7_75t_L g129 ( .A(n_90), .B(n_115), .Y(n_129) );
AND2x2_ASAP7_75t_L g90 ( .A(n_91), .B(n_94), .Y(n_90) );
AND2x2_ASAP7_75t_L g116 ( .A(n_91), .B(n_95), .Y(n_116) );
AND2x2_ASAP7_75t_L g123 ( .A(n_91), .B(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g175 ( .A(n_91), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g98 ( .A(n_92), .B(n_99), .Y(n_98) );
INVx2_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
NAND2xp33_ASAP7_75t_L g96 ( .A(n_93), .B(n_97), .Y(n_96) );
INVx3_ASAP7_75t_L g104 ( .A(n_93), .Y(n_104) );
NAND2xp33_ASAP7_75t_L g110 ( .A(n_93), .B(n_111), .Y(n_110) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_93), .Y(n_121) );
INVx1_ASAP7_75t_L g126 ( .A(n_93), .Y(n_126) );
AND2x4_ASAP7_75t_L g174 ( .A(n_94), .B(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
NAND2xp5_ASAP7_75t_L g95 ( .A(n_96), .B(n_98), .Y(n_95) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_97), .B(n_136), .Y(n_135) );
INVxp67_ASAP7_75t_L g206 ( .A(n_97), .Y(n_206) );
OAI21xp5_ASAP7_75t_L g124 ( .A1(n_99), .A2(n_125), .B(n_126), .Y(n_124) );
AND2x4_ASAP7_75t_L g131 ( .A(n_100), .B(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g140 ( .A(n_100), .B(n_116), .Y(n_140) );
AND2x2_ASAP7_75t_L g180 ( .A(n_100), .B(n_174), .Y(n_180) );
AND2x4_ASAP7_75t_L g100 ( .A(n_101), .B(n_106), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x4_ASAP7_75t_L g115 ( .A(n_102), .B(n_106), .Y(n_115) );
AND2x2_ASAP7_75t_L g119 ( .A(n_102), .B(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g158 ( .A(n_102), .B(n_159), .Y(n_158) );
AND2x4_ASAP7_75t_L g167 ( .A(n_102), .B(n_168), .Y(n_167) );
AND2x4_ASAP7_75t_L g102 ( .A(n_103), .B(n_105), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_104), .B(n_109), .Y(n_108) );
INVxp67_ASAP7_75t_L g134 ( .A(n_104), .Y(n_134) );
NAND3xp33_ASAP7_75t_L g150 ( .A(n_105), .B(n_133), .C(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g159 ( .A(n_107), .Y(n_159) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
AND2x4_ASAP7_75t_L g182 ( .A(n_115), .B(n_174), .Y(n_182) );
AND2x4_ASAP7_75t_L g161 ( .A(n_116), .B(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_L g170 ( .A(n_116), .B(n_167), .Y(n_170) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x4_ASAP7_75t_L g118 ( .A(n_119), .B(n_123), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
INVx1_ASAP7_75t_L g146 ( .A(n_121), .Y(n_146) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_122), .Y(n_203) );
BUFx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x4_ASAP7_75t_L g156 ( .A(n_132), .B(n_157), .Y(n_156) );
AND2x4_ASAP7_75t_L g166 ( .A(n_132), .B(n_167), .Y(n_166) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_137), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_136), .Y(n_207) );
BUFx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AO21x2_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_150), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
NAND4xp25_ASAP7_75t_L g152 ( .A(n_153), .B(n_163), .C(n_171), .D(n_178), .Y(n_152) );
INVx5_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx6_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x4_ASAP7_75t_L g173 ( .A(n_157), .B(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g162 ( .A(n_158), .Y(n_162) );
INVx1_ASAP7_75t_L g168 ( .A(n_159), .Y(n_168) );
BUFx12f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx8_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AND2x4_ASAP7_75t_L g177 ( .A(n_167), .B(n_174), .Y(n_177) );
BUFx4f_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
BUFx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
BUFx12f_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
OAI22xp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B1(n_190), .B2(n_191), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_185), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B1(n_188), .B2(n_189), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_186), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_187), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_191), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B1(n_194), .B2(n_195), .Y(n_191) );
CKINVDCx16_ASAP7_75t_R g192 ( .A(n_193), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_195), .Y(n_194) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
BUFx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_200), .B(n_208), .Y(n_199) );
INVxp67_ASAP7_75t_SL g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g649 ( .A(n_201), .B(n_208), .Y(n_649) );
AOI211xp5_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_203), .B(n_204), .C(n_207), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_209), .B(n_212), .Y(n_208) );
OR2x2_ASAP7_75t_L g653 ( .A(n_209), .B(n_213), .Y(n_653) );
INVx1_ASAP7_75t_L g656 ( .A(n_209), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_209), .B(n_212), .Y(n_657) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_217), .Y(n_214) );
OAI21x1_ASAP7_75t_L g294 ( .A1(n_215), .A2(n_295), .B(n_304), .Y(n_294) );
AO31x2_ASAP7_75t_L g334 ( .A1(n_215), .A2(n_335), .A3(n_345), .B(n_348), .Y(n_334) );
AO31x2_ASAP7_75t_L g389 ( .A1(n_215), .A2(n_335), .A3(n_345), .B(n_348), .Y(n_389) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx3_ASAP7_75t_L g243 ( .A(n_216), .Y(n_243) );
INVx1_ASAP7_75t_L g266 ( .A(n_216), .Y(n_266) );
INVx3_ASAP7_75t_L g356 ( .A(n_216), .Y(n_356) );
OA21x2_ASAP7_75t_L g655 ( .A1(n_217), .A2(n_656), .B(n_657), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_218), .B(n_222), .Y(n_217) );
HB1xp67_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_219), .B(n_299), .Y(n_298) );
OAI22x1_ASAP7_75t_L g335 ( .A1(n_219), .A2(n_336), .B1(n_341), .B2(n_343), .Y(n_335) );
INVx4_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g295 ( .A1(n_220), .A2(n_296), .B1(n_298), .B2(n_301), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_220), .B(n_355), .Y(n_354) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_220), .A2(n_376), .B(n_377), .Y(n_375) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx4_ASAP7_75t_L g238 ( .A(n_221), .Y(n_238) );
INVx3_ASAP7_75t_L g260 ( .A(n_221), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_221), .B(n_270), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_221), .B(n_277), .Y(n_276) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_221), .Y(n_308) );
INVxp67_ASAP7_75t_L g318 ( .A(n_221), .Y(n_318) );
INVx1_ASAP7_75t_L g342 ( .A(n_221), .Y(n_342) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g275 ( .A(n_224), .Y(n_275) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx3_ASAP7_75t_L g250 ( .A(n_225), .Y(n_250) );
INVx6_ASAP7_75t_L g273 ( .A(n_225), .Y(n_273) );
INVx2_ASAP7_75t_L g303 ( .A(n_225), .Y(n_303) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NAND2x1p5_ASAP7_75t_L g229 ( .A(n_230), .B(n_518), .Y(n_229) );
NOR4xp75_ASAP7_75t_L g230 ( .A(n_231), .B(n_431), .C(n_449), .D(n_475), .Y(n_230) );
AO21x1_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_287), .B(n_395), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_234), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g439 ( .A(n_234), .B(n_405), .Y(n_439) );
INVx2_ASAP7_75t_L g501 ( .A(n_234), .Y(n_501) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_262), .Y(n_234) );
INVx1_ASAP7_75t_L g366 ( .A(n_235), .Y(n_366) );
INVx1_ASAP7_75t_L g394 ( .A(n_235), .Y(n_394) );
AND2x2_ASAP7_75t_L g421 ( .A(n_235), .B(n_263), .Y(n_421) );
INVx1_ASAP7_75t_L g452 ( .A(n_235), .Y(n_452) );
INVx2_ASAP7_75t_L g484 ( .A(n_235), .Y(n_484) );
NOR2x1_ASAP7_75t_L g526 ( .A(n_235), .B(n_527), .Y(n_526) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_235), .Y(n_541) );
AND2x2_ASAP7_75t_L g590 ( .A(n_235), .B(n_370), .Y(n_590) );
OR2x6_ASAP7_75t_L g235 ( .A(n_236), .B(n_257), .Y(n_235) );
OAI21x1_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_244), .B(n_251), .Y(n_236) );
NAND3xp33_ASAP7_75t_SL g237 ( .A(n_238), .B(n_239), .C(n_242), .Y(n_237) );
NOR2xp33_ASAP7_75t_SL g279 ( .A(n_238), .B(n_280), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_238), .B(n_282), .Y(n_281) );
NAND3xp33_ASAP7_75t_L g258 ( .A(n_239), .B(n_242), .C(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g265 ( .A(n_239), .Y(n_265) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g347 ( .A(n_240), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_240), .B(n_356), .Y(n_355) );
AOI21xp33_ASAP7_75t_SL g327 ( .A1(n_242), .A2(n_328), .B(n_330), .Y(n_327) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NOR2x1_ASAP7_75t_L g384 ( .A(n_243), .B(n_373), .Y(n_384) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g283 ( .A(n_247), .Y(n_283) );
INVx2_ASAP7_75t_L g297 ( .A(n_247), .Y(n_297) );
INVx2_ASAP7_75t_L g382 ( .A(n_247), .Y(n_382) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g361 ( .A(n_249), .Y(n_361) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g380 ( .A(n_250), .Y(n_380) );
INVx1_ASAP7_75t_L g417 ( .A(n_250), .Y(n_417) );
OR2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
INVx1_ASAP7_75t_L g311 ( .A(n_253), .Y(n_311) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx3_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g329 ( .A(n_255), .Y(n_329) );
INVx4_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g286 ( .A(n_256), .Y(n_286) );
BUFx3_ASAP7_75t_L g309 ( .A(n_256), .Y(n_309) );
NOR2xp67_ASAP7_75t_L g257 ( .A(n_258), .B(n_261), .Y(n_257) );
INVx3_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g483 ( .A(n_262), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g488 ( .A(n_263), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g508 ( .A(n_263), .Y(n_508) );
INVx1_ASAP7_75t_L g527 ( .A(n_263), .Y(n_527) );
AND2x2_ASAP7_75t_L g589 ( .A(n_263), .B(n_454), .Y(n_589) );
INVxp67_ASAP7_75t_L g619 ( .A(n_263), .Y(n_619) );
AO21x2_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_267), .B(n_284), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
OR2x2_ASAP7_75t_L g407 ( .A(n_266), .B(n_311), .Y(n_407) );
NAND3xp33_ASAP7_75t_SL g267 ( .A(n_268), .B(n_274), .C(n_278), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g317 ( .A(n_273), .Y(n_317) );
INVx1_ASAP7_75t_L g323 ( .A(n_273), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g278 ( .A1(n_275), .A2(n_279), .B1(n_281), .B2(n_283), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx3_ASAP7_75t_L g373 ( .A(n_286), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_363), .B1(n_385), .B2(n_392), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x4_ASAP7_75t_L g289 ( .A(n_290), .B(n_331), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g560 ( .A(n_291), .Y(n_560) );
OR2x2_ASAP7_75t_L g642 ( .A(n_291), .B(n_474), .Y(n_642) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g473 ( .A(n_292), .B(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_312), .Y(n_292) );
AND2x2_ASAP7_75t_L g386 ( .A(n_293), .B(n_387), .Y(n_386) );
NAND2x1_ASAP7_75t_L g435 ( .A(n_293), .B(n_333), .Y(n_435) );
AND2x2_ASAP7_75t_L g570 ( .A(n_293), .B(n_352), .Y(n_570) );
OA21x2_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_309), .B(n_310), .Y(n_293) );
OA21x2_ASAP7_75t_L g401 ( .A1(n_294), .A2(n_309), .B(n_310), .Y(n_401) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_306), .B(n_307), .Y(n_304) );
INVxp67_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_SL g326 ( .A(n_308), .Y(n_326) );
INVx1_ASAP7_75t_L g383 ( .A(n_308), .Y(n_383) );
INVx1_ASAP7_75t_L g409 ( .A(n_308), .Y(n_409) );
INVx3_ASAP7_75t_L g350 ( .A(n_309), .Y(n_350) );
AND2x2_ASAP7_75t_L g396 ( .A(n_312), .B(n_389), .Y(n_396) );
AND2x4_ASAP7_75t_L g424 ( .A(n_312), .B(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g543 ( .A(n_312), .B(n_389), .Y(n_543) );
AO21x2_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_319), .B(n_327), .Y(n_312) );
AO21x2_ASAP7_75t_L g391 ( .A1(n_313), .A2(n_319), .B(n_327), .Y(n_391) );
OAI21x1_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_315), .B(n_318), .Y(n_313) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g344 ( .A(n_317), .Y(n_344) );
OAI21x1_ASAP7_75t_SL g319 ( .A1(n_320), .A2(n_321), .B(n_325), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_324), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g330 ( .A(n_324), .Y(n_330) );
AOI21x1_ASAP7_75t_L g414 ( .A1(n_326), .A2(n_415), .B(n_416), .Y(n_414) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_351), .Y(n_331) );
INVx2_ASAP7_75t_L g426 ( .A(n_332), .Y(n_426) );
INVx1_ASAP7_75t_L g458 ( .A(n_332), .Y(n_458) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g448 ( .A(n_333), .B(n_391), .Y(n_448) );
INVx1_ASAP7_75t_L g462 ( .A(n_333), .Y(n_462) );
AND2x2_ASAP7_75t_L g602 ( .A(n_333), .B(n_402), .Y(n_602) );
INVx3_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx3_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g413 ( .A(n_340), .Y(n_413) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_342), .B(n_355), .Y(n_359) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NOR2xp67_ASAP7_75t_SL g348 ( .A(n_349), .B(n_350), .Y(n_348) );
OR2x2_ASAP7_75t_L g418 ( .A(n_350), .B(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g474 ( .A(n_351), .Y(n_474) );
OR2x2_ASAP7_75t_L g586 ( .A(n_351), .B(n_435), .Y(n_586) );
INVx2_ASAP7_75t_L g594 ( .A(n_351), .Y(n_594) );
INVx2_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_358), .Y(n_352) );
NAND2x1p5_ASAP7_75t_L g387 ( .A(n_353), .B(n_358), .Y(n_387) );
OR2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_357), .Y(n_353) );
OA21x2_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_360), .B(n_362), .Y(n_358) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_367), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g509 ( .A(n_366), .B(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g534 ( .A(n_368), .B(n_494), .Y(n_534) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OR2x2_ASAP7_75t_L g468 ( .A(n_369), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g405 ( .A(n_370), .B(n_406), .Y(n_405) );
INVx3_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g430 ( .A(n_371), .Y(n_430) );
AND2x2_ASAP7_75t_L g453 ( .A(n_371), .B(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g465 ( .A(n_371), .B(n_406), .Y(n_465) );
AND2x4_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
OAI21x1_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_378), .B(n_384), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_381), .B(n_383), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_388), .Y(n_385) );
AND2x2_ASAP7_75t_L g490 ( .A(n_386), .B(n_434), .Y(n_490) );
INVx1_ASAP7_75t_L g603 ( .A(n_386), .Y(n_603) );
AND2x2_ASAP7_75t_L g635 ( .A(n_386), .B(n_462), .Y(n_635) );
INVx2_ASAP7_75t_L g402 ( .A(n_387), .Y(n_402) );
AND2x2_ASAP7_75t_L g445 ( .A(n_387), .B(n_400), .Y(n_445) );
INVx1_ASAP7_75t_L g495 ( .A(n_387), .Y(n_495) );
INVx1_ASAP7_75t_L g547 ( .A(n_387), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_387), .B(n_514), .Y(n_555) );
BUFx3_ASAP7_75t_L g442 ( .A(n_388), .Y(n_442) );
NOR2xp67_ASAP7_75t_L g562 ( .A(n_388), .B(n_444), .Y(n_562) );
AND2x4_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx1_ASAP7_75t_L g472 ( .A(n_389), .Y(n_472) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVxp67_ASAP7_75t_L g434 ( .A(n_391), .Y(n_434) );
INVx1_ASAP7_75t_L g514 ( .A(n_391), .Y(n_514) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g464 ( .A(n_393), .B(n_465), .Y(n_464) );
OR2x2_ASAP7_75t_L g467 ( .A(n_393), .B(n_468), .Y(n_467) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_393), .Y(n_496) );
OR2x2_ASAP7_75t_L g623 ( .A(n_393), .B(n_500), .Y(n_623) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g486 ( .A(n_394), .B(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_394), .B(n_552), .Y(n_551) );
OAI32xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .A3(n_403), .B1(n_422), .B2(n_427), .Y(n_395) );
INVx2_ASAP7_75t_L g558 ( .A(n_396), .Y(n_558) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g585 ( .A(n_398), .Y(n_585) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVxp67_ASAP7_75t_L g505 ( .A(n_399), .Y(n_505) );
OR2x2_ASAP7_75t_L g512 ( .A(n_399), .B(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_402), .Y(n_399) );
INVx1_ASAP7_75t_L g597 ( .A(n_400), .Y(n_597) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g425 ( .A(n_401), .Y(n_425) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_401), .Y(n_553) );
INVx1_ASAP7_75t_L g447 ( .A(n_402), .Y(n_447) );
INVx2_ASAP7_75t_L g437 ( .A(n_403), .Y(n_437) );
OR2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_420), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AND2x4_ASAP7_75t_L g525 ( .A(n_405), .B(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g612 ( .A(n_405), .B(n_483), .Y(n_612) );
INVx2_ASAP7_75t_SL g454 ( .A(n_406), .Y(n_454) );
OAI21x1_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_408), .B(n_418), .Y(n_406) );
OAI21xp5_ASAP7_75t_L g489 ( .A1(n_407), .A2(n_408), .B(n_418), .Y(n_489) );
AOI21x1_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B(n_414), .Y(n_408) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g561 ( .A(n_421), .B(n_465), .Y(n_561) );
NAND2x1_ASAP7_75t_SL g583 ( .A(n_421), .B(n_453), .Y(n_583) );
AND2x2_ASAP7_75t_L g592 ( .A(n_421), .B(n_481), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_421), .B(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g636 ( .A(n_423), .B(n_494), .Y(n_636) );
AND2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_426), .Y(n_423) );
AND2x4_ASAP7_75t_SL g461 ( .A(n_424), .B(n_462), .Y(n_461) );
BUFx3_ASAP7_75t_L g537 ( .A(n_424), .Y(n_537) );
INVxp67_ASAP7_75t_SL g530 ( .A(n_425), .Y(n_530) );
INVx1_ASAP7_75t_L g563 ( .A(n_427), .Y(n_563) );
AOI211xp5_ASAP7_75t_SL g550 ( .A1(n_428), .A2(n_462), .B(n_551), .C(n_553), .Y(n_550) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g507 ( .A(n_429), .B(n_508), .Y(n_507) );
OR2x2_ASAP7_75t_L g565 ( .A(n_429), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g632 ( .A(n_429), .B(n_483), .Y(n_632) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g516 ( .A(n_430), .B(n_452), .Y(n_516) );
OR2x2_ASAP7_75t_L g531 ( .A(n_430), .B(n_488), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_430), .B(n_619), .Y(n_618) );
OAI22xp5_ASAP7_75t_SL g431 ( .A1(n_432), .A2(n_436), .B1(n_438), .B2(n_440), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_435), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_434), .Y(n_529) );
AND3x2_ASAP7_75t_L g609 ( .A(n_434), .B(n_594), .C(n_597), .Y(n_609) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OA21x2_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_443), .B(n_446), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g628 ( .A(n_443), .Y(n_628) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g459 ( .A(n_445), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
BUFx3_ASAP7_75t_L g523 ( .A(n_448), .Y(n_523) );
AND2x2_ASAP7_75t_L g593 ( .A(n_448), .B(n_594), .Y(n_593) );
OAI21xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_455), .B(n_463), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
AND2x2_ASAP7_75t_L g573 ( .A(n_453), .B(n_483), .Y(n_573) );
INVx2_ASAP7_75t_L g581 ( .A(n_453), .Y(n_581) );
INVx1_ASAP7_75t_L g469 ( .A(n_454), .Y(n_469) );
INVx1_ASAP7_75t_L g498 ( .A(n_454), .Y(n_498) );
INVxp67_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_457), .B(n_460), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_457), .A2(n_478), .B1(n_493), .B2(n_499), .Y(n_492) );
OR2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
OR2x2_ASAP7_75t_L g568 ( .A(n_458), .B(n_569), .Y(n_568) );
INVx2_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g478 ( .A(n_461), .Y(n_478) );
OAI21xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_466), .B(n_470), .Y(n_463) );
INVx2_ASAP7_75t_L g500 ( .A(n_465), .Y(n_500) );
AND2x2_ASAP7_75t_L g545 ( .A(n_465), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g595 ( .A1(n_467), .A2(n_568), .B1(n_596), .B2(n_598), .Y(n_595) );
INVxp67_ASAP7_75t_SL g481 ( .A(n_469), .Y(n_481) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_473), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_471), .B(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_471), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NAND3x1_ASAP7_75t_L g475 ( .A(n_476), .B(n_491), .C(n_502), .Y(n_475) );
AOI21x1_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_479), .B(n_485), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_480), .A2(n_565), .B1(n_642), .B2(n_643), .Y(n_641) );
OR2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_490), .Y(n_485) );
INVx1_ASAP7_75t_L g535 ( .A(n_487), .Y(n_535) );
AND2x2_ASAP7_75t_L g615 ( .A(n_487), .B(n_541), .Y(n_615) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g517 ( .A(n_488), .Y(n_517) );
BUFx2_ASAP7_75t_L g510 ( .A(n_489), .Y(n_510) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NAND3xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_496), .C(n_497), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g549 ( .A(n_498), .B(n_508), .Y(n_549) );
OR2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
INVxp67_ASAP7_75t_L g539 ( .A(n_501), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_506), .B1(n_511), .B2(n_515), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NAND3xp33_ASAP7_75t_SL g557 ( .A(n_504), .B(n_558), .C(n_559), .Y(n_557) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_509), .Y(n_506) );
AND2x2_ASAP7_75t_L g617 ( .A(n_509), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_509), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g552 ( .A(n_510), .Y(n_552) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_513), .B(n_547), .Y(n_643) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_514), .A2(n_539), .B1(n_540), .B2(n_542), .Y(n_538) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
NAND2x2_ASAP7_75t_L g626 ( .A(n_516), .B(n_627), .Y(n_626) );
NOR2x1_ASAP7_75t_L g518 ( .A(n_519), .B(n_604), .Y(n_518) );
NAND4xp25_ASAP7_75t_L g519 ( .A(n_520), .B(n_556), .C(n_571), .D(n_591), .Y(n_519) );
NOR2xp67_ASAP7_75t_L g520 ( .A(n_521), .B(n_532), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_524), .B1(n_528), .B2(n_531), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AOI21xp33_ASAP7_75t_L g613 ( .A1(n_524), .A2(n_536), .B(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g566 ( .A(n_526), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
OAI211xp5_ASAP7_75t_SL g548 ( .A1(n_530), .A2(n_549), .B(n_550), .C(n_554), .Y(n_548) );
INVx1_ASAP7_75t_L g575 ( .A(n_530), .Y(n_575) );
AOI21xp33_ASAP7_75t_L g600 ( .A1(n_531), .A2(n_601), .B(n_603), .Y(n_600) );
OAI321xp33_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_535), .A3(n_536), .B1(n_538), .B2(n_544), .C(n_548), .Y(n_532) );
INVx2_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
OR2x2_ASAP7_75t_L g598 ( .A(n_535), .B(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_537), .B(n_578), .Y(n_577) );
NOR2x1_ASAP7_75t_R g620 ( .A(n_537), .B(n_601), .Y(n_620) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g621 ( .A(n_542), .B(n_570), .Y(n_621) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
OR2x2_ASAP7_75t_L g596 ( .A(n_543), .B(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g608 ( .A(n_543), .Y(n_608) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g578 ( .A(n_547), .Y(n_578) );
INVxp67_ASAP7_75t_L g634 ( .A(n_552), .Y(n_634) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AOI222xp33_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_561), .B1(n_562), .B2(n_563), .C1(n_564), .C2(n_567), .Y(n_556) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g625 ( .A(n_560), .Y(n_625) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g580 ( .A(n_566), .B(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AOI221x1_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_574), .B1(n_576), .B2(n_579), .C(n_582), .Y(n_571) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OAI22xp33_ASAP7_75t_SL g582 ( .A1(n_583), .A2(n_584), .B1(n_586), .B2(n_587), .Y(n_582) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x4_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
BUFx3_ASAP7_75t_L g627 ( .A(n_589), .Y(n_627) );
INVx2_ASAP7_75t_L g599 ( .A(n_590), .Y(n_599) );
AOI211xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_593), .B(n_595), .C(n_600), .Y(n_591) );
NAND2x1_ASAP7_75t_L g607 ( .A(n_594), .B(n_608), .Y(n_607) );
OAI22xp5_ASAP7_75t_SL g624 ( .A1(n_598), .A2(n_625), .B1(n_626), .B2(n_628), .Y(n_624) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND3xp33_ASAP7_75t_SL g604 ( .A(n_605), .B(n_616), .C(n_629), .Y(n_604) );
O2A1O1Ixp33_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_609), .B(n_610), .C(n_613), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AOI221xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_620), .B1(n_621), .B2(n_622), .C(n_624), .Y(n_616) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_619), .Y(n_640) );
INVxp67_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_635), .B1(n_636), .B2(n_637), .C(n_641), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVxp67_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI222xp33_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_646), .B1(n_648), .B2(n_650), .C1(n_652), .C2(n_654), .Y(n_644) );
CKINVDCx5p33_ASAP7_75t_R g646 ( .A(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
BUFx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
endmodule