module fake_jpeg_24321_n_307 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_307);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_307;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx4f_ASAP7_75t_SL g42 ( 
.A(n_26),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_42),
.Y(n_54)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_35),
.B1(n_32),
.B2(n_23),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_47),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_18),
.A2(n_0),
.B(n_1),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_48),
.B(n_37),
.C(n_21),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_18),
.B(n_19),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_57),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_23),
.B1(n_32),
.B2(n_35),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_55),
.A2(n_58),
.B1(n_65),
.B2(n_81),
.Y(n_111)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_23),
.B1(n_32),
.B2(n_35),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_42),
.B(n_46),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_48),
.C(n_27),
.Y(n_82)
);

NAND2x2_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_37),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_63),
.A2(n_67),
.B1(n_68),
.B2(n_72),
.Y(n_93)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_66),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_19),
.B1(n_22),
.B2(n_24),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_44),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_43),
.A2(n_19),
.B1(n_22),
.B2(n_24),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_22),
.B1(n_34),
.B2(n_24),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_40),
.A2(n_34),
.B1(n_25),
.B2(n_29),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_76),
.Y(n_97)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g102 ( 
.A(n_75),
.Y(n_102)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g103 ( 
.A(n_77),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_SL g78 ( 
.A(n_45),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

XNOR2x1_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_80),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_40),
.A2(n_34),
.B1(n_25),
.B2(n_29),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_47),
.A2(n_33),
.B1(n_31),
.B2(n_28),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_82),
.B(n_116),
.Y(n_129)
);

AO22x1_ASAP7_75t_SL g83 ( 
.A1(n_62),
.A2(n_37),
.B1(n_21),
.B2(n_45),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_83),
.A2(n_90),
.B1(n_99),
.B2(n_105),
.Y(n_125)
);

AOI32xp33_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_36),
.A3(n_30),
.B1(n_47),
.B2(n_37),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_85),
.B(n_41),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_21),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_95),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_63),
.B1(n_51),
.B2(n_33),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_21),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_113),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_18),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_98),
.B(n_111),
.C(n_88),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_63),
.A2(n_31),
.B1(n_36),
.B2(n_38),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_53),
.Y(n_100)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_57),
.B(n_18),
.Y(n_104)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_51),
.A2(n_38),
.B1(n_27),
.B2(n_30),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_3),
.B(n_5),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_50),
.B(n_0),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_109),
.B(n_110),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_30),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_18),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_112),
.B(n_114),
.Y(n_135)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_1),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_50),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_5),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_52),
.B(n_2),
.Y(n_116)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_119),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_94),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_120),
.Y(n_164)
);

OAI32xp33_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_54),
.A3(n_41),
.B1(n_59),
.B2(n_77),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_140),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_82),
.B(n_2),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_126),
.B(n_138),
.Y(n_153)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_131),
.Y(n_152)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_95),
.A2(n_54),
.B(n_59),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_132),
.A2(n_147),
.B(n_148),
.Y(n_182)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_134),
.Y(n_156)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_83),
.Y(n_134)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_137),
.A2(n_116),
.B(n_84),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_111),
.B(n_5),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_75),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_118),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_141),
.Y(n_165)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_144),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_143),
.A2(n_150),
.B1(n_129),
.B2(n_147),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_6),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_106),
.B(n_6),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_149),
.Y(n_163)
);

O2A1O1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_88),
.A2(n_41),
.B(n_8),
.C(n_9),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_41),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_96),
.B(n_7),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_118),
.C(n_103),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_154),
.A2(n_126),
.B(n_129),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_134),
.A2(n_93),
.B1(n_84),
.B2(n_116),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_155),
.A2(n_177),
.B1(n_157),
.B2(n_156),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_142),
.A2(n_102),
.B1(n_103),
.B2(n_108),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_158),
.A2(n_173),
.B1(n_179),
.B2(n_123),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_92),
.Y(n_160)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_92),
.Y(n_161)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_139),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_167),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_182),
.Y(n_185)
);

A2O1A1O1Ixp25_ASAP7_75t_L g169 ( 
.A1(n_137),
.A2(n_148),
.B(n_150),
.C(n_151),
.D(n_124),
.Y(n_169)
);

MAJx2_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_12),
.C(n_13),
.Y(n_201)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_170),
.B(n_172),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_108),
.Y(n_171)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_L g173 ( 
.A1(n_140),
.A2(n_118),
.B1(n_102),
.B2(n_87),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_135),
.B(n_7),
.Y(n_174)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_138),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_175),
.B(n_176),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_135),
.B(n_9),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_10),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_177),
.A2(n_180),
.B(n_122),
.Y(n_189)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_181),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_121),
.B(n_12),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_121),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_125),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_13),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_185),
.B(n_199),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_186),
.B(n_191),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_159),
.A2(n_125),
.B1(n_129),
.B2(n_122),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_187),
.A2(n_192),
.B1(n_197),
.B2(n_198),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_188),
.A2(n_201),
.B(n_209),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_180),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_165),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_159),
.A2(n_128),
.B1(n_120),
.B2(n_130),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_178),
.A2(n_182),
.B(n_156),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_193),
.A2(n_171),
.B(n_169),
.Y(n_227)
);

BUFx24_ASAP7_75t_SL g194 ( 
.A(n_181),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_202),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_183),
.A2(n_128),
.B1(n_131),
.B2(n_123),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_141),
.Y(n_199)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_203),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_155),
.A2(n_146),
.B1(n_91),
.B2(n_87),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_204),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_165),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_205),
.A2(n_191),
.B1(n_170),
.B2(n_172),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_154),
.A2(n_14),
.B(n_15),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_153),
.A2(n_14),
.B(n_15),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_210),
.A2(n_211),
.B(n_163),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_153),
.A2(n_15),
.B(n_16),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_206),
.B(n_175),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_213),
.Y(n_245)
);

NAND3xp33_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_174),
.C(n_176),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_215),
.B(n_218),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_216),
.A2(n_219),
.B(n_221),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_161),
.Y(n_217)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_217),
.Y(n_247)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_206),
.B(n_157),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_202),
.B(n_160),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_192),
.B(n_179),
.Y(n_225)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_225),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_226),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_227),
.A2(n_222),
.B(n_231),
.Y(n_248)
);

XOR2x1_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_209),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_184),
.B(n_164),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_197),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_199),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_234),
.A2(n_196),
.B1(n_186),
.B2(n_189),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_230),
.B(n_227),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_235),
.B(n_241),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_185),
.C(n_193),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_240),
.C(n_246),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_221),
.A2(n_214),
.B1(n_220),
.B2(n_232),
.Y(n_237)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_237),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_214),
.A2(n_187),
.B1(n_195),
.B2(n_184),
.Y(n_238)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_195),
.C(n_188),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_233),
.A2(n_225),
.B1(n_216),
.B2(n_217),
.Y(n_243)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_244),
.B(n_250),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_208),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_248),
.A2(n_213),
.B(n_229),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_223),
.A2(n_158),
.B1(n_190),
.B2(n_164),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_167),
.Y(n_253)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_253),
.Y(n_271)
);

NOR2xp67_ASAP7_75t_SL g254 ( 
.A(n_241),
.B(n_224),
.Y(n_254)
);

XNOR2x1_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_261),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_212),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_260),
.B(n_268),
.Y(n_273)
);

OAI21xp33_ASAP7_75t_L g261 ( 
.A1(n_252),
.A2(n_218),
.B(n_219),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_228),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_263),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_239),
.A2(n_162),
.B(n_166),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_265),
.A2(n_266),
.B(n_248),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_252),
.A2(n_211),
.B(n_210),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_162),
.C(n_166),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_235),
.C(n_246),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_212),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_255),
.A2(n_237),
.B1(n_245),
.B2(n_251),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_269),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_261),
.B(n_249),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_275),
.B(n_278),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_279),
.C(n_280),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_257),
.A2(n_247),
.B1(n_251),
.B2(n_242),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_277),
.A2(n_256),
.B1(n_263),
.B2(n_265),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_267),
.B(n_152),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_242),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_247),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_287),
.Y(n_290)
);

INVx11_ASAP7_75t_L g286 ( 
.A(n_270),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_272),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_259),
.C(n_264),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_266),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_272),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_288),
.B(n_271),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_291),
.Y(n_297)
);

AOI31xp33_ASAP7_75t_L g291 ( 
.A1(n_284),
.A2(n_270),
.A3(n_277),
.B(n_274),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_293),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_280),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_294),
.B(n_284),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_290),
.Y(n_295)
);

AOI322xp5_ASAP7_75t_L g302 ( 
.A1(n_295),
.A2(n_296),
.A3(n_283),
.B1(n_262),
.B2(n_285),
.C1(n_286),
.C2(n_276),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_281),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_299),
.A2(n_281),
.B(n_283),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_298),
.B(n_282),
.C(n_287),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_301),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_302),
.A2(n_286),
.B1(n_297),
.B2(n_259),
.Y(n_304)
);

AOI21x1_ASAP7_75t_L g305 ( 
.A1(n_304),
.A2(n_163),
.B(n_16),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_146),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_303),
.Y(n_307)
);


endmodule