module fake_jpeg_13454_n_390 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_390);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_390;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_2),
.B(n_6),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_SL g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_16),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_55),
.B(n_58),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_53),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_56),
.Y(n_124)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_13),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_59),
.B(n_62),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_60),
.Y(n_161)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_61),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_63),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_13),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_64),
.B(n_66),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_65),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_10),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_67),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_33),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_69),
.B(n_77),
.Y(n_114)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_70),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_71),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_10),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_72),
.B(n_82),
.Y(n_131)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

BUFx24_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

CKINVDCx6p67_ASAP7_75t_R g127 ( 
.A(n_74),
.Y(n_127)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_33),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_79),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_80),
.Y(n_162)
);

BUFx16f_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_81),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_43),
.B(n_0),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_0),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_84),
.B(n_87),
.Y(n_153)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_86),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_46),
.B(n_0),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_88),
.Y(n_167)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

BUFx10_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_98),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_1),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_92),
.B(n_97),
.Y(n_168)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_17),
.Y(n_94)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_96),
.Y(n_150)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_26),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_100),
.Y(n_123)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_102),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_30),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_49),
.B(n_2),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_103),
.B(n_104),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_25),
.B(n_3),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_42),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_106),
.Y(n_149)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

CKINVDCx11_ASAP7_75t_R g132 ( 
.A(n_107),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_57),
.A2(n_21),
.B1(n_35),
.B2(n_28),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_110),
.A2(n_142),
.B1(n_145),
.B2(n_152),
.Y(n_191)
);

CKINVDCx12_ASAP7_75t_R g116 ( 
.A(n_74),
.Y(n_116)
);

INVx4_ASAP7_75t_SL g173 ( 
.A(n_116),
.Y(n_173)
);

OR2x2_ASAP7_75t_SL g117 ( 
.A(n_74),
.B(n_19),
.Y(n_117)
);

OR2x4_ASAP7_75t_L g176 ( 
.A(n_117),
.B(n_4),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_60),
.A2(n_21),
.B1(n_35),
.B2(n_28),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_120),
.A2(n_144),
.B1(n_164),
.B2(n_113),
.Y(n_203)
);

AOI21xp33_ASAP7_75t_SL g122 ( 
.A1(n_81),
.A2(n_51),
.B(n_50),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_122),
.B(n_124),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_86),
.B(n_32),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_133),
.B(n_167),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_56),
.A2(n_22),
.B1(n_48),
.B2(n_28),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_135),
.A2(n_146),
.B1(n_166),
.B2(n_162),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_65),
.A2(n_35),
.B1(n_48),
.B2(n_32),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_67),
.A2(n_48),
.B1(n_23),
.B2(n_25),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_L g145 ( 
.A1(n_68),
.A2(n_71),
.B1(n_101),
.B2(n_78),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_90),
.A2(n_23),
.B1(n_52),
.B2(n_31),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_63),
.A2(n_29),
.B1(n_45),
.B2(n_40),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_91),
.B(n_40),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_154),
.B(n_155),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_91),
.B(n_29),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_83),
.B(n_20),
.C(n_45),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_4),
.C(n_6),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_102),
.B(n_20),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_158),
.B(n_163),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_102),
.A2(n_52),
.B1(n_39),
.B2(n_31),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_159),
.A2(n_127),
.B(n_124),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_105),
.B(n_39),
.Y(n_163)
);

OA22x2_ASAP7_75t_L g164 ( 
.A1(n_85),
.A2(n_51),
.B1(n_4),
.B2(n_5),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_105),
.A2(n_89),
.B1(n_107),
.B2(n_5),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_114),
.B(n_3),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_169),
.B(n_175),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_170),
.B(n_180),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_108),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_171),
.B(n_207),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_161),
.Y(n_172)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_172),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_127),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_174),
.B(n_188),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_4),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_176),
.B(n_184),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_119),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_177),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_115),
.B(n_7),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_178),
.B(n_186),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_159),
.A2(n_144),
.B1(n_156),
.B2(n_164),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_179),
.A2(n_185),
.B1(n_201),
.B2(n_203),
.Y(n_235)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_182),
.Y(n_236)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_137),
.Y(n_183)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_183),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_164),
.A2(n_145),
.B1(n_117),
.B2(n_133),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_129),
.B(n_131),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_187),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_168),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_137),
.Y(n_189)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_189),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_127),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_194),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_109),
.B(n_139),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_192),
.B(n_196),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_142),
.A2(n_164),
.B1(n_123),
.B2(n_167),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_193),
.A2(n_217),
.B1(n_199),
.B2(n_204),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_126),
.B(n_128),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_111),
.B(n_147),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_126),
.B(n_128),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_197),
.B(n_204),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_127),
.B(n_149),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_198),
.B(n_208),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_157),
.A2(n_121),
.B1(n_161),
.B2(n_148),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_199),
.A2(n_191),
.B1(n_190),
.B2(n_197),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_121),
.A2(n_157),
.B1(n_148),
.B2(n_136),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_138),
.Y(n_202)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_202),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_150),
.B(n_118),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_138),
.Y(n_205)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_205),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_130),
.B(n_125),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_206),
.B(n_211),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_112),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_132),
.B(n_141),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_113),
.A2(n_162),
.B1(n_112),
.B2(n_160),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_209),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_136),
.Y(n_210)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_210),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_125),
.B(n_160),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_112),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_212),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_162),
.B(n_141),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_215),
.Y(n_244)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_118),
.Y(n_214)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_112),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_143),
.Y(n_216)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_143),
.A2(n_151),
.B1(n_134),
.B2(n_140),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_140),
.B(n_143),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_218),
.B(n_220),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_134),
.A2(n_151),
.B1(n_120),
.B2(n_133),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_219),
.A2(n_203),
.B1(n_174),
.B2(n_201),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_151),
.B(n_133),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_133),
.B(n_69),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_206),
.Y(n_233)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_137),
.Y(n_222)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_222),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_218),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_230),
.B(n_234),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_233),
.B(n_231),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_218),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_237),
.A2(n_258),
.B1(n_261),
.B2(n_265),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_238),
.A2(n_260),
.B1(n_232),
.B2(n_255),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_184),
.B(n_180),
.C(n_220),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_241),
.B(n_248),
.C(n_260),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_191),
.A2(n_190),
.B1(n_221),
.B2(n_219),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_242),
.A2(n_183),
.B1(n_215),
.B2(n_212),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_204),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_246),
.B(n_247),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_194),
.B(n_170),
.Y(n_248)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_210),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_177),
.A2(n_187),
.B1(n_211),
.B2(n_214),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_176),
.A2(n_195),
.B1(n_181),
.B2(n_222),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_243),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_181),
.A2(n_195),
.B1(n_202),
.B2(n_189),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_266),
.B(n_275),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_236),
.Y(n_267)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_267),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_235),
.A2(n_237),
.B1(n_223),
.B2(n_242),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_268),
.A2(n_270),
.B1(n_280),
.B2(n_286),
.Y(n_298)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_228),
.Y(n_269)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_269),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_235),
.A2(n_171),
.B1(n_172),
.B2(n_213),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_271),
.A2(n_281),
.B1(n_252),
.B2(n_278),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_223),
.A2(n_173),
.B(n_207),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_273),
.A2(n_289),
.B(n_295),
.Y(n_306)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_225),
.Y(n_274)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_274),
.Y(n_307)
);

AND2x6_ASAP7_75t_L g275 ( 
.A(n_227),
.B(n_173),
.Y(n_275)
);

INVx13_ASAP7_75t_L g277 ( 
.A(n_236),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_277),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_227),
.A2(n_182),
.B(n_173),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_278),
.A2(n_226),
.B(n_257),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_240),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_283),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_263),
.A2(n_172),
.B1(n_210),
.B2(n_205),
.Y(n_280)
);

OAI32xp33_ASAP7_75t_L g282 ( 
.A1(n_255),
.A2(n_243),
.A3(n_263),
.B1(n_238),
.B2(n_262),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_282),
.B(n_287),
.Y(n_319)
);

INVx13_ASAP7_75t_L g284 ( 
.A(n_229),
.Y(n_284)
);

INVxp33_ASAP7_75t_L g318 ( 
.A(n_284),
.Y(n_318)
);

INVx13_ASAP7_75t_L g285 ( 
.A(n_245),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_285),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_231),
.B(n_233),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_293),
.C(n_254),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_260),
.A2(n_239),
.B(n_232),
.Y(n_289)
);

A2O1A1Ixp33_ASAP7_75t_L g290 ( 
.A1(n_241),
.A2(n_261),
.B(n_244),
.C(n_248),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_291),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_224),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_249),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_292),
.A2(n_294),
.B1(n_274),
.B2(n_286),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_265),
.B(n_251),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_254),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_259),
.B(n_253),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_289),
.A2(n_239),
.B(n_250),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_296),
.B(n_316),
.Y(n_329)
);

AO22x1_ASAP7_75t_SL g299 ( 
.A1(n_268),
.A2(n_257),
.B1(n_226),
.B2(n_225),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_299),
.B(n_302),
.Y(n_321)
);

MAJx2_ASAP7_75t_L g327 ( 
.A(n_304),
.B(n_305),
.C(n_319),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_256),
.C(n_245),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_305),
.B(n_276),
.C(n_271),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_312),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_270),
.A2(n_252),
.B1(n_276),
.B2(n_286),
.Y(n_310)
);

OAI21xp33_ASAP7_75t_L g336 ( 
.A1(n_310),
.A2(n_284),
.B(n_285),
.Y(n_336)
);

OAI21xp33_ASAP7_75t_SL g312 ( 
.A1(n_279),
.A2(n_275),
.B(n_273),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_269),
.Y(n_313)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_313),
.Y(n_324)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_314),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_272),
.A2(n_275),
.B(n_283),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_280),
.Y(n_317)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_317),
.Y(n_330)
);

NOR3xp33_ASAP7_75t_SL g322 ( 
.A(n_315),
.B(n_266),
.C(n_287),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_322),
.B(n_331),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_301),
.A2(n_298),
.B1(n_310),
.B2(n_314),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_325),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_326),
.B(n_327),
.C(n_328),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_304),
.B(n_293),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_299),
.B(n_282),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_298),
.A2(n_290),
.B1(n_272),
.B2(n_292),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_332),
.A2(n_336),
.B1(n_308),
.B2(n_320),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_304),
.B(n_319),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_333),
.B(n_334),
.C(n_335),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_305),
.B(n_294),
.C(n_295),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_303),
.B(n_306),
.C(n_315),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_307),
.Y(n_337)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_337),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_332),
.B(n_301),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_338),
.B(n_344),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_303),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_339),
.B(n_349),
.Y(n_363)
);

BUFx4f_ASAP7_75t_SL g340 ( 
.A(n_323),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_340),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_329),
.A2(n_302),
.B(n_312),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_335),
.A2(n_306),
.B(n_316),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_345),
.B(n_346),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_334),
.B(n_318),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_347),
.B(n_351),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_333),
.B(n_299),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_323),
.A2(n_296),
.B(n_309),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_350),
.A2(n_320),
.B(n_330),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_321),
.Y(n_351)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_341),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_353),
.B(n_355),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_351),
.B(n_324),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_342),
.B(n_327),
.C(n_326),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_356),
.B(n_364),
.C(n_322),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_340),
.A2(n_321),
.B(n_331),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_357),
.B(n_352),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_359),
.B(n_347),
.Y(n_366)
);

BUFx24_ASAP7_75t_SL g361 ( 
.A(n_343),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_361),
.B(n_300),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_342),
.B(n_348),
.C(n_339),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_354),
.A2(n_352),
.B1(n_317),
.B2(n_330),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_365),
.B(n_368),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_366),
.B(n_369),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_364),
.B(n_348),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_356),
.B(n_349),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_370),
.B(n_363),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_371),
.B(n_372),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_360),
.B(n_340),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_373),
.B(n_357),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_377),
.A2(n_366),
.B(n_363),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_378),
.A2(n_369),
.B(n_362),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_373),
.B(n_358),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_379),
.B(n_370),
.C(n_367),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_380),
.A2(n_374),
.B1(n_309),
.B2(n_311),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_381),
.B(n_382),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_376),
.A2(n_362),
.B1(n_337),
.B2(n_307),
.Y(n_383)
);

OA21x2_ASAP7_75t_SL g385 ( 
.A1(n_383),
.A2(n_384),
.B(n_299),
.Y(n_385)
);

NOR2xp67_ASAP7_75t_L g384 ( 
.A(n_374),
.B(n_375),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_385),
.A2(n_297),
.B1(n_300),
.B2(n_267),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_388),
.B(n_387),
.C(n_386),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_389),
.B(n_285),
.Y(n_390)
);


endmodule