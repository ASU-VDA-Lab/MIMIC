module real_jpeg_6572_n_30 (n_17, n_8, n_0, n_21, n_168, n_2, n_29, n_10, n_9, n_12, n_24, n_165, n_166, n_170, n_6, n_28, n_171, n_169, n_162, n_167, n_23, n_11, n_14, n_25, n_163, n_7, n_22, n_18, n_3, n_5, n_4, n_1, n_26, n_27, n_20, n_19, n_164, n_16, n_15, n_13, n_30);

input n_17;
input n_8;
input n_0;
input n_21;
input n_168;
input n_2;
input n_29;
input n_10;
input n_9;
input n_12;
input n_24;
input n_165;
input n_166;
input n_170;
input n_6;
input n_28;
input n_171;
input n_169;
input n_162;
input n_167;
input n_23;
input n_11;
input n_14;
input n_25;
input n_163;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_164;
input n_16;
input n_15;
input n_13;

output n_30;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_64;
wire n_47;
wire n_131;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_150;
wire n_41;
wire n_74;
wire n_32;
wire n_80;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

INVx5_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_0),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_0),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_0),
.B(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_1),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_2),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_2),
.B(n_33),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_2),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_3),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_5),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_5),
.B(n_58),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_6),
.B(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_7),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_9),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_9),
.B(n_50),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_10),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_10),
.B(n_54),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_11),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_11),
.B(n_145),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_12),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_12),
.B(n_148),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_13),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_14),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_14),
.B(n_44),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_15),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_16),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_18),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_18),
.B(n_93),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_19),
.Y(n_135)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_21),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_21),
.B(n_106),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_22),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_23),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_24),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_24),
.B(n_121),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_25),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_25),
.B(n_70),
.Y(n_99)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_28),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_28),
.B(n_67),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_29),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_29),
.B(n_130),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_154),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_39),
.B(n_153),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_35),
.B(n_102),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_35),
.B(n_158),
.Y(n_157)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_143),
.B(n_150),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_123),
.B(n_137),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_62),
.B(n_111),
.C(n_120),
.Y(n_41)
);

NOR4xp25_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_49),
.C(n_53),
.D(n_57),
.Y(n_42)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_43),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_49),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_52),
.B(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_53),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_105),
.B(n_110),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_100),
.B(n_104),
.Y(n_63)
);

AO221x1_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_76),
.B1(n_97),
.B2(n_98),
.C(n_99),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_75),
.B(n_94),
.Y(n_93)
);

AO21x1_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_82),
.B(n_96),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_81),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_92),
.B(n_95),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_87),
.B(n_91),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_90),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_90),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_103),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_103),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_122),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_149),
.Y(n_148)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

A2O1A1O1Ixp25_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B(n_117),
.C(n_118),
.D(n_119),
.Y(n_112)
);

NAND3xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.C(n_133),
.Y(n_123)
);

A2O1A1O1Ixp25_ASAP7_75t_L g137 ( 
.A1(n_124),
.A2(n_133),
.B(n_138),
.C(n_141),
.D(n_142),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_126),
.Y(n_142)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_129),
.A2(n_139),
.B(n_140),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_136),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_147),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_160),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_159),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_162),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_163),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_164),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_165),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_166),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_167),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_168),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_169),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_170),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_171),
.Y(n_107)
);


endmodule