module real_jpeg_32037_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx3_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_0),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_0),
.Y(n_179)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_0),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_1),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_1),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_1),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_1),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_1),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_1),
.B(n_255),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_1),
.Y(n_279)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_2),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_2),
.B(n_66),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_2),
.B(n_272),
.Y(n_271)
);

NAND2xp33_ASAP7_75t_SL g302 ( 
.A(n_2),
.B(n_303),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_3),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_3),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_3),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_3),
.B(n_188),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_4),
.Y(n_160)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_5),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_5),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_5),
.B(n_159),
.Y(n_158)
);

AND2x2_ASAP7_75t_SL g270 ( 
.A(n_5),
.B(n_157),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_5),
.B(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_5),
.B(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_6),
.B(n_117),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_6),
.B(n_157),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_6),
.Y(n_180)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_7),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_8),
.B(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_8),
.B(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_8),
.B(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_8),
.B(n_123),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_8),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_8),
.B(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_9),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_10),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_10),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_10),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_12),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_13),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_13),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_13),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_13),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_13),
.B(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_13),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_13),
.B(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_13),
.B(n_319),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_14),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_14),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_14),
.Y(n_197)
);

NAND2x1_ASAP7_75t_L g54 ( 
.A(n_15),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_15),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_15),
.B(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_15),
.B(n_152),
.Y(n_151)
);

AND2x2_ASAP7_75t_SL g165 ( 
.A(n_15),
.B(n_166),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g184 ( 
.A(n_15),
.B(n_185),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_203),
.Y(n_16)
);

NAND2xp33_ASAP7_75t_R g17 ( 
.A(n_18),
.B(n_202),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_167),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_19),
.B(n_167),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_97),
.Y(n_19)
);

MAJx2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_44),
.C(n_59),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_21),
.B(n_44),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_34),
.B2(n_43),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_24),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_26),
.Y(n_307)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_27),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_28),
.Y(n_334)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_29),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_32),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_32),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_33),
.B(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

MAJx2_ASAP7_75t_L g100 ( 
.A(n_34),
.B(n_101),
.C(n_102),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_36),
.Y(n_280)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OA21x2_ASAP7_75t_SL g171 ( 
.A1(n_43),
.A2(n_172),
.B(n_177),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_54),
.B2(n_58),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_46)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_48),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_50),
.B(n_53),
.C(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_50),
.B(n_184),
.Y(n_183)
);

OA21x2_ASAP7_75t_L g257 ( 
.A1(n_50),
.A2(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_50),
.B(n_258),
.Y(n_259)
);

OAI21xp33_ASAP7_75t_L g290 ( 
.A1(n_50),
.A2(n_258),
.B(n_259),
.Y(n_290)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_52),
.Y(n_316)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_57),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_59),
.B(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_74),
.C(n_81),
.Y(n_59)
);

XOR2x2_ASAP7_75t_L g231 ( 
.A(n_60),
.B(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_61),
.B(n_65),
.C(n_73),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_63),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_68),
.B1(n_72),
.B2(n_73),
.Y(n_64)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_68),
.Y(n_73)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_74),
.B(n_82),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_80),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_75),
.B(n_80),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NOR2x1_ASAP7_75t_L g138 ( 
.A(n_79),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_79),
.B(n_253),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_79),
.B(n_331),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_80),
.B(n_165),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.C(n_91),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_83),
.A2(n_87),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_83),
.Y(n_215)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_86),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_87),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_89),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_90),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_91),
.B(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_94),
.Y(n_268)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_96),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_144),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_113),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_106),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_109),
.B1(n_111),
.B2(n_112),
.Y(n_106)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_109),
.Y(n_112)
);

MAJx2_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_131),
.C(n_132),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_114),
.B(n_131),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_121),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_125),
.C(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_120),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_120),
.Y(n_253)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_120),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_125),
.B1(n_129),
.B2(n_130),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

XOR2x2_ASAP7_75t_L g200 ( 
.A(n_132),
.B(n_201),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_138),
.C(n_140),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_133),
.B(n_140),
.Y(n_199)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2x2_ASAP7_75t_L g198 ( 
.A(n_138),
.B(n_199),
.Y(n_198)
);

OR2x2_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_143),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2x1_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_161),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_149),
.B2(n_150),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_155),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_165),
.B(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_165),
.B(n_251),
.Y(n_286)
);

INVx8_ASAP7_75t_L g328 ( 
.A(n_166),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.C(n_200),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_168),
.B(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_170),
.B(n_200),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_181),
.C(n_198),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_198),
.Y(n_209)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

BUFx4f_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_181),
.B(n_209),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_186),
.C(n_191),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_182),
.A2(n_183),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_184),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_186),
.A2(n_187),
.B1(n_191),
.B2(n_192),
.Y(n_247)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_235),
.B(n_354),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_233),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g354 ( 
.A(n_207),
.B(n_233),
.Y(n_354)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.C(n_231),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_239),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_231),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_217),
.C(n_218),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_243),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_217),
.A2(n_218),
.B1(n_219),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_225),
.C(n_227),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_220),
.A2(n_221),
.B1(n_225),
.B2(n_226),
.Y(n_294)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_227),
.B(n_294),
.Y(n_293)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVxp67_ASAP7_75t_SL g235 ( 
.A(n_236),
.Y(n_235)
);

AO21x2_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_260),
.B(n_353),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_238),
.B(n_240),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_245),
.C(n_248),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_241),
.A2(n_242),
.B1(n_351),
.B2(n_352),
.Y(n_350)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_242),
.B(n_347),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_245),
.B(n_248),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_245),
.B(n_248),
.Y(n_352)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_254),
.C(n_257),
.Y(n_248)
);

XNOR2x1_ASAP7_75t_L g288 ( 
.A(n_249),
.B(n_289),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_254),
.A2(n_257),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_254),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_345),
.B(n_349),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_296),
.B(n_344),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_287),
.Y(n_262)
);

NOR2x1_ASAP7_75t_L g344 ( 
.A(n_263),
.B(n_287),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_276),
.C(n_286),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_265),
.B(n_341),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_269),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_266),
.B(n_270),
.C(n_275),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_267),
.B(n_326),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_274),
.B2(n_275),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_270),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_271),
.Y(n_275)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

AO22x1_ASAP7_75t_L g341 ( 
.A1(n_276),
.A2(n_277),
.B1(n_286),
.B2(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_281),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_278),
.A2(n_281),
.B1(n_282),
.B2(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_278),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_286),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_292),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_288),
.B(n_293),
.C(n_295),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_295),
.Y(n_292)
);

OAI21x1_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_338),
.B(n_343),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_322),
.B(n_337),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_311),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_299),
.B(n_311),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_308),
.B2(n_309),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_305),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_302),
.B(n_305),
.C(n_308),
.Y(n_339)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_317),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_312),
.A2(n_313),
.B1(n_317),
.B2(n_318),
.Y(n_335)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx3_ASAP7_75t_SL g314 ( 
.A(n_315),
.Y(n_314)
);

INVx8_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

OAI21x1_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_329),
.B(n_336),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_335),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_330),
.B(n_335),
.Y(n_336)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_339),
.B(n_340),
.Y(n_343)
);

NOR2x1p5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_348),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);


endmodule