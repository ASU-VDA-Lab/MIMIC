module fake_jpeg_8610_n_113 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_113);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_113;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx11_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_62),
.B(n_1),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_66),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g64 ( 
.A(n_50),
.B(n_1),
.Y(n_64)
);

OA22x2_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_53),
.B1(n_2),
.B2(n_3),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_69),
.Y(n_84)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_51),
.B1(n_49),
.B2(n_58),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_71),
.A2(n_72),
.B1(n_81),
.B2(n_82),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_68),
.A2(n_58),
.B1(n_52),
.B2(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_78),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_67),
.B(n_46),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_75),
.Y(n_92)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

OR2x2_ASAP7_75t_SL g88 ( 
.A(n_76),
.B(n_83),
.Y(n_88)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_85),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_55),
.B1(n_54),
.B2(n_3),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_70),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_4),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_70),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_87),
.A2(n_21),
.B1(n_22),
.B2(n_25),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_90),
.B1(n_91),
.B2(n_93),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_17),
.B1(n_18),
.B2(n_20),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_79),
.B(n_27),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

AND2x6_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_86),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_100),
.A2(n_95),
.B1(n_99),
.B2(n_92),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_101),
.B(n_92),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_97),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_103),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

NOR2xp67_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_88),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_96),
.B1(n_97),
.B2(n_84),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

AOI322xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_28),
.A3(n_29),
.B1(n_30),
.B2(n_32),
.C1(n_33),
.C2(n_38),
.Y(n_109)
);

INVxp33_ASAP7_75t_L g110 ( 
.A(n_109),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_110),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_39),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_40),
.Y(n_113)
);


endmodule