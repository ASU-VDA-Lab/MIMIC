module fake_aes_6686_n_1311 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_272, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_270, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_1311);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_272;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
output n_1311;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_613;
wire n_648;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1079;
wire n_315;
wire n_409;
wire n_295;
wire n_677;
wire n_1242;
wire n_283;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_281;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_280;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_275;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1117;
wire n_1007;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_287;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_596;
wire n_1215;
wire n_286;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_282;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_285;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_290;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_288;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_274;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_276;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_335;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_819;
wire n_772;
wire n_405;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g273 ( .A(n_190), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_235), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_37), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_84), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_26), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_72), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_202), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_173), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_60), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_30), .Y(n_282) );
OR2x2_ASAP7_75t_L g283 ( .A(n_49), .B(n_161), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_56), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_167), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_237), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g287 ( .A(n_35), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_205), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_139), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_238), .Y(n_290) );
BUFx2_ASAP7_75t_L g291 ( .A(n_270), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_192), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_197), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_31), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_60), .Y(n_295) );
INVx1_ASAP7_75t_SL g296 ( .A(n_162), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_79), .Y(n_297) );
INVx1_ASAP7_75t_SL g298 ( .A(n_102), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_31), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_216), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_128), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_142), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_116), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_99), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_105), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_154), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_165), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_61), .Y(n_308) );
BUFx2_ASAP7_75t_L g309 ( .A(n_172), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_8), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_84), .B(n_245), .Y(n_311) );
CKINVDCx14_ASAP7_75t_R g312 ( .A(n_175), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_196), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_258), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_232), .Y(n_315) );
CKINVDCx16_ASAP7_75t_R g316 ( .A(n_20), .Y(n_316) );
CKINVDCx20_ASAP7_75t_R g317 ( .A(n_179), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_33), .Y(n_318) );
NOR2xp67_ASAP7_75t_L g319 ( .A(n_83), .B(n_77), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_217), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_184), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_231), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_261), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_4), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_45), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_164), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_2), .Y(n_327) );
CKINVDCx20_ASAP7_75t_R g328 ( .A(n_272), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_158), .Y(n_329) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_195), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_121), .Y(n_331) );
INVx1_ASAP7_75t_SL g332 ( .A(n_57), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_86), .Y(n_333) );
CKINVDCx20_ASAP7_75t_R g334 ( .A(n_252), .Y(n_334) );
CKINVDCx20_ASAP7_75t_R g335 ( .A(n_185), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_255), .Y(n_336) );
CKINVDCx20_ASAP7_75t_R g337 ( .A(n_104), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_57), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_138), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_95), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_250), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_187), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_49), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_135), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_101), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_123), .Y(n_346) );
CKINVDCx20_ASAP7_75t_R g347 ( .A(n_126), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_213), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_159), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_117), .Y(n_350) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_153), .Y(n_351) );
INVxp67_ASAP7_75t_SL g352 ( .A(n_78), .Y(n_352) );
CKINVDCx20_ASAP7_75t_R g353 ( .A(n_91), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_193), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_207), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_80), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_249), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_111), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_44), .Y(n_359) );
CKINVDCx20_ASAP7_75t_R g360 ( .A(n_247), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_157), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_204), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_91), .Y(n_363) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_109), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_41), .Y(n_365) );
CKINVDCx20_ASAP7_75t_R g366 ( .A(n_146), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_27), .Y(n_367) );
INVxp67_ASAP7_75t_SL g368 ( .A(n_36), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_143), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_51), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_30), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_2), .Y(n_372) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_66), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_13), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_83), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_125), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_110), .Y(n_377) );
INVx1_ASAP7_75t_SL g378 ( .A(n_65), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_118), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_92), .Y(n_380) );
BUFx2_ASAP7_75t_SL g381 ( .A(n_0), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_4), .Y(n_382) );
BUFx3_ASAP7_75t_L g383 ( .A(n_156), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_37), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_144), .Y(n_385) );
CKINVDCx20_ASAP7_75t_R g386 ( .A(n_150), .Y(n_386) );
INVx1_ASAP7_75t_SL g387 ( .A(n_224), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_79), .Y(n_388) );
BUFx10_ASAP7_75t_L g389 ( .A(n_1), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_14), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_74), .Y(n_391) );
BUFx5_ASAP7_75t_L g392 ( .A(n_229), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_262), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_48), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_67), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_65), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_191), .Y(n_397) );
CKINVDCx16_ASAP7_75t_R g398 ( .A(n_140), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_119), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_13), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_152), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_233), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_263), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_264), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_70), .Y(n_405) );
BUFx8_ASAP7_75t_SL g406 ( .A(n_194), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_97), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_171), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_254), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_52), .Y(n_410) );
CKINVDCx20_ASAP7_75t_R g411 ( .A(n_9), .Y(n_411) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_68), .Y(n_412) );
CKINVDCx14_ASAP7_75t_R g413 ( .A(n_137), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_259), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_246), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_115), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_32), .Y(n_417) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_90), .Y(n_418) );
INVxp67_ASAP7_75t_L g419 ( .A(n_176), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_160), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_225), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_130), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_188), .Y(n_423) );
CKINVDCx5p33_ASAP7_75t_R g424 ( .A(n_34), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_6), .Y(n_425) );
CKINVDCx5p33_ASAP7_75t_R g426 ( .A(n_17), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_198), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_278), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_392), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_392), .Y(n_430) );
BUFx3_ASAP7_75t_L g431 ( .A(n_320), .Y(n_431) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_279), .Y(n_432) );
BUFx8_ASAP7_75t_L g433 ( .A(n_291), .Y(n_433) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_278), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_320), .B(n_0), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_281), .Y(n_436) );
BUFx3_ASAP7_75t_L g437 ( .A(n_383), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_316), .A2(n_5), .B1(n_1), .B2(n_3), .Y(n_438) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_279), .Y(n_439) );
INVx5_ASAP7_75t_L g440 ( .A(n_279), .Y(n_440) );
INVxp67_ASAP7_75t_L g441 ( .A(n_309), .Y(n_441) );
BUFx2_ASAP7_75t_L g442 ( .A(n_406), .Y(n_442) );
AND2x4_ASAP7_75t_L g443 ( .A(n_281), .B(n_3), .Y(n_443) );
AND2x4_ASAP7_75t_L g444 ( .A(n_382), .B(n_5), .Y(n_444) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_279), .Y(n_445) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_330), .Y(n_446) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_330), .Y(n_447) );
BUFx2_ASAP7_75t_L g448 ( .A(n_406), .Y(n_448) );
OA21x2_ASAP7_75t_L g449 ( .A1(n_303), .A2(n_100), .B(n_98), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_392), .Y(n_450) );
INVx3_ASAP7_75t_L g451 ( .A(n_303), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_382), .B(n_6), .Y(n_452) );
OAI21x1_ASAP7_75t_L g453 ( .A1(n_321), .A2(n_106), .B(n_103), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_395), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_395), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_400), .Y(n_456) );
BUFx2_ASAP7_75t_L g457 ( .A(n_312), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_351), .B(n_7), .Y(n_458) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_330), .Y(n_459) );
BUFx2_ASAP7_75t_L g460 ( .A(n_312), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_400), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_419), .B(n_7), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_273), .Y(n_463) );
BUFx3_ASAP7_75t_L g464 ( .A(n_383), .Y(n_464) );
OA21x2_ASAP7_75t_L g465 ( .A1(n_321), .A2(n_108), .B(n_107), .Y(n_465) );
INVx3_ASAP7_75t_L g466 ( .A(n_345), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_280), .Y(n_467) );
INVx2_ASAP7_75t_SL g468 ( .A(n_389), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_443), .Y(n_469) );
AO22x2_ASAP7_75t_L g470 ( .A1(n_438), .A2(n_381), .B1(n_283), .B2(n_368), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_429), .Y(n_471) );
AND3x1_ASAP7_75t_L g472 ( .A(n_468), .B(n_294), .C(n_282), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g473 ( .A1(n_441), .A2(n_398), .B1(n_335), .B2(n_337), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_457), .B(n_274), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_443), .A2(n_297), .B1(n_299), .B2(n_295), .Y(n_475) );
INVx3_ASAP7_75t_L g476 ( .A(n_435), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_430), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_457), .B(n_413), .Y(n_478) );
OAI22xp33_ASAP7_75t_L g479 ( .A1(n_442), .A2(n_353), .B1(n_418), .B2(n_287), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_430), .Y(n_480) );
NAND2xp33_ASAP7_75t_R g481 ( .A(n_442), .B(n_275), .Y(n_481) );
INVx3_ASAP7_75t_L g482 ( .A(n_435), .Y(n_482) );
AO21x1_ASAP7_75t_L g483 ( .A1(n_435), .A2(n_311), .B(n_286), .Y(n_483) );
INVx2_ASAP7_75t_SL g484 ( .A(n_457), .Y(n_484) );
INVx8_ASAP7_75t_L g485 ( .A(n_435), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_443), .A2(n_310), .B1(n_327), .B2(n_308), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_443), .A2(n_333), .B1(n_340), .B2(n_338), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_443), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_444), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_430), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_450), .Y(n_491) );
BUFx3_ASAP7_75t_L g492 ( .A(n_460), .Y(n_492) );
OR2x6_ASAP7_75t_L g493 ( .A(n_442), .B(n_319), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_460), .B(n_413), .Y(n_494) );
INVx2_ASAP7_75t_SL g495 ( .A(n_460), .Y(n_495) );
AND2x6_ASAP7_75t_L g496 ( .A(n_435), .B(n_285), .Y(n_496) );
INVx5_ASAP7_75t_L g497 ( .A(n_440), .Y(n_497) );
NAND3xp33_ASAP7_75t_L g498 ( .A(n_458), .B(n_433), .C(n_463), .Y(n_498) );
NAND2xp33_ASAP7_75t_SL g499 ( .A(n_448), .B(n_334), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_450), .Y(n_500) );
AND3x2_ASAP7_75t_L g501 ( .A(n_448), .B(n_352), .C(n_343), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_450), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_444), .A2(n_356), .B1(n_367), .B2(n_359), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_468), .B(n_290), .Y(n_504) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_432), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_448), .Y(n_506) );
NAND2xp33_ASAP7_75t_SL g507 ( .A(n_468), .B(n_334), .Y(n_507) );
OAI21xp33_ASAP7_75t_SL g508 ( .A1(n_463), .A2(n_372), .B(n_371), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_440), .Y(n_509) );
BUFx6f_ASAP7_75t_SL g510 ( .A(n_444), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_467), .B(n_292), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_431), .B(n_276), .Y(n_512) );
INVx8_ASAP7_75t_L g513 ( .A(n_444), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_452), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_476), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_484), .B(n_433), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_483), .B(n_433), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_484), .B(n_433), .Y(n_518) );
BUFx5_ASAP7_75t_L g519 ( .A(n_496), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_495), .B(n_433), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_492), .B(n_431), .Y(n_521) );
BUFx3_ASAP7_75t_L g522 ( .A(n_492), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_478), .B(n_431), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_476), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_476), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_498), .B(n_458), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_482), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_494), .B(n_462), .Y(n_528) );
BUFx3_ASAP7_75t_L g529 ( .A(n_506), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_506), .B(n_434), .Y(n_530) );
NOR3xp33_ASAP7_75t_L g531 ( .A(n_479), .B(n_438), .C(n_378), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_482), .A2(n_452), .B(n_453), .C(n_451), .Y(n_532) );
NOR2xp67_ASAP7_75t_L g533 ( .A(n_473), .B(n_434), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_482), .Y(n_534) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_485), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_474), .B(n_455), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_493), .B(n_455), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_512), .B(n_464), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_485), .B(n_452), .Y(n_539) );
NAND3xp33_ASAP7_75t_SL g540 ( .A(n_475), .B(n_284), .C(n_277), .Y(n_540) );
AND3x1_ASAP7_75t_L g541 ( .A(n_486), .B(n_394), .C(n_390), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_485), .Y(n_542) );
INVx2_ASAP7_75t_SL g543 ( .A(n_501), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_485), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_510), .A2(n_452), .B1(n_337), .B2(n_347), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_513), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_513), .B(n_437), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_513), .B(n_437), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_504), .B(n_437), .Y(n_549) );
OAI21xp5_ASAP7_75t_L g550 ( .A1(n_477), .A2(n_453), .B(n_449), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_469), .B(n_293), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_488), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_487), .B(n_437), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_503), .B(n_451), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_493), .B(n_335), .Y(n_555) );
OAI22xp33_ASAP7_75t_L g556 ( .A1(n_489), .A2(n_347), .B1(n_366), .B2(n_360), .Y(n_556) );
BUFx3_ASAP7_75t_L g557 ( .A(n_477), .Y(n_557) );
AND2x2_ASAP7_75t_SL g558 ( .A(n_472), .B(n_449), .Y(n_558) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_496), .Y(n_559) );
NOR2x1p5_ASAP7_75t_L g560 ( .A(n_481), .B(n_318), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_499), .B(n_332), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_510), .A2(n_366), .B1(n_386), .B2(n_360), .Y(n_562) );
NOR2x1_ASAP7_75t_L g563 ( .A(n_493), .B(n_317), .Y(n_563) );
INVxp67_ASAP7_75t_SL g564 ( .A(n_514), .Y(n_564) );
AOI22xp33_ASAP7_75t_SL g565 ( .A1(n_470), .A2(n_353), .B1(n_418), .B2(n_287), .Y(n_565) );
INVxp67_ASAP7_75t_L g566 ( .A(n_510), .Y(n_566) );
A2O1A1Ixp33_ASAP7_75t_L g567 ( .A1(n_511), .A2(n_453), .B(n_466), .C(n_451), .Y(n_567) );
INVxp67_ASAP7_75t_SL g568 ( .A(n_491), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_500), .B(n_300), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_508), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_493), .B(n_470), .Y(n_571) );
INVxp67_ASAP7_75t_L g572 ( .A(n_496), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_500), .B(n_304), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_471), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_507), .A2(n_386), .B1(n_328), .B2(n_363), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_507), .B(n_288), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_480), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_480), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_490), .B(n_451), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_502), .B(n_428), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_470), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_470), .B(n_466), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_509), .B(n_436), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_497), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_499), .A2(n_365), .B1(n_370), .B2(n_325), .Y(n_585) );
NAND2x1_ASAP7_75t_L g586 ( .A(n_505), .B(n_449), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_497), .B(n_454), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_497), .B(n_305), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_505), .B(n_456), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_505), .B(n_456), .Y(n_590) );
BUFx3_ASAP7_75t_L g591 ( .A(n_492), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_485), .A2(n_465), .B(n_449), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_484), .B(n_461), .Y(n_593) );
INVxp67_ASAP7_75t_L g594 ( .A(n_492), .Y(n_594) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_492), .Y(n_595) );
OR2x6_ASAP7_75t_L g596 ( .A(n_485), .B(n_410), .Y(n_596) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_485), .Y(n_597) );
BUFx2_ASAP7_75t_L g598 ( .A(n_492), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_568), .B(n_373), .Y(n_599) );
AOI21xp5_ASAP7_75t_L g600 ( .A1(n_592), .A2(n_465), .B(n_449), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_568), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_594), .B(n_374), .Y(n_602) );
BUFx2_ASAP7_75t_L g603 ( .A(n_596), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_532), .A2(n_465), .B(n_313), .Y(n_604) );
AOI21xp5_ASAP7_75t_L g605 ( .A1(n_586), .A2(n_465), .B(n_314), .Y(n_605) );
AOI21xp5_ASAP7_75t_L g606 ( .A1(n_526), .A2(n_465), .B(n_323), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_533), .A2(n_380), .B1(n_384), .B2(n_375), .Y(n_607) );
INVxp67_ASAP7_75t_L g608 ( .A(n_529), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_535), .B(n_289), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_557), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_530), .B(n_389), .Y(n_611) );
NAND2x1p5_ASAP7_75t_L g612 ( .A(n_535), .B(n_324), .Y(n_612) );
NAND2x1p5_ASAP7_75t_L g613 ( .A(n_535), .B(n_324), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_541), .A2(n_391), .B1(n_396), .B2(n_388), .Y(n_614) );
BUFx2_ASAP7_75t_L g615 ( .A(n_596), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_594), .B(n_417), .Y(n_616) );
NAND3xp33_ASAP7_75t_SL g617 ( .A(n_565), .B(n_411), .C(n_405), .Y(n_617) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_597), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_550), .A2(n_326), .B(n_307), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_515), .Y(n_620) );
A2O1A1Ixp33_ASAP7_75t_L g621 ( .A1(n_570), .A2(n_331), .B(n_341), .C(n_339), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_540), .A2(n_424), .B1(n_426), .B2(n_425), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g623 ( .A1(n_538), .A2(n_355), .B(n_349), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_595), .B(n_389), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_598), .B(n_296), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_595), .B(n_301), .Y(n_626) );
BUFx8_ASAP7_75t_L g627 ( .A(n_555), .Y(n_627) );
O2A1O1Ixp33_ASAP7_75t_L g628 ( .A1(n_581), .A2(n_358), .B(n_369), .C(n_357), .Y(n_628) );
NOR3xp33_ASAP7_75t_L g629 ( .A(n_556), .B(n_387), .C(n_298), .Y(n_629) );
CKINVDCx20_ASAP7_75t_R g630 ( .A(n_562), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_593), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_523), .A2(n_385), .B(n_379), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_564), .B(n_302), .Y(n_633) );
NAND2x1_ASAP7_75t_L g634 ( .A(n_596), .B(n_345), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_567), .A2(n_397), .B(n_393), .Y(n_635) );
CKINVDCx20_ASAP7_75t_R g636 ( .A(n_575), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_545), .A2(n_412), .B1(n_401), .B2(n_402), .Y(n_637) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_549), .A2(n_404), .B(n_399), .Y(n_638) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_597), .B(n_306), .Y(n_639) );
AOI21xp5_ASAP7_75t_L g640 ( .A1(n_539), .A2(n_408), .B(n_407), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_524), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_552), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_525), .Y(n_643) );
INVx3_ASAP7_75t_L g644 ( .A(n_542), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_564), .B(n_315), .Y(n_645) );
NAND3xp33_ASAP7_75t_L g646 ( .A(n_517), .B(n_415), .C(n_414), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_527), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_528), .A2(n_420), .B(n_416), .Y(n_648) );
BUFx3_ASAP7_75t_L g649 ( .A(n_522), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_534), .Y(n_650) );
AND2x4_ASAP7_75t_L g651 ( .A(n_591), .B(n_422), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g652 ( .A1(n_547), .A2(n_427), .B(n_421), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_516), .B(n_322), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_559), .A2(n_336), .B1(n_342), .B2(n_329), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_536), .B(n_344), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_536), .B(n_346), .Y(n_656) );
O2A1O1Ixp33_ASAP7_75t_L g657 ( .A1(n_582), .A2(n_10), .B(n_8), .C(n_9), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_540), .A2(n_348), .B1(n_354), .B2(n_350), .Y(n_658) );
AOI21xp5_ASAP7_75t_L g659 ( .A1(n_548), .A2(n_440), .B(n_362), .Y(n_659) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_566), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_544), .B(n_361), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_537), .B(n_10), .Y(n_662) );
NOR2xp67_ASAP7_75t_L g663 ( .A(n_543), .B(n_11), .Y(n_663) );
O2A1O1Ixp33_ASAP7_75t_L g664 ( .A1(n_531), .A2(n_554), .B(n_553), .C(n_561), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_580), .Y(n_665) );
INVx11_ASAP7_75t_L g666 ( .A(n_565), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_546), .B(n_376), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_518), .B(n_377), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_574), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_577), .Y(n_670) );
INVx3_ASAP7_75t_L g671 ( .A(n_559), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_520), .B(n_403), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_571), .A2(n_392), .B1(n_423), .B2(n_409), .Y(n_673) );
AO21x2_ASAP7_75t_L g674 ( .A1(n_569), .A2(n_392), .B(n_364), .Y(n_674) );
OA22x2_ASAP7_75t_L g675 ( .A1(n_555), .A2(n_14), .B1(n_11), .B2(n_12), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_585), .B(n_12), .Y(n_676) );
NAND3xp33_ASAP7_75t_L g677 ( .A(n_558), .B(n_440), .C(n_364), .Y(n_677) );
BUFx4f_ASAP7_75t_L g678 ( .A(n_558), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_578), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_572), .A2(n_566), .B1(n_521), .B2(n_551), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_551), .B(n_576), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_583), .Y(n_682) );
OR2x2_ASAP7_75t_L g683 ( .A(n_531), .B(n_560), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_519), .B(n_432), .Y(n_684) );
OA22x2_ASAP7_75t_L g685 ( .A1(n_563), .A2(n_18), .B1(n_15), .B2(n_16), .Y(n_685) );
OAI22xp33_ASAP7_75t_L g686 ( .A1(n_579), .A2(n_439), .B1(n_445), .B2(n_432), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_573), .B(n_18), .Y(n_687) );
CKINVDCx20_ASAP7_75t_R g688 ( .A(n_519), .Y(n_688) );
OA22x2_ASAP7_75t_L g689 ( .A1(n_588), .A2(n_21), .B1(n_19), .B2(n_20), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_590), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_587), .B(n_22), .Y(n_691) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_584), .B(n_445), .Y(n_692) );
OAI21x1_ASAP7_75t_L g693 ( .A1(n_589), .A2(n_113), .B(n_112), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_568), .B(n_23), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_568), .A2(n_447), .B1(n_459), .B2(n_446), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_568), .B(n_24), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_568), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_530), .B(n_25), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_568), .B(n_27), .Y(n_699) );
A2O1A1Ixp33_ASAP7_75t_L g700 ( .A1(n_570), .A2(n_459), .B(n_447), .C(n_32), .Y(n_700) );
A2O1A1Ixp33_ASAP7_75t_L g701 ( .A1(n_570), .A2(n_459), .B(n_447), .C(n_33), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_530), .B(n_28), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_568), .A2(n_28), .B1(n_29), .B2(n_36), .Y(n_703) );
AND2x4_ASAP7_75t_L g704 ( .A(n_596), .B(n_29), .Y(n_704) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_535), .B(n_38), .Y(n_705) );
AOI21xp5_ASAP7_75t_L g706 ( .A1(n_592), .A2(n_120), .B(n_114), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_533), .A2(n_38), .B1(n_39), .B2(n_40), .Y(n_707) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_531), .A2(n_39), .B1(n_40), .B2(n_41), .C(n_42), .Y(n_708) );
INVx3_ASAP7_75t_L g709 ( .A(n_535), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_530), .B(n_42), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_592), .A2(n_124), .B(n_122), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_568), .B(n_43), .Y(n_712) );
A2O1A1Ixp33_ASAP7_75t_L g713 ( .A1(n_570), .A2(n_43), .B(n_44), .C(n_45), .Y(n_713) );
BUFx3_ASAP7_75t_L g714 ( .A(n_522), .Y(n_714) );
NAND2xp5_ASAP7_75t_SL g715 ( .A(n_535), .B(n_46), .Y(n_715) );
NOR3xp33_ASAP7_75t_L g716 ( .A(n_556), .B(n_46), .C(n_47), .Y(n_716) );
O2A1O1Ixp33_ASAP7_75t_L g717 ( .A1(n_581), .A2(n_47), .B(n_48), .C(n_50), .Y(n_717) );
OAI21xp33_ASAP7_75t_SL g718 ( .A1(n_568), .A2(n_50), .B(n_52), .Y(n_718) );
A2O1A1Ixp33_ASAP7_75t_L g719 ( .A1(n_570), .A2(n_53), .B(n_54), .C(n_55), .Y(n_719) );
NAND2x1p5_ASAP7_75t_L g720 ( .A(n_535), .B(n_53), .Y(n_720) );
O2A1O1Ixp33_ASAP7_75t_L g721 ( .A1(n_581), .A2(n_54), .B(n_55), .C(n_56), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_631), .B(n_58), .Y(n_722) );
AOI21xp5_ASAP7_75t_L g723 ( .A1(n_600), .A2(n_129), .B(n_127), .Y(n_723) );
NAND2xp5_ASAP7_75t_SL g724 ( .A(n_603), .B(n_58), .Y(n_724) );
OAI21xp5_ASAP7_75t_L g725 ( .A1(n_604), .A2(n_132), .B(n_131), .Y(n_725) );
BUFx2_ASAP7_75t_L g726 ( .A(n_704), .Y(n_726) );
OAI22x1_ASAP7_75t_L g727 ( .A1(n_704), .A2(n_59), .B1(n_61), .B2(n_62), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_642), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g729 ( .A(n_615), .B(n_59), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_675), .Y(n_730) );
BUFx6f_ASAP7_75t_L g731 ( .A(n_618), .Y(n_731) );
OAI21xp5_ASAP7_75t_L g732 ( .A1(n_635), .A2(n_134), .B(n_133), .Y(n_732) );
CKINVDCx11_ASAP7_75t_R g733 ( .A(n_630), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_601), .B(n_62), .Y(n_734) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_605), .A2(n_141), .B(n_136), .Y(n_735) );
OAI21xp5_ASAP7_75t_L g736 ( .A1(n_619), .A2(n_646), .B(n_677), .Y(n_736) );
BUFx6f_ASAP7_75t_L g737 ( .A(n_618), .Y(n_737) );
INVx6_ASAP7_75t_L g738 ( .A(n_627), .Y(n_738) );
AO21x1_ASAP7_75t_L g739 ( .A1(n_720), .A2(n_147), .B(n_145), .Y(n_739) );
BUFx6f_ASAP7_75t_L g740 ( .A(n_612), .Y(n_740) );
BUFx8_ASAP7_75t_L g741 ( .A(n_649), .Y(n_741) );
AOI21xp5_ASAP7_75t_L g742 ( .A1(n_681), .A2(n_149), .B(n_148), .Y(n_742) );
AND2x4_ASAP7_75t_L g743 ( .A(n_714), .B(n_63), .Y(n_743) );
OAI21x1_ASAP7_75t_L g744 ( .A1(n_693), .A2(n_155), .B(n_151), .Y(n_744) );
AO31x2_ASAP7_75t_L g745 ( .A1(n_700), .A2(n_64), .A3(n_67), .B(n_68), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_627), .Y(n_746) );
NOR2xp67_ASAP7_75t_SL g747 ( .A(n_660), .B(n_69), .Y(n_747) );
NOR2x1_ASAP7_75t_L g748 ( .A(n_617), .B(n_69), .Y(n_748) );
OR2x6_ASAP7_75t_L g749 ( .A(n_608), .B(n_70), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_697), .B(n_71), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_710), .B(n_71), .Y(n_751) );
NAND2x1p5_ASAP7_75t_L g752 ( .A(n_709), .B(n_72), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_698), .B(n_73), .Y(n_753) );
OAI21xp5_ASAP7_75t_L g754 ( .A1(n_646), .A2(n_212), .B(n_269), .Y(n_754) );
AO21x1_ASAP7_75t_L g755 ( .A1(n_720), .A2(n_211), .B(n_268), .Y(n_755) );
OAI21x1_ASAP7_75t_L g756 ( .A1(n_706), .A2(n_210), .B(n_267), .Y(n_756) );
OAI21xp5_ASAP7_75t_SL g757 ( .A1(n_629), .A2(n_75), .B(n_76), .Y(n_757) );
AOI21xp5_ASAP7_75t_L g758 ( .A1(n_659), .A2(n_209), .B(n_266), .Y(n_758) );
NAND2xp5_ASAP7_75t_SL g759 ( .A(n_654), .B(n_75), .Y(n_759) );
AOI21xp33_ASAP7_75t_L g760 ( .A1(n_664), .A2(n_77), .B(n_78), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_702), .B(n_80), .Y(n_761) );
AOI21xp5_ASAP7_75t_L g762 ( .A1(n_680), .A2(n_214), .B(n_265), .Y(n_762) );
INVx4_ASAP7_75t_L g763 ( .A(n_709), .Y(n_763) );
BUFx2_ASAP7_75t_L g764 ( .A(n_636), .Y(n_764) );
AND2x4_ASAP7_75t_L g765 ( .A(n_682), .B(n_81), .Y(n_765) );
OAI21x1_ASAP7_75t_L g766 ( .A1(n_711), .A2(n_208), .B(n_260), .Y(n_766) );
BUFx3_ASAP7_75t_L g767 ( .A(n_651), .Y(n_767) );
O2A1O1Ixp5_ASAP7_75t_L g768 ( .A1(n_678), .A2(n_206), .B(n_257), .C(n_256), .Y(n_768) );
OR2x2_ASAP7_75t_L g769 ( .A(n_611), .B(n_82), .Y(n_769) );
A2O1A1Ixp33_ASAP7_75t_L g770 ( .A1(n_628), .A2(n_82), .B(n_85), .C(n_86), .Y(n_770) );
AOI21xp5_ASAP7_75t_L g771 ( .A1(n_638), .A2(n_215), .B(n_253), .Y(n_771) );
AO31x2_ASAP7_75t_L g772 ( .A1(n_701), .A2(n_85), .A3(n_87), .B(n_88), .Y(n_772) );
AOI21xp5_ASAP7_75t_L g773 ( .A1(n_632), .A2(n_203), .B(n_251), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_599), .B(n_87), .Y(n_774) );
NOR2xp33_ASAP7_75t_L g775 ( .A(n_683), .B(n_88), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_669), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_675), .Y(n_777) );
NOR2xp33_ASAP7_75t_L g778 ( .A(n_607), .B(n_89), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g779 ( .A(n_666), .B(n_92), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_662), .B(n_93), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_665), .B(n_93), .Y(n_781) );
AOI21xp5_ASAP7_75t_L g782 ( .A1(n_684), .A2(n_623), .B(n_633), .Y(n_782) );
NAND3xp33_ASAP7_75t_SL g783 ( .A(n_716), .B(n_94), .C(n_95), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_670), .Y(n_784) );
OAI22x1_ASAP7_75t_L g785 ( .A1(n_707), .A2(n_96), .B1(n_163), .B2(n_166), .Y(n_785) );
AND2x6_ASAP7_75t_SL g786 ( .A(n_676), .B(n_168), .Y(n_786) );
INVx2_ASAP7_75t_SL g787 ( .A(n_651), .Y(n_787) );
O2A1O1Ixp5_ASAP7_75t_L g788 ( .A1(n_678), .A2(n_169), .B(n_170), .C(n_174), .Y(n_788) );
AOI21xp5_ASAP7_75t_L g789 ( .A1(n_645), .A2(n_177), .B(n_178), .Y(n_789) );
NAND2xp33_ASAP7_75t_R g790 ( .A(n_671), .B(n_180), .Y(n_790) );
AOI21xp5_ASAP7_75t_SL g791 ( .A1(n_694), .A2(n_181), .B(n_182), .Y(n_791) );
OAI21xp5_ASAP7_75t_L g792 ( .A1(n_652), .A2(n_183), .B(n_186), .Y(n_792) );
CKINVDCx5p33_ASAP7_75t_R g793 ( .A(n_614), .Y(n_793) );
CKINVDCx11_ASAP7_75t_R g794 ( .A(n_688), .Y(n_794) );
CKINVDCx5p33_ASAP7_75t_R g795 ( .A(n_637), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_679), .Y(n_796) );
OR2x6_ASAP7_75t_L g797 ( .A(n_685), .B(n_189), .Y(n_797) );
INVx4_ASAP7_75t_L g798 ( .A(n_612), .Y(n_798) );
BUFx5_ASAP7_75t_L g799 ( .A(n_647), .Y(n_799) );
A2O1A1Ixp33_ASAP7_75t_L g800 ( .A1(n_718), .A2(n_199), .B(n_200), .C(n_201), .Y(n_800) );
NAND2xp5_ASAP7_75t_SL g801 ( .A(n_625), .B(n_610), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_621), .B(n_622), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_696), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_699), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_712), .Y(n_805) );
AOI21xp5_ASAP7_75t_SL g806 ( .A1(n_613), .A2(n_271), .B(n_218), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_602), .B(n_219), .Y(n_807) );
INVx2_ASAP7_75t_L g808 ( .A(n_620), .Y(n_808) );
OR2x2_ASAP7_75t_L g809 ( .A(n_624), .B(n_220), .Y(n_809) );
INVx2_ASAP7_75t_SL g810 ( .A(n_634), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_616), .B(n_221), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_655), .B(n_222), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_690), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_656), .B(n_223), .Y(n_814) );
AO32x2_ASAP7_75t_L g815 ( .A1(n_703), .A2(n_226), .A3(n_227), .B1(n_228), .B2(n_230), .Y(n_815) );
AO21x1_ASAP7_75t_L g816 ( .A1(n_657), .A2(n_234), .B(n_236), .Y(n_816) );
OAI21xp5_ASAP7_75t_L g817 ( .A1(n_640), .A2(n_239), .B(n_240), .Y(n_817) );
OAI21xp5_ASAP7_75t_L g818 ( .A1(n_650), .A2(n_241), .B(n_242), .Y(n_818) );
AND2x2_ASAP7_75t_L g819 ( .A(n_658), .B(n_243), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_644), .B(n_244), .Y(n_820) );
INVx2_ASAP7_75t_L g821 ( .A(n_641), .Y(n_821) );
AND2x4_ASAP7_75t_L g822 ( .A(n_609), .B(n_248), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_643), .Y(n_823) );
AND2x2_ASAP7_75t_L g824 ( .A(n_626), .B(n_685), .Y(n_824) );
OR2x2_ASAP7_75t_L g825 ( .A(n_661), .B(n_667), .Y(n_825) );
NAND3xp33_ASAP7_75t_L g826 ( .A(n_653), .B(n_672), .C(n_668), .Y(n_826) );
BUFx3_ASAP7_75t_L g827 ( .A(n_687), .Y(n_827) );
AO22x2_ASAP7_75t_L g828 ( .A1(n_705), .A2(n_715), .B1(n_689), .B2(n_721), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_717), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_691), .Y(n_830) );
O2A1O1Ixp33_ASAP7_75t_L g831 ( .A1(n_713), .A2(n_719), .B(n_708), .C(n_639), .Y(n_831) );
AND2x2_ASAP7_75t_L g832 ( .A(n_663), .B(n_673), .Y(n_832) );
INVx5_ASAP7_75t_L g833 ( .A(n_686), .Y(n_833) );
AND2x2_ASAP7_75t_L g834 ( .A(n_674), .B(n_695), .Y(n_834) );
NAND3xp33_ASAP7_75t_SL g835 ( .A(n_692), .B(n_448), .C(n_442), .Y(n_835) );
AOI211x1_ASAP7_75t_L g836 ( .A1(n_648), .A2(n_581), .B(n_517), .C(n_483), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_631), .B(n_581), .Y(n_837) );
AO31x2_ASAP7_75t_L g838 ( .A1(n_604), .A2(n_567), .A3(n_532), .B(n_635), .Y(n_838) );
OR2x2_ASAP7_75t_L g839 ( .A(n_617), .B(n_556), .Y(n_839) );
OAI22x1_ASAP7_75t_L g840 ( .A1(n_704), .A2(n_473), .B1(n_562), .B2(n_575), .Y(n_840) );
INVx2_ASAP7_75t_L g841 ( .A(n_669), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_642), .Y(n_842) );
AOI21xp5_ASAP7_75t_L g843 ( .A1(n_600), .A2(n_592), .B(n_606), .Y(n_843) );
AO21x1_ASAP7_75t_L g844 ( .A1(n_635), .A2(n_604), .B(n_619), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_631), .B(n_581), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_642), .Y(n_846) );
BUFx2_ASAP7_75t_SL g847 ( .A(n_704), .Y(n_847) );
NOR4xp25_ASAP7_75t_L g848 ( .A(n_718), .B(n_617), .C(n_664), .D(n_717), .Y(n_848) );
INVx2_ASAP7_75t_L g849 ( .A(n_669), .Y(n_849) );
NOR2xp67_ASAP7_75t_L g850 ( .A(n_617), .B(n_562), .Y(n_850) );
BUFx6f_ASAP7_75t_L g851 ( .A(n_618), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_601), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_631), .B(n_581), .Y(n_853) );
OAI21x1_ASAP7_75t_L g854 ( .A1(n_600), .A2(n_605), .B(n_586), .Y(n_854) );
NAND2xp5_ASAP7_75t_SL g855 ( .A(n_603), .B(n_535), .Y(n_855) );
AND2x4_ASAP7_75t_L g856 ( .A(n_631), .B(n_603), .Y(n_856) );
NOR2x1_ASAP7_75t_SL g857 ( .A(n_631), .B(n_596), .Y(n_857) );
AOI21xp5_ASAP7_75t_L g858 ( .A1(n_600), .A2(n_592), .B(n_606), .Y(n_858) );
NOR3xp33_ASAP7_75t_SL g859 ( .A(n_617), .B(n_499), .C(n_479), .Y(n_859) );
BUFx2_ASAP7_75t_L g860 ( .A(n_746), .Y(n_860) );
OA21x2_ASAP7_75t_L g861 ( .A1(n_843), .A2(n_858), .B(n_854), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_852), .B(n_813), .Y(n_862) );
AO31x2_ASAP7_75t_L g863 ( .A1(n_844), .A2(n_816), .A3(n_755), .B(n_739), .Y(n_863) );
HB1xp67_ASAP7_75t_L g864 ( .A(n_765), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_852), .B(n_813), .Y(n_865) );
OA21x2_ASAP7_75t_L g866 ( .A1(n_736), .A2(n_725), .B(n_744), .Y(n_866) );
INVx3_ASAP7_75t_L g867 ( .A(n_798), .Y(n_867) );
NOR2xp67_ASAP7_75t_L g868 ( .A(n_840), .B(n_839), .Y(n_868) );
AND2x4_ASAP7_75t_L g869 ( .A(n_857), .B(n_856), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_728), .B(n_842), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_846), .B(n_803), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_784), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_784), .Y(n_873) );
INVx3_ASAP7_75t_L g874 ( .A(n_798), .Y(n_874) );
BUFx3_ASAP7_75t_L g875 ( .A(n_741), .Y(n_875) );
NOR2xp33_ASAP7_75t_L g876 ( .A(n_793), .B(n_726), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_796), .Y(n_877) );
OR2x2_ASAP7_75t_L g878 ( .A(n_764), .B(n_847), .Y(n_878) );
BUFx6f_ASAP7_75t_L g879 ( .A(n_731), .Y(n_879) );
BUFx3_ASAP7_75t_L g880 ( .A(n_741), .Y(n_880) );
INVx2_ASAP7_75t_L g881 ( .A(n_776), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_804), .B(n_805), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_830), .B(n_837), .Y(n_883) );
CKINVDCx6p67_ASAP7_75t_R g884 ( .A(n_749), .Y(n_884) );
OA21x2_ASAP7_75t_L g885 ( .A1(n_732), .A2(n_754), .B(n_834), .Y(n_885) );
A2O1A1Ixp33_ASAP7_75t_L g886 ( .A1(n_831), .A2(n_826), .B(n_829), .C(n_730), .Y(n_886) );
NOR2x1_ASAP7_75t_SL g887 ( .A(n_797), .B(n_749), .Y(n_887) );
OAI21xp5_ASAP7_75t_L g888 ( .A1(n_777), .A2(n_802), .B(n_782), .Y(n_888) );
OAI22xp5_ASAP7_75t_L g889 ( .A1(n_765), .A2(n_797), .B1(n_853), .B2(n_845), .Y(n_889) );
BUFx2_ASAP7_75t_SL g890 ( .A(n_856), .Y(n_890) );
INVx3_ASAP7_75t_L g891 ( .A(n_763), .Y(n_891) );
INVx1_ASAP7_75t_L g892 ( .A(n_841), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_849), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_830), .B(n_824), .Y(n_894) );
INVx2_ASAP7_75t_SL g895 ( .A(n_738), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_734), .Y(n_896) );
OA21x2_ASAP7_75t_L g897 ( .A1(n_723), .A2(n_792), .B(n_818), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_750), .Y(n_898) );
OA21x2_ASAP7_75t_L g899 ( .A1(n_735), .A2(n_766), .B(n_756), .Y(n_899) );
OR2x6_ASAP7_75t_L g900 ( .A(n_738), .B(n_743), .Y(n_900) );
AOI21xp5_ASAP7_75t_L g901 ( .A1(n_814), .A2(n_807), .B(n_811), .Y(n_901) );
A2O1A1Ixp33_ASAP7_75t_L g902 ( .A1(n_775), .A2(n_757), .B(n_760), .C(n_812), .Y(n_902) );
OR2x2_ASAP7_75t_L g903 ( .A(n_769), .B(n_787), .Y(n_903) );
INVx1_ASAP7_75t_SL g904 ( .A(n_767), .Y(n_904) );
AOI21xp33_ASAP7_75t_SL g905 ( .A1(n_779), .A2(n_727), .B(n_778), .Y(n_905) );
AND2x4_ASAP7_75t_L g906 ( .A(n_827), .B(n_825), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_722), .Y(n_907) );
OA21x2_ASAP7_75t_L g908 ( .A1(n_800), .A2(n_788), .B(n_768), .Y(n_908) );
BUFx2_ASAP7_75t_L g909 ( .A(n_743), .Y(n_909) );
INVx4_ASAP7_75t_L g910 ( .A(n_794), .Y(n_910) );
OAI22xp33_ASAP7_75t_SL g911 ( .A1(n_752), .A2(n_748), .B1(n_795), .B2(n_724), .Y(n_911) );
OAI21x1_ASAP7_75t_L g912 ( .A1(n_758), .A2(n_762), .B(n_820), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_848), .B(n_823), .Y(n_913) );
AND2x4_ASAP7_75t_L g914 ( .A(n_822), .B(n_763), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_823), .B(n_836), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_781), .Y(n_916) );
BUFx3_ASAP7_75t_L g917 ( .A(n_733), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_808), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_821), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_850), .B(n_774), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_747), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_799), .B(n_832), .Y(n_922) );
AO31x2_ASAP7_75t_L g923 ( .A1(n_785), .A2(n_770), .A3(n_789), .B(n_742), .Y(n_923) );
INVx2_ASAP7_75t_SL g924 ( .A(n_855), .Y(n_924) );
OR2x2_ASAP7_75t_L g925 ( .A(n_751), .B(n_780), .Y(n_925) );
OA21x2_ASAP7_75t_L g926 ( .A1(n_817), .A2(n_771), .B(n_773), .Y(n_926) );
INVx2_ASAP7_75t_SL g927 ( .A(n_729), .Y(n_927) );
INVxp67_ASAP7_75t_L g928 ( .A(n_790), .Y(n_928) );
BUFx2_ASAP7_75t_R g929 ( .A(n_801), .Y(n_929) );
AO21x1_ASAP7_75t_L g930 ( .A1(n_759), .A2(n_761), .B(n_753), .Y(n_930) );
OAI21x1_ASAP7_75t_L g931 ( .A1(n_806), .A2(n_791), .B(n_809), .Y(n_931) );
OAI21x1_ASAP7_75t_L g932 ( .A1(n_838), .A2(n_819), .B(n_783), .Y(n_932) );
AND2x4_ASAP7_75t_L g933 ( .A(n_822), .B(n_810), .Y(n_933) );
NOR2x1_ASAP7_75t_SL g934 ( .A(n_737), .B(n_851), .Y(n_934) );
CKINVDCx6p67_ASAP7_75t_R g935 ( .A(n_799), .Y(n_935) );
INVx2_ASAP7_75t_SL g936 ( .A(n_737), .Y(n_936) );
OAI21x1_ASAP7_75t_L g937 ( .A1(n_838), .A2(n_851), .B(n_740), .Y(n_937) );
OAI21xp5_ASAP7_75t_L g938 ( .A1(n_859), .A2(n_833), .B(n_835), .Y(n_938) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_828), .B(n_786), .Y(n_939) );
OAI21xp33_ASAP7_75t_SL g940 ( .A1(n_815), .A2(n_833), .B(n_745), .Y(n_940) );
INVx1_ASAP7_75t_L g941 ( .A(n_745), .Y(n_941) );
NOR2xp33_ASAP7_75t_R g942 ( .A(n_772), .B(n_746), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_772), .Y(n_943) );
AND2x4_ASAP7_75t_L g944 ( .A(n_772), .B(n_857), .Y(n_944) );
INVx3_ASAP7_75t_L g945 ( .A(n_798), .Y(n_945) );
INVx1_ASAP7_75t_L g946 ( .A(n_728), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_852), .B(n_631), .Y(n_947) );
NOR2xp33_ASAP7_75t_L g948 ( .A(n_839), .B(n_555), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_728), .Y(n_949) );
NAND3xp33_ASAP7_75t_L g950 ( .A(n_800), .B(n_757), .C(n_760), .Y(n_950) );
BUFx2_ASAP7_75t_L g951 ( .A(n_746), .Y(n_951) );
NAND2xp5_ASAP7_75t_SL g952 ( .A(n_765), .B(n_704), .Y(n_952) );
A2O1A1Ixp33_ASAP7_75t_L g953 ( .A1(n_831), .A2(n_826), .B(n_664), .C(n_829), .Y(n_953) );
INVxp67_ASAP7_75t_L g954 ( .A(n_765), .Y(n_954) );
BUFx3_ASAP7_75t_L g955 ( .A(n_741), .Y(n_955) );
AO31x2_ASAP7_75t_L g956 ( .A1(n_844), .A2(n_843), .A3(n_858), .B(n_567), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g957 ( .A(n_852), .B(n_631), .Y(n_957) );
HB1xp67_ASAP7_75t_L g958 ( .A(n_765), .Y(n_958) );
HB1xp67_ASAP7_75t_L g959 ( .A(n_856), .Y(n_959) );
NAND2x1p5_ASAP7_75t_L g960 ( .A(n_765), .B(n_704), .Y(n_960) );
OR2x2_ASAP7_75t_L g961 ( .A(n_764), .B(n_530), .Y(n_961) );
AO31x2_ASAP7_75t_L g962 ( .A1(n_844), .A2(n_843), .A3(n_858), .B(n_567), .Y(n_962) );
AND2x2_ASAP7_75t_L g963 ( .A(n_856), .B(n_530), .Y(n_963) );
INVx3_ASAP7_75t_L g964 ( .A(n_798), .Y(n_964) );
INVx3_ASAP7_75t_L g965 ( .A(n_798), .Y(n_965) );
INVx3_ASAP7_75t_L g966 ( .A(n_798), .Y(n_966) );
AO31x2_ASAP7_75t_L g967 ( .A1(n_844), .A2(n_843), .A3(n_858), .B(n_567), .Y(n_967) );
INVx2_ASAP7_75t_SL g968 ( .A(n_741), .Y(n_968) );
NAND2xp5_ASAP7_75t_SL g969 ( .A(n_765), .B(n_704), .Y(n_969) );
HB1xp67_ASAP7_75t_L g970 ( .A(n_856), .Y(n_970) );
INVx2_ASAP7_75t_L g971 ( .A(n_852), .Y(n_971) );
BUFx2_ASAP7_75t_L g972 ( .A(n_746), .Y(n_972) );
CKINVDCx5p33_ASAP7_75t_R g973 ( .A(n_746), .Y(n_973) );
AOI22xp5_ASAP7_75t_L g974 ( .A1(n_850), .A2(n_617), .B1(n_556), .B2(n_479), .Y(n_974) );
AND2x2_ASAP7_75t_L g975 ( .A(n_856), .B(n_530), .Y(n_975) );
AOI22xp5_ASAP7_75t_L g976 ( .A1(n_850), .A2(n_617), .B1(n_556), .B2(n_479), .Y(n_976) );
BUFx3_ASAP7_75t_L g977 ( .A(n_935), .Y(n_977) );
OR2x6_ASAP7_75t_L g978 ( .A(n_889), .B(n_960), .Y(n_978) );
HB1xp67_ASAP7_75t_L g979 ( .A(n_906), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_915), .Y(n_980) );
BUFx2_ASAP7_75t_L g981 ( .A(n_960), .Y(n_981) );
AND2x2_ASAP7_75t_L g982 ( .A(n_971), .B(n_862), .Y(n_982) );
HB1xp67_ASAP7_75t_L g983 ( .A(n_906), .Y(n_983) );
INVx1_ASAP7_75t_L g984 ( .A(n_915), .Y(n_984) );
HB1xp67_ASAP7_75t_L g985 ( .A(n_900), .Y(n_985) );
OR2x2_ASAP7_75t_L g986 ( .A(n_862), .B(n_865), .Y(n_986) );
AND2x2_ASAP7_75t_L g987 ( .A(n_865), .B(n_872), .Y(n_987) );
INVx2_ASAP7_75t_L g988 ( .A(n_861), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_913), .Y(n_989) );
OR2x2_ASAP7_75t_L g990 ( .A(n_889), .B(n_894), .Y(n_990) );
AND2x2_ASAP7_75t_L g991 ( .A(n_873), .B(n_877), .Y(n_991) );
BUFx2_ASAP7_75t_L g992 ( .A(n_864), .Y(n_992) );
INVx1_ASAP7_75t_SL g993 ( .A(n_860), .Y(n_993) );
AND2x2_ASAP7_75t_L g994 ( .A(n_894), .B(n_881), .Y(n_994) );
AND2x2_ASAP7_75t_L g995 ( .A(n_887), .B(n_886), .Y(n_995) );
INVx1_ASAP7_75t_L g996 ( .A(n_941), .Y(n_996) );
OAI21xp33_ASAP7_75t_L g997 ( .A1(n_942), .A2(n_976), .B(n_974), .Y(n_997) );
OR2x2_ASAP7_75t_L g998 ( .A(n_864), .B(n_958), .Y(n_998) );
OR2x2_ASAP7_75t_L g999 ( .A(n_958), .B(n_947), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_943), .Y(n_1000) );
INVx2_ASAP7_75t_L g1001 ( .A(n_956), .Y(n_1001) );
CKINVDCx6p67_ASAP7_75t_R g1002 ( .A(n_875), .Y(n_1002) );
HB1xp67_ASAP7_75t_L g1003 ( .A(n_900), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_963), .B(n_975), .Y(n_1004) );
BUFx2_ASAP7_75t_SL g1005 ( .A(n_869), .Y(n_1005) );
BUFx2_ASAP7_75t_L g1006 ( .A(n_937), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_892), .B(n_893), .Y(n_1007) );
INVx2_ASAP7_75t_L g1008 ( .A(n_956), .Y(n_1008) );
OR2x2_ASAP7_75t_L g1009 ( .A(n_947), .B(n_957), .Y(n_1009) );
BUFx2_ASAP7_75t_L g1010 ( .A(n_909), .Y(n_1010) );
HB1xp67_ASAP7_75t_L g1011 ( .A(n_900), .Y(n_1011) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_957), .B(n_882), .Y(n_1012) );
NAND2x1p5_ASAP7_75t_L g1013 ( .A(n_914), .B(n_952), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_948), .B(n_882), .Y(n_1014) );
HB1xp67_ASAP7_75t_L g1015 ( .A(n_959), .Y(n_1015) );
HB1xp67_ASAP7_75t_L g1016 ( .A(n_970), .Y(n_1016) );
INVx3_ASAP7_75t_L g1017 ( .A(n_879), .Y(n_1017) );
INVx1_ASAP7_75t_L g1018 ( .A(n_888), .Y(n_1018) );
INVx2_ASAP7_75t_L g1019 ( .A(n_962), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g1020 ( .A(n_871), .B(n_946), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_870), .Y(n_1021) );
HB1xp67_ASAP7_75t_L g1022 ( .A(n_903), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g1023 ( .A(n_871), .B(n_949), .Y(n_1023) );
INVxp67_ASAP7_75t_L g1024 ( .A(n_890), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_870), .Y(n_1025) );
HB1xp67_ASAP7_75t_L g1026 ( .A(n_904), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_918), .B(n_919), .Y(n_1027) );
CKINVDCx6p67_ASAP7_75t_R g1028 ( .A(n_880), .Y(n_1028) );
HB1xp67_ASAP7_75t_L g1029 ( .A(n_904), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_922), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_922), .Y(n_1031) );
INVx1_ASAP7_75t_L g1032 ( .A(n_967), .Y(n_1032) );
OR2x2_ASAP7_75t_L g1033 ( .A(n_939), .B(n_883), .Y(n_1033) );
HB1xp67_ASAP7_75t_L g1034 ( .A(n_954), .Y(n_1034) );
INVx1_ASAP7_75t_L g1035 ( .A(n_883), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_953), .B(n_907), .Y(n_1036) );
AOI21x1_ASAP7_75t_L g1037 ( .A1(n_866), .A2(n_901), .B(n_897), .Y(n_1037) );
HB1xp67_ASAP7_75t_L g1038 ( .A(n_954), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_944), .Y(n_1039) );
NOR2xp33_ASAP7_75t_L g1040 ( .A(n_905), .B(n_884), .Y(n_1040) );
INVx2_ASAP7_75t_SL g1041 ( .A(n_867), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_944), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_932), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_896), .B(n_898), .Y(n_1044) );
OAI22xp5_ASAP7_75t_L g1045 ( .A1(n_969), .A2(n_928), .B1(n_939), .B2(n_929), .Y(n_1045) );
OR2x2_ASAP7_75t_L g1046 ( .A(n_868), .B(n_961), .Y(n_1046) );
AOI21x1_ASAP7_75t_L g1047 ( .A1(n_866), .A2(n_901), .B(n_897), .Y(n_1047) );
AOI21xp33_ASAP7_75t_L g1048 ( .A1(n_920), .A2(n_902), .B(n_950), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_869), .B(n_920), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_940), .Y(n_1050) );
OR2x2_ASAP7_75t_L g1051 ( .A(n_1033), .B(n_928), .Y(n_1051) );
AND2x2_ASAP7_75t_L g1052 ( .A(n_1030), .B(n_885), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g1053 ( .A1(n_997), .A2(n_921), .B1(n_938), .B2(n_927), .Y(n_1053) );
INVx1_ASAP7_75t_L g1054 ( .A(n_996), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_996), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_997), .A2(n_938), .B1(n_933), .B2(n_911), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_1030), .B(n_885), .Y(n_1057) );
OAI22xp5_ASAP7_75t_L g1058 ( .A1(n_978), .A2(n_929), .B1(n_914), .B2(n_933), .Y(n_1058) );
NOR2x1_ASAP7_75t_L g1059 ( .A(n_977), .B(n_945), .Y(n_1059) );
INVx1_ASAP7_75t_L g1060 ( .A(n_1000), .Y(n_1060) );
NAND2xp5_ASAP7_75t_L g1061 ( .A(n_1012), .B(n_916), .Y(n_1061) );
NAND2xp5_ASAP7_75t_L g1062 ( .A(n_1012), .B(n_876), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1000), .Y(n_1063) );
BUFx2_ASAP7_75t_L g1064 ( .A(n_978), .Y(n_1064) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_1044), .B(n_911), .Y(n_1065) );
AND2x2_ASAP7_75t_L g1066 ( .A(n_1031), .B(n_982), .Y(n_1066) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_978), .A2(n_925), .B1(n_930), .B2(n_910), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_1031), .B(n_863), .Y(n_1068) );
BUFx3_ASAP7_75t_L g1069 ( .A(n_977), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_1044), .B(n_878), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_982), .B(n_863), .Y(n_1071) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_980), .B(n_863), .Y(n_1072) );
INVx2_ASAP7_75t_L g1073 ( .A(n_988), .Y(n_1073) );
AOI22xp5_ASAP7_75t_L g1074 ( .A1(n_1036), .A2(n_867), .B1(n_874), .B2(n_945), .Y(n_1074) );
NAND3xp33_ASAP7_75t_L g1075 ( .A(n_1048), .B(n_924), .C(n_964), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_984), .B(n_874), .Y(n_1076) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_984), .B(n_966), .Y(n_1077) );
AND2x2_ASAP7_75t_L g1078 ( .A(n_987), .B(n_966), .Y(n_1078) );
BUFx12f_ASAP7_75t_L g1079 ( .A(n_977), .Y(n_1079) );
NAND2xp5_ASAP7_75t_L g1080 ( .A(n_1035), .B(n_965), .Y(n_1080) );
BUFx2_ASAP7_75t_SL g1081 ( .A(n_1041), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_987), .B(n_965), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_994), .B(n_964), .Y(n_1083) );
BUFx2_ASAP7_75t_L g1084 ( .A(n_978), .Y(n_1084) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_994), .B(n_923), .Y(n_1085) );
OR2x2_ASAP7_75t_L g1086 ( .A(n_1033), .B(n_891), .Y(n_1086) );
AOI21xp5_ASAP7_75t_SL g1087 ( .A1(n_978), .A2(n_934), .B(n_926), .Y(n_1087) );
HB1xp67_ASAP7_75t_L g1088 ( .A(n_1026), .Y(n_1088) );
HB1xp67_ASAP7_75t_L g1089 ( .A(n_1029), .Y(n_1089) );
HB1xp67_ASAP7_75t_L g1090 ( .A(n_1015), .Y(n_1090) );
NAND2xp5_ASAP7_75t_L g1091 ( .A(n_1035), .B(n_895), .Y(n_1091) );
OR2x2_ASAP7_75t_L g1092 ( .A(n_989), .B(n_891), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_989), .B(n_936), .Y(n_1093) );
NAND2xp5_ASAP7_75t_L g1094 ( .A(n_1036), .B(n_972), .Y(n_1094) );
AOI21xp33_ASAP7_75t_L g1095 ( .A1(n_1046), .A2(n_908), .B(n_926), .Y(n_1095) );
NAND2xp5_ASAP7_75t_L g1096 ( .A(n_1009), .B(n_1021), .Y(n_1096) );
OAI222xp33_ASAP7_75t_L g1097 ( .A1(n_1045), .A2(n_910), .B1(n_968), .B2(n_951), .C1(n_973), .C2(n_917), .Y(n_1097) );
OR2x2_ASAP7_75t_L g1098 ( .A(n_990), .B(n_955), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_991), .B(n_931), .Y(n_1099) );
OR2x2_ASAP7_75t_L g1100 ( .A(n_990), .B(n_899), .Y(n_1100) );
BUFx2_ASAP7_75t_L g1101 ( .A(n_1039), .Y(n_1101) );
NAND2xp5_ASAP7_75t_L g1102 ( .A(n_1009), .B(n_1021), .Y(n_1102) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1032), .Y(n_1103) );
AND2x4_ASAP7_75t_L g1104 ( .A(n_1039), .B(n_912), .Y(n_1104) );
INVx1_ASAP7_75t_SL g1105 ( .A(n_1002), .Y(n_1105) );
INVxp67_ASAP7_75t_SL g1106 ( .A(n_986), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_991), .B(n_899), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1085), .B(n_1050), .Y(n_1108) );
INVx3_ASAP7_75t_SL g1109 ( .A(n_1105), .Y(n_1109) );
NAND2xp5_ASAP7_75t_L g1110 ( .A(n_1106), .B(n_1025), .Y(n_1110) );
INVxp67_ASAP7_75t_L g1111 ( .A(n_1090), .Y(n_1111) );
INVx1_ASAP7_75t_SL g1112 ( .A(n_1079), .Y(n_1112) );
INVx1_ASAP7_75t_L g1113 ( .A(n_1054), .Y(n_1113) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_1066), .B(n_1025), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1054), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1085), .B(n_1050), .Y(n_1116) );
INVx2_ASAP7_75t_L g1117 ( .A(n_1073), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_1071), .B(n_1042), .Y(n_1118) );
AND2x4_ASAP7_75t_L g1119 ( .A(n_1099), .B(n_1042), .Y(n_1119) );
AND2x4_ASAP7_75t_L g1120 ( .A(n_1099), .B(n_1043), .Y(n_1120) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1055), .Y(n_1121) );
AND2x2_ASAP7_75t_SL g1122 ( .A(n_1064), .B(n_995), .Y(n_1122) );
INVx2_ASAP7_75t_SL g1123 ( .A(n_1059), .Y(n_1123) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1055), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1060), .Y(n_1125) );
HB1xp67_ASAP7_75t_L g1126 ( .A(n_1088), .Y(n_1126) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1060), .Y(n_1127) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_1071), .B(n_1001), .Y(n_1128) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1063), .Y(n_1129) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1063), .Y(n_1130) );
INVx4_ASAP7_75t_L g1131 ( .A(n_1069), .Y(n_1131) );
INVxp67_ASAP7_75t_L g1132 ( .A(n_1089), .Y(n_1132) );
AND2x2_ASAP7_75t_SL g1133 ( .A(n_1084), .B(n_995), .Y(n_1133) );
AND2x2_ASAP7_75t_L g1134 ( .A(n_1107), .B(n_1008), .Y(n_1134) );
INVxp67_ASAP7_75t_SL g1135 ( .A(n_1086), .Y(n_1135) );
NOR2xp33_ASAP7_75t_L g1136 ( .A(n_1097), .B(n_993), .Y(n_1136) );
HB1xp67_ASAP7_75t_L g1137 ( .A(n_1078), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_1107), .B(n_1008), .Y(n_1138) );
OR2x2_ASAP7_75t_L g1139 ( .A(n_1066), .B(n_1018), .Y(n_1139) );
BUFx6f_ASAP7_75t_L g1140 ( .A(n_1104), .Y(n_1140) );
NAND2xp5_ASAP7_75t_SL g1141 ( .A(n_1059), .B(n_1041), .Y(n_1141) );
AND2x4_ASAP7_75t_L g1142 ( .A(n_1104), .B(n_1006), .Y(n_1142) );
NAND2xp5_ASAP7_75t_L g1143 ( .A(n_1096), .B(n_1049), .Y(n_1143) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_1102), .B(n_1049), .Y(n_1144) );
BUFx3_ASAP7_75t_L g1145 ( .A(n_1069), .Y(n_1145) );
BUFx2_ASAP7_75t_L g1146 ( .A(n_1101), .Y(n_1146) );
NAND2xp5_ASAP7_75t_L g1147 ( .A(n_1061), .B(n_999), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_1052), .B(n_1019), .Y(n_1148) );
AND2x4_ASAP7_75t_L g1149 ( .A(n_1140), .B(n_1104), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1113), .Y(n_1150) );
HB1xp67_ASAP7_75t_L g1151 ( .A(n_1126), .Y(n_1151) );
OR2x2_ASAP7_75t_L g1152 ( .A(n_1139), .B(n_1100), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_1108), .B(n_1052), .Y(n_1153) );
OR2x2_ASAP7_75t_L g1154 ( .A(n_1139), .B(n_1100), .Y(n_1154) );
INVx2_ASAP7_75t_L g1155 ( .A(n_1117), .Y(n_1155) );
HB1xp67_ASAP7_75t_L g1156 ( .A(n_1146), .Y(n_1156) );
OR2x2_ASAP7_75t_L g1157 ( .A(n_1137), .B(n_1051), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1113), .Y(n_1158) );
HB1xp67_ASAP7_75t_L g1159 ( .A(n_1146), .Y(n_1159) );
NAND2xp5_ASAP7_75t_L g1160 ( .A(n_1108), .B(n_1072), .Y(n_1160) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1115), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1116), .B(n_1057), .Y(n_1162) );
INVx2_ASAP7_75t_SL g1163 ( .A(n_1145), .Y(n_1163) );
OAI21x1_ASAP7_75t_L g1164 ( .A1(n_1141), .A2(n_1037), .B(n_1047), .Y(n_1164) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1115), .Y(n_1165) );
AND2x4_ASAP7_75t_SL g1166 ( .A(n_1131), .B(n_1078), .Y(n_1166) );
BUFx2_ASAP7_75t_L g1167 ( .A(n_1131), .Y(n_1167) );
OR2x2_ASAP7_75t_L g1168 ( .A(n_1116), .B(n_1051), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1118), .B(n_1057), .Y(n_1169) );
NOR2xp33_ASAP7_75t_L g1170 ( .A(n_1109), .B(n_1040), .Y(n_1170) );
NAND2xp5_ASAP7_75t_L g1171 ( .A(n_1121), .B(n_1072), .Y(n_1171) );
NAND2xp5_ASAP7_75t_L g1172 ( .A(n_1121), .B(n_1068), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1124), .Y(n_1173) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1124), .Y(n_1174) );
INVx2_ASAP7_75t_SL g1175 ( .A(n_1145), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1118), .B(n_1068), .Y(n_1176) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1125), .Y(n_1177) );
NAND2xp5_ASAP7_75t_L g1178 ( .A(n_1125), .B(n_1103), .Y(n_1178) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1127), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1128), .B(n_1101), .Y(n_1180) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1127), .Y(n_1181) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1129), .Y(n_1182) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_1130), .B(n_1103), .Y(n_1183) );
OR2x2_ASAP7_75t_L g1184 ( .A(n_1135), .B(n_1092), .Y(n_1184) );
INVx1_ASAP7_75t_SL g1185 ( .A(n_1131), .Y(n_1185) );
INVx4_ASAP7_75t_L g1186 ( .A(n_1109), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1153), .B(n_1134), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1150), .Y(n_1188) );
INVx2_ASAP7_75t_L g1189 ( .A(n_1155), .Y(n_1189) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1150), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1153), .B(n_1134), .Y(n_1191) );
NAND2xp5_ASAP7_75t_L g1192 ( .A(n_1176), .B(n_1111), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1162), .B(n_1169), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1162), .B(n_1138), .Y(n_1194) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1158), .Y(n_1195) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1158), .Y(n_1196) );
NOR2xp67_ASAP7_75t_SL g1197 ( .A(n_1167), .B(n_1081), .Y(n_1197) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1161), .Y(n_1198) );
INVx2_ASAP7_75t_L g1199 ( .A(n_1155), .Y(n_1199) );
HB1xp67_ASAP7_75t_L g1200 ( .A(n_1159), .Y(n_1200) );
NAND2x1_ASAP7_75t_L g1201 ( .A(n_1186), .B(n_1087), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1161), .Y(n_1202) );
AND2x4_ASAP7_75t_L g1203 ( .A(n_1167), .B(n_1142), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1204 ( .A(n_1169), .B(n_1138), .Y(n_1204) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1165), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1165), .Y(n_1206) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1173), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1176), .B(n_1120), .Y(n_1208) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1173), .Y(n_1209) );
INVx2_ASAP7_75t_SL g1210 ( .A(n_1166), .Y(n_1210) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_1151), .B(n_1160), .Y(n_1211) );
INVxp67_ASAP7_75t_L g1212 ( .A(n_1170), .Y(n_1212) );
OR2x2_ASAP7_75t_L g1213 ( .A(n_1152), .B(n_1132), .Y(n_1213) );
NAND2xp5_ASAP7_75t_L g1214 ( .A(n_1160), .B(n_1114), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1180), .B(n_1120), .Y(n_1215) );
HB1xp67_ASAP7_75t_L g1216 ( .A(n_1159), .Y(n_1216) );
NAND2xp5_ASAP7_75t_L g1217 ( .A(n_1168), .B(n_1110), .Y(n_1217) );
OR2x2_ASAP7_75t_L g1218 ( .A(n_1152), .B(n_1148), .Y(n_1218) );
NOR2xp33_ASAP7_75t_L g1219 ( .A(n_1186), .B(n_1112), .Y(n_1219) );
INVx2_ASAP7_75t_SL g1220 ( .A(n_1210), .Y(n_1220) );
OR2x2_ASAP7_75t_L g1221 ( .A(n_1218), .B(n_1154), .Y(n_1221) );
A2O1A1Ixp33_ASAP7_75t_L g1222 ( .A1(n_1219), .A2(n_1166), .B(n_1136), .C(n_1069), .Y(n_1222) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1213), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1213), .Y(n_1224) );
AOI222xp33_ASAP7_75t_L g1225 ( .A1(n_1212), .A2(n_1062), .B1(n_1079), .B2(n_1094), .C1(n_1186), .C2(n_1070), .Y(n_1225) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1218), .Y(n_1226) );
NAND2xp5_ASAP7_75t_L g1227 ( .A(n_1193), .B(n_1156), .Y(n_1227) );
AOI22xp5_ASAP7_75t_L g1228 ( .A1(n_1210), .A2(n_1186), .B1(n_1122), .B2(n_1133), .Y(n_1228) );
AOI221xp5_ASAP7_75t_L g1229 ( .A1(n_1211), .A2(n_1065), .B1(n_1172), .B2(n_1171), .C(n_1056), .Y(n_1229) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1188), .Y(n_1230) );
OAI21xp5_ASAP7_75t_L g1231 ( .A1(n_1197), .A2(n_1185), .B(n_1075), .Y(n_1231) );
OR2x2_ASAP7_75t_L g1232 ( .A(n_1217), .B(n_1154), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g1233 ( .A(n_1193), .B(n_1168), .Y(n_1233) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1188), .Y(n_1234) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1190), .Y(n_1235) );
AOI21xp33_ASAP7_75t_L g1236 ( .A1(n_1201), .A2(n_1046), .B(n_1098), .Y(n_1236) );
OR2x2_ASAP7_75t_L g1237 ( .A(n_1187), .B(n_1157), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1208), .B(n_1166), .Y(n_1238) );
OAI21xp5_ASAP7_75t_L g1239 ( .A1(n_1197), .A2(n_1185), .B(n_1067), .Y(n_1239) );
A2O1A1Ixp33_ASAP7_75t_L g1240 ( .A1(n_1201), .A2(n_1175), .B(n_1163), .C(n_1133), .Y(n_1240) );
OAI32xp33_ASAP7_75t_L g1241 ( .A1(n_1200), .A2(n_1184), .A3(n_1157), .B1(n_1175), .B2(n_1163), .Y(n_1241) );
AOI22xp5_ASAP7_75t_L g1242 ( .A1(n_1192), .A2(n_1122), .B1(n_1058), .B2(n_1180), .Y(n_1242) );
OAI22xp5_ASAP7_75t_L g1243 ( .A1(n_1203), .A2(n_1163), .B1(n_1175), .B2(n_1184), .Y(n_1243) );
NOR3xp33_ASAP7_75t_L g1244 ( .A(n_1241), .B(n_1075), .C(n_1024), .Y(n_1244) );
OAI22xp5_ASAP7_75t_L g1245 ( .A1(n_1228), .A2(n_1203), .B1(n_1208), .B2(n_1214), .Y(n_1245) );
AOI22xp5_ASAP7_75t_L g1246 ( .A1(n_1242), .A2(n_1203), .B1(n_1215), .B2(n_1216), .Y(n_1246) );
AOI22xp5_ASAP7_75t_L g1247 ( .A1(n_1225), .A2(n_1215), .B1(n_1187), .B2(n_1204), .Y(n_1247) );
NOR3xp33_ASAP7_75t_L g1248 ( .A(n_1231), .B(n_1091), .C(n_1098), .Y(n_1248) );
OAI32xp33_ASAP7_75t_L g1249 ( .A1(n_1243), .A2(n_1191), .A3(n_1194), .B1(n_1204), .B2(n_1172), .Y(n_1249) );
OAI221xp5_ASAP7_75t_L g1250 ( .A1(n_1240), .A2(n_1053), .B1(n_1171), .B2(n_1206), .C(n_1207), .Y(n_1250) );
OAI22xp5_ASAP7_75t_L g1251 ( .A1(n_1222), .A2(n_1194), .B1(n_1191), .B2(n_1081), .Y(n_1251) );
AOI22xp5_ASAP7_75t_L g1252 ( .A1(n_1225), .A2(n_1119), .B1(n_1120), .B2(n_1209), .Y(n_1252) );
OAI322xp33_ASAP7_75t_L g1253 ( .A1(n_1223), .A2(n_1209), .A3(n_1207), .B1(n_1206), .B2(n_1205), .C1(n_1202), .C2(n_1195), .Y(n_1253) );
OAI221xp5_ASAP7_75t_L g1254 ( .A1(n_1239), .A2(n_1205), .B1(n_1196), .B2(n_1202), .C(n_1198), .Y(n_1254) );
OAI22xp5_ASAP7_75t_L g1255 ( .A1(n_1220), .A2(n_1123), .B1(n_1028), .B2(n_1002), .Y(n_1255) );
A2O1A1Ixp33_ASAP7_75t_L g1256 ( .A1(n_1238), .A2(n_1005), .B(n_1123), .C(n_1074), .Y(n_1256) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1221), .Y(n_1257) );
AOI22xp5_ASAP7_75t_L g1258 ( .A1(n_1229), .A2(n_1119), .B1(n_1190), .B2(n_1198), .Y(n_1258) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1237), .Y(n_1259) );
A2O1A1Ixp33_ASAP7_75t_L g1260 ( .A1(n_1236), .A2(n_1231), .B(n_1233), .C(n_1227), .Y(n_1260) );
OAI22xp5_ASAP7_75t_L g1261 ( .A1(n_1247), .A2(n_1224), .B1(n_1226), .B2(n_1232), .Y(n_1261) );
NAND4xp25_ASAP7_75t_L g1262 ( .A(n_1255), .B(n_1074), .C(n_1014), .D(n_1086), .Y(n_1262) );
AOI22xp5_ASAP7_75t_L g1263 ( .A1(n_1252), .A2(n_1235), .B1(n_1230), .B2(n_1234), .Y(n_1263) );
NAND3xp33_ASAP7_75t_L g1264 ( .A(n_1260), .B(n_1196), .C(n_1195), .Y(n_1264) );
NOR4xp25_ASAP7_75t_L g1265 ( .A(n_1254), .B(n_1023), .C(n_1020), .D(n_1004), .Y(n_1265) );
AOI21xp5_ASAP7_75t_L g1266 ( .A1(n_1249), .A2(n_1087), .B(n_1178), .Y(n_1266) );
AOI222xp33_ASAP7_75t_L g1267 ( .A1(n_1245), .A2(n_1010), .B1(n_1022), .B2(n_1147), .C1(n_1181), .C2(n_1179), .Y(n_1267) );
OAI211xp5_ASAP7_75t_L g1268 ( .A1(n_1246), .A2(n_1003), .B(n_1011), .C(n_985), .Y(n_1268) );
OAI21xp5_ASAP7_75t_L g1269 ( .A1(n_1244), .A2(n_1080), .B(n_1083), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1259), .B(n_1149), .Y(n_1270) );
OAI221xp5_ASAP7_75t_L g1271 ( .A1(n_1258), .A2(n_1178), .B1(n_1183), .B2(n_1182), .C(n_1174), .Y(n_1271) );
AOI21xp5_ASAP7_75t_L g1272 ( .A1(n_1251), .A2(n_1183), .B(n_1189), .Y(n_1272) );
NOR2x1_ASAP7_75t_L g1273 ( .A(n_1264), .B(n_1268), .Y(n_1273) );
OAI221xp5_ASAP7_75t_L g1274 ( .A1(n_1265), .A2(n_1248), .B1(n_1250), .B2(n_1256), .C(n_1257), .Y(n_1274) );
NOR3xp33_ASAP7_75t_L g1275 ( .A(n_1261), .B(n_1253), .C(n_1010), .Y(n_1275) );
A2O1A1Ixp33_ASAP7_75t_L g1276 ( .A1(n_1263), .A2(n_1266), .B(n_1272), .C(n_1269), .Y(n_1276) );
NAND4xp25_ASAP7_75t_L g1277 ( .A(n_1267), .B(n_981), .C(n_1082), .D(n_1083), .Y(n_1277) );
AOI21xp5_ASAP7_75t_L g1278 ( .A1(n_1271), .A2(n_1199), .B(n_1189), .Y(n_1278) );
NOR4xp25_ASAP7_75t_L g1279 ( .A(n_1262), .B(n_1027), .C(n_1007), .D(n_1028), .Y(n_1279) );
O2A1O1Ixp33_ASAP7_75t_L g1280 ( .A1(n_1270), .A2(n_1034), .B(n_1038), .C(n_1016), .Y(n_1280) );
NAND4xp75_ASAP7_75t_L g1281 ( .A(n_1273), .B(n_1093), .C(n_1076), .D(n_1077), .Y(n_1281) );
NAND4xp25_ASAP7_75t_L g1282 ( .A(n_1276), .B(n_1277), .C(n_1274), .D(n_1275), .Y(n_1282) );
NOR2x1_ASAP7_75t_L g1283 ( .A(n_1279), .B(n_1005), .Y(n_1283) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1280), .Y(n_1284) );
NOR3xp33_ASAP7_75t_L g1285 ( .A(n_1278), .B(n_981), .C(n_1017), .Y(n_1285) );
NAND3xp33_ASAP7_75t_L g1286 ( .A(n_1273), .B(n_1177), .C(n_1174), .Y(n_1286) );
INVx2_ASAP7_75t_L g1287 ( .A(n_1281), .Y(n_1287) );
NAND2xp5_ASAP7_75t_L g1288 ( .A(n_1284), .B(n_1177), .Y(n_1288) );
INVx2_ASAP7_75t_L g1289 ( .A(n_1283), .Y(n_1289) );
AND4x1_ASAP7_75t_L g1290 ( .A(n_1286), .B(n_1082), .C(n_1143), .D(n_1144), .Y(n_1290) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1288), .Y(n_1291) );
NOR2xp67_ASAP7_75t_L g1292 ( .A(n_1289), .B(n_1282), .Y(n_1292) );
HB1xp67_ASAP7_75t_L g1293 ( .A(n_1287), .Y(n_1293) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1290), .Y(n_1294) );
AOI22xp5_ASAP7_75t_L g1295 ( .A1(n_1292), .A2(n_1285), .B1(n_983), .B2(n_979), .Y(n_1295) );
NOR2xp33_ASAP7_75t_L g1296 ( .A(n_1293), .B(n_1013), .Y(n_1296) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1291), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1297), .Y(n_1298) );
INVx2_ASAP7_75t_L g1299 ( .A(n_1296), .Y(n_1299) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1295), .Y(n_1300) );
OA21x2_ASAP7_75t_L g1301 ( .A1(n_1298), .A2(n_1291), .B(n_1294), .Y(n_1301) );
AOI22xp5_ASAP7_75t_L g1302 ( .A1(n_1300), .A2(n_1013), .B1(n_1007), .B2(n_1027), .Y(n_1302) );
AOI22x1_ASAP7_75t_L g1303 ( .A1(n_1299), .A2(n_1013), .B1(n_992), .B2(n_1017), .Y(n_1303) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_1301), .B(n_1299), .Y(n_1304) );
BUFx2_ASAP7_75t_L g1305 ( .A(n_1302), .Y(n_1305) );
OAI22xp5_ASAP7_75t_L g1306 ( .A1(n_1303), .A2(n_1092), .B1(n_999), .B2(n_998), .Y(n_1306) );
AO21x2_ASAP7_75t_L g1307 ( .A1(n_1304), .A2(n_1095), .B(n_1179), .Y(n_1307) );
AO21x2_ASAP7_75t_L g1308 ( .A1(n_1305), .A2(n_1181), .B(n_1182), .Y(n_1308) );
OAI21xp5_ASAP7_75t_L g1309 ( .A1(n_1306), .A2(n_998), .B(n_1164), .Y(n_1309) );
OAI21xp5_ASAP7_75t_L g1310 ( .A1(n_1309), .A2(n_1077), .B(n_1076), .Y(n_1310) );
AOI22xp33_ASAP7_75t_L g1311 ( .A1(n_1310), .A2(n_1307), .B1(n_1308), .B2(n_1149), .Y(n_1311) );
endmodule