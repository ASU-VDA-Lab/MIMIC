module fake_jpeg_31995_n_138 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_138);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_138;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_6),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_8),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_28),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_61),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_1),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_62),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_2),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_2),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_55),
.A2(n_45),
.B1(n_48),
.B2(n_40),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_42),
.B1(n_43),
.B2(n_54),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_66),
.B1(n_68),
.B2(n_71),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_67),
.B(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_59),
.B(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_62),
.B(n_52),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_74),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_48),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_62),
.B(n_47),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_76),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_39),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_74),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_79),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_63),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_72),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_81),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_83),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_44),
.B(n_38),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_89),
.Y(n_99)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_45),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_45),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_94),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_3),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_88),
.A2(n_18),
.B1(n_36),
.B2(n_35),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_95),
.A2(n_97),
.B1(n_100),
.B2(n_7),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_88),
.A2(n_17),
.B1(n_32),
.B2(n_30),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_14),
.C(n_29),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_107),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_86),
.B(n_4),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_105),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_81),
.B(n_5),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_6),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_96),
.A2(n_82),
.B1(n_8),
.B2(n_7),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_109),
.A2(n_110),
.B1(n_116),
.B2(n_95),
.Y(n_121)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_111),
.B(n_112),
.Y(n_126)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_99),
.B(n_9),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_114),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_103),
.B(n_37),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_97),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_106),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_100),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_121),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_110),
.A2(n_108),
.B1(n_98),
.B2(n_23),
.Y(n_122)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_124),
.A2(n_109),
.B1(n_116),
.B2(n_115),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_129),
.A2(n_123),
.B1(n_126),
.B2(n_124),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_130),
.A2(n_131),
.B(n_128),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_118),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_132),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_125),
.C(n_117),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_13),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_15),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);


endmodule