module fake_jpeg_13047_n_517 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_517);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_517;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_293;
wire n_38;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_352;
wire n_350;
wire n_150;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_3),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx4f_ASAP7_75t_SL g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_52),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_22),
.B(n_15),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_53),
.B(n_63),
.Y(n_113)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_26),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_54),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx11_ASAP7_75t_L g150 ( 
.A(n_57),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_62),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_22),
.B(n_13),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_67),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_68),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_28),
.B(n_13),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_69),
.B(n_83),
.Y(n_139)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_72),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_73),
.Y(n_111)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_74),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_76),
.Y(n_149)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_16),
.Y(n_77)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_16),
.Y(n_78)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_18),
.B(n_12),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_27),
.Y(n_104)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_16),
.Y(n_81)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_31),
.B(n_12),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_35),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_89),
.A2(n_30),
.B1(n_23),
.B2(n_46),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_90),
.A2(n_27),
.B1(n_30),
.B2(n_34),
.Y(n_124)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_91),
.Y(n_151)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_93),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_97),
.B(n_98),
.Y(n_145)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_21),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_18),
.B(n_0),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_99),
.B(n_1),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_104),
.B(n_109),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_61),
.A2(n_21),
.B1(n_19),
.B2(n_39),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_105),
.A2(n_118),
.B1(n_133),
.B2(n_134),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_31),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_86),
.B(n_40),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_131),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_60),
.A2(n_19),
.B1(n_39),
.B2(n_48),
.Y(n_118)
);

NAND2x1_ASAP7_75t_L g194 ( 
.A(n_124),
.B(n_41),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_72),
.B(n_42),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_132),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_88),
.B(n_40),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_73),
.B(n_42),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_93),
.A2(n_19),
.B1(n_39),
.B2(n_48),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_76),
.B(n_49),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_143),
.Y(n_175)
);

AND2x4_ASAP7_75t_L g141 ( 
.A(n_89),
.B(n_50),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_51),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_87),
.B(n_49),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_147),
.B(n_153),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_52),
.B(n_34),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_159),
.B(n_190),
.Y(n_218)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_160),
.B(n_165),
.Y(n_226)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_115),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_164),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_145),
.Y(n_165)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_166),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_120),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_167),
.Y(n_221)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_103),
.Y(n_168)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_168),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_134),
.A2(n_79),
.B1(n_62),
.B2(n_141),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_169),
.A2(n_97),
.B1(n_50),
.B2(n_142),
.Y(n_237)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_170),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_81),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_171),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_121),
.A2(n_59),
.B1(n_70),
.B2(n_48),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_172),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_145),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_173),
.B(n_177),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_121),
.A2(n_50),
.B1(n_96),
.B2(n_94),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_174),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_122),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_176),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_110),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_113),
.B(n_46),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_178),
.B(n_192),
.Y(n_234)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_123),
.Y(n_180)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_77),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_181),
.Y(n_209)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_123),
.Y(n_182)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_182),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_129),
.Y(n_183)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_149),
.Y(n_185)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_186),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_136),
.Y(n_187)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_187),
.Y(n_240)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_119),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_188),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_125),
.Y(n_189)
);

INVx4_ASAP7_75t_SL g211 ( 
.A(n_189),
.Y(n_211)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_148),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_191),
.B(n_193),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_139),
.B(n_44),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_194),
.B(n_205),
.Y(n_231)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_196),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_102),
.B(n_44),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_197),
.B(n_206),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_107),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_137),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_125),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_137),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_201),
.B(n_202),
.Y(n_235)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_157),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_141),
.A2(n_64),
.B1(n_84),
.B2(n_82),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_203),
.A2(n_65),
.B1(n_55),
.B2(n_56),
.Y(n_228)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_138),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_118),
.Y(n_206)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_152),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_207),
.B(n_106),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_206),
.A2(n_141),
.B(n_117),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_216),
.A2(n_100),
.B(n_142),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_194),
.A2(n_105),
.B1(n_133),
.B2(n_108),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_219),
.A2(n_237),
.B1(n_239),
.B2(n_242),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_195),
.B(n_57),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_241),
.C(n_175),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_228),
.A2(n_126),
.B1(n_200),
.B2(n_166),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_229),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_159),
.A2(n_108),
.B1(n_75),
.B2(n_67),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_163),
.B(n_128),
.C(n_130),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_159),
.A2(n_112),
.B1(n_144),
.B2(n_155),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_161),
.A2(n_112),
.B1(n_144),
.B2(n_155),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_243),
.A2(n_126),
.B1(n_167),
.B2(n_189),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_248),
.B(n_213),
.Y(n_318)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_249),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_181),
.C(n_171),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_250),
.B(n_254),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_251),
.A2(n_233),
.B1(n_228),
.B2(n_209),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_216),
.A2(n_164),
.B(n_183),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_252),
.A2(n_267),
.B(n_273),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_178),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_192),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_255),
.B(n_261),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_256),
.A2(n_246),
.B1(n_221),
.B2(n_240),
.Y(n_299)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_235),
.Y(n_257)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_257),
.Y(n_288)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_236),
.Y(n_258)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_258),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_236),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_259),
.B(n_269),
.Y(n_305)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_260),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_158),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_214),
.B(n_204),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_262),
.B(n_264),
.Y(n_310)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_236),
.Y(n_263)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_263),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_214),
.B(n_205),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_208),
.Y(n_265)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_265),
.Y(n_306)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_230),
.Y(n_266)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_266),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_219),
.A2(n_171),
.B1(n_181),
.B2(n_129),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_231),
.B(n_193),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_268),
.B(n_279),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_229),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_231),
.A2(n_101),
.B1(n_156),
.B2(n_162),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_270),
.A2(n_242),
.B1(n_239),
.B2(n_243),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_226),
.B(n_202),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_271),
.B(n_278),
.Y(n_303)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_211),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_272),
.B(n_280),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_225),
.A2(n_185),
.B(n_187),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_230),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_275),
.B(n_276),
.Y(n_314)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_224),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_277),
.A2(n_282),
.B(n_273),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_241),
.B(n_196),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_218),
.B(n_168),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_224),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_218),
.B(n_170),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_281),
.B(n_284),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_238),
.A2(n_23),
.B(n_176),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_244),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_283),
.B(n_213),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_218),
.B(n_188),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_271),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_285),
.B(n_291),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_286),
.A2(n_298),
.B1(n_299),
.B2(n_302),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_253),
.A2(n_247),
.B1(n_218),
.B2(n_209),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_289),
.A2(n_277),
.B(n_267),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_268),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_295),
.A2(n_309),
.B1(n_317),
.B2(n_256),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_283),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_297),
.B(n_300),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_249),
.A2(n_237),
.B1(n_247),
.B2(n_232),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_282),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_257),
.A2(n_232),
.B1(n_217),
.B2(n_210),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_252),
.A2(n_217),
.B1(n_210),
.B2(n_246),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_304),
.A2(n_307),
.B1(n_212),
.B2(n_215),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_252),
.A2(n_246),
.B1(n_240),
.B2(n_244),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_274),
.A2(n_226),
.B1(n_245),
.B2(n_221),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_284),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_311),
.B(n_272),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_315),
.A2(n_266),
.B(n_272),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_274),
.A2(n_245),
.B1(n_221),
.B2(n_101),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_278),
.C(n_250),
.Y(n_326)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_319),
.Y(n_321)
);

OAI21xp33_ASAP7_75t_L g320 ( 
.A1(n_289),
.A2(n_262),
.B(n_264),
.Y(n_320)
);

NAND3xp33_ASAP7_75t_L g381 ( 
.A(n_320),
.B(n_343),
.C(n_335),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_313),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_322),
.B(n_328),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_301),
.B(n_248),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_323),
.B(n_326),
.C(n_327),
.Y(n_361)
);

AND2x2_ASAP7_75t_SL g325 ( 
.A(n_304),
.B(n_248),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_325),
.A2(n_351),
.B(n_222),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_301),
.B(n_254),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_313),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_314),
.Y(n_329)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_329),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_254),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_330),
.B(n_337),
.C(n_338),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_314),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_331),
.B(n_345),
.Y(n_370)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_319),
.Y(n_333)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_333),
.Y(n_367)
);

OAI221xp5_ASAP7_75t_L g334 ( 
.A1(n_294),
.A2(n_261),
.B1(n_255),
.B2(n_259),
.C(n_263),
.Y(n_334)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_334),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_335),
.B(n_336),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_294),
.B(n_250),
.C(n_277),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_310),
.B(n_260),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_310),
.B(n_269),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_339),
.B(n_287),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_308),
.B(n_312),
.C(n_292),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_340),
.B(n_344),
.C(n_346),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_309),
.A2(n_253),
.B1(n_256),
.B2(n_274),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_342),
.B(n_349),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_305),
.B(n_275),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_308),
.B(n_258),
.C(n_267),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_313),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_312),
.B(n_281),
.C(n_279),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_305),
.B(n_270),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_347),
.B(n_348),
.C(n_223),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_287),
.B(n_270),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_317),
.A2(n_273),
.B1(n_282),
.B2(n_251),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_300),
.A2(n_251),
.B1(n_276),
.B2(n_280),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_350),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_352),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_292),
.A2(n_265),
.B1(n_215),
.B2(n_212),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_353),
.B(n_296),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_354),
.A2(n_324),
.B1(n_295),
.B2(n_293),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_355),
.B(n_339),
.Y(n_393)
);

OA21x2_ASAP7_75t_L g356 ( 
.A1(n_332),
.A2(n_307),
.B(n_315),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_356),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_357),
.A2(n_360),
.B1(n_362),
.B2(n_366),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_332),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_359),
.B(n_374),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_325),
.A2(n_291),
.B1(n_288),
.B2(n_303),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_325),
.A2(n_288),
.B1(n_303),
.B2(n_311),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_321),
.A2(n_285),
.B1(n_293),
.B2(n_290),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_327),
.B(n_296),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_368),
.B(n_375),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_321),
.B(n_297),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_372),
.B(n_347),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_323),
.B(n_290),
.Y(n_375)
);

NOR2xp67_ASAP7_75t_L g376 ( 
.A(n_333),
.B(n_302),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_376),
.B(n_381),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_329),
.A2(n_316),
.B1(n_286),
.B2(n_298),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_377),
.A2(n_378),
.B1(n_371),
.B2(n_373),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_352),
.A2(n_316),
.B1(n_306),
.B2(n_222),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_341),
.B(n_306),
.Y(n_379)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_379),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_382),
.B(n_346),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_330),
.B(n_326),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_383),
.B(n_384),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_340),
.B(n_149),
.Y(n_384)
);

XOR2x2_ASAP7_75t_L g389 ( 
.A(n_385),
.B(n_353),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_338),
.B(n_223),
.Y(n_386)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_386),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_367),
.Y(n_388)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_388),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_389),
.A2(n_403),
.B(n_363),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_390),
.B(n_412),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_369),
.A2(n_336),
.B1(n_342),
.B2(n_344),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_391),
.A2(n_400),
.B1(n_365),
.B2(n_358),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_393),
.B(n_414),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_361),
.B(n_384),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_394),
.B(n_405),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g397 ( 
.A(n_366),
.B(n_350),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_397),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_361),
.B(n_383),
.C(n_364),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_398),
.B(n_406),
.C(n_382),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_357),
.A2(n_349),
.B1(n_337),
.B2(n_351),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_402),
.B(n_404),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_363),
.B(n_348),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_387),
.B(n_222),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_364),
.B(n_220),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_380),
.B(n_220),
.C(n_208),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_370),
.B(n_201),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_407),
.B(n_411),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_408),
.A2(n_358),
.B1(n_363),
.B2(n_356),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_371),
.A2(n_100),
.B1(n_199),
.B2(n_182),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_410),
.A2(n_377),
.B1(n_378),
.B2(n_385),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_380),
.B(n_207),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_375),
.B(n_128),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_413),
.B(n_415),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_368),
.B(n_190),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_355),
.B(n_211),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_417),
.B(n_420),
.C(n_437),
.Y(n_447)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_418),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_412),
.B(n_362),
.C(n_360),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_421),
.A2(n_41),
.B1(n_47),
.B2(n_16),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_422),
.B(n_431),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_401),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_425),
.B(n_435),
.Y(n_457)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_427),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_416),
.B(n_356),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_430),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_397),
.A2(n_211),
.B1(n_17),
.B2(n_180),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_432),
.B(n_433),
.Y(n_453)
);

OAI22x1_ASAP7_75t_L g433 ( 
.A1(n_399),
.A2(n_156),
.B1(n_130),
.B2(n_150),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_433),
.A2(n_439),
.B1(n_17),
.B2(n_41),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_398),
.B(n_111),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_434),
.B(n_436),
.Y(n_440)
);

FAx1_ASAP7_75t_SL g435 ( 
.A(n_393),
.B(n_399),
.CI(n_415),
.CON(n_435),
.SN(n_435)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_394),
.B(n_111),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_405),
.B(n_150),
.C(n_37),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_392),
.A2(n_389),
.B1(n_403),
.B2(n_414),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_419),
.B(n_409),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_SL g464 ( 
.A(n_441),
.B(n_424),
.Y(n_464)
);

OAI221xp5_ASAP7_75t_L g443 ( 
.A1(n_423),
.A2(n_396),
.B1(n_406),
.B2(n_390),
.C(n_395),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_443),
.A2(n_446),
.B1(n_33),
.B2(n_4),
.Y(n_472)
);

OAI221xp5_ASAP7_75t_L g446 ( 
.A1(n_438),
.A2(n_395),
.B1(n_409),
.B2(n_413),
.C(n_410),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_417),
.B(n_37),
.C(n_38),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_448),
.B(n_450),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_421),
.A2(n_136),
.B(n_38),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_449),
.A2(n_451),
.B(n_452),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_428),
.B(n_74),
.C(n_45),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_439),
.A2(n_33),
.B(n_54),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_420),
.A2(n_418),
.B(n_435),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_SL g465 ( 
.A1(n_453),
.A2(n_436),
.B1(n_429),
.B2(n_434),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_428),
.B(n_74),
.C(n_47),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_454),
.B(n_441),
.C(n_419),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_455),
.A2(n_458),
.B1(n_432),
.B2(n_426),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_459),
.A2(n_462),
.B1(n_465),
.B2(n_475),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_424),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_460),
.B(n_466),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_442),
.A2(n_437),
.B1(n_435),
.B2(n_429),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_463),
.B(n_464),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_444),
.B(n_47),
.Y(n_466)
);

OAI21xp33_ASAP7_75t_SL g467 ( 
.A1(n_442),
.A2(n_33),
.B(n_4),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_467),
.B(n_451),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_444),
.B(n_47),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_469),
.B(n_471),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_447),
.B(n_47),
.C(n_4),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_470),
.B(n_448),
.C(n_440),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_456),
.B(n_3),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_472),
.A2(n_458),
.B1(n_450),
.B2(n_449),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_445),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_473),
.B(n_5),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_457),
.A2(n_3),
.B(n_5),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_474),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_453),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g496 ( 
.A(n_476),
.B(n_11),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_477),
.B(n_479),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_460),
.B(n_456),
.C(n_452),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_481),
.B(n_482),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_464),
.B(n_440),
.C(n_454),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_483),
.A2(n_463),
.B(n_461),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_459),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_485),
.B(n_487),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_475),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_486),
.B(n_489),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_461),
.B(n_6),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_491),
.A2(n_492),
.B(n_499),
.Y(n_507)
);

OAI21x1_ASAP7_75t_L g492 ( 
.A1(n_488),
.A2(n_468),
.B(n_474),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_481),
.B(n_462),
.C(n_470),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_493),
.B(n_495),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_480),
.B(n_6),
.C(n_7),
.Y(n_495)
);

INVxp33_ASAP7_75t_L g503 ( 
.A(n_496),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_498),
.A2(n_500),
.B(n_476),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_478),
.B(n_6),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_483),
.A2(n_7),
.B(n_8),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_494),
.A2(n_484),
.B(n_477),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_501),
.A2(n_506),
.B(n_496),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_497),
.B(n_487),
.C(n_489),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_502),
.B(n_495),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_505),
.Y(n_510)
);

OAI21xp33_ASAP7_75t_L g506 ( 
.A1(n_493),
.A2(n_479),
.B(n_9),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_508),
.B(n_509),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_507),
.B(n_490),
.C(n_8),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_511),
.A2(n_503),
.B(n_504),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_512),
.A2(n_510),
.B(n_8),
.Y(n_514)
);

BUFx24_ASAP7_75t_SL g515 ( 
.A(n_514),
.Y(n_515)
);

AOI21x1_ASAP7_75t_L g516 ( 
.A1(n_515),
.A2(n_513),
.B(n_11),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_11),
.Y(n_517)
);


endmodule