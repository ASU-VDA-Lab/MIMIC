module fake_jpeg_14425_n_601 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_601);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_601;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_2),
.B(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_15),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_15),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

BUFx4f_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_57),
.Y(n_147)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_58),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_22),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_59),
.B(n_71),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

AND2x4_ASAP7_75t_SL g63 ( 
.A(n_21),
.B(n_1),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_63),
.B(n_87),
.Y(n_130)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx11_ASAP7_75t_L g171 ( 
.A(n_64),
.Y(n_171)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_65),
.Y(n_191)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_66),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_67),
.Y(n_127)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_27),
.B(n_10),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_69),
.B(n_75),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g175 ( 
.A(n_70),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_22),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_73),
.B(n_78),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_27),
.B(n_10),
.Y(n_75)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_76),
.Y(n_169)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_22),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_25),
.B(n_14),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_79),
.B(n_110),
.Y(n_150)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_80),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_22),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_81),
.B(n_84),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_82),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_85),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_22),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_86),
.B(n_89),
.Y(n_166)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_47),
.B(n_2),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g185 ( 
.A(n_88),
.Y(n_185)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_40),
.A2(n_9),
.B1(n_3),
.B2(n_4),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_90),
.A2(n_49),
.B1(n_51),
.B2(n_45),
.Y(n_161)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_23),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_91),
.B(n_92),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_21),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_21),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_93),
.B(n_94),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_25),
.B(n_36),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

BUFx12_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_51),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_97),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_98),
.Y(n_187)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_99),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_100),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_102),
.Y(n_193)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_24),
.Y(n_103)
);

INVx3_ASAP7_75t_SL g181 ( 
.A(n_103),
.Y(n_181)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

BUFx4f_ASAP7_75t_SL g105 ( 
.A(n_48),
.Y(n_105)
);

INVx5_ASAP7_75t_SL g179 ( 
.A(n_105),
.Y(n_179)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_21),
.Y(n_106)
);

INVx11_ASAP7_75t_L g194 ( 
.A(n_106),
.Y(n_194)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

INVx3_ASAP7_75t_SL g108 ( 
.A(n_16),
.Y(n_108)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_108),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_33),
.Y(n_109)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_29),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_37),
.Y(n_112)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_112),
.Y(n_168)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_28),
.Y(n_113)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_114),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_37),
.Y(n_115)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_115),
.Y(n_197)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_24),
.Y(n_116)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_47),
.B(n_11),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_2),
.Y(n_153)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_24),
.Y(n_118)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_119),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_29),
.Y(n_120)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_76),
.A2(n_41),
.B1(n_50),
.B2(n_16),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_124),
.A2(n_135),
.B1(n_70),
.B2(n_31),
.Y(n_251)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_129),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_97),
.A2(n_51),
.B1(n_41),
.B2(n_50),
.Y(n_135)
);

AND2x2_ASAP7_75t_SL g136 ( 
.A(n_117),
.B(n_37),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_136),
.B(n_115),
.Y(n_227)
);

BUFx10_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

INVxp67_ASAP7_75t_SL g206 ( 
.A(n_137),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_90),
.A2(n_16),
.B1(n_55),
.B2(n_41),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_141),
.A2(n_161),
.B1(n_182),
.B2(n_49),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_106),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_151),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_153),
.B(n_53),
.Y(n_240)
);

AOI21xp33_ASAP7_75t_L g160 ( 
.A1(n_63),
.A2(n_38),
.B(n_36),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_160),
.B(n_184),
.Y(n_219)
);

BUFx2_ASAP7_75t_R g164 ( 
.A(n_62),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_164),
.B(n_83),
.Y(n_266)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_67),
.Y(n_165)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_104),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_167),
.B(n_105),
.Y(n_207)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_72),
.Y(n_172)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_172),
.Y(n_217)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_68),
.Y(n_173)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_173),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_87),
.B(n_35),
.C(n_42),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_174),
.B(n_35),
.C(n_30),
.Y(n_249)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_95),
.Y(n_177)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_108),
.A2(n_63),
.B1(n_114),
.B2(n_109),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_74),
.Y(n_183)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_183),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_96),
.Y(n_184)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_121),
.Y(n_188)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_188),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_107),
.Y(n_189)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_189),
.Y(n_226)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_80),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g230 ( 
.A(n_195),
.Y(n_230)
);

INVx11_ASAP7_75t_L g199 ( 
.A(n_120),
.Y(n_199)
);

INVx11_ASAP7_75t_L g260 ( 
.A(n_199),
.Y(n_260)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_77),
.Y(n_200)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_200),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_201),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_204),
.A2(n_228),
.B1(n_241),
.B2(n_268),
.Y(n_294)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_155),
.Y(n_205)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_205),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_207),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_182),
.A2(n_87),
.B1(n_103),
.B2(n_98),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_208),
.A2(n_229),
.B1(n_247),
.B2(n_100),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_42),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_210),
.B(n_222),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_170),
.A2(n_31),
.B1(n_29),
.B2(n_54),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_211),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_186),
.Y(n_213)
);

INVx6_ASAP7_75t_L g292 ( 
.A(n_213),
.Y(n_292)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_162),
.Y(n_214)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_214),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_187),
.Y(n_215)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_215),
.Y(n_277)
);

NAND2x1p5_ASAP7_75t_L g216 ( 
.A(n_130),
.B(n_88),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_216),
.B(n_239),
.C(n_249),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_136),
.B(n_53),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_220),
.B(n_261),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_124),
.A2(n_85),
.B1(n_102),
.B2(n_116),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_221),
.A2(n_231),
.B1(n_251),
.B2(n_258),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_146),
.B(n_43),
.Y(n_222)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_122),
.Y(n_224)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_224),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_187),
.Y(n_225)
);

INVx8_ASAP7_75t_L g321 ( 
.A(n_225),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_227),
.B(n_257),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_193),
.A2(n_119),
.B1(n_118),
.B2(n_45),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_130),
.A2(n_99),
.B1(n_55),
.B2(n_50),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_150),
.A2(n_55),
.B1(n_112),
.B2(n_101),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_190),
.B(n_43),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_232),
.B(n_237),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_179),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_234),
.Y(n_320)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_147),
.Y(n_235)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_235),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_166),
.B(n_46),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_152),
.B(n_163),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_238),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_138),
.B(n_82),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_240),
.B(n_246),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_193),
.A2(n_38),
.B1(n_26),
.B2(n_52),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_156),
.Y(n_242)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_242),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_179),
.A2(n_31),
.B1(n_28),
.B2(n_54),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_243),
.A2(n_267),
.B1(n_133),
.B2(n_159),
.Y(n_276)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_181),
.Y(n_244)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_244),
.Y(n_303)
);

INVx6_ASAP7_75t_L g245 ( 
.A(n_140),
.Y(n_245)
);

INVx3_ASAP7_75t_SL g297 ( 
.A(n_245),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_131),
.B(n_52),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_181),
.A2(n_169),
.B1(n_198),
.B2(n_180),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_191),
.B(n_46),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_248),
.B(n_252),
.Y(n_315)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_129),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_250),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_189),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_169),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_253),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_126),
.Y(n_254)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_139),
.Y(n_255)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_255),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_158),
.B(n_175),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_256),
.B(n_259),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_144),
.B(n_96),
.C(n_39),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_135),
.A2(n_30),
.B1(n_39),
.B2(n_32),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_142),
.B(n_26),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_149),
.B(n_32),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_137),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_262),
.B(n_264),
.Y(n_323)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_165),
.Y(n_263)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_263),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_175),
.B(n_105),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_126),
.Y(n_265)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_265),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_266),
.B(n_185),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_123),
.A2(n_111),
.B1(n_100),
.B2(n_60),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_154),
.A2(n_56),
.B1(n_4),
.B2(n_8),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_176),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_269),
.Y(n_327)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_172),
.Y(n_270)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_270),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_175),
.B(n_111),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_271),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_239),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_274),
.B(n_300),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_221),
.A2(n_128),
.B1(n_132),
.B2(n_178),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_275),
.A2(n_282),
.B1(n_293),
.B2(n_244),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_276),
.A2(n_317),
.B1(n_234),
.B2(n_230),
.Y(n_331)
);

AOI32xp33_ASAP7_75t_L g279 ( 
.A1(n_216),
.A2(n_137),
.A3(n_194),
.B1(n_171),
.B2(n_167),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_SL g340 ( 
.A(n_279),
.B(n_195),
.C(n_143),
.Y(n_340)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_224),
.Y(n_280)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_280),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_231),
.A2(n_196),
.B1(n_151),
.B2(n_134),
.Y(n_282)
);

INVx13_ASAP7_75t_L g283 ( 
.A(n_230),
.Y(n_283)
);

INVx13_ASAP7_75t_L g329 ( 
.A(n_283),
.Y(n_329)
);

OAI22x1_ASAP7_75t_SL g284 ( 
.A1(n_204),
.A2(n_133),
.B1(n_159),
.B2(n_199),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_284),
.A2(n_314),
.B1(n_325),
.B2(n_266),
.Y(n_339)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_205),
.Y(n_287)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_287),
.Y(n_358)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_214),
.Y(n_289)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_289),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_227),
.A2(n_194),
.B1(n_171),
.B2(n_178),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_239),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_261),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_301),
.B(n_226),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_220),
.B(n_168),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_306),
.B(n_313),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_208),
.A2(n_132),
.B1(n_128),
.B2(n_127),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_311),
.B(n_312),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_227),
.B(n_197),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_219),
.A2(n_127),
.B1(n_125),
.B2(n_148),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_257),
.B(n_2),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_318),
.B(n_4),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_229),
.A2(n_125),
.B1(n_157),
.B2(n_56),
.Y(n_325)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_218),
.Y(n_328)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_328),
.Y(n_370)
);

BUFx24_ASAP7_75t_SL g330 ( 
.A(n_278),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_330),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_331),
.A2(n_308),
.B1(n_321),
.B2(n_277),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_315),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_332),
.B(n_346),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_309),
.B(n_216),
.C(n_249),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_333),
.B(n_348),
.C(n_353),
.Y(n_390)
);

INVx13_ASAP7_75t_L g334 ( 
.A(n_283),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_334),
.Y(n_395)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_295),
.Y(n_335)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_335),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_299),
.B(n_209),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_336),
.B(n_363),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_339),
.A2(n_349),
.B1(n_365),
.B2(n_312),
.Y(n_373)
);

OR2x2_ASAP7_75t_L g392 ( 
.A(n_340),
.B(n_145),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_310),
.A2(n_206),
.B1(n_230),
.B2(n_260),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_341),
.A2(n_344),
.B(n_350),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_310),
.A2(n_260),
.B1(n_236),
.B2(n_245),
.Y(n_344)
);

BUFx24_ASAP7_75t_L g345 ( 
.A(n_320),
.Y(n_345)
);

INVxp33_ASAP7_75t_L g408 ( 
.A(n_345),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_323),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_347),
.B(n_357),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_309),
.B(n_223),
.Y(n_348)
);

OAI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_281),
.A2(n_247),
.B1(n_236),
.B2(n_263),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_312),
.A2(n_233),
.B(n_212),
.Y(n_350)
);

AND2x6_ASAP7_75t_L g351 ( 
.A(n_285),
.B(n_143),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_351),
.B(n_354),
.Y(n_401)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_295),
.Y(n_352)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_352),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_285),
.B(n_318),
.C(n_299),
.Y(n_353)
);

AND2x6_ASAP7_75t_L g355 ( 
.A(n_285),
.B(n_157),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_355),
.B(n_361),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_L g372 ( 
.A1(n_356),
.A2(n_317),
.B1(n_284),
.B2(n_294),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_319),
.B(n_255),
.Y(n_357)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_288),
.Y(n_360)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_360),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_316),
.Y(n_361)
);

INVx13_ASAP7_75t_L g362 ( 
.A(n_307),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_362),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_290),
.B(n_242),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_327),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_364),
.B(n_366),
.Y(n_393)
);

OAI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_281),
.A2(n_270),
.B1(n_217),
.B2(n_203),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_306),
.B(n_202),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_288),
.Y(n_367)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_367),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_291),
.B(n_202),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_368),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_326),
.B(n_217),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_369),
.A2(n_371),
.B(n_302),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_326),
.B(n_203),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_372),
.A2(n_399),
.B1(n_335),
.B2(n_303),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_373),
.B(n_375),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_350),
.B(n_313),
.Y(n_375)
);

XNOR2x1_ASAP7_75t_L g376 ( 
.A(n_348),
.B(n_282),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_376),
.B(n_280),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_378),
.B(n_352),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_353),
.A2(n_293),
.B1(n_302),
.B2(n_253),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_383),
.A2(n_386),
.B1(n_400),
.B2(n_402),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_337),
.A2(n_336),
.B1(n_333),
.B2(n_366),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_342),
.A2(n_328),
.B(n_327),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_388),
.A2(n_392),
.B(n_334),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_338),
.A2(n_356),
.B1(n_337),
.B2(n_355),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_389),
.A2(n_394),
.B1(n_359),
.B2(n_358),
.Y(n_418)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_370),
.Y(n_391)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_391),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_338),
.A2(n_286),
.B1(n_297),
.B2(n_273),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_345),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_397),
.B(n_406),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_354),
.B(n_327),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_398),
.B(n_340),
.C(n_359),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_L g399 ( 
.A1(n_338),
.A2(n_346),
.B1(n_364),
.B2(n_332),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_351),
.A2(n_297),
.B1(n_225),
.B2(n_215),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_361),
.A2(n_213),
.B1(n_201),
.B2(n_273),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_403),
.B(n_394),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_345),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_363),
.B(n_298),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_407),
.B(n_324),
.C(n_289),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_384),
.B(n_371),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_412),
.B(n_413),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_405),
.B(n_369),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_384),
.B(n_370),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_415),
.B(n_419),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_416),
.B(n_443),
.Y(n_468)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_417),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_418),
.A2(n_427),
.B1(n_433),
.B2(n_439),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_380),
.B(n_345),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_393),
.B(n_358),
.Y(n_420)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_420),
.Y(n_469)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_393),
.Y(n_421)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_421),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_380),
.B(n_343),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_422),
.B(n_423),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_405),
.B(n_343),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_391),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_424),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_377),
.A2(n_334),
.B(n_329),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_425),
.A2(n_436),
.B(n_392),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_397),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_426),
.B(n_428),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_389),
.A2(n_272),
.B1(n_292),
.B2(n_308),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_385),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_406),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_429),
.B(n_432),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_430),
.B(n_431),
.Y(n_467)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_385),
.Y(n_432)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_387),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_434),
.B(n_435),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_382),
.B(n_360),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_377),
.A2(n_401),
.B(n_396),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_408),
.B(n_367),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_437),
.B(n_440),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_438),
.B(n_376),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_373),
.A2(n_292),
.B1(n_321),
.B2(n_272),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_401),
.A2(n_277),
.B1(n_296),
.B2(n_265),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_387),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_441),
.B(n_442),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_396),
.A2(n_296),
.B1(n_254),
.B2(n_287),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_444),
.A2(n_460),
.B(n_461),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_410),
.A2(n_392),
.B1(n_390),
.B2(n_376),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_445),
.A2(n_464),
.B1(n_411),
.B2(n_418),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_422),
.B(n_386),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_451),
.B(n_413),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_409),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_452),
.B(n_454),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_409),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_431),
.B(n_375),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_455),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_420),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_458),
.B(n_379),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_459),
.B(n_465),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_411),
.A2(n_375),
.B(n_378),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_411),
.B(n_400),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_425),
.A2(n_402),
.B(n_388),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_462),
.A2(n_463),
.B(n_471),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_411),
.A2(n_383),
.B(n_382),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_410),
.A2(n_390),
.B1(n_407),
.B2(n_381),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_438),
.B(n_398),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_416),
.B(n_374),
.C(n_381),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_466),
.B(n_443),
.C(n_426),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_436),
.A2(n_395),
.B(n_374),
.Y(n_471)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_446),
.Y(n_475)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_475),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_476),
.B(n_485),
.C(n_487),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_479),
.B(n_480),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_468),
.B(n_435),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_446),
.Y(n_481)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_481),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_482),
.A2(n_483),
.B1(n_486),
.B2(n_447),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_461),
.A2(n_433),
.B1(n_440),
.B2(n_427),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_449),
.A2(n_421),
.B1(n_417),
.B2(n_430),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_484),
.A2(n_489),
.B1(n_494),
.B2(n_500),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_466),
.B(n_429),
.C(n_414),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_449),
.A2(n_439),
.B1(n_442),
.B2(n_415),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_468),
.B(n_414),
.C(n_424),
.Y(n_487)
);

INVx4_ASAP7_75t_L g488 ( 
.A(n_452),
.Y(n_488)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_488),
.Y(n_505)
);

AOI211xp5_ASAP7_75t_L g489 ( 
.A1(n_463),
.A2(n_412),
.B(n_419),
.C(n_423),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_453),
.Y(n_490)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_490),
.Y(n_510)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_453),
.Y(n_491)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_491),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_464),
.B(n_441),
.C(n_428),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_493),
.B(n_467),
.C(n_454),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_469),
.A2(n_434),
.B1(n_432),
.B2(n_437),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_456),
.A2(n_379),
.B1(n_395),
.B2(n_403),
.Y(n_495)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_495),
.Y(n_517)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_498),
.Y(n_523)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_450),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_499),
.B(n_502),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_469),
.A2(n_395),
.B1(n_305),
.B2(n_307),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_459),
.B(n_445),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_501),
.B(n_465),
.Y(n_503)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_470),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_503),
.B(n_511),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_487),
.B(n_444),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_512),
.B(n_516),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_485),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_513),
.B(n_479),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_480),
.B(n_471),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_478),
.B(n_460),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_518),
.B(n_478),
.C(n_501),
.Y(n_526)
);

OAI21xp33_ASAP7_75t_L g519 ( 
.A1(n_477),
.A2(n_467),
.B(n_455),
.Y(n_519)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_519),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_520),
.A2(n_472),
.B1(n_524),
.B2(n_508),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_492),
.B(n_404),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_521),
.B(n_448),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_476),
.B(n_455),
.C(n_473),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_522),
.B(n_524),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_493),
.B(n_473),
.C(n_462),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_488),
.B(n_456),
.Y(n_525)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_525),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_526),
.B(n_530),
.Y(n_547)
);

AO221x1_ASAP7_75t_L g527 ( 
.A1(n_513),
.A2(n_450),
.B1(n_491),
.B2(n_490),
.C(n_502),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_527),
.A2(n_542),
.B(n_541),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_523),
.A2(n_486),
.B1(n_447),
.B2(n_483),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_528),
.B(n_534),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_517),
.A2(n_489),
.B1(n_484),
.B2(n_461),
.Y(n_529)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_529),
.Y(n_551)
);

BUFx2_ASAP7_75t_L g532 ( 
.A(n_505),
.Y(n_532)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_532),
.Y(n_552)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_533),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_514),
.A2(n_458),
.B1(n_474),
.B2(n_472),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_514),
.A2(n_497),
.B1(n_496),
.B2(n_474),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_536),
.A2(n_509),
.B1(n_522),
.B2(n_500),
.Y(n_553)
);

A2O1A1Ixp33_ASAP7_75t_SL g538 ( 
.A1(n_519),
.A2(n_496),
.B(n_497),
.C(n_470),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_538),
.B(n_515),
.C(n_510),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_540),
.B(n_542),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_506),
.B(n_494),
.C(n_457),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_507),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_543),
.B(n_506),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_511),
.B(n_448),
.Y(n_544)
);

CKINVDCx16_ASAP7_75t_R g548 ( 
.A(n_544),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_545),
.B(n_550),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_526),
.B(n_518),
.Y(n_550)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_553),
.Y(n_564)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_555),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_539),
.B(n_537),
.Y(n_556)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_556),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_537),
.B(n_504),
.C(n_512),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_557),
.A2(n_305),
.B(n_322),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_536),
.A2(n_516),
.B1(n_504),
.B2(n_503),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g566 ( 
.A(n_558),
.B(n_559),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_SL g559 ( 
.A(n_531),
.B(n_457),
.Y(n_559)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_560),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_557),
.B(n_533),
.C(n_530),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_561),
.B(n_562),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_556),
.B(n_549),
.C(n_550),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_SL g563 ( 
.A1(n_551),
.A2(n_535),
.B(n_538),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_SL g577 ( 
.A1(n_563),
.A2(n_571),
.B(n_552),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_SL g567 ( 
.A(n_548),
.B(n_529),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_567),
.B(n_569),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_L g568 ( 
.A1(n_558),
.A2(n_538),
.B(n_532),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_568),
.A2(n_545),
.B(n_546),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_553),
.B(n_538),
.C(n_322),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g585 ( 
.A1(n_574),
.A2(n_575),
.B(n_581),
.Y(n_585)
);

NOR2x1_ASAP7_75t_L g575 ( 
.A(n_572),
.B(n_554),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_577),
.B(n_582),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_562),
.B(n_547),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_579),
.B(n_580),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_565),
.B(n_547),
.C(n_559),
.Y(n_580)
);

NOR2xp67_ASAP7_75t_L g581 ( 
.A(n_570),
.B(n_329),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_565),
.B(n_304),
.C(n_362),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_573),
.B(n_304),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_583),
.B(n_8),
.Y(n_589)
);

AOI322xp5_ASAP7_75t_L g586 ( 
.A1(n_576),
.A2(n_564),
.A3(n_563),
.B1(n_569),
.B2(n_561),
.C1(n_566),
.C2(n_362),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_586),
.A2(n_589),
.B1(n_582),
.B2(n_575),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_578),
.A2(n_329),
.B1(n_250),
.B2(n_60),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_587),
.B(n_588),
.C(n_11),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_580),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_591),
.B(n_592),
.Y(n_596)
);

OAI21xp5_ASAP7_75t_L g592 ( 
.A1(n_585),
.A2(n_11),
.B(n_12),
.Y(n_592)
);

AOI21xp5_ASAP7_75t_SL g593 ( 
.A1(n_584),
.A2(n_11),
.B(n_13),
.Y(n_593)
);

BUFx24_ASAP7_75t_SL g595 ( 
.A(n_593),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_596),
.B(n_590),
.C(n_595),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_597),
.B(n_594),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g599 ( 
.A1(n_598),
.A2(n_586),
.B1(n_14),
.B2(n_56),
.Y(n_599)
);

BUFx24_ASAP7_75t_SL g600 ( 
.A(n_599),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_600),
.B(n_14),
.Y(n_601)
);


endmodule