module fake_jpeg_1528_n_148 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_148);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx8_ASAP7_75t_SL g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_14),
.B(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_21),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_53),
.B(n_55),
.Y(n_59)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_42),
.B(n_1),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_36),
.Y(n_56)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_1),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_35),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_37),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_72),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_64),
.B(n_37),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_64),
.A2(n_50),
.B1(n_47),
.B2(n_48),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_73),
.A2(n_84),
.B1(n_2),
.B2(n_3),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_77),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_43),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_60),
.A2(n_50),
.B1(n_45),
.B2(n_39),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_82),
.B1(n_47),
.B2(n_68),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_64),
.B(n_44),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_81),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_50),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_62),
.A2(n_48),
.B(n_3),
.C(n_4),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_45),
.B1(n_39),
.B2(n_38),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_71),
.A2(n_63),
.B1(n_66),
.B2(n_69),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_20),
.Y(n_108)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_94),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_2),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_95),
.B(n_98),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_96),
.Y(n_105)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_5),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_19),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_88),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_109),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_93),
.A2(n_83),
.B(n_6),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_104),
.A2(n_112),
.B(n_10),
.Y(n_120)
);

XOR2x2_ASAP7_75t_SL g106 ( 
.A(n_97),
.B(n_5),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_12),
.C(n_13),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_108),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_34),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_92),
.B(n_6),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_114),
.Y(n_121)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_111),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_85),
.A2(n_7),
.B(n_8),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_7),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_115),
.B(n_116),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_8),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_119),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_9),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_120),
.A2(n_122),
.B1(n_126),
.B2(n_129),
.Y(n_133)
);

OAI22x1_ASAP7_75t_L g122 ( 
.A1(n_113),
.A2(n_25),
.B1(n_30),
.B2(n_16),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_106),
.C(n_105),
.Y(n_135)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_125),
.Y(n_131)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_104),
.A2(n_18),
.B(n_22),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_112),
.B(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_31),
.Y(n_129)
);

BUFx24_ASAP7_75t_SL g132 ( 
.A(n_121),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_134),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_123),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_131),
.A2(n_122),
.B(n_118),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_138),
.Y(n_140)
);

NOR2xp67_ASAP7_75t_SL g139 ( 
.A(n_130),
.B(n_120),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_139),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_140),
.B(n_136),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_141),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_143),
.A2(n_127),
.B(n_133),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_124),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_145),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_108),
.C(n_26),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_24),
.Y(n_148)
);


endmodule