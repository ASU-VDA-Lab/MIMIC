module real_jpeg_7351_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_38;
wire n_33;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_44;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_40;
wire n_36;
wire n_39;
wire n_41;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_26;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

BUFx10_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

AND2x2_ASAP7_75t_SL g29 ( 
.A(n_1),
.B(n_5),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_1),
.B(n_19),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_3),
.B(n_12),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_4),
.B(n_11),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_4),
.B(n_11),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_4),
.B(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

AOI221xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_16),
.B1(n_23),
.B2(n_29),
.C(n_30),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_8),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_SL g8 ( 
.A(n_9),
.B(n_15),
.Y(n_8)
);

AND2x2_ASAP7_75t_SL g28 ( 
.A(n_9),
.B(n_15),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g9 ( 
.A1(n_10),
.A2(n_13),
.B(n_14),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_11),
.B(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_12),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_27),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_15),
.B(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_15),
.B(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_21),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_20),
.Y(n_18)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

OR2x4_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_27),
.A2(n_38),
.B(n_40),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_33),
.B1(n_41),
.B2(n_42),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);


endmodule