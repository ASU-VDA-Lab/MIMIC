module fake_netlist_1_5705_n_514 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_514);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_514;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_141;
wire n_119;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_493;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_SL g77 ( .A(n_44), .Y(n_77) );
CKINVDCx5p33_ASAP7_75t_R g78 ( .A(n_52), .Y(n_78) );
CKINVDCx16_ASAP7_75t_R g79 ( .A(n_51), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_58), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_30), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_20), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_35), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_17), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_48), .Y(n_85) );
INVxp33_ASAP7_75t_L g86 ( .A(n_69), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_76), .Y(n_87) );
BUFx5_ASAP7_75t_L g88 ( .A(n_65), .Y(n_88) );
CKINVDCx20_ASAP7_75t_R g89 ( .A(n_39), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_71), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_19), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_42), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_68), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_14), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_49), .Y(n_95) );
INVx2_ASAP7_75t_SL g96 ( .A(n_36), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_28), .Y(n_97) );
INVxp67_ASAP7_75t_SL g98 ( .A(n_9), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_59), .Y(n_99) );
INVxp33_ASAP7_75t_L g100 ( .A(n_41), .Y(n_100) );
NOR2xp33_ASAP7_75t_L g101 ( .A(n_37), .B(n_21), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_72), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_43), .Y(n_103) );
CKINVDCx16_ASAP7_75t_R g104 ( .A(n_54), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_40), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_57), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_26), .Y(n_107) );
INVxp67_ASAP7_75t_L g108 ( .A(n_55), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_50), .Y(n_109) );
INVxp33_ASAP7_75t_SL g110 ( .A(n_45), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g111 ( .A(n_73), .B(n_18), .Y(n_111) );
BUFx10_ASAP7_75t_L g112 ( .A(n_70), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_80), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_81), .Y(n_114) );
INVx3_ASAP7_75t_L g115 ( .A(n_112), .Y(n_115) );
BUFx2_ASAP7_75t_L g116 ( .A(n_79), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_82), .Y(n_117) );
OR2x6_ASAP7_75t_L g118 ( .A(n_84), .B(n_0), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_96), .B(n_0), .Y(n_119) );
AND2x2_ASAP7_75t_L g120 ( .A(n_86), .B(n_1), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_96), .B(n_1), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_86), .B(n_2), .Y(n_122) );
INVx3_ASAP7_75t_L g123 ( .A(n_112), .Y(n_123) );
AND2x2_ASAP7_75t_L g124 ( .A(n_100), .B(n_2), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_93), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_100), .B(n_3), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_94), .B(n_3), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_104), .B(n_4), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_83), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_85), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_90), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_91), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_92), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_88), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_93), .B(n_4), .Y(n_135) );
AO21x2_ASAP7_75t_L g136 ( .A1(n_135), .A2(n_102), .B(n_97), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_134), .Y(n_137) );
BUFx2_ASAP7_75t_L g138 ( .A(n_116), .Y(n_138) );
AND2x6_ASAP7_75t_L g139 ( .A(n_120), .B(n_107), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_134), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_113), .B(n_105), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_113), .B(n_106), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_114), .B(n_95), .Y(n_143) );
OAI22xp33_ASAP7_75t_L g144 ( .A1(n_118), .A2(n_98), .B1(n_89), .B2(n_110), .Y(n_144) );
INVx1_ASAP7_75t_SL g145 ( .A(n_116), .Y(n_145) );
INVxp33_ASAP7_75t_L g146 ( .A(n_128), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_125), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_114), .B(n_103), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_125), .Y(n_149) );
AND2x2_ASAP7_75t_L g150 ( .A(n_115), .B(n_112), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_134), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_117), .B(n_109), .Y(n_152) );
INVx4_ASAP7_75t_L g153 ( .A(n_118), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_125), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_115), .B(n_123), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_125), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_115), .B(n_99), .Y(n_157) );
NAND2x1p5_ASAP7_75t_L g158 ( .A(n_120), .B(n_111), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_115), .B(n_108), .Y(n_159) );
AND2x6_ASAP7_75t_L g160 ( .A(n_124), .B(n_101), .Y(n_160) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_145), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_137), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_151), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_151), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_145), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_137), .Y(n_166) );
INVx2_ASAP7_75t_SL g167 ( .A(n_153), .Y(n_167) );
INVx5_ASAP7_75t_L g168 ( .A(n_153), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_140), .Y(n_169) );
AND2x2_ASAP7_75t_L g170 ( .A(n_153), .B(n_124), .Y(n_170) );
BUFx4f_ASAP7_75t_L g171 ( .A(n_139), .Y(n_171) );
HB1xp67_ASAP7_75t_L g172 ( .A(n_138), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_151), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_139), .A2(n_118), .B1(n_128), .B2(n_131), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_151), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_153), .B(n_118), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_150), .B(n_123), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_150), .B(n_123), .Y(n_178) );
BUFx4f_ASAP7_75t_L g179 ( .A(n_139), .Y(n_179) );
BUFx3_ASAP7_75t_L g180 ( .A(n_139), .Y(n_180) );
INVx2_ASAP7_75t_SL g181 ( .A(n_159), .Y(n_181) );
NAND2xp33_ASAP7_75t_L g182 ( .A(n_139), .B(n_88), .Y(n_182) );
BUFx4f_ASAP7_75t_L g183 ( .A(n_139), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_140), .Y(n_184) );
AND2x6_ASAP7_75t_L g185 ( .A(n_157), .B(n_123), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_136), .Y(n_186) );
BUFx2_ASAP7_75t_L g187 ( .A(n_138), .Y(n_187) );
INVx5_ASAP7_75t_L g188 ( .A(n_139), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_147), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_147), .Y(n_190) );
INVx1_ASAP7_75t_SL g191 ( .A(n_159), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_184), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_188), .B(n_180), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_184), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_186), .A2(n_155), .B(n_157), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_170), .B(n_139), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_168), .B(n_174), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_174), .A2(n_146), .B1(n_144), .B2(n_118), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_170), .B(n_159), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_185), .B(n_159), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_185), .B(n_157), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_185), .B(n_157), .Y(n_202) );
INVx3_ASAP7_75t_L g203 ( .A(n_184), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_188), .B(n_136), .Y(n_204) );
INVx3_ASAP7_75t_L g205 ( .A(n_168), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_168), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_162), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_162), .Y(n_208) );
INVxp67_ASAP7_75t_L g209 ( .A(n_161), .Y(n_209) );
A2O1A1Ixp33_ASAP7_75t_L g210 ( .A1(n_186), .A2(n_141), .B(n_142), .C(n_143), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_168), .Y(n_211) );
OAI22xp33_ASAP7_75t_L g212 ( .A1(n_165), .A2(n_89), .B1(n_126), .B2(n_122), .Y(n_212) );
AND2x4_ASAP7_75t_L g213 ( .A(n_188), .B(n_136), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_187), .B(n_152), .Y(n_214) );
HB1xp67_ASAP7_75t_L g215 ( .A(n_187), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_172), .B(n_152), .Y(n_216) );
INVx4_ASAP7_75t_L g217 ( .A(n_171), .Y(n_217) );
OR2x6_ASAP7_75t_L g218 ( .A(n_180), .B(n_158), .Y(n_218) );
INVx4_ASAP7_75t_L g219 ( .A(n_171), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_166), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_168), .Y(n_221) );
NAND2x1p5_ASAP7_75t_L g222 ( .A(n_188), .B(n_131), .Y(n_222) );
INVx4_ASAP7_75t_SL g223 ( .A(n_185), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_209), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_192), .Y(n_225) );
BUFx10_ASAP7_75t_L g226 ( .A(n_193), .Y(n_226) );
INVx3_ASAP7_75t_L g227 ( .A(n_211), .Y(n_227) );
INVx3_ASAP7_75t_L g228 ( .A(n_211), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_214), .B(n_166), .Y(n_229) );
OAI221xp5_ASAP7_75t_L g230 ( .A1(n_198), .A2(n_178), .B1(n_177), .B2(n_191), .C(n_148), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_207), .B(n_181), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_215), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_192), .Y(n_233) );
NAND2xp33_ASAP7_75t_L g234 ( .A(n_211), .B(n_168), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_214), .A2(n_185), .B1(n_181), .B2(n_136), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_216), .B(n_169), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_207), .B(n_169), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_216), .B(n_141), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g239 ( .A1(n_210), .A2(n_179), .B1(n_171), .B2(n_183), .Y(n_239) );
INVxp67_ASAP7_75t_SL g240 ( .A(n_192), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_207), .B(n_185), .Y(n_241) );
INVx2_ASAP7_75t_SL g242 ( .A(n_211), .Y(n_242) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_208), .A2(n_179), .B1(n_183), .B2(n_180), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_208), .B(n_176), .Y(n_244) );
CKINVDCx20_ASAP7_75t_R g245 ( .A(n_223), .Y(n_245) );
OAI221xp5_ASAP7_75t_L g246 ( .A1(n_199), .A2(n_142), .B1(n_143), .B2(n_148), .C(n_127), .Y(n_246) );
AOI21x1_ASAP7_75t_L g247 ( .A1(n_195), .A2(n_156), .B(n_154), .Y(n_247) );
OR2x2_ASAP7_75t_L g248 ( .A(n_212), .B(n_158), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_194), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g250 ( .A1(n_248), .A2(n_185), .B1(n_218), .B2(n_160), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_236), .B(n_194), .Y(n_251) );
AO31x2_ASAP7_75t_L g252 ( .A1(n_239), .A2(n_208), .A3(n_220), .B(n_194), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_233), .Y(n_253) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_226), .Y(n_254) );
AND4x1_ASAP7_75t_L g255 ( .A(n_235), .B(n_176), .C(n_119), .D(n_121), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_233), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_236), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_230), .A2(n_218), .B1(n_220), .B2(n_179), .Y(n_258) );
AOI21xp33_ASAP7_75t_SL g259 ( .A1(n_224), .A2(n_110), .B(n_77), .Y(n_259) );
NAND2x1p5_ASAP7_75t_L g260 ( .A(n_227), .B(n_203), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_236), .B(n_203), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_237), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g263 ( .A1(n_248), .A2(n_218), .B1(n_160), .B2(n_197), .Y(n_263) );
BUFx2_ASAP7_75t_L g264 ( .A(n_240), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_230), .A2(n_218), .B1(n_160), .B2(n_182), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_229), .Y(n_266) );
AOI221x1_ASAP7_75t_L g267 ( .A1(n_239), .A2(n_204), .B1(n_213), .B2(n_125), .C(n_196), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_229), .B(n_203), .Y(n_268) );
OR2x6_ASAP7_75t_L g269 ( .A(n_229), .B(n_218), .Y(n_269) );
AOI221xp5_ASAP7_75t_L g270 ( .A1(n_246), .A2(n_132), .B1(n_117), .B2(n_133), .C(n_129), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_246), .A2(n_183), .B1(n_203), .B2(n_200), .Y(n_271) );
BUFx2_ASAP7_75t_L g272 ( .A(n_264), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_264), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_253), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_253), .Y(n_275) );
OAI33xp33_ASAP7_75t_L g276 ( .A1(n_257), .A2(n_133), .A3(n_129), .B1(n_130), .B2(n_132), .B3(n_232), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_251), .B(n_240), .Y(n_277) );
AOI33xp33_ASAP7_75t_L g278 ( .A1(n_266), .A2(n_130), .A3(n_235), .B1(n_244), .B2(n_156), .B3(n_154), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_251), .B(n_249), .Y(n_279) );
OAI221xp5_ASAP7_75t_L g280 ( .A1(n_255), .A2(n_238), .B1(n_158), .B2(n_202), .C(n_201), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_256), .Y(n_281) );
OR2x2_ASAP7_75t_L g282 ( .A(n_256), .B(n_238), .Y(n_282) );
AOI221xp5_ASAP7_75t_L g283 ( .A1(n_259), .A2(n_270), .B1(n_262), .B2(n_271), .C(n_258), .Y(n_283) );
OAI21xp33_ASAP7_75t_L g284 ( .A1(n_265), .A2(n_237), .B(n_225), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_262), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_261), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g287 ( .A1(n_269), .A2(n_244), .B1(n_231), .B2(n_249), .Y(n_287) );
AOI221xp5_ASAP7_75t_L g288 ( .A1(n_261), .A2(n_244), .B1(n_77), .B2(n_231), .C(n_241), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_268), .B(n_249), .Y(n_289) );
NAND3xp33_ASAP7_75t_L g290 ( .A(n_267), .B(n_225), .C(n_125), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_268), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_252), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_269), .A2(n_160), .B1(n_243), .B2(n_241), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_272), .B(n_269), .Y(n_294) );
AOI211xp5_ASAP7_75t_L g295 ( .A1(n_280), .A2(n_254), .B(n_78), .C(n_87), .Y(n_295) );
NAND3xp33_ASAP7_75t_L g296 ( .A(n_283), .B(n_267), .C(n_78), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_277), .B(n_252), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_274), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_272), .B(n_269), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_282), .B(n_254), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_277), .B(n_252), .Y(n_301) );
AOI22xp5_ASAP7_75t_L g302 ( .A1(n_288), .A2(n_250), .B1(n_263), .B2(n_254), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_274), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_282), .B(n_225), .Y(n_304) );
INVx2_ASAP7_75t_SL g305 ( .A(n_273), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_273), .B(n_252), .Y(n_306) );
A2O1A1Ixp33_ASAP7_75t_L g307 ( .A1(n_278), .A2(n_254), .B(n_213), .C(n_204), .Y(n_307) );
AOI33xp33_ASAP7_75t_L g308 ( .A1(n_286), .A2(n_154), .A3(n_149), .B1(n_7), .B2(n_8), .B3(n_9), .Y(n_308) );
OAI211xp5_ASAP7_75t_SL g309 ( .A1(n_287), .A2(n_281), .B(n_286), .C(n_293), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_281), .Y(n_310) );
INVx2_ASAP7_75t_SL g311 ( .A(n_273), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_275), .Y(n_312) );
INVx2_ASAP7_75t_SL g313 ( .A(n_285), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_275), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_279), .B(n_252), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_285), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_292), .Y(n_317) );
AOI211xp5_ASAP7_75t_L g318 ( .A1(n_276), .A2(n_87), .B(n_254), .C(n_243), .Y(n_318) );
NAND4xp25_ASAP7_75t_L g319 ( .A(n_287), .B(n_149), .C(n_213), .D(n_204), .Y(n_319) );
BUFx2_ASAP7_75t_L g320 ( .A(n_292), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_279), .B(n_260), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_291), .Y(n_322) );
OAI221xp5_ASAP7_75t_SL g323 ( .A1(n_291), .A2(n_205), .B1(n_206), .B2(n_242), .C(n_227), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_309), .B(n_284), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_310), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_317), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_310), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_322), .B(n_289), .Y(n_328) );
NAND4xp25_ASAP7_75t_L g329 ( .A(n_295), .B(n_290), .C(n_289), .D(n_284), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_312), .Y(n_330) );
OAI22xp33_ASAP7_75t_L g331 ( .A1(n_319), .A2(n_290), .B1(n_245), .B2(n_260), .Y(n_331) );
INVx1_ASAP7_75t_SL g332 ( .A(n_305), .Y(n_332) );
NAND2x1_ASAP7_75t_L g333 ( .A(n_313), .B(n_227), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_322), .B(n_5), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_300), .B(n_5), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_317), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_315), .B(n_88), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_315), .B(n_88), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_297), .B(n_88), .Y(n_339) );
INVx1_ASAP7_75t_SL g340 ( .A(n_305), .Y(n_340) );
AND2x4_ASAP7_75t_L g341 ( .A(n_306), .B(n_242), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_298), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_297), .B(n_88), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_301), .B(n_88), .Y(n_344) );
INVxp67_ASAP7_75t_SL g345 ( .A(n_313), .Y(n_345) );
INVx4_ASAP7_75t_L g346 ( .A(n_311), .Y(n_346) );
NOR3xp33_ASAP7_75t_L g347 ( .A(n_308), .B(n_149), .C(n_227), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_298), .Y(n_348) );
AOI22xp5_ASAP7_75t_L g349 ( .A1(n_295), .A2(n_160), .B1(n_213), .B2(n_204), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_301), .B(n_247), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_304), .B(n_6), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_316), .B(n_6), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_303), .B(n_247), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_303), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_311), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_314), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_320), .B(n_260), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_294), .B(n_7), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_314), .Y(n_359) );
NOR2xp67_ASAP7_75t_SL g360 ( .A(n_296), .B(n_188), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_306), .B(n_8), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_316), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_306), .B(n_242), .Y(n_363) );
AOI32xp33_ASAP7_75t_L g364 ( .A1(n_318), .A2(n_10), .A3(n_11), .B1(n_12), .B2(n_13), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_306), .B(n_10), .Y(n_365) );
NOR3xp33_ASAP7_75t_SL g366 ( .A(n_307), .B(n_11), .C(n_12), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_337), .B(n_320), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_337), .B(n_294), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_338), .B(n_299), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_325), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_338), .B(n_299), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_339), .B(n_343), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_335), .B(n_323), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_326), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_339), .B(n_321), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_343), .B(n_302), .Y(n_376) );
OAI211xp5_ASAP7_75t_L g377 ( .A1(n_364), .A2(n_302), .B(n_228), .C(n_205), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_336), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_344), .B(n_13), .Y(n_379) );
NOR3xp33_ASAP7_75t_L g380 ( .A(n_344), .B(n_228), .C(n_205), .Y(n_380) );
NAND3xp33_ASAP7_75t_L g381 ( .A(n_324), .B(n_234), .C(n_228), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_361), .B(n_14), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_345), .B(n_328), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_350), .B(n_15), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_361), .B(n_15), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_358), .B(n_16), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_354), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_350), .B(n_16), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_327), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_332), .B(n_17), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_330), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_365), .B(n_160), .Y(n_392) );
INVx2_ASAP7_75t_SL g393 ( .A(n_346), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_342), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_340), .B(n_22), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_324), .A2(n_351), .B1(n_334), .B2(n_355), .C(n_352), .Y(n_396) );
OAI21xp5_ASAP7_75t_L g397 ( .A1(n_366), .A2(n_222), .B(n_205), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_346), .B(n_362), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_348), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_356), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_341), .B(n_23), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_346), .B(n_226), .Y(n_402) );
NAND4xp25_ASAP7_75t_L g403 ( .A(n_349), .B(n_206), .C(n_219), .D(n_217), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_329), .B(n_24), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_359), .Y(n_405) );
OA21x2_ASAP7_75t_L g406 ( .A1(n_353), .A2(n_173), .B(n_164), .Y(n_406) );
INVx1_ASAP7_75t_SL g407 ( .A(n_357), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_354), .Y(n_408) );
CKINVDCx6p67_ASAP7_75t_R g409 ( .A(n_357), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_353), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_341), .B(n_25), .Y(n_411) );
INVxp67_ASAP7_75t_L g412 ( .A(n_333), .Y(n_412) );
AO22x1_ASAP7_75t_L g413 ( .A1(n_393), .A2(n_363), .B1(n_341), .B2(n_347), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_370), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_383), .B(n_363), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_389), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_384), .B(n_360), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_410), .B(n_27), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_384), .B(n_29), .Y(n_419) );
XOR2x2_ASAP7_75t_L g420 ( .A(n_386), .B(n_31), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_388), .B(n_32), .Y(n_421) );
INVx2_ASAP7_75t_SL g422 ( .A(n_393), .Y(n_422) );
OAI221xp5_ASAP7_75t_L g423 ( .A1(n_396), .A2(n_206), .B1(n_222), .B2(n_221), .C(n_211), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_391), .Y(n_424) );
INVx1_ASAP7_75t_SL g425 ( .A(n_409), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_409), .B(n_33), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_407), .B(n_34), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_394), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g429 ( .A(n_412), .B(n_223), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_368), .B(n_38), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_399), .Y(n_431) );
XNOR2x1_ASAP7_75t_L g432 ( .A(n_390), .B(n_46), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_388), .B(n_47), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_368), .B(n_53), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_400), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_374), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_371), .B(n_56), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_373), .B(n_60), .Y(n_438) );
NAND3xp33_ASAP7_75t_SL g439 ( .A(n_377), .B(n_222), .C(n_219), .Y(n_439) );
OA211x2_ASAP7_75t_L g440 ( .A1(n_386), .A2(n_61), .B(n_62), .C(n_63), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_405), .Y(n_441) );
OAI221xp5_ASAP7_75t_SL g442 ( .A1(n_373), .A2(n_206), .B1(n_226), .B2(n_223), .C(n_167), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_398), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_406), .Y(n_444) );
NOR2xp33_ASAP7_75t_SL g445 ( .A(n_379), .B(n_221), .Y(n_445) );
NAND2xp33_ASAP7_75t_SL g446 ( .A(n_401), .B(n_221), .Y(n_446) );
XNOR2x2_ASAP7_75t_L g447 ( .A(n_379), .B(n_223), .Y(n_447) );
NAND2x1_ASAP7_75t_L g448 ( .A(n_406), .B(n_221), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_371), .B(n_64), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_408), .Y(n_450) );
AOI221x1_ASAP7_75t_SL g451 ( .A1(n_382), .A2(n_66), .B1(n_67), .B2(n_74), .C(n_75), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_376), .B(n_164), .Y(n_452) );
OAI21xp5_ASAP7_75t_SL g453 ( .A1(n_404), .A2(n_193), .B(n_223), .Y(n_453) );
AOI211xp5_ASAP7_75t_L g454 ( .A1(n_404), .A2(n_193), .B(n_173), .C(n_175), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_367), .B(n_173), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_380), .A2(n_188), .B1(n_219), .B2(n_217), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_385), .B(n_219), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_378), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_372), .B(n_163), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_406), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g461 ( .A1(n_402), .A2(n_217), .B1(n_193), .B2(n_167), .Y(n_461) );
XNOR2xp5_ASAP7_75t_L g462 ( .A(n_375), .B(n_163), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_369), .B(n_175), .Y(n_463) );
INVxp67_ASAP7_75t_L g464 ( .A(n_387), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_395), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_401), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_411), .A2(n_217), .B1(n_189), .B2(n_190), .Y(n_467) );
INVx1_ASAP7_75t_SL g468 ( .A(n_411), .Y(n_468) );
AOI222xp33_ASAP7_75t_L g469 ( .A1(n_392), .A2(n_189), .B1(n_190), .B2(n_381), .C1(n_397), .C2(n_403), .Y(n_469) );
INVxp67_ASAP7_75t_L g470 ( .A(n_398), .Y(n_470) );
AOI211xp5_ASAP7_75t_L g471 ( .A1(n_377), .A2(n_190), .B(n_331), .C(n_373), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_370), .Y(n_472) );
NOR2x1_ASAP7_75t_L g473 ( .A(n_390), .B(n_190), .Y(n_473) );
AOI222xp33_ASAP7_75t_L g474 ( .A1(n_386), .A2(n_190), .B1(n_396), .B2(n_344), .C1(n_343), .C2(n_339), .Y(n_474) );
AOI221xp5_ASAP7_75t_L g475 ( .A1(n_396), .A2(n_386), .B1(n_373), .B2(n_385), .C(n_382), .Y(n_475) );
INVxp67_ASAP7_75t_L g476 ( .A(n_425), .Y(n_476) );
AOI221xp5_ASAP7_75t_L g477 ( .A1(n_475), .A2(n_470), .B1(n_443), .B2(n_416), .C(n_414), .Y(n_477) );
CKINVDCx16_ASAP7_75t_R g478 ( .A(n_445), .Y(n_478) );
OAI221xp5_ASAP7_75t_L g479 ( .A1(n_471), .A2(n_451), .B1(n_470), .B2(n_423), .C(n_453), .Y(n_479) );
OAI21xp5_ASAP7_75t_SL g480 ( .A1(n_432), .A2(n_439), .B(n_474), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_436), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_424), .Y(n_482) );
AOI221xp5_ASAP7_75t_L g483 ( .A1(n_472), .A2(n_441), .B1(n_431), .B2(n_435), .C(n_428), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_468), .A2(n_438), .B1(n_432), .B2(n_420), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_422), .A2(n_415), .B1(n_462), .B2(n_417), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_450), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_464), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_438), .A2(n_420), .B1(n_466), .B2(n_469), .Y(n_488) );
OAI211xp5_ASAP7_75t_SL g489 ( .A1(n_454), .A2(n_473), .B(n_419), .C(n_421), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_413), .A2(n_446), .B(n_422), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_464), .Y(n_491) );
AOI31xp33_ASAP7_75t_L g492 ( .A1(n_484), .A2(n_426), .A3(n_446), .B(n_429), .Y(n_492) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_487), .Y(n_493) );
OAI211xp5_ASAP7_75t_L g494 ( .A1(n_480), .A2(n_433), .B(n_467), .C(n_457), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_490), .A2(n_429), .B1(n_460), .B2(n_444), .Y(n_495) );
OAI311xp33_ASAP7_75t_L g496 ( .A1(n_480), .A2(n_427), .A3(n_437), .B1(n_459), .C1(n_452), .Y(n_496) );
AOI211xp5_ASAP7_75t_SL g497 ( .A1(n_479), .A2(n_442), .B(n_437), .C(n_434), .Y(n_497) );
OA22x2_ASAP7_75t_L g498 ( .A1(n_476), .A2(n_447), .B1(n_465), .B2(n_430), .Y(n_498) );
AOI21xp33_ASAP7_75t_SL g499 ( .A1(n_478), .A2(n_460), .B(n_444), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_477), .B(n_458), .Y(n_500) );
AOI221xp5_ASAP7_75t_L g501 ( .A1(n_499), .A2(n_485), .B1(n_483), .B2(n_482), .C(n_491), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_L g502 ( .A1(n_495), .A2(n_489), .B(n_486), .C(n_461), .Y(n_502) );
NAND4xp25_ASAP7_75t_L g503 ( .A(n_497), .B(n_488), .C(n_440), .D(n_449), .Y(n_503) );
NAND3xp33_ASAP7_75t_SL g504 ( .A(n_494), .B(n_456), .C(n_448), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_493), .B(n_481), .Y(n_505) );
OAI221xp5_ASAP7_75t_R g506 ( .A1(n_504), .A2(n_498), .B1(n_492), .B2(n_496), .C(n_500), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_505), .Y(n_507) );
AOI211xp5_ASAP7_75t_L g508 ( .A1(n_503), .A2(n_498), .B(n_418), .C(n_455), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_508), .B(n_501), .Y(n_509) );
OAI211xp5_ASAP7_75t_SL g510 ( .A1(n_507), .A2(n_506), .B(n_502), .C(n_456), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_510), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_511), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_512), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_513), .A2(n_509), .B(n_463), .Y(n_514) );
endmodule