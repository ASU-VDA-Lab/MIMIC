module real_aes_7534_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_733;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g441 ( .A(n_0), .Y(n_441) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_1), .A2(n_120), .B(n_124), .C(n_205), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_2), .A2(n_154), .B(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g510 ( .A(n_3), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_4), .B(n_221), .Y(n_240) );
AOI21xp33_ASAP7_75t_L g475 ( .A1(n_5), .A2(n_154), .B(n_476), .Y(n_475) );
AND2x6_ASAP7_75t_L g120 ( .A(n_6), .B(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g195 ( .A(n_7), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_8), .B(n_41), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_9), .A2(n_153), .B(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_10), .B(n_132), .Y(n_207) );
INVx1_ASAP7_75t_L g480 ( .A(n_11), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_12), .B(n_235), .Y(n_535) );
INVx1_ASAP7_75t_L g140 ( .A(n_13), .Y(n_140) );
INVx1_ASAP7_75t_L g547 ( .A(n_14), .Y(n_547) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_15), .A2(n_130), .B(n_217), .C(n_219), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_16), .B(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_17), .B(n_498), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_18), .B(n_154), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_19), .B(n_166), .Y(n_165) );
A2O1A1Ixp33_ASAP7_75t_L g249 ( .A1(n_20), .A2(n_235), .B(n_250), .C(n_252), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_21), .B(n_221), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_22), .B(n_132), .Y(n_177) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_23), .A2(n_162), .B(n_219), .C(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g131 ( .A(n_24), .B(n_132), .Y(n_131) );
CKINVDCx16_ASAP7_75t_R g171 ( .A(n_25), .Y(n_171) );
INVx1_ASAP7_75t_L g128 ( .A(n_26), .Y(n_128) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_27), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_28), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_29), .B(n_132), .Y(n_511) );
OAI22xp5_ASAP7_75t_SL g744 ( .A1(n_30), .A2(n_31), .B1(n_745), .B2(n_746), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_30), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_31), .Y(n_745) );
INVx1_ASAP7_75t_L g160 ( .A(n_32), .Y(n_160) );
INVx1_ASAP7_75t_L g489 ( .A(n_33), .Y(n_489) );
INVx2_ASAP7_75t_L g118 ( .A(n_34), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g209 ( .A(n_35), .Y(n_209) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_36), .A2(n_235), .B(n_236), .C(n_238), .Y(n_234) );
INVxp67_ASAP7_75t_L g161 ( .A(n_37), .Y(n_161) );
A2O1A1Ixp33_ASAP7_75t_L g123 ( .A1(n_38), .A2(n_124), .B(n_127), .C(n_135), .Y(n_123) );
CKINVDCx14_ASAP7_75t_R g233 ( .A(n_39), .Y(n_233) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_40), .A2(n_120), .B(n_124), .C(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g488 ( .A(n_42), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_43), .A2(n_179), .B(n_193), .C(n_194), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_44), .B(n_132), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g742 ( .A1(n_45), .A2(n_743), .B1(n_744), .B2(n_747), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_45), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g142 ( .A(n_46), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_47), .Y(n_156) );
INVx1_ASAP7_75t_L g248 ( .A(n_48), .Y(n_248) );
CKINVDCx16_ASAP7_75t_R g490 ( .A(n_49), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_50), .B(n_154), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_51), .B(n_444), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_52), .A2(n_124), .B1(n_252), .B2(n_487), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_53), .Y(n_526) );
CKINVDCx16_ASAP7_75t_R g507 ( .A(n_54), .Y(n_507) );
CKINVDCx14_ASAP7_75t_R g191 ( .A(n_55), .Y(n_191) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_56), .A2(n_193), .B(n_238), .C(n_479), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g563 ( .A(n_57), .Y(n_563) );
INVx1_ASAP7_75t_L g477 ( .A(n_58), .Y(n_477) );
AOI22xp5_ASAP7_75t_L g433 ( .A1(n_59), .A2(n_88), .B1(n_434), .B2(n_435), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_59), .Y(n_435) );
INVx1_ASAP7_75t_L g121 ( .A(n_60), .Y(n_121) );
INVx1_ASAP7_75t_L g139 ( .A(n_61), .Y(n_139) );
INVx1_ASAP7_75t_SL g237 ( .A(n_62), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_63), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_64), .B(n_221), .Y(n_254) );
INVx1_ASAP7_75t_L g174 ( .A(n_65), .Y(n_174) );
A2O1A1Ixp33_ASAP7_75t_SL g497 ( .A1(n_66), .A2(n_238), .B(n_498), .C(n_499), .Y(n_497) );
INVxp67_ASAP7_75t_L g500 ( .A(n_67), .Y(n_500) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_68), .A2(n_103), .B1(n_446), .B2(n_454), .C1(n_457), .C2(n_754), .Y(n_102) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_68), .A2(n_105), .B1(n_106), .B2(n_107), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_68), .Y(n_105) );
INVx1_ASAP7_75t_L g453 ( .A(n_69), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_70), .A2(n_154), .B(n_190), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_71), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_72), .A2(n_154), .B(n_214), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_73), .Y(n_492) );
INVx1_ASAP7_75t_L g557 ( .A(n_74), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_75), .A2(n_153), .B(n_155), .Y(n_152) );
CKINVDCx16_ASAP7_75t_R g122 ( .A(n_76), .Y(n_122) );
INVx1_ASAP7_75t_L g215 ( .A(n_77), .Y(n_215) );
A2O1A1Ixp33_ASAP7_75t_L g558 ( .A1(n_78), .A2(n_120), .B(n_124), .C(n_559), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_79), .A2(n_154), .B(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g218 ( .A(n_80), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_81), .B(n_129), .Y(n_523) );
INVx2_ASAP7_75t_L g137 ( .A(n_82), .Y(n_137) );
INVx1_ASAP7_75t_L g206 ( .A(n_83), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_84), .B(n_498), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_85), .A2(n_120), .B(n_124), .C(n_509), .Y(n_508) );
OR2x2_ASAP7_75t_L g438 ( .A(n_86), .B(n_439), .Y(n_438) );
OR2x2_ASAP7_75t_L g462 ( .A(n_86), .B(n_440), .Y(n_462) );
INVx2_ASAP7_75t_L g466 ( .A(n_86), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g172 ( .A1(n_87), .A2(n_124), .B(n_173), .C(n_181), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_88), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_89), .B(n_136), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_90), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_91), .A2(n_120), .B(n_124), .C(n_533), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_92), .Y(n_539) );
INVx1_ASAP7_75t_L g496 ( .A(n_93), .Y(n_496) );
CKINVDCx16_ASAP7_75t_R g544 ( .A(n_94), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_95), .B(n_129), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_96), .B(n_144), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_97), .B(n_144), .Y(n_548) );
INVx2_ASAP7_75t_L g251 ( .A(n_98), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_99), .B(n_453), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_100), .A2(n_154), .B(n_495), .Y(n_494) );
AOI222xp33_ASAP7_75t_L g458 ( .A1(n_101), .A2(n_459), .B1(n_741), .B2(n_742), .C1(n_748), .C2(n_751), .Y(n_458) );
OAI21xp5_ASAP7_75t_SL g103 ( .A1(n_104), .A2(n_436), .B(n_443), .Y(n_103) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
XOR2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_433), .Y(n_107) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_108), .A2(n_460), .B1(n_463), .B2(n_467), .Y(n_459) );
INVx1_ASAP7_75t_L g749 ( .A(n_108), .Y(n_749) );
OR4x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_323), .C(n_370), .D(n_410), .Y(n_108) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_110), .B(n_269), .C(n_298), .Y(n_109) );
AOI211xp5_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_184), .B(n_222), .C(n_262), .Y(n_110) );
O2A1O1Ixp33_ASAP7_75t_L g298 ( .A1(n_111), .A2(n_282), .B(n_299), .C(n_303), .Y(n_298) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_146), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_113), .B(n_261), .Y(n_260) );
INVx3_ASAP7_75t_SL g265 ( .A(n_113), .Y(n_265) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_113), .Y(n_277) );
AND2x4_ASAP7_75t_L g281 ( .A(n_113), .B(n_229), .Y(n_281) );
AND2x2_ASAP7_75t_L g292 ( .A(n_113), .B(n_169), .Y(n_292) );
OR2x2_ASAP7_75t_L g316 ( .A(n_113), .B(n_225), .Y(n_316) );
AND2x2_ASAP7_75t_L g329 ( .A(n_113), .B(n_230), .Y(n_329) );
AND2x2_ASAP7_75t_L g369 ( .A(n_113), .B(n_355), .Y(n_369) );
AND2x2_ASAP7_75t_L g376 ( .A(n_113), .B(n_339), .Y(n_376) );
AND2x2_ASAP7_75t_L g406 ( .A(n_113), .B(n_147), .Y(n_406) );
OR2x6_ASAP7_75t_L g113 ( .A(n_114), .B(n_141), .Y(n_113) );
O2A1O1Ixp33_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_122), .B(n_123), .C(n_136), .Y(n_114) );
OAI21xp5_ASAP7_75t_L g170 ( .A1(n_115), .A2(n_171), .B(n_172), .Y(n_170) );
OAI21xp5_ASAP7_75t_L g202 ( .A1(n_115), .A2(n_203), .B(n_204), .Y(n_202) );
OAI22xp33_ASAP7_75t_L g485 ( .A1(n_115), .A2(n_164), .B1(n_486), .B2(n_490), .Y(n_485) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_115), .A2(n_507), .B(n_508), .Y(n_506) );
OAI21xp5_ASAP7_75t_L g556 ( .A1(n_115), .A2(n_557), .B(n_558), .Y(n_556) );
NAND2x1p5_ASAP7_75t_L g115 ( .A(n_116), .B(n_120), .Y(n_115) );
AND2x4_ASAP7_75t_L g154 ( .A(n_116), .B(n_120), .Y(n_154) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_119), .Y(n_116) );
INVx1_ASAP7_75t_L g134 ( .A(n_117), .Y(n_134) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g125 ( .A(n_118), .Y(n_125) );
INVx1_ASAP7_75t_L g253 ( .A(n_118), .Y(n_253) );
INVx1_ASAP7_75t_L g126 ( .A(n_119), .Y(n_126) );
INVx3_ASAP7_75t_L g130 ( .A(n_119), .Y(n_130) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_119), .Y(n_132) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_119), .Y(n_163) );
INVx1_ASAP7_75t_L g498 ( .A(n_119), .Y(n_498) );
BUFx3_ASAP7_75t_L g135 ( .A(n_120), .Y(n_135) );
INVx4_ASAP7_75t_SL g164 ( .A(n_120), .Y(n_164) );
INVx5_ASAP7_75t_L g157 ( .A(n_124), .Y(n_157) );
AND2x6_ASAP7_75t_L g124 ( .A(n_125), .B(n_126), .Y(n_124) );
BUFx3_ASAP7_75t_L g180 ( .A(n_125), .Y(n_180) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_125), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_129), .B(n_131), .C(n_133), .Y(n_127) );
OAI22xp33_ASAP7_75t_L g159 ( .A1(n_129), .A2(n_160), .B1(n_161), .B2(n_162), .Y(n_159) );
O2A1O1Ixp33_ASAP7_75t_L g509 ( .A1(n_129), .A2(n_510), .B(n_511), .C(n_512), .Y(n_509) );
INVx5_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_130), .B(n_195), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_130), .B(n_480), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_130), .B(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g193 ( .A(n_132), .Y(n_193) );
INVx4_ASAP7_75t_L g235 ( .A(n_132), .Y(n_235) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_134), .B(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g167 ( .A(n_136), .Y(n_167) );
OA21x2_ASAP7_75t_L g188 ( .A1(n_136), .A2(n_189), .B(n_196), .Y(n_188) );
INVx1_ASAP7_75t_L g201 ( .A(n_136), .Y(n_201) );
OA21x2_ASAP7_75t_L g541 ( .A1(n_136), .A2(n_542), .B(n_548), .Y(n_541) );
AND2x2_ASAP7_75t_SL g136 ( .A(n_137), .B(n_138), .Y(n_136) );
AND2x2_ASAP7_75t_L g145 ( .A(n_137), .B(n_138), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
AO21x2_ASAP7_75t_L g169 ( .A1(n_143), .A2(n_170), .B(n_182), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_143), .B(n_209), .Y(n_208) );
INVx3_ASAP7_75t_L g221 ( .A(n_143), .Y(n_221) );
NOR2xp33_ASAP7_75t_SL g525 ( .A(n_143), .B(n_526), .Y(n_525) );
INVx4_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_144), .Y(n_212) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_144), .A2(n_494), .B(n_501), .Y(n_493) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g151 ( .A(n_145), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_146), .B(n_333), .Y(n_345) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_168), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_147), .B(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g283 ( .A(n_147), .B(n_168), .Y(n_283) );
BUFx3_ASAP7_75t_L g291 ( .A(n_147), .Y(n_291) );
OR2x2_ASAP7_75t_L g312 ( .A(n_147), .B(n_187), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_147), .B(n_333), .Y(n_423) );
OA21x2_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_152), .B(n_165), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_149), .A2(n_226), .B(n_227), .Y(n_225) );
AO21x2_ASAP7_75t_L g555 ( .A1(n_149), .A2(n_556), .B(n_562), .Y(n_555) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AOI21xp5_ASAP7_75t_SL g519 ( .A1(n_150), .A2(n_520), .B(n_521), .Y(n_519) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AO21x2_ASAP7_75t_L g484 ( .A1(n_151), .A2(n_485), .B(n_491), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_151), .B(n_492), .Y(n_491) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_151), .A2(n_506), .B(n_513), .Y(n_505) );
INVx1_ASAP7_75t_L g226 ( .A(n_152), .Y(n_226) );
BUFx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
O2A1O1Ixp33_ASAP7_75t_SL g155 ( .A1(n_156), .A2(n_157), .B(n_158), .C(n_164), .Y(n_155) );
O2A1O1Ixp33_ASAP7_75t_SL g190 ( .A1(n_157), .A2(n_164), .B(n_191), .C(n_192), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_SL g214 ( .A1(n_157), .A2(n_164), .B(n_215), .C(n_216), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_157), .A2(n_164), .B(n_233), .C(n_234), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_SL g247 ( .A1(n_157), .A2(n_164), .B(n_248), .C(n_249), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_157), .A2(n_164), .B(n_477), .C(n_478), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g495 ( .A1(n_157), .A2(n_164), .B(n_496), .C(n_497), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_L g543 ( .A1(n_157), .A2(n_164), .B(n_544), .C(n_545), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_162), .B(n_218), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_162), .B(n_251), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_162), .B(n_547), .Y(n_546) );
INVx4_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g176 ( .A(n_163), .Y(n_176) );
OAI22xp5_ASAP7_75t_SL g487 ( .A1(n_163), .A2(n_176), .B1(n_488), .B2(n_489), .Y(n_487) );
INVx1_ASAP7_75t_L g181 ( .A(n_164), .Y(n_181) );
INVx1_ASAP7_75t_L g227 ( .A(n_165), .Y(n_227) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_167), .B(n_183), .Y(n_182) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_167), .A2(n_531), .B(n_538), .Y(n_530) );
AND2x2_ASAP7_75t_L g228 ( .A(n_168), .B(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g276 ( .A(n_168), .Y(n_276) );
AND2x2_ASAP7_75t_L g339 ( .A(n_168), .B(n_230), .Y(n_339) );
AOI221xp5_ASAP7_75t_L g341 ( .A1(n_168), .A2(n_342), .B1(n_344), .B2(n_346), .C(n_347), .Y(n_341) );
AND2x2_ASAP7_75t_L g355 ( .A(n_168), .B(n_225), .Y(n_355) );
AND2x2_ASAP7_75t_L g381 ( .A(n_168), .B(n_265), .Y(n_381) );
INVx2_ASAP7_75t_SL g168 ( .A(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_L g261 ( .A(n_169), .B(n_230), .Y(n_261) );
BUFx2_ASAP7_75t_L g395 ( .A(n_169), .Y(n_395) );
O2A1O1Ixp33_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_177), .C(n_178), .Y(n_173) );
O2A1O1Ixp5_ASAP7_75t_L g205 ( .A1(n_175), .A2(n_178), .B(n_206), .C(n_207), .Y(n_205) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_178), .A2(n_523), .B(n_524), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_178), .A2(n_560), .B(n_561), .Y(n_559) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g219 ( .A(n_180), .Y(n_219) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
OAI32xp33_ASAP7_75t_L g361 ( .A1(n_185), .A2(n_322), .A3(n_336), .B1(n_362), .B2(n_363), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_186), .B(n_197), .Y(n_185) );
AND2x2_ASAP7_75t_L g302 ( .A(n_186), .B(n_244), .Y(n_302) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
OR2x2_ASAP7_75t_L g284 ( .A(n_187), .B(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_187), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g356 ( .A(n_187), .B(n_244), .Y(n_356) );
AND2x2_ASAP7_75t_L g367 ( .A(n_187), .B(n_259), .Y(n_367) );
BUFx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
OR2x2_ASAP7_75t_L g268 ( .A(n_188), .B(n_245), .Y(n_268) );
AND2x2_ASAP7_75t_L g272 ( .A(n_188), .B(n_245), .Y(n_272) );
AND2x2_ASAP7_75t_L g307 ( .A(n_188), .B(n_258), .Y(n_307) );
AND2x2_ASAP7_75t_L g314 ( .A(n_188), .B(n_210), .Y(n_314) );
OAI211xp5_ASAP7_75t_L g319 ( .A1(n_188), .A2(n_265), .B(n_276), .C(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g373 ( .A(n_188), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_188), .B(n_199), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_197), .B(n_256), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_197), .B(n_272), .Y(n_362) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
OR2x2_ASAP7_75t_L g267 ( .A(n_198), .B(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_199), .B(n_210), .Y(n_198) );
AND2x2_ASAP7_75t_L g259 ( .A(n_199), .B(n_211), .Y(n_259) );
OR2x2_ASAP7_75t_L g274 ( .A(n_199), .B(n_211), .Y(n_274) );
AND2x2_ASAP7_75t_L g297 ( .A(n_199), .B(n_258), .Y(n_297) );
INVx1_ASAP7_75t_L g301 ( .A(n_199), .Y(n_301) );
AND2x2_ASAP7_75t_L g320 ( .A(n_199), .B(n_257), .Y(n_320) );
OAI22xp33_ASAP7_75t_L g330 ( .A1(n_199), .A2(n_285), .B1(n_331), .B2(n_332), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_199), .B(n_373), .Y(n_397) );
AND2x2_ASAP7_75t_L g412 ( .A(n_199), .B(n_272), .Y(n_412) );
INVx4_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
BUFx3_ASAP7_75t_L g242 ( .A(n_200), .Y(n_242) );
AND2x2_ASAP7_75t_L g286 ( .A(n_200), .B(n_211), .Y(n_286) );
AND2x2_ASAP7_75t_L g288 ( .A(n_200), .B(n_244), .Y(n_288) );
AND3x2_ASAP7_75t_L g350 ( .A(n_200), .B(n_314), .C(n_351), .Y(n_350) );
AO21x2_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_202), .B(n_208), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_201), .B(n_514), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_201), .B(n_539), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_201), .B(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g385 ( .A(n_210), .B(n_257), .Y(n_385) );
INVx1_ASAP7_75t_SL g210 ( .A(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g244 ( .A(n_211), .B(n_245), .Y(n_244) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_211), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_211), .B(n_256), .Y(n_318) );
NAND3xp33_ASAP7_75t_L g425 ( .A(n_211), .B(n_297), .C(n_373), .Y(n_425) );
OA21x2_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_220), .Y(n_211) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_212), .A2(n_231), .B(n_240), .Y(n_230) );
OA21x2_ASAP7_75t_L g245 ( .A1(n_212), .A2(n_246), .B(n_254), .Y(n_245) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_221), .A2(n_475), .B(n_481), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_241), .B1(n_255), .B2(n_260), .Y(n_222) );
INVx1_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_228), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_225), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_SL g337 ( .A(n_225), .Y(n_337) );
OAI31xp33_ASAP7_75t_L g353 ( .A1(n_228), .A2(n_354), .A3(n_355), .B(n_356), .Y(n_353) );
AND2x2_ASAP7_75t_L g378 ( .A(n_228), .B(n_265), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_228), .B(n_291), .Y(n_424) );
AND2x2_ASAP7_75t_L g333 ( .A(n_229), .B(n_265), .Y(n_333) );
AND2x2_ASAP7_75t_L g394 ( .A(n_229), .B(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g264 ( .A(n_230), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g322 ( .A(n_230), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_235), .B(n_237), .Y(n_236) );
INVx3_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_239), .Y(n_536) );
OR2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
CKINVDCx16_ASAP7_75t_R g343 ( .A(n_242), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_243), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
AOI221x1_ASAP7_75t_SL g310 ( .A1(n_244), .A2(n_311), .B1(n_313), .B2(n_315), .C(n_317), .Y(n_310) );
INVx2_ASAP7_75t_L g258 ( .A(n_245), .Y(n_258) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_245), .Y(n_352) );
INVx2_ASAP7_75t_L g512 ( .A(n_252), .Y(n_512) );
INVx3_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g340 ( .A(n_255), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_259), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_256), .B(n_273), .Y(n_365) );
INVx1_ASAP7_75t_SL g428 ( .A(n_256), .Y(n_428) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g346 ( .A(n_259), .B(n_272), .Y(n_346) );
INVx1_ASAP7_75t_L g414 ( .A(n_260), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_260), .B(n_343), .Y(n_427) );
INVx2_ASAP7_75t_SL g266 ( .A(n_261), .Y(n_266) );
AND2x2_ASAP7_75t_L g309 ( .A(n_261), .B(n_265), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_261), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_261), .B(n_336), .Y(n_363) );
AOI21xp33_ASAP7_75t_SL g262 ( .A1(n_263), .A2(n_266), .B(n_267), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_264), .B(n_336), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_264), .B(n_291), .Y(n_432) );
OR2x2_ASAP7_75t_L g304 ( .A(n_265), .B(n_283), .Y(n_304) );
AND2x2_ASAP7_75t_L g403 ( .A(n_265), .B(n_394), .Y(n_403) );
OAI22xp5_ASAP7_75t_SL g278 ( .A1(n_266), .A2(n_279), .B1(n_284), .B2(n_287), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_266), .B(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g326 ( .A(n_268), .B(n_274), .Y(n_326) );
INVx1_ASAP7_75t_L g390 ( .A(n_268), .Y(n_390) );
AOI311xp33_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_275), .A3(n_277), .B(n_278), .C(n_289), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_273), .A2(n_405), .B1(n_417), .B2(n_420), .C(n_422), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_273), .B(n_428), .Y(n_430) );
INVx2_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g327 ( .A(n_275), .Y(n_327) );
AOI211xp5_ASAP7_75t_L g317 ( .A1(n_276), .A2(n_318), .B(n_319), .C(n_321), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
O2A1O1Ixp33_ASAP7_75t_SL g386 ( .A1(n_280), .A2(n_282), .B(n_387), .C(n_388), .Y(n_386) );
INVx3_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_281), .B(n_355), .Y(n_421) );
INVx1_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
OAI221xp5_ASAP7_75t_L g303 ( .A1(n_284), .A2(n_304), .B1(n_305), .B2(n_308), .C(n_310), .Y(n_303) );
INVx1_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g306 ( .A(n_286), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g389 ( .A(n_286), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_290), .B(n_293), .Y(n_289) );
A2O1A1Ixp33_ASAP7_75t_L g347 ( .A1(n_290), .A2(n_348), .B(n_349), .C(n_353), .Y(n_347) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_291), .B(n_292), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_291), .B(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_291), .B(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
INVxp67_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g313 ( .A(n_297), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_301), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g415 ( .A(n_304), .Y(n_415) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_307), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g342 ( .A(n_307), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_SL g419 ( .A(n_307), .Y(n_419) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g360 ( .A(n_309), .B(n_336), .Y(n_360) );
INVx1_ASAP7_75t_SL g354 ( .A(n_316), .Y(n_354) );
INVx1_ASAP7_75t_L g331 ( .A(n_322), .Y(n_331) );
NAND3xp33_ASAP7_75t_SL g323 ( .A(n_324), .B(n_341), .C(n_357), .Y(n_323) );
AOI322xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_327), .A3(n_328), .B1(n_330), .B2(n_334), .C1(n_338), .C2(n_340), .Y(n_324) );
AOI211xp5_ASAP7_75t_L g377 ( .A1(n_325), .A2(n_378), .B(n_379), .C(n_386), .Y(n_377) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_328), .A2(n_349), .B1(n_380), .B2(n_382), .Y(n_379) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g338 ( .A(n_336), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g375 ( .A(n_336), .B(n_376), .Y(n_375) );
AOI32xp33_ASAP7_75t_L g426 ( .A1(n_336), .A2(n_427), .A3(n_428), .B1(n_429), .B2(n_431), .Y(n_426) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g348 ( .A(n_339), .Y(n_348) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_339), .A2(n_392), .B1(n_396), .B2(n_398), .C(n_401), .Y(n_391) );
AND2x2_ASAP7_75t_L g405 ( .A(n_339), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g408 ( .A(n_343), .B(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g418 ( .A(n_343), .B(n_419), .Y(n_418) );
INVxp67_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
INVxp67_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g409 ( .A(n_352), .B(n_373), .Y(n_409) );
AOI211xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_360), .B(n_361), .C(n_364), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AOI21xp33_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_366), .B(n_368), .Y(n_364) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OAI211xp5_ASAP7_75t_SL g370 ( .A1(n_371), .A2(n_374), .B(n_377), .C(n_391), .Y(n_370) );
INVxp67_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_385), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g400 ( .A(n_397), .Y(n_400) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AOI21xp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_404), .B(n_407), .Y(n_401) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI211xp5_ASAP7_75t_SL g410 ( .A1(n_411), .A2(n_413), .B(n_416), .C(n_426), .Y(n_410) );
CKINVDCx20_ASAP7_75t_R g411 ( .A(n_412), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
INVx1_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AOI21xp33_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_424), .B(n_425), .Y(n_422) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_438), .Y(n_445) );
BUFx2_ASAP7_75t_L g456 ( .A(n_438), .Y(n_456) );
INVx1_ASAP7_75t_SL g758 ( .A(n_438), .Y(n_758) );
NOR2x2_ASAP7_75t_L g753 ( .A(n_439), .B(n_466), .Y(n_753) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OR2x2_ASAP7_75t_L g465 ( .A(n_440), .B(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_451), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OA21x2_ASAP7_75t_L g455 ( .A1(n_450), .A2(n_451), .B(n_456), .Y(n_455) );
NOR2xp33_ASAP7_75t_SL g756 ( .A(n_450), .B(n_452), .Y(n_756) );
INVx1_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
INVxp67_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OAI22x1_ASAP7_75t_L g748 ( .A1(n_460), .A2(n_463), .B1(n_749), .B2(n_750), .Y(n_748) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVxp67_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx2_ASAP7_75t_L g750 ( .A(n_468), .Y(n_750) );
BUFx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND3x1_ASAP7_75t_L g469 ( .A(n_470), .B(n_663), .C(n_708), .Y(n_469) );
NOR4xp25_ASAP7_75t_L g470 ( .A(n_471), .B(n_586), .C(n_627), .D(n_644), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_502), .B(n_516), .C(n_549), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_482), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_473), .B(n_503), .Y(n_502) );
NOR4xp25_ASAP7_75t_L g610 ( .A(n_473), .B(n_604), .C(n_611), .D(n_617), .Y(n_610) );
AND2x2_ASAP7_75t_L g683 ( .A(n_473), .B(n_572), .Y(n_683) );
AND2x2_ASAP7_75t_L g702 ( .A(n_473), .B(n_648), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_473), .B(n_697), .Y(n_711) );
AND2x2_ASAP7_75t_L g724 ( .A(n_473), .B(n_515), .Y(n_724) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_SL g569 ( .A(n_474), .Y(n_569) );
AND2x2_ASAP7_75t_L g576 ( .A(n_474), .B(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g626 ( .A(n_474), .B(n_483), .Y(n_626) );
AND2x2_ASAP7_75t_SL g637 ( .A(n_474), .B(n_572), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_474), .B(n_483), .Y(n_641) );
AND2x2_ASAP7_75t_L g650 ( .A(n_474), .B(n_575), .Y(n_650) );
BUFx2_ASAP7_75t_L g673 ( .A(n_474), .Y(n_673) );
AND2x2_ASAP7_75t_L g677 ( .A(n_474), .B(n_493), .Y(n_677) );
OR2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_493), .Y(n_482) );
AND2x2_ASAP7_75t_L g515 ( .A(n_483), .B(n_493), .Y(n_515) );
BUFx2_ASAP7_75t_L g579 ( .A(n_483), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_483), .A2(n_612), .B1(n_614), .B2(n_615), .Y(n_611) );
OR2x2_ASAP7_75t_L g633 ( .A(n_483), .B(n_505), .Y(n_633) );
AND2x2_ASAP7_75t_L g697 ( .A(n_483), .B(n_575), .Y(n_697) );
INVx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g565 ( .A(n_484), .B(n_505), .Y(n_565) );
AND2x2_ASAP7_75t_L g572 ( .A(n_484), .B(n_493), .Y(n_572) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_484), .Y(n_614) );
OR2x2_ASAP7_75t_L g649 ( .A(n_484), .B(n_504), .Y(n_649) );
INVx1_ASAP7_75t_L g568 ( .A(n_493), .Y(n_568) );
INVx3_ASAP7_75t_L g577 ( .A(n_493), .Y(n_577) );
BUFx2_ASAP7_75t_L g601 ( .A(n_493), .Y(n_601) );
AND2x2_ASAP7_75t_L g634 ( .A(n_493), .B(n_569), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_502), .A2(n_720), .B1(n_721), .B2(n_722), .Y(n_719) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_515), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_504), .B(n_577), .Y(n_581) );
INVx1_ASAP7_75t_L g609 ( .A(n_504), .Y(n_609) );
INVx3_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx3_ASAP7_75t_L g575 ( .A(n_505), .Y(n_575) );
INVx1_ASAP7_75t_L g587 ( .A(n_515), .Y(n_587) );
NAND2x1_ASAP7_75t_SL g516 ( .A(n_517), .B(n_527), .Y(n_516) );
AND2x2_ASAP7_75t_L g585 ( .A(n_517), .B(n_540), .Y(n_585) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_517), .Y(n_659) );
AND2x2_ASAP7_75t_L g686 ( .A(n_517), .B(n_606), .Y(n_686) );
AND2x2_ASAP7_75t_L g694 ( .A(n_517), .B(n_656), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_517), .B(n_552), .Y(n_721) );
INVx3_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g553 ( .A(n_518), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g570 ( .A(n_518), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g591 ( .A(n_518), .Y(n_591) );
INVx1_ASAP7_75t_L g597 ( .A(n_518), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_518), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g630 ( .A(n_518), .B(n_555), .Y(n_630) );
OR2x2_ASAP7_75t_L g668 ( .A(n_518), .B(n_623), .Y(n_668) );
AOI32xp33_ASAP7_75t_L g680 ( .A1(n_518), .A2(n_681), .A3(n_684), .B1(n_685), .B2(n_686), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_518), .B(n_656), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_518), .B(n_616), .Y(n_731) );
OR2x6_ASAP7_75t_L g518 ( .A(n_519), .B(n_525), .Y(n_518) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OR2x2_ASAP7_75t_L g642 ( .A(n_528), .B(n_643), .Y(n_642) );
OR2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_540), .Y(n_528) );
INVx1_ASAP7_75t_L g604 ( .A(n_529), .Y(n_604) );
AND2x2_ASAP7_75t_L g606 ( .A(n_529), .B(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_529), .B(n_554), .Y(n_623) );
AND2x2_ASAP7_75t_L g656 ( .A(n_529), .B(n_632), .Y(n_656) );
AND2x2_ASAP7_75t_L g693 ( .A(n_529), .B(n_555), .Y(n_693) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g552 ( .A(n_530), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_530), .B(n_554), .Y(n_583) );
AND2x2_ASAP7_75t_L g590 ( .A(n_530), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g631 ( .A(n_530), .B(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_537), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_535), .B(n_536), .Y(n_533) );
INVx2_ASAP7_75t_L g607 ( .A(n_540), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_540), .B(n_554), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_540), .B(n_598), .Y(n_679) );
INVx1_ASAP7_75t_L g701 ( .A(n_540), .Y(n_701) );
INVx1_ASAP7_75t_L g718 ( .A(n_540), .Y(n_718) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g571 ( .A(n_541), .B(n_554), .Y(n_571) );
AND2x2_ASAP7_75t_L g593 ( .A(n_541), .B(n_555), .Y(n_593) );
INVx1_ASAP7_75t_L g632 ( .A(n_541), .Y(n_632) );
AOI221x1_ASAP7_75t_SL g549 ( .A1(n_550), .A2(n_564), .B1(n_570), .B2(n_572), .C(n_573), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_550), .A2(n_637), .B1(n_704), .B2(n_705), .Y(n_703) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_553), .Y(n_550) );
AND2x2_ASAP7_75t_L g595 ( .A(n_551), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g690 ( .A(n_551), .B(n_570), .Y(n_690) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g646 ( .A(n_552), .B(n_571), .Y(n_646) );
INVx1_ASAP7_75t_L g658 ( .A(n_553), .Y(n_658) );
AND2x2_ASAP7_75t_L g669 ( .A(n_553), .B(n_656), .Y(n_669) );
AND2x2_ASAP7_75t_L g736 ( .A(n_553), .B(n_631), .Y(n_736) );
INVx2_ASAP7_75t_L g598 ( .A(n_554), .Y(n_598) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_565), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g688 ( .A(n_565), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_566), .B(n_649), .Y(n_652) );
INVx3_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g732 ( .A1(n_567), .A2(n_688), .B(n_733), .Y(n_732) );
AND2x4_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NOR2xp33_ASAP7_75t_SL g710 ( .A(n_570), .B(n_596), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_571), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g662 ( .A(n_571), .B(n_590), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_571), .B(n_597), .Y(n_739) );
AND2x2_ASAP7_75t_L g608 ( .A(n_572), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g675 ( .A(n_572), .Y(n_675) );
AOI21xp33_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_578), .B(n_582), .Y(n_573) );
NAND2x1_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_575), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g624 ( .A(n_575), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_SL g636 ( .A(n_575), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_575), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g660 ( .A(n_576), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_576), .B(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_576), .B(n_579), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
AOI211xp5_ASAP7_75t_L g647 ( .A1(n_579), .A2(n_618), .B(n_648), .C(n_650), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g665 ( .A1(n_579), .A2(n_666), .B1(n_669), .B2(n_670), .C(n_674), .Y(n_665) );
AND2x2_ASAP7_75t_L g661 ( .A(n_580), .B(n_614), .Y(n_661) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g621 ( .A(n_585), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g692 ( .A(n_585), .B(n_693), .Y(n_692) );
OAI211xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_588), .B(n_594), .C(n_619), .Y(n_586) );
NAND3xp33_ASAP7_75t_SL g705 ( .A(n_587), .B(n_706), .C(n_707), .Y(n_705) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_592), .Y(n_588) );
OR2x2_ASAP7_75t_L g678 ( .A(n_589), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AOI221xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_599), .B1(n_602), .B2(n_608), .C(n_610), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_596), .B(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_596), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g618 ( .A(n_601), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_601), .A2(n_658), .B1(n_659), .B2(n_660), .Y(n_657) );
OR2x2_ASAP7_75t_L g738 ( .A(n_601), .B(n_649), .Y(n_738) );
NAND2xp5_ASAP7_75t_SL g602 ( .A(n_603), .B(n_605), .Y(n_602) );
INVxp67_ASAP7_75t_L g712 ( .A(n_604), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_606), .B(n_727), .Y(n_726) );
INVxp67_ASAP7_75t_L g613 ( .A(n_607), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_609), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_609), .B(n_656), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_609), .B(n_676), .Y(n_715) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_613), .Y(n_639) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OR2x2_ASAP7_75t_L g729 ( .A(n_618), .B(n_649), .Y(n_729) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_624), .Y(n_620) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_SL g707 ( .A(n_624), .Y(n_707) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OAI322xp33_ASAP7_75t_SL g627 ( .A1(n_628), .A2(n_633), .A3(n_634), .B1(n_635), .B2(n_638), .C1(n_640), .C2(n_642), .Y(n_627) );
OAI322xp33_ASAP7_75t_L g709 ( .A1(n_628), .A2(n_710), .A3(n_711), .B1(n_712), .B2(n_713), .C1(n_714), .C2(n_716), .Y(n_709) );
CKINVDCx16_ASAP7_75t_R g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
INVx4_ASAP7_75t_L g643 ( .A(n_630), .Y(n_643) );
AND2x2_ASAP7_75t_L g704 ( .A(n_630), .B(n_656), .Y(n_704) );
AND2x2_ASAP7_75t_L g717 ( .A(n_630), .B(n_718), .Y(n_717) );
CKINVDCx16_ASAP7_75t_R g728 ( .A(n_633), .Y(n_728) );
INVx1_ASAP7_75t_L g706 ( .A(n_634), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
OR2x2_ASAP7_75t_L g640 ( .A(n_636), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g723 ( .A(n_636), .B(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_636), .B(n_677), .Y(n_734) );
OR2x2_ASAP7_75t_L g667 ( .A(n_639), .B(n_668), .Y(n_667) );
INVxp33_ASAP7_75t_L g684 ( .A(n_639), .Y(n_684) );
OAI221xp5_ASAP7_75t_SL g644 ( .A1(n_643), .A2(n_645), .B1(n_647), .B2(n_651), .C(n_653), .Y(n_644) );
NOR2xp67_ASAP7_75t_L g700 ( .A(n_643), .B(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g727 ( .A(n_643), .Y(n_727) );
INVx1_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
INVx3_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
AOI322xp5_ASAP7_75t_L g691 ( .A1(n_650), .A2(n_675), .A3(n_692), .B1(n_694), .B2(n_695), .C1(n_698), .C2(n_702), .Y(n_691) );
INVxp67_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_657), .B1(n_661), .B2(n_662), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_687), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_665), .B(n_680), .Y(n_664) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g698 ( .A(n_668), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
NAND2xp33_ASAP7_75t_SL g685 ( .A(n_671), .B(n_682), .Y(n_685) );
INVx1_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
OAI322xp33_ASAP7_75t_L g725 ( .A1(n_673), .A2(n_726), .A3(n_728), .B1(n_729), .B2(n_730), .C1(n_732), .C2(n_735), .Y(n_725) );
AOI21xp33_ASAP7_75t_SL g674 ( .A1(n_675), .A2(n_676), .B(n_678), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_683), .B(n_731), .Y(n_740) );
OAI211xp5_ASAP7_75t_SL g687 ( .A1(n_688), .A2(n_689), .B(n_691), .C(n_703), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NOR4xp25_ASAP7_75t_L g708 ( .A(n_709), .B(n_719), .C(n_725), .D(n_737), .Y(n_708) );
INVxp67_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
INVxp67_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
CKINVDCx14_ASAP7_75t_R g735 ( .A(n_736), .Y(n_735) );
OAI21xp5_ASAP7_75t_SL g737 ( .A1(n_738), .A2(n_739), .B(n_740), .Y(n_737) );
CKINVDCx16_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
INVx3_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
NAND2xp33_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
endmodule