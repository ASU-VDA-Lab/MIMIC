module fake_jpeg_12985_n_647 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_647);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_647;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_3),
.B(n_18),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_13),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_13),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_59),
.Y(n_162)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_60),
.Y(n_139)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_61),
.Y(n_153)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_62),
.Y(n_164)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_46),
.Y(n_63)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_63),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_28),
.B(n_8),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_64),
.B(n_68),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_28),
.B(n_8),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_65),
.B(n_75),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_22),
.B(n_31),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_67),
.B(n_109),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_19),
.B(n_7),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_70),
.Y(n_152)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_74),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_30),
.B(n_7),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_76),
.Y(n_167)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_77),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_79),
.Y(n_146)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_80),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_30),
.B(n_51),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_81),
.B(n_91),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_82),
.Y(n_182)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_83),
.Y(n_158)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

INVx6_ASAP7_75t_SL g86 ( 
.A(n_46),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_86),
.B(n_101),
.Y(n_142)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_87),
.Y(n_154)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_88),
.Y(n_157)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_89),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_22),
.B(n_9),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_90),
.B(n_0),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_32),
.B(n_35),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_92),
.Y(n_165)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g171 ( 
.A(n_93),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_94),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_32),
.B(n_9),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_95),
.B(n_52),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_96),
.Y(n_218)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_97),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_98),
.Y(n_198)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_99),
.Y(n_173)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_100),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_35),
.B(n_9),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_102),
.Y(n_211)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_25),
.Y(n_103)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_25),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_104),
.Y(n_219)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_105),
.Y(n_205)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_43),
.Y(n_106)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_106),
.Y(n_215)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_108),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_22),
.B(n_18),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_111),
.Y(n_190)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_40),
.Y(n_112)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_112),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_25),
.Y(n_113)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_113),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_54),
.Y(n_114)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_19),
.Y(n_115)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_34),
.Y(n_117)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_117),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_34),
.Y(n_118)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_119),
.Y(n_221)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_120),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_34),
.Y(n_121)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_121),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_22),
.B(n_6),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_122),
.B(n_124),
.Y(n_185)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_21),
.Y(n_123)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_123),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_41),
.B(n_6),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_34),
.Y(n_125)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_125),
.Y(n_207)
);

INVx3_ASAP7_75t_SL g126 ( 
.A(n_42),
.Y(n_126)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_126),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_38),
.Y(n_127)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_127),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_41),
.B(n_6),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_128),
.B(n_16),
.Y(n_189)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_38),
.Y(n_129)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_L g133 ( 
.A1(n_89),
.A2(n_21),
.B1(n_42),
.B2(n_55),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_133),
.A2(n_156),
.B1(n_200),
.B2(n_113),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_72),
.A2(n_21),
.B1(n_59),
.B2(n_42),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_137),
.A2(n_166),
.B1(n_204),
.B2(n_206),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_68),
.B(n_53),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_147),
.B(n_155),
.Y(n_273)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_151),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_90),
.B(n_53),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_66),
.A2(n_55),
.B1(n_48),
.B2(n_26),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_114),
.B(n_44),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_160),
.B(n_176),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_61),
.B(n_57),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_163),
.B(n_217),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_73),
.A2(n_55),
.B1(n_48),
.B2(n_50),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_60),
.A2(n_48),
.B1(n_57),
.B2(n_45),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_169),
.A2(n_213),
.B1(n_98),
.B2(n_85),
.Y(n_265)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_110),
.Y(n_175)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_175),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_78),
.B(n_52),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_177),
.B(n_178),
.Y(n_280)
);

AND2x2_ASAP7_75t_SL g178 ( 
.A(n_80),
.B(n_12),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_111),
.Y(n_180)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_180),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_197),
.Y(n_228)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_116),
.Y(n_191)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_191),
.Y(n_255)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_99),
.Y(n_195)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_195),
.Y(n_262)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_102),
.Y(n_196)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_196),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_70),
.A2(n_48),
.B1(n_26),
.B2(n_39),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_120),
.B(n_51),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_208),
.Y(n_230)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_62),
.Y(n_203)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_203),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_73),
.A2(n_49),
.B1(n_45),
.B2(n_36),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_126),
.A2(n_74),
.B1(n_129),
.B2(n_100),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_119),
.B(n_44),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_76),
.B(n_50),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_222),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_83),
.B(n_49),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_210),
.B(n_0),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_93),
.A2(n_36),
.B1(n_24),
.B2(n_39),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_106),
.B(n_24),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_82),
.B(n_10),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_173),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_223),
.B(n_270),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_161),
.Y(n_224)
);

NAND3xp33_ASAP7_75t_L g311 ( 
.A(n_224),
.B(n_295),
.C(n_139),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_159),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_225),
.B(n_227),
.Y(n_325)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_162),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_226),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_159),
.Y(n_227)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_144),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_229),
.Y(n_358)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_165),
.Y(n_231)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_231),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_216),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_232),
.Y(n_323)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_170),
.Y(n_233)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_233),
.Y(n_307)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_183),
.Y(n_236)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_236),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_133),
.A2(n_125),
.B1(n_121),
.B2(n_118),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_237),
.A2(n_267),
.B1(n_274),
.B2(n_288),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_238),
.A2(n_249),
.B1(n_212),
.B2(n_150),
.Y(n_312)
);

AO22x2_ASAP7_75t_L g240 ( 
.A1(n_178),
.A2(n_104),
.B1(n_96),
.B2(n_94),
.Y(n_240)
);

OA22x2_ASAP7_75t_L g339 ( 
.A1(n_240),
.A2(n_132),
.B1(n_152),
.B2(n_167),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_173),
.Y(n_241)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_241),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_130),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_242),
.Y(n_334)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_187),
.Y(n_243)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_243),
.Y(n_342)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_162),
.Y(n_244)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_244),
.Y(n_308)
);

INVx4_ASAP7_75t_SL g245 ( 
.A(n_161),
.Y(n_245)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_245),
.Y(n_353)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_162),
.Y(n_246)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_246),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_185),
.A2(n_98),
.B1(n_85),
.B2(n_77),
.Y(n_249)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_141),
.Y(n_250)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_250),
.Y(n_322)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_201),
.Y(n_251)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_251),
.Y(n_324)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_136),
.Y(n_254)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_254),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_214),
.Y(n_256)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_256),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_216),
.Y(n_257)
);

INVx8_ASAP7_75t_L g318 ( 
.A(n_257),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_135),
.Y(n_258)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_258),
.Y(n_360)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_198),
.Y(n_259)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_259),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_174),
.B(n_12),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_260),
.B(n_286),
.Y(n_336)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_221),
.Y(n_261)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_261),
.Y(n_335)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_220),
.Y(n_264)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_264),
.Y(n_347)
);

OA21x2_ASAP7_75t_L g331 ( 
.A1(n_265),
.A2(n_277),
.B(n_3),
.Y(n_331)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_214),
.Y(n_266)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_266),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_156),
.A2(n_37),
.B1(n_10),
.B2(n_12),
.Y(n_267)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_221),
.Y(n_268)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_268),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_138),
.A2(n_5),
.B1(n_17),
.B2(n_16),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_269),
.A2(n_271),
.B1(n_293),
.B2(n_297),
.Y(n_346)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_157),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_135),
.A2(n_13),
.B1(n_5),
.B2(n_37),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_200),
.A2(n_37),
.B1(n_5),
.B2(n_2),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_192),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_275),
.B(n_278),
.Y(n_315)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_172),
.Y(n_276)
);

INVx3_ASAP7_75t_SL g305 ( 
.A(n_276),
.Y(n_305)
);

O2A1O1Ixp33_ASAP7_75t_SL g277 ( 
.A1(n_163),
.A2(n_37),
.B(n_5),
.C(n_2),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_172),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_218),
.Y(n_279)
);

BUFx4f_ASAP7_75t_L g348 ( 
.A(n_279),
.Y(n_348)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_184),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_281),
.B(n_284),
.Y(n_316)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_184),
.Y(n_282)
);

BUFx24_ASAP7_75t_L g356 ( 
.A(n_282),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_217),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_283),
.Y(n_332)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_131),
.Y(n_284)
);

AND2x2_ASAP7_75t_SL g285 ( 
.A(n_143),
.B(n_177),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_158),
.C(n_204),
.Y(n_306)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_134),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_287),
.A2(n_205),
.B1(n_153),
.B2(n_188),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_194),
.A2(n_37),
.B1(n_1),
.B2(n_3),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_179),
.B(n_0),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_289),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_140),
.B(n_1),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_290),
.B(n_292),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_211),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_291),
.B(n_298),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_142),
.B(n_1),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_211),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_146),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_294),
.Y(n_310)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_145),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_148),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_296),
.Y(n_321)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_190),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_215),
.B(n_1),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_149),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_299),
.A2(n_219),
.B1(n_171),
.B2(n_4),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_207),
.A2(n_3),
.B1(n_4),
.B2(n_210),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_300),
.A2(n_166),
.B1(n_206),
.B2(n_137),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_154),
.B(n_3),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_301),
.B(n_4),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_239),
.B(n_230),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_302),
.B(n_320),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_303),
.A2(n_313),
.B1(n_331),
.B2(n_339),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_306),
.B(n_317),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_247),
.A2(n_186),
.B(n_164),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_309),
.A2(n_317),
.B(n_333),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_311),
.B(n_353),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_312),
.A2(n_337),
.B1(n_300),
.B2(n_288),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_234),
.A2(n_193),
.B1(n_181),
.B2(n_168),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_280),
.A2(n_199),
.B(n_190),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_285),
.B(n_199),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_327),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_280),
.B(n_150),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_328),
.B(n_329),
.C(n_293),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_253),
.B(n_193),
.C(n_132),
.Y(n_329)
);

O2A1O1Ixp33_ASAP7_75t_L g333 ( 
.A1(n_277),
.A2(n_283),
.B(n_234),
.C(n_245),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_240),
.A2(n_168),
.B1(n_181),
.B2(n_152),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_287),
.B(n_240),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_338),
.B(n_351),
.Y(n_389)
);

OAI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_269),
.A2(n_167),
.B1(n_182),
.B2(n_218),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_344),
.A2(n_258),
.B1(n_358),
.B2(n_353),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_289),
.B(n_182),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_355),
.B(n_263),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_359),
.A2(n_256),
.B1(n_242),
.B2(n_299),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g426 ( 
.A1(n_362),
.A2(n_372),
.B1(n_392),
.B2(n_396),
.Y(n_426)
);

MAJx2_ASAP7_75t_L g363 ( 
.A(n_328),
.B(n_228),
.C(n_272),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_363),
.B(n_375),
.C(n_393),
.Y(n_418)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_304),
.Y(n_364)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_364),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_306),
.A2(n_271),
.B(n_266),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_366),
.A2(n_346),
.B(n_312),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_356),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_367),
.B(n_369),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_338),
.A2(n_237),
.B1(n_274),
.B2(n_267),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_368),
.A2(n_377),
.B1(n_398),
.B2(n_326),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_356),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_360),
.Y(n_371)
);

BUFx4f_ASAP7_75t_SL g446 ( 
.A(n_371),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_L g372 ( 
.A1(n_313),
.A2(n_219),
.B1(n_252),
.B2(n_235),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_318),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_373),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_309),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_374),
.B(n_382),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_320),
.B(n_273),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_378),
.A2(n_331),
.B(n_357),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_302),
.B(n_248),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_379),
.B(n_387),
.Y(n_411)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_348),
.Y(n_380)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_380),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_333),
.A2(n_241),
.B(n_262),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_381),
.A2(n_400),
.B(n_350),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_340),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_347),
.Y(n_383)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_383),
.Y(n_416)
);

CKINVDCx14_ASAP7_75t_R g384 ( 
.A(n_325),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_384),
.Y(n_421)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_347),
.Y(n_385)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_385),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_327),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_386),
.B(n_391),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_356),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_314),
.Y(n_388)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_388),
.Y(n_425)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_307),
.Y(n_390)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_390),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_318),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_329),
.B(n_255),
.C(n_261),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_351),
.B(n_282),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_394),
.B(n_402),
.Y(n_428)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_330),
.Y(n_395)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_395),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_L g396 ( 
.A1(n_303),
.A2(n_276),
.B1(n_232),
.B2(n_257),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_361),
.B(n_268),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_397),
.B(n_408),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_337),
.A2(n_279),
.B1(n_250),
.B2(n_259),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_319),
.A2(n_226),
.B1(n_244),
.B2(n_246),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_399),
.A2(n_358),
.B1(n_305),
.B2(n_314),
.Y(n_415)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_348),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_336),
.B(n_343),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_403),
.B(n_407),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_404),
.B(n_315),
.C(n_321),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_405),
.B(n_406),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_323),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_316),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_332),
.B(n_310),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_410),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_381),
.B(n_339),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_412),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_414),
.B(n_437),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_415),
.A2(n_443),
.B1(n_398),
.B2(n_377),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_374),
.A2(n_386),
.B1(n_365),
.B2(n_364),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_417),
.A2(n_438),
.B(n_441),
.Y(n_459)
);

OAI21xp33_ASAP7_75t_SL g419 ( 
.A1(n_381),
.A2(n_331),
.B(n_339),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_419),
.B(n_376),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_408),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_422),
.B(n_433),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_401),
.B(n_339),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_424),
.B(n_442),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_432),
.B(n_434),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_367),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_375),
.B(n_404),
.C(n_393),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_370),
.B(n_342),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_401),
.A2(n_326),
.B(n_308),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_440),
.A2(n_413),
.B1(n_426),
.B2(n_421),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_382),
.A2(n_360),
.B1(n_322),
.B2(n_349),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_376),
.A2(n_323),
.B1(n_335),
.B2(n_352),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_363),
.B(n_335),
.C(n_352),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_444),
.B(n_407),
.Y(n_450)
);

XOR2x2_ASAP7_75t_SL g445 ( 
.A(n_389),
.B(n_305),
.Y(n_445)
);

A2O1A1Ixp33_ASAP7_75t_L g470 ( 
.A1(n_445),
.A2(n_395),
.B(n_390),
.C(n_350),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g494 ( 
.A(n_448),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_450),
.B(n_418),
.Y(n_488)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_420),
.Y(n_451)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_451),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_440),
.A2(n_389),
.B1(n_366),
.B2(n_370),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_452),
.A2(n_461),
.B1(n_462),
.B2(n_466),
.Y(n_486)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_420),
.Y(n_454)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_454),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_428),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_455),
.B(n_456),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_428),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_410),
.A2(n_400),
.B1(n_378),
.B2(n_399),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_427),
.A2(n_378),
.B1(n_403),
.B2(n_394),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_463),
.A2(n_476),
.B1(n_477),
.B2(n_480),
.Y(n_497)
);

OAI32xp33_ASAP7_75t_L g464 ( 
.A1(n_436),
.A2(n_427),
.A3(n_429),
.B1(n_445),
.B2(n_411),
.Y(n_464)
);

AOI221xp5_ASAP7_75t_L g513 ( 
.A1(n_464),
.A2(n_446),
.B1(n_341),
.B2(n_345),
.C(n_334),
.Y(n_513)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_416),
.Y(n_465)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_465),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_417),
.A2(n_379),
.B1(n_368),
.B2(n_397),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_436),
.A2(n_363),
.B1(n_391),
.B2(n_385),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_467),
.A2(n_473),
.B1(n_415),
.B2(n_409),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_411),
.B(n_383),
.Y(n_468)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_468),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_437),
.B(n_369),
.Y(n_469)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_469),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_470),
.A2(n_438),
.B(n_412),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_422),
.B(n_387),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_471),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_430),
.B(n_371),
.Y(n_472)
);

CKINVDCx14_ASAP7_75t_R g484 ( 
.A(n_472),
.Y(n_484)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_416),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_474),
.B(n_475),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_433),
.B(n_373),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_443),
.A2(n_392),
.B1(n_373),
.B2(n_406),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_419),
.A2(n_412),
.B1(n_424),
.B2(n_414),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_430),
.Y(n_478)
);

INVxp33_ASAP7_75t_L g499 ( 
.A(n_478),
.Y(n_499)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_423),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_412),
.A2(n_392),
.B1(n_406),
.B2(n_402),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_481),
.A2(n_482),
.B1(n_447),
.B2(n_380),
.Y(n_502)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_423),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_409),
.Y(n_483)
);

CKINVDCx16_ASAP7_75t_R g493 ( 
.A(n_483),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_478),
.B(n_413),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_487),
.B(n_507),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_488),
.B(n_513),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_SL g490 ( 
.A(n_458),
.B(n_434),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_490),
.B(n_495),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_458),
.B(n_418),
.C(n_432),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_492),
.B(n_500),
.C(n_510),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_450),
.B(n_444),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_496),
.A2(n_515),
.B(n_470),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_448),
.A2(n_445),
.B1(n_429),
.B2(n_442),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_498),
.A2(n_501),
.B1(n_459),
.B2(n_460),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_452),
.B(n_424),
.C(n_425),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_479),
.A2(n_421),
.B1(n_441),
.B2(n_425),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_502),
.B(n_482),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_463),
.A2(n_409),
.B1(n_435),
.B2(n_439),
.Y(n_504)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_504),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_506),
.A2(n_477),
.B1(n_457),
.B2(n_459),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_467),
.B(n_439),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_461),
.A2(n_431),
.B1(n_435),
.B2(n_447),
.Y(n_508)
);

XOR2x1_ASAP7_75t_L g526 ( 
.A(n_508),
.B(n_471),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_464),
.B(n_324),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_462),
.B(n_324),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_512),
.B(n_514),
.C(n_517),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_451),
.B(n_322),
.C(n_349),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_460),
.A2(n_308),
.B(n_354),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_466),
.B(n_354),
.Y(n_517)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_489),
.Y(n_519)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_519),
.Y(n_549)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_489),
.Y(n_520)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_520),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_521),
.A2(n_532),
.B1(n_533),
.B2(n_543),
.Y(n_570)
);

CKINVDCx16_ASAP7_75t_R g522 ( 
.A(n_491),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_522),
.B(n_535),
.Y(n_548)
);

NOR3xp33_ASAP7_75t_L g524 ( 
.A(n_503),
.B(n_449),
.C(n_454),
.Y(n_524)
);

CKINVDCx14_ASAP7_75t_R g567 ( 
.A(n_524),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_526),
.B(n_547),
.Y(n_550)
);

AOI22x1_ASAP7_75t_L g527 ( 
.A1(n_494),
.A2(n_460),
.B1(n_457),
.B2(n_498),
.Y(n_527)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_527),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_515),
.B(n_457),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_528),
.Y(n_551)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_503),
.Y(n_529)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_529),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_511),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_511),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_505),
.Y(n_534)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_534),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_493),
.B(n_449),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_536),
.A2(n_544),
.B1(n_508),
.B2(n_494),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_490),
.B(n_460),
.C(n_483),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_537),
.B(n_540),
.Y(n_561)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_538),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_492),
.B(n_468),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_539),
.B(n_542),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_488),
.B(n_469),
.C(n_456),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g564 ( 
.A1(n_541),
.A2(n_496),
.B(n_499),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_495),
.B(n_455),
.C(n_472),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_486),
.A2(n_453),
.B1(n_481),
.B2(n_470),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_497),
.A2(n_473),
.B1(n_453),
.B2(n_475),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_485),
.B(n_480),
.Y(n_545)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_545),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_500),
.B(n_474),
.C(n_465),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_539),
.B(n_510),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g577 ( 
.A(n_554),
.B(n_569),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_520),
.B(n_485),
.Y(n_555)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_555),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_525),
.B(n_509),
.Y(n_556)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_556),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_538),
.B(n_516),
.Y(n_558)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_558),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_SL g562 ( 
.A(n_540),
.B(n_499),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_562),
.A2(n_560),
.B1(n_559),
.B2(n_556),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_564),
.B(n_521),
.Y(n_579)
);

OAI22xp33_ASAP7_75t_SL g565 ( 
.A1(n_544),
.A2(n_516),
.B1(n_509),
.B2(n_506),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_565),
.B(n_566),
.Y(n_582)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_518),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_543),
.B(n_484),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_568),
.B(n_517),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_563),
.B(n_530),
.C(n_547),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_572),
.B(n_575),
.Y(n_596)
);

FAx1_ASAP7_75t_SL g573 ( 
.A(n_564),
.B(n_537),
.CI(n_542),
.CON(n_573),
.SN(n_573)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_573),
.B(n_560),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_567),
.B(n_563),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_SL g595 ( 
.A(n_574),
.B(n_580),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_561),
.B(n_530),
.C(n_546),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_SL g576 ( 
.A1(n_570),
.A2(n_486),
.B1(n_536),
.B2(n_541),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_576),
.A2(n_578),
.B1(n_589),
.B2(n_501),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_SL g578 ( 
.A1(n_568),
.A2(n_531),
.B1(n_526),
.B2(n_523),
.Y(n_578)
);

XOR2xp5_ASAP7_75t_L g592 ( 
.A(n_579),
.B(n_558),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_562),
.B(n_514),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_550),
.B(n_546),
.C(n_554),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_581),
.B(n_587),
.Y(n_600)
);

XOR2xp5_ASAP7_75t_L g583 ( 
.A(n_550),
.B(n_531),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_583),
.B(n_566),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_586),
.B(n_588),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_569),
.B(n_523),
.C(n_527),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_559),
.A2(n_527),
.B1(n_512),
.B2(n_476),
.Y(n_589)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_592),
.B(n_593),
.Y(n_609)
);

OAI21xp5_ASAP7_75t_SL g594 ( 
.A1(n_582),
.A2(n_571),
.B(n_551),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_594),
.A2(n_584),
.B(n_585),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_582),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_SL g614 ( 
.A(n_597),
.B(n_599),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_572),
.B(n_551),
.C(n_571),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_598),
.B(n_601),
.C(n_577),
.Y(n_608)
);

CKINVDCx16_ASAP7_75t_R g599 ( 
.A(n_588),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_583),
.B(n_555),
.C(n_528),
.Y(n_601)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_602),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_590),
.B(n_548),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_603),
.B(n_604),
.Y(n_612)
);

INVxp33_ASAP7_75t_SL g604 ( 
.A(n_578),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_573),
.B(n_553),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_SL g620 ( 
.A(n_605),
.B(n_600),
.Y(n_620)
);

XOR2xp5_ASAP7_75t_L g606 ( 
.A(n_579),
.B(n_528),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_606),
.B(n_573),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_SL g617 ( 
.A1(n_607),
.A2(n_587),
.B1(n_577),
.B2(n_581),
.Y(n_617)
);

XNOR2x1_ASAP7_75t_L g629 ( 
.A(n_608),
.B(n_617),
.Y(n_629)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_611),
.Y(n_627)
);

A2O1A1Ixp33_ASAP7_75t_SL g630 ( 
.A1(n_613),
.A2(n_610),
.B(n_614),
.C(n_615),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_591),
.A2(n_585),
.B1(n_576),
.B2(n_589),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_615),
.B(n_618),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_SL g616 ( 
.A1(n_591),
.A2(n_552),
.B1(n_553),
.B2(n_549),
.Y(n_616)
);

XOR2xp5_ASAP7_75t_L g625 ( 
.A(n_616),
.B(n_552),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_596),
.B(n_598),
.C(n_593),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_595),
.B(n_575),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_619),
.B(n_620),
.Y(n_626)
);

XOR2xp5_ASAP7_75t_L g621 ( 
.A(n_617),
.B(n_601),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_621),
.B(n_628),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_L g622 ( 
.A1(n_612),
.A2(n_594),
.B(n_607),
.Y(n_622)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_622),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_608),
.B(n_592),
.C(n_606),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_624),
.B(n_618),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_625),
.B(n_446),
.Y(n_636)
);

XOR2xp5_ASAP7_75t_L g628 ( 
.A(n_609),
.B(n_549),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g633 ( 
.A(n_630),
.B(n_609),
.C(n_557),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g640 ( 
.A(n_631),
.B(n_636),
.C(n_621),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_SL g632 ( 
.A1(n_626),
.A2(n_612),
.B(n_613),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_632),
.A2(n_633),
.B(n_634),
.Y(n_641)
);

A2O1A1Ixp33_ASAP7_75t_L g634 ( 
.A1(n_627),
.A2(n_505),
.B(n_557),
.C(n_446),
.Y(n_634)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g638 ( 
.A1(n_635),
.A2(n_630),
.B(n_628),
.C(n_629),
.D(n_623),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_638),
.B(n_639),
.Y(n_643)
);

OAI21xp33_ASAP7_75t_L g639 ( 
.A1(n_637),
.A2(n_630),
.B(n_629),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_640),
.B(n_631),
.Y(n_642)
);

OAI21xp5_ASAP7_75t_L g644 ( 
.A1(n_642),
.A2(n_641),
.B(n_446),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_SL g645 ( 
.A1(n_644),
.A2(n_643),
.B(n_345),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_SL g646 ( 
.A1(n_645),
.A2(n_334),
.B(n_348),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_646),
.B(n_341),
.Y(n_647)
);


endmodule