module real_jpeg_13950_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_288, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_288;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_249;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_281;
wire n_131;
wire n_276;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_200;
wire n_164;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_267;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_285;
wire n_160;
wire n_45;
wire n_211;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_278;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_0),
.A2(n_23),
.B1(n_26),
.B2(n_36),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_0),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_0),
.A2(n_36),
.B1(n_45),
.B2(n_46),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_0),
.A2(n_8),
.B(n_32),
.C(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_0),
.A2(n_36),
.B1(n_56),
.B2(n_57),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_0),
.B(n_37),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_0),
.B(n_54),
.C(n_57),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_0),
.B(n_44),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_0),
.B(n_29),
.C(n_33),
.Y(n_165)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_3),
.Y(n_98)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_40),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_6),
.A2(n_23),
.B1(n_26),
.B2(n_40),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_6),
.A2(n_40),
.B1(n_56),
.B2(n_57),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_6),
.A2(n_40),
.B1(n_45),
.B2(n_46),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

AO22x1_ASAP7_75t_L g44 ( 
.A1(n_8),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_10),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_10),
.A2(n_23),
.B1(n_26),
.B2(n_48),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_10),
.A2(n_48),
.B1(n_56),
.B2(n_57),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_11),
.A2(n_15),
.B(n_284),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_11),
.B(n_285),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_12),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_12),
.A2(n_25),
.B1(n_32),
.B2(n_33),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_12),
.A2(n_25),
.B1(n_45),
.B2(n_46),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_12),
.A2(n_25),
.B1(n_56),
.B2(n_57),
.Y(n_112)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_13),
.Y(n_285)
);

AOI21xp33_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_280),
.B(n_282),
.Y(n_15)
);

AO21x1_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_72),
.B(n_279),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_69),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_18),
.B(n_69),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_62),
.C(n_66),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_19),
.B(n_276),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_38),
.C(n_49),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_20),
.A2(n_105),
.B1(n_115),
.B2(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_20),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_20),
.B(n_115),
.C(n_178),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_20),
.A2(n_81),
.B1(n_82),
.B2(n_180),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_20),
.A2(n_180),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_27),
.B1(n_35),
.B2(n_37),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OA21x2_ASAP7_75t_L g168 ( 
.A1(n_22),
.A2(n_31),
.B(n_68),
.Y(n_168)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_26),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_27),
.B(n_35),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_27),
.B(n_37),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_29),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_31),
.A2(n_67),
.B(n_68),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_31),
.A2(n_67),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_42),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

INVxp33_ASAP7_75t_L g236 ( 
.A(n_35),
.Y(n_236)
);

OAI21xp33_ASAP7_75t_SL g94 ( 
.A1(n_36),
.A2(n_42),
.B(n_45),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_36),
.B(n_101),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_36),
.B(n_60),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_38),
.A2(n_49),
.B1(n_254),
.B2(n_268),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_38),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_41),
.B1(n_44),
.B2(n_47),
.Y(n_38)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_39),
.Y(n_256)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_41),
.B(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_46),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_46),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_49),
.A2(n_254),
.B1(n_255),
.B2(n_257),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_49),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_49),
.B(n_168),
.C(n_255),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_60),
.B(n_61),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_50),
.A2(n_60),
.B(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_90),
.Y(n_89)
);

AO22x1_ASAP7_75t_SL g120 ( 
.A1(n_51),
.A2(n_55),
.B1(n_88),
.B2(n_90),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_51),
.A2(n_55),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

NOR2x1_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

AO22x1_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_56),
.B(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_57),
.B(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OA21x2_ASAP7_75t_L g86 ( 
.A1(n_60),
.A2(n_87),
.B(n_89),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_60),
.A2(n_89),
.B(n_220),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_61),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_62),
.B(n_66),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_64),
.A2(n_65),
.B1(n_83),
.B2(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_64),
.A2(n_65),
.B(n_106),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_83),
.B(n_84),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_65),
.A2(n_84),
.B(n_256),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_69),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_69),
.B(n_281),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_71),
.B(n_237),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_274),
.B(n_278),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_246),
.B(n_271),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_224),
.B(n_245),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_207),
.B(n_223),
.Y(n_75)
);

OAI321xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_175),
.A3(n_202),
.B1(n_205),
.B2(n_206),
.C(n_288),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_157),
.B(n_174),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_123),
.B(n_156),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_102),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_80),
.B(n_102),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_86),
.C(n_91),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_81),
.A2(n_82),
.B1(n_86),
.B2(n_140),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_81),
.A2(n_82),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_82),
.B(n_167),
.C(n_172),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_82),
.B(n_180),
.C(n_212),
.Y(n_244)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_86),
.B(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_86),
.A2(n_127),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_86),
.A2(n_140),
.B1(n_182),
.B2(n_184),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_90),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_91),
.A2(n_92),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_95),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_96),
.A2(n_100),
.B1(n_101),
.B2(n_112),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_97),
.B(n_200),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_100),
.A2(n_101),
.B1(n_183),
.B2(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_112),
.B(n_113),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_101),
.A2(n_113),
.B(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_117),
.B2(n_118),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_103),
.B(n_120),
.C(n_121),
.Y(n_158)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_107),
.B1(n_115),
.B2(n_116),
.Y(n_104)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_105),
.B(n_108),
.C(n_111),
.Y(n_161)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_110),
.B(n_138),
.Y(n_148)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_111),
.B(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_115),
.A2(n_240),
.B(n_243),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_115),
.B(n_240),
.Y(n_243)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_119),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_120),
.A2(n_122),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_132),
.C(n_134),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_120),
.A2(n_122),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_120),
.B(n_199),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_150),
.B(n_155),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_136),
.B(n_149),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_126),
.B(n_129),
.Y(n_149)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_129)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_130),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_131),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_133),
.A2(n_134),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_134),
.B(n_146),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_163),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_141),
.B(n_148),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_140),
.B(n_182),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_145),
.B(n_147),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_151),
.B(n_152),
.Y(n_155)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_158),
.B(n_159),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_166),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_162),
.C(n_166),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_167),
.A2(n_168),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_167),
.B(n_190),
.C(n_195),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_167),
.A2(n_168),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_167),
.A2(n_168),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_168),
.B(n_265),
.C(n_269),
.Y(n_277)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_186),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_186),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_181),
.C(n_185),
.Y(n_176)
);

FAx1_ASAP7_75t_SL g204 ( 
.A(n_177),
.B(n_181),
.CI(n_185),
.CON(n_204),
.SN(n_204)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_182),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_201),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_196),
.B2(n_197),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_197),
.C(n_201),
.Y(n_222)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_203),
.B(n_204),
.Y(n_205)
);

BUFx24_ASAP7_75t_SL g287 ( 
.A(n_204),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_222),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_222),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_211),
.C(n_216),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_216),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_219),
.B2(n_221),
.Y(n_216)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_217),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_219),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_217),
.A2(n_221),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_221),
.A2(n_230),
.B(n_235),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_226),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_244),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_238),
.B2(n_239),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_238),
.C(n_244),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_243),
.A2(n_250),
.B1(n_251),
.B2(n_258),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_243),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_261),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_260),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_260),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_259),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_258),
.C(n_259),
.Y(n_270)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_255),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_261),
.A2(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_270),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_270),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_269),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_277),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_277),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);


endmodule