module fake_netlist_6_387_n_1621 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1621);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1621;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_544;
wire n_250;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_107),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_108),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_60),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_76),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_1),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_112),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_25),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_44),
.Y(n_159)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_75),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_110),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_46),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_65),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_13),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_79),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_42),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_25),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_13),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_100),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_1),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_37),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_36),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_118),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_30),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_142),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_94),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_135),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_81),
.Y(n_181)
);

BUFx2_ASAP7_75t_SL g182 ( 
.A(n_126),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_35),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_63),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_50),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_23),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_123),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_138),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_136),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_117),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_36),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_8),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_23),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_45),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_18),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_143),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_34),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_35),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_12),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_61),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_124),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_55),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_5),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_146),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_16),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_19),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_99),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_70),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_27),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_140),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_2),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_82),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_15),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_33),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_103),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_91),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_109),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_121),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_73),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_137),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_132),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_38),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_15),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_104),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_74),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_12),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_53),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_4),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_28),
.Y(n_229)
);

BUFx2_ASAP7_75t_SL g230 ( 
.A(n_148),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_57),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_125),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_88),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_42),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_89),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_86),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_68),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_69),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_19),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_113),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_102),
.Y(n_241)
);

BUFx10_ASAP7_75t_L g242 ( 
.A(n_9),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_17),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_78),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_38),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_120),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_0),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_128),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_84),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_3),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_27),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_80),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_48),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_83),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_98),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_28),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_115),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_114),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_105),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_116),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_2),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_144),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_134),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_9),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_52),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_47),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_64),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_85),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_39),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_34),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_3),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_14),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_97),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_29),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_11),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_37),
.Y(n_276)
);

INVxp67_ASAP7_75t_SL g277 ( 
.A(n_141),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_32),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_45),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_133),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_58),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_67),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_56),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_92),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_24),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_5),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_127),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_26),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_20),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_122),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_39),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_10),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_44),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_17),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_6),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_8),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_129),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_29),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_87),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_59),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_18),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_192),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_285),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_183),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_200),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_292),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_0),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_292),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_225),
.B(n_4),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_177),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_244),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_164),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_191),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_169),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_193),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_180),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_195),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_177),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_169),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_176),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_176),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_223),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_L g323 ( 
.A(n_160),
.B(n_6),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_189),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_197),
.Y(n_325)
);

NOR2xp67_ASAP7_75t_L g326 ( 
.A(n_160),
.B(n_7),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_158),
.Y(n_327)
);

INVxp33_ASAP7_75t_L g328 ( 
.A(n_155),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_282),
.B(n_7),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_200),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_159),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_265),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_284),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_163),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_255),
.Y(n_335)
);

NOR2xp67_ASAP7_75t_L g336 ( 
.A(n_160),
.B(n_10),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_190),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_186),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_198),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_263),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_242),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_194),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_228),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_243),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_251),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_199),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_227),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_274),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_223),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_227),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_229),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_151),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_282),
.B(n_11),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_229),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_264),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_264),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_205),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_275),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_206),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_242),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_294),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_252),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_252),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_153),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_301),
.Y(n_365)
);

INVxp33_ASAP7_75t_L g366 ( 
.A(n_301),
.Y(n_366)
);

INVxp33_ASAP7_75t_SL g367 ( 
.A(n_158),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_242),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_185),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_150),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_187),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_150),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_156),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_156),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_209),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_211),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_181),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_370),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_305),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_327),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_377),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_369),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_310),
.Y(n_383)
);

NAND2xp33_ASAP7_75t_L g384 ( 
.A(n_303),
.B(n_168),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_305),
.Y(n_385)
);

NOR2xp67_ASAP7_75t_L g386 ( 
.A(n_318),
.B(n_232),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_371),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_318),
.B(n_152),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_330),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_377),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_330),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_304),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_304),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_372),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_303),
.B(n_152),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_310),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_372),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_312),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_313),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_316),
.B(n_170),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_373),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_313),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_318),
.B(n_154),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_373),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_374),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_315),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_374),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_314),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_363),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_314),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_319),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_363),
.B(n_154),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_319),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_320),
.Y(n_414)
);

INVx6_ASAP7_75t_L g415 ( 
.A(n_337),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_315),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_320),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_321),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_321),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_317),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_362),
.B(n_181),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_317),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_322),
.Y(n_423)
);

INVx5_ASAP7_75t_L g424 ( 
.A(n_363),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_322),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_349),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_325),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_349),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_324),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_351),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_351),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_354),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_325),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_364),
.B(n_161),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_339),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_347),
.B(n_161),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_350),
.B(n_249),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_306),
.B(n_157),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_332),
.Y(n_439)
);

OA21x2_ASAP7_75t_L g440 ( 
.A1(n_354),
.A2(n_356),
.B(n_355),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_339),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_355),
.Y(n_442)
);

AND2x2_ASAP7_75t_SL g443 ( 
.A(n_307),
.B(n_216),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_356),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_365),
.Y(n_445)
);

AND2x6_ASAP7_75t_L g446 ( 
.A(n_353),
.B(n_216),
.Y(n_446)
);

NOR2xp67_ASAP7_75t_L g447 ( 
.A(n_365),
.B(n_290),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_346),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g449 ( 
.A(n_436),
.B(n_368),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_409),
.B(n_308),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_409),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_436),
.B(n_367),
.Y(n_452)
);

OR2x2_ASAP7_75t_L g453 ( 
.A(n_380),
.B(n_311),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_420),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_379),
.B(n_323),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_409),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_383),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_413),
.Y(n_458)
);

INVx4_ASAP7_75t_SL g459 ( 
.A(n_446),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_383),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_379),
.B(n_326),
.Y(n_461)
);

BUFx8_ASAP7_75t_SL g462 ( 
.A(n_398),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_400),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_379),
.B(n_336),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_437),
.B(n_352),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_396),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_396),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_385),
.B(n_335),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_443),
.A2(n_340),
.B1(n_375),
.B2(n_359),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_395),
.B(n_346),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_443),
.A2(n_329),
.B1(n_309),
.B2(n_366),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_440),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_440),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_440),
.Y(n_474)
);

INVx2_ASAP7_75t_SL g475 ( 
.A(n_415),
.Y(n_475)
);

NAND2x1p5_ASAP7_75t_L g476 ( 
.A(n_443),
.B(n_262),
.Y(n_476)
);

AND2x6_ASAP7_75t_L g477 ( 
.A(n_438),
.B(n_216),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_440),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_437),
.B(n_357),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_440),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_378),
.Y(n_481)
);

OR2x2_ASAP7_75t_L g482 ( 
.A(n_380),
.B(n_357),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_415),
.Y(n_483)
);

INVxp67_ASAP7_75t_SL g484 ( 
.A(n_385),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_413),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_385),
.B(n_200),
.Y(n_486)
);

OR2x2_ASAP7_75t_SL g487 ( 
.A(n_415),
.B(n_166),
.Y(n_487)
);

AND2x6_ASAP7_75t_L g488 ( 
.A(n_438),
.B(n_216),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_378),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_424),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_381),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_400),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_388),
.B(n_359),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_388),
.B(n_375),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_389),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_415),
.Y(n_496)
);

AND2x6_ASAP7_75t_L g497 ( 
.A(n_438),
.B(n_216),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_415),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_403),
.B(n_376),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_389),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_392),
.B(n_376),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_389),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_429),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_391),
.B(n_446),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_391),
.B(n_200),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_391),
.B(n_200),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_446),
.B(n_200),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_413),
.Y(n_508)
);

AND2x6_ASAP7_75t_L g509 ( 
.A(n_421),
.B(n_219),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_403),
.B(n_302),
.Y(n_510)
);

INVxp33_ASAP7_75t_SL g511 ( 
.A(n_382),
.Y(n_511)
);

AND2x6_ASAP7_75t_L g512 ( 
.A(n_421),
.B(n_219),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_412),
.B(n_341),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_446),
.B(n_200),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_390),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_393),
.B(n_360),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_446),
.B(n_200),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_446),
.B(n_277),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_420),
.B(n_328),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_399),
.B(n_162),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_434),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_387),
.Y(n_522)
);

CKINVDCx6p67_ASAP7_75t_R g523 ( 
.A(n_439),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_422),
.B(n_331),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_421),
.B(n_334),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_441),
.A2(n_203),
.B1(n_276),
.B2(n_261),
.Y(n_526)
);

INVx1_ASAP7_75t_SL g527 ( 
.A(n_422),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_441),
.B(n_338),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_394),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_446),
.A2(n_361),
.B1(n_358),
.B2(n_348),
.Y(n_530)
);

INVxp33_ASAP7_75t_SL g531 ( 
.A(n_402),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_446),
.B(n_184),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_446),
.B(n_204),
.Y(n_533)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_424),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_394),
.Y(n_535)
);

NAND2xp33_ASAP7_75t_L g536 ( 
.A(n_412),
.B(n_219),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_413),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_434),
.B(n_342),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_384),
.A2(n_333),
.B1(n_241),
.B2(n_179),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_386),
.B(n_343),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_406),
.B(n_162),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_424),
.B(n_218),
.Y(n_542)
);

BUFx4f_ASAP7_75t_L g543 ( 
.A(n_413),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_416),
.B(n_167),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_401),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_427),
.B(n_167),
.Y(n_546)
);

OR2x2_ASAP7_75t_L g547 ( 
.A(n_433),
.B(n_165),
.Y(n_547)
);

BUFx10_ASAP7_75t_L g548 ( 
.A(n_435),
.Y(n_548)
);

NAND3xp33_ASAP7_75t_L g549 ( 
.A(n_448),
.B(n_345),
.C(n_344),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_401),
.Y(n_550)
);

BUFx10_ASAP7_75t_L g551 ( 
.A(n_408),
.Y(n_551)
);

OR2x6_ASAP7_75t_L g552 ( 
.A(n_447),
.B(n_182),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_413),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_425),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_407),
.B(n_171),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_410),
.A2(n_219),
.B1(n_237),
.B2(n_254),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_425),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_425),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_386),
.B(n_171),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_424),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_410),
.A2(n_219),
.B1(n_237),
.B2(n_221),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_407),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_447),
.B(n_175),
.Y(n_563)
);

AND2x6_ASAP7_75t_L g564 ( 
.A(n_445),
.B(n_237),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_408),
.A2(n_300),
.B1(n_299),
.B2(n_175),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_425),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_411),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_411),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_425),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_418),
.B(n_178),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_424),
.B(n_178),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_424),
.B(n_410),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_424),
.B(n_179),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_L g574 ( 
.A1(n_410),
.A2(n_237),
.B1(n_253),
.B2(n_231),
.Y(n_574)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_418),
.B(n_172),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_419),
.B(n_212),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_419),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_425),
.B(n_212),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_423),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_423),
.A2(n_241),
.B1(n_300),
.B2(n_299),
.Y(n_580)
);

NAND2xp33_ASAP7_75t_R g581 ( 
.A(n_426),
.B(n_246),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_426),
.A2(n_237),
.B1(n_248),
.B2(n_240),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_428),
.B(n_222),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_430),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_430),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_430),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_428),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_426),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_430),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_430),
.Y(n_590)
);

OR2x2_ASAP7_75t_L g591 ( 
.A(n_432),
.B(n_278),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_430),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_426),
.B(n_246),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_519),
.B(n_524),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_521),
.B(n_430),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_452),
.B(n_257),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_521),
.B(n_279),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_493),
.B(n_397),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_494),
.B(n_397),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_513),
.B(n_257),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_499),
.B(n_397),
.Y(n_601)
);

OAI22xp33_ASAP7_75t_L g602 ( 
.A1(n_476),
.A2(n_583),
.B1(n_591),
.B2(n_575),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_452),
.B(n_259),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_588),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_538),
.B(n_404),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_510),
.B(n_404),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_528),
.B(n_432),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_450),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_495),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_510),
.B(n_404),
.Y(n_610)
);

NOR3x1_ASAP7_75t_L g611 ( 
.A(n_526),
.B(n_266),
.C(n_280),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_484),
.B(n_405),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_450),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_484),
.B(n_471),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_481),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_471),
.B(n_405),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_593),
.B(n_405),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_593),
.B(n_235),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_500),
.Y(n_619)
);

AND2x6_ASAP7_75t_SL g620 ( 
.A(n_470),
.B(n_238),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_476),
.B(n_451),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g622 ( 
.A(n_453),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_551),
.B(n_469),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_456),
.B(n_472),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_502),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_473),
.B(n_258),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_489),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_518),
.B(n_268),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_474),
.B(n_273),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_551),
.B(n_259),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_479),
.B(n_449),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_457),
.B(n_260),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_491),
.Y(n_633)
);

NAND2xp33_ASAP7_75t_L g634 ( 
.A(n_556),
.B(n_188),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_467),
.B(n_460),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_478),
.B(n_480),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_527),
.B(n_442),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_515),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_466),
.B(n_260),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_529),
.Y(n_640)
);

NOR3xp33_ASAP7_75t_L g641 ( 
.A(n_465),
.B(n_267),
.C(n_214),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_454),
.B(n_442),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_535),
.Y(n_643)
);

AO22x1_ASAP7_75t_L g644 ( 
.A1(n_475),
.A2(n_174),
.B1(n_298),
.B2(n_296),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_547),
.B(n_267),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_545),
.B(n_414),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_468),
.B(n_213),
.Y(n_647)
);

NAND2xp33_ASAP7_75t_SL g648 ( 
.A(n_568),
.B(n_168),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_468),
.B(n_226),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_550),
.B(n_414),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_520),
.B(n_234),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_462),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_562),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_503),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_567),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_577),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_579),
.Y(n_657)
);

OR2x6_ASAP7_75t_L g658 ( 
.A(n_483),
.B(n_230),
.Y(n_658)
);

AND2x6_ASAP7_75t_SL g659 ( 
.A(n_552),
.B(n_173),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_587),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_455),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_570),
.B(n_414),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_525),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_576),
.B(n_417),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_525),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_555),
.B(n_417),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_455),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_482),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_556),
.A2(n_173),
.B1(n_174),
.B2(n_245),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_555),
.B(n_417),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_461),
.B(n_431),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_461),
.B(n_431),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_464),
.B(n_431),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_581),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_464),
.B(n_444),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_540),
.B(n_444),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_541),
.B(n_239),
.Y(n_677)
);

AND2x4_ASAP7_75t_SL g678 ( 
.A(n_523),
.B(n_445),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_486),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_544),
.B(n_272),
.Y(n_680)
);

INVxp67_ASAP7_75t_L g681 ( 
.A(n_549),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_522),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_539),
.B(n_196),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_546),
.B(n_286),
.Y(n_684)
);

NAND2xp33_ASAP7_75t_L g685 ( 
.A(n_561),
.B(n_201),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_561),
.B(n_202),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_486),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_505),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_565),
.B(n_288),
.Y(n_689)
);

INVx8_ASAP7_75t_L g690 ( 
.A(n_552),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_580),
.B(n_289),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_574),
.B(n_207),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_496),
.B(n_498),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_574),
.B(n_208),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_501),
.B(n_559),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_458),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_582),
.B(n_210),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_554),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_505),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_531),
.B(n_215),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_485),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_582),
.B(n_530),
.Y(n_702)
);

A2O1A1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_504),
.A2(n_217),
.B(n_220),
.C(n_224),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_516),
.B(n_291),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_548),
.B(n_298),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_530),
.B(n_233),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_506),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_548),
.B(n_296),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_506),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_552),
.B(n_563),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_487),
.B(n_295),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_518),
.B(n_532),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_526),
.B(n_295),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_578),
.Y(n_714)
);

BUFx5_ASAP7_75t_L g715 ( 
.A(n_509),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_532),
.B(n_236),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_533),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_533),
.B(n_293),
.Y(n_718)
);

INVxp67_ASAP7_75t_L g719 ( 
.A(n_507),
.Y(n_719)
);

OR2x6_ASAP7_75t_L g720 ( 
.A(n_507),
.B(n_14),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_459),
.B(n_511),
.Y(n_721)
);

A2O1A1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_514),
.A2(n_517),
.B(n_536),
.C(n_542),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_514),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_571),
.B(n_293),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_573),
.B(n_269),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_584),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_459),
.B(n_287),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_584),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_485),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_477),
.B(n_283),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_517),
.B(n_256),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_592),
.B(n_256),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_508),
.Y(n_733)
);

INVx2_ASAP7_75t_SL g734 ( 
.A(n_542),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_477),
.B(n_281),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_543),
.A2(n_270),
.B(n_269),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_463),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_477),
.A2(n_488),
.B1(n_497),
.B2(n_509),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_572),
.Y(n_739)
);

NAND2x1_ASAP7_75t_L g740 ( 
.A(n_592),
.B(n_71),
.Y(n_740)
);

OR2x6_ASAP7_75t_L g741 ( 
.A(n_572),
.B(n_16),
.Y(n_741)
);

NAND2x1_ASAP7_75t_L g742 ( 
.A(n_590),
.B(n_72),
.Y(n_742)
);

NAND2xp33_ASAP7_75t_L g743 ( 
.A(n_477),
.B(n_271),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_537),
.Y(n_744)
);

INVxp67_ASAP7_75t_L g745 ( 
.A(n_509),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_553),
.A2(n_569),
.B1(n_589),
.B2(n_586),
.Y(n_746)
);

AND2x6_ASAP7_75t_L g747 ( 
.A(n_459),
.B(n_66),
.Y(n_747)
);

NOR3xp33_ASAP7_75t_L g748 ( 
.A(n_492),
.B(n_271),
.C(n_270),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_488),
.B(n_250),
.Y(n_749)
);

AO221x1_ASAP7_75t_L g750 ( 
.A1(n_485),
.A2(n_250),
.B1(n_247),
.B2(n_245),
.C(n_24),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_557),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_488),
.B(n_247),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_488),
.B(n_62),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_497),
.B(n_54),
.Y(n_754)
);

NAND3xp33_ASAP7_75t_L g755 ( 
.A(n_600),
.B(n_597),
.C(n_689),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_615),
.Y(n_756)
);

OR2x2_ASAP7_75t_L g757 ( 
.A(n_594),
.B(n_20),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_712),
.A2(n_543),
.B(n_590),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_627),
.Y(n_759)
);

A2O1A1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_600),
.A2(n_585),
.B(n_566),
.C(n_558),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_633),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_661),
.B(n_497),
.Y(n_762)
);

AO21x1_ASAP7_75t_L g763 ( 
.A1(n_618),
.A2(n_497),
.B(n_509),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_667),
.B(n_497),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_712),
.A2(n_560),
.B(n_534),
.Y(n_765)
);

NAND2x1p5_ASAP7_75t_L g766 ( 
.A(n_742),
.B(n_490),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_719),
.B(n_512),
.Y(n_767)
);

O2A1O1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_614),
.A2(n_509),
.B(n_512),
.C(n_26),
.Y(n_768)
);

OR2x6_ASAP7_75t_L g769 ( 
.A(n_690),
.B(n_490),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_638),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_656),
.Y(n_771)
);

BUFx4f_ASAP7_75t_L g772 ( 
.A(n_690),
.Y(n_772)
);

BUFx6f_ASAP7_75t_SL g773 ( 
.A(n_652),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_606),
.B(n_512),
.Y(n_774)
);

AO32x1_ASAP7_75t_L g775 ( 
.A1(n_746),
.A2(n_734),
.A3(n_657),
.B1(n_714),
.B2(n_640),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_636),
.A2(n_512),
.B(n_564),
.Y(n_776)
);

OAI21xp5_ASAP7_75t_L g777 ( 
.A1(n_723),
.A2(n_564),
.B(n_77),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_665),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_602),
.B(n_564),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_597),
.B(n_21),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_637),
.B(n_21),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_612),
.A2(n_564),
.B(n_90),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_605),
.A2(n_564),
.B(n_93),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_642),
.B(n_22),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_635),
.Y(n_785)
);

INVx11_ASAP7_75t_L g786 ( 
.A(n_747),
.Y(n_786)
);

INVx3_ASAP7_75t_L g787 ( 
.A(n_696),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_610),
.B(n_22),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_598),
.B(n_30),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_607),
.B(n_31),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_599),
.B(n_31),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_622),
.B(n_32),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_617),
.A2(n_702),
.B(n_624),
.Y(n_793)
);

OAI21xp5_ASAP7_75t_L g794 ( 
.A1(n_722),
.A2(n_96),
.B(n_139),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_665),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_595),
.A2(n_51),
.B(n_131),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_643),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_601),
.A2(n_49),
.B(n_119),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_653),
.Y(n_799)
);

O2A1O1Ixp33_ASAP7_75t_L g800 ( 
.A1(n_616),
.A2(n_33),
.B(n_40),
.C(n_41),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_647),
.B(n_40),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_647),
.B(n_41),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_701),
.Y(n_803)
);

OAI21xp5_ASAP7_75t_L g804 ( 
.A1(n_679),
.A2(n_106),
.B(n_111),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_655),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_660),
.Y(n_806)
);

AOI21x1_ASAP7_75t_L g807 ( 
.A1(n_629),
.A2(n_147),
.B(n_43),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_622),
.B(n_43),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_609),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_649),
.B(n_46),
.Y(n_810)
);

OAI21x1_ASAP7_75t_L g811 ( 
.A1(n_739),
.A2(n_744),
.B(n_733),
.Y(n_811)
);

OAI22xp5_ASAP7_75t_L g812 ( 
.A1(n_669),
.A2(n_689),
.B1(n_691),
.B2(n_720),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_602),
.B(n_631),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_646),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_631),
.B(n_596),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_687),
.A2(n_699),
.B(n_709),
.Y(n_816)
);

INVxp67_ASAP7_75t_L g817 ( 
.A(n_632),
.Y(n_817)
);

CKINVDCx10_ASAP7_75t_R g818 ( 
.A(n_737),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_SL g819 ( 
.A(n_747),
.B(n_690),
.Y(n_819)
);

NOR2x1_ASAP7_75t_L g820 ( 
.A(n_721),
.B(n_682),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_663),
.B(n_608),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_671),
.A2(n_673),
.B(n_672),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_695),
.B(n_649),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_688),
.A2(n_707),
.B(n_717),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_650),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_613),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_621),
.A2(n_670),
.B(n_666),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_L g828 ( 
.A1(n_669),
.A2(n_691),
.B1(n_720),
.B2(n_681),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_675),
.B(n_731),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_731),
.B(n_662),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_604),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_676),
.Y(n_832)
);

NOR2x1_ASAP7_75t_L g833 ( 
.A(n_623),
.B(n_700),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_664),
.B(n_718),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_718),
.B(n_732),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_701),
.Y(n_836)
);

NOR2x1_ASAP7_75t_L g837 ( 
.A(n_693),
.B(n_695),
.Y(n_837)
);

BUFx2_ASAP7_75t_L g838 ( 
.A(n_668),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_732),
.B(n_724),
.Y(n_839)
);

AOI21x1_ASAP7_75t_L g840 ( 
.A1(n_628),
.A2(n_716),
.B(n_727),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_619),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_729),
.A2(n_727),
.B(n_728),
.Y(n_842)
);

AND2x6_ASAP7_75t_L g843 ( 
.A(n_738),
.B(n_710),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_625),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_628),
.B(n_681),
.Y(n_845)
);

O2A1O1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_603),
.A2(n_683),
.B(n_685),
.C(n_634),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_645),
.B(n_704),
.Y(n_847)
);

NOR2x1p5_ASAP7_75t_SL g848 ( 
.A(n_715),
.B(n_751),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_729),
.Y(n_849)
);

OAI21xp33_ASAP7_75t_L g850 ( 
.A1(n_704),
.A2(n_680),
.B(n_651),
.Y(n_850)
);

BUFx4f_ASAP7_75t_L g851 ( 
.A(n_678),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_710),
.A2(n_680),
.B1(n_651),
.B2(n_684),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_724),
.B(n_725),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_725),
.B(n_677),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_729),
.A2(n_698),
.B(n_726),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_741),
.Y(n_856)
);

INVx4_ASAP7_75t_L g857 ( 
.A(n_747),
.Y(n_857)
);

INVx1_ASAP7_75t_SL g858 ( 
.A(n_648),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_654),
.Y(n_859)
);

OR2x2_ASAP7_75t_L g860 ( 
.A(n_713),
.B(n_708),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_730),
.A2(n_735),
.B(n_703),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_745),
.A2(n_694),
.B(n_692),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_720),
.Y(n_863)
);

AOI21x1_ASAP7_75t_L g864 ( 
.A1(n_706),
.A2(n_749),
.B(n_752),
.Y(n_864)
);

OAI21xp5_ASAP7_75t_L g865 ( 
.A1(n_745),
.A2(n_697),
.B(n_686),
.Y(n_865)
);

CKINVDCx10_ASAP7_75t_R g866 ( 
.A(n_658),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_677),
.B(n_684),
.Y(n_867)
);

O2A1O1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_743),
.A2(n_741),
.B(n_711),
.C(n_641),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_632),
.B(n_639),
.Y(n_869)
);

AO22x1_ASAP7_75t_L g870 ( 
.A1(n_611),
.A2(n_641),
.B1(n_748),
.B2(n_711),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_753),
.A2(n_754),
.B(n_740),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_705),
.B(n_639),
.Y(n_872)
);

INVx4_ASAP7_75t_L g873 ( 
.A(n_747),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_741),
.A2(n_658),
.B1(n_630),
.B2(n_736),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_658),
.A2(n_715),
.B(n_644),
.Y(n_875)
);

AO21x1_ASAP7_75t_L g876 ( 
.A1(n_748),
.A2(n_750),
.B(n_620),
.Y(n_876)
);

NAND2xp33_ASAP7_75t_L g877 ( 
.A(n_715),
.B(n_659),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_715),
.B(n_674),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_712),
.A2(n_719),
.B(n_636),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_712),
.A2(n_719),
.B(n_636),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_615),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_661),
.B(n_667),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_615),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_661),
.B(n_667),
.Y(n_884)
);

BUFx2_ASAP7_75t_L g885 ( 
.A(n_594),
.Y(n_885)
);

AND3x2_ASAP7_75t_L g886 ( 
.A(n_600),
.B(n_691),
.C(n_689),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_L g887 ( 
.A1(n_702),
.A2(n_471),
.B1(n_476),
.B2(n_614),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_674),
.B(n_602),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_674),
.B(n_600),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_712),
.A2(n_719),
.B(n_636),
.Y(n_890)
);

NOR2x1_ASAP7_75t_L g891 ( 
.A(n_721),
.B(n_496),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_615),
.Y(n_892)
);

CKINVDCx10_ASAP7_75t_R g893 ( 
.A(n_652),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_712),
.A2(n_719),
.B(n_636),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_661),
.B(n_667),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_637),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_615),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_615),
.Y(n_898)
);

OAI22xp5_ASAP7_75t_L g899 ( 
.A1(n_702),
.A2(n_471),
.B1(n_476),
.B2(n_614),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_712),
.A2(n_719),
.B(n_636),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_712),
.A2(n_719),
.B(n_636),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_719),
.B(n_712),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_594),
.Y(n_903)
);

O2A1O1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_614),
.A2(n_521),
.B(n_616),
.C(n_600),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_719),
.B(n_712),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_719),
.B(n_712),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_712),
.A2(n_719),
.B(n_636),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_674),
.B(n_600),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_661),
.B(n_667),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_615),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_615),
.Y(n_911)
);

AND2x2_ASAP7_75t_SL g912 ( 
.A(n_600),
.B(n_454),
.Y(n_912)
);

NAND3xp33_ASAP7_75t_L g913 ( 
.A(n_600),
.B(n_597),
.C(n_689),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_682),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_627),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_661),
.B(n_667),
.Y(n_916)
);

AOI22xp5_ASAP7_75t_L g917 ( 
.A1(n_600),
.A2(n_631),
.B1(n_521),
.B2(n_452),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_615),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_729),
.Y(n_919)
);

AO21x1_ASAP7_75t_L g920 ( 
.A1(n_618),
.A2(n_476),
.B(n_600),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_615),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_729),
.Y(n_922)
);

AOI21x1_ASAP7_75t_L g923 ( 
.A1(n_624),
.A2(n_629),
.B(n_626),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_696),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_594),
.B(n_519),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_729),
.Y(n_926)
);

O2A1O1Ixp5_ASAP7_75t_L g927 ( 
.A1(n_600),
.A2(n_628),
.B(n_618),
.C(n_716),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_661),
.B(n_667),
.Y(n_928)
);

NOR2xp67_ASAP7_75t_L g929 ( 
.A(n_674),
.B(n_522),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_661),
.B(n_667),
.Y(n_930)
);

NAND2x1p5_ASAP7_75t_L g931 ( 
.A(n_742),
.B(n_740),
.Y(n_931)
);

CKINVDCx16_ASAP7_75t_R g932 ( 
.A(n_682),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_674),
.B(n_600),
.Y(n_933)
);

NAND3xp33_ASAP7_75t_L g934 ( 
.A(n_755),
.B(n_913),
.C(n_852),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_879),
.A2(n_890),
.B(n_880),
.Y(n_935)
);

A2O1A1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_850),
.A2(n_867),
.B(n_854),
.C(n_853),
.Y(n_936)
);

AO21x1_ASAP7_75t_L g937 ( 
.A1(n_835),
.A2(n_853),
.B(n_839),
.Y(n_937)
);

BUFx8_ASAP7_75t_L g938 ( 
.A(n_773),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_902),
.B(n_905),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_812),
.A2(n_917),
.B1(n_902),
.B2(n_906),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_849),
.Y(n_941)
);

OAI21x1_ASAP7_75t_L g942 ( 
.A1(n_864),
.A2(n_855),
.B(n_758),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_793),
.A2(n_900),
.B(n_894),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_905),
.B(n_906),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_901),
.A2(n_907),
.B(n_822),
.Y(n_945)
);

AOI21x1_ASAP7_75t_SL g946 ( 
.A1(n_801),
.A2(n_810),
.B(n_802),
.Y(n_946)
);

OA21x2_ASAP7_75t_L g947 ( 
.A1(n_794),
.A2(n_816),
.B(n_760),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_820),
.B(n_821),
.Y(n_948)
);

NAND2xp33_ASAP7_75t_L g949 ( 
.A(n_812),
.B(n_869),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_889),
.B(n_908),
.Y(n_950)
);

OAI21x1_ASAP7_75t_L g951 ( 
.A1(n_840),
.A2(n_923),
.B(n_931),
.Y(n_951)
);

AO21x1_ASAP7_75t_L g952 ( 
.A1(n_813),
.A2(n_823),
.B(n_887),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_756),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_834),
.B(n_829),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_821),
.B(n_785),
.Y(n_955)
);

OR2x6_ASAP7_75t_L g956 ( 
.A(n_859),
.B(n_857),
.Y(n_956)
);

AOI21x1_ASAP7_75t_L g957 ( 
.A1(n_827),
.A2(n_779),
.B(n_774),
.Y(n_957)
);

OAI21x1_ASAP7_75t_L g958 ( 
.A1(n_862),
.A2(n_765),
.B(n_865),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_824),
.A2(n_830),
.B(n_816),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_846),
.A2(n_884),
.B(n_882),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_933),
.B(n_895),
.Y(n_961)
);

AO31x2_ASAP7_75t_L g962 ( 
.A1(n_920),
.A2(n_887),
.A3(n_899),
.B(n_763),
.Y(n_962)
);

INVx2_ASAP7_75t_SL g963 ( 
.A(n_838),
.Y(n_963)
);

OAI21xp5_ASAP7_75t_L g964 ( 
.A1(n_899),
.A2(n_904),
.B(n_927),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_914),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_925),
.B(n_863),
.Y(n_966)
);

OAI21xp5_ASAP7_75t_L g967 ( 
.A1(n_794),
.A2(n_828),
.B(n_845),
.Y(n_967)
);

A2O1A1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_847),
.A2(n_815),
.B(n_780),
.C(n_828),
.Y(n_968)
);

INVxp67_ASAP7_75t_L g969 ( 
.A(n_831),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_909),
.B(n_916),
.Y(n_970)
);

AOI21x1_ASAP7_75t_L g971 ( 
.A1(n_767),
.A2(n_764),
.B(n_762),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_817),
.B(n_886),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_814),
.B(n_825),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_826),
.B(n_770),
.Y(n_974)
);

INVxp67_ASAP7_75t_L g975 ( 
.A(n_885),
.Y(n_975)
);

OAI21x1_ASAP7_75t_L g976 ( 
.A1(n_766),
.A2(n_776),
.B(n_803),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_896),
.B(n_903),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_928),
.B(n_930),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_778),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_868),
.A2(n_845),
.B(n_832),
.C(n_833),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_843),
.B(n_888),
.Y(n_981)
);

INVx4_ASAP7_75t_L g982 ( 
.A(n_849),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_912),
.B(n_929),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_837),
.A2(n_875),
.B(n_872),
.C(n_804),
.Y(n_984)
);

INVx5_ASAP7_75t_L g985 ( 
.A(n_857),
.Y(n_985)
);

OA21x2_ASAP7_75t_L g986 ( 
.A1(n_777),
.A2(n_788),
.B(n_789),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_860),
.B(n_795),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_893),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_771),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_791),
.A2(n_768),
.B(n_878),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_790),
.A2(n_843),
.B(n_757),
.Y(n_991)
);

OAI21x1_ASAP7_75t_L g992 ( 
.A1(n_787),
.A2(n_924),
.B(n_836),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_781),
.B(n_897),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_856),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_873),
.A2(n_819),
.B(n_891),
.Y(n_995)
);

INVx1_ASAP7_75t_SL g996 ( 
.A(n_818),
.Y(n_996)
);

OAI211xp5_ASAP7_75t_L g997 ( 
.A1(n_792),
.A2(n_808),
.B(n_784),
.C(n_858),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_843),
.B(n_881),
.Y(n_998)
);

OAI21x1_ASAP7_75t_L g999 ( 
.A1(n_798),
.A2(n_783),
.B(n_782),
.Y(n_999)
);

OAI21x1_ASAP7_75t_L g1000 ( 
.A1(n_796),
.A2(n_807),
.B(n_841),
.Y(n_1000)
);

AOI21x1_ASAP7_75t_L g1001 ( 
.A1(n_874),
.A2(n_911),
.B(n_910),
.Y(n_1001)
);

AO21x2_ASAP7_75t_L g1002 ( 
.A1(n_775),
.A2(n_898),
.B(n_892),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_919),
.A2(n_922),
.B(n_926),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_843),
.B(n_883),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_858),
.B(n_932),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_870),
.B(n_876),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_851),
.Y(n_1007)
);

AO31x2_ASAP7_75t_L g1008 ( 
.A1(n_775),
.A2(n_918),
.A3(n_921),
.B(n_761),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_851),
.B(n_759),
.Y(n_1009)
);

NAND2x1p5_ASAP7_75t_L g1010 ( 
.A(n_919),
.B(n_926),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_844),
.Y(n_1011)
);

NAND3xp33_ASAP7_75t_SL g1012 ( 
.A(n_800),
.B(n_805),
.C(n_806),
.Y(n_1012)
);

AO21x1_ASAP7_75t_L g1013 ( 
.A1(n_877),
.A2(n_775),
.B(n_915),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_797),
.B(n_799),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_919),
.A2(n_922),
.B(n_769),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_922),
.B(n_848),
.Y(n_1016)
);

OAI22x1_ASAP7_75t_L g1017 ( 
.A1(n_866),
.A2(n_772),
.B1(n_773),
.B2(n_786),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_769),
.A2(n_880),
.B(n_879),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_769),
.A2(n_880),
.B(n_879),
.Y(n_1019)
);

OAI21x1_ASAP7_75t_SL g1020 ( 
.A1(n_794),
.A2(n_816),
.B(n_804),
.Y(n_1020)
);

AO31x2_ASAP7_75t_L g1021 ( 
.A1(n_920),
.A2(n_899),
.A3(n_887),
.B(n_760),
.Y(n_1021)
);

AO31x2_ASAP7_75t_L g1022 ( 
.A1(n_920),
.A2(n_899),
.A3(n_887),
.B(n_760),
.Y(n_1022)
);

OR2x2_ASAP7_75t_L g1023 ( 
.A(n_860),
.B(n_737),
.Y(n_1023)
);

AOI21x1_ASAP7_75t_L g1024 ( 
.A1(n_861),
.A2(n_864),
.B(n_923),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_879),
.A2(n_890),
.B(n_880),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_879),
.A2(n_890),
.B(n_880),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_902),
.B(n_905),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_902),
.B(n_905),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_879),
.A2(n_890),
.B(n_880),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_914),
.Y(n_1030)
);

AOI211x1_ASAP7_75t_L g1031 ( 
.A1(n_755),
.A2(n_913),
.B(n_812),
.C(n_850),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_902),
.B(n_905),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_914),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_809),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_879),
.A2(n_890),
.B(n_880),
.Y(n_1035)
);

AO31x2_ASAP7_75t_L g1036 ( 
.A1(n_920),
.A2(n_899),
.A3(n_887),
.B(n_760),
.Y(n_1036)
);

AOI21x1_ASAP7_75t_SL g1037 ( 
.A1(n_867),
.A2(n_802),
.B(n_801),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_755),
.A2(n_913),
.B(n_850),
.C(n_867),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_902),
.B(n_905),
.Y(n_1039)
);

OAI21x1_ASAP7_75t_L g1040 ( 
.A1(n_811),
.A2(n_842),
.B(n_871),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_812),
.A2(n_913),
.B1(n_755),
.B2(n_852),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_879),
.A2(n_890),
.B(n_880),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_793),
.A2(n_880),
.B(n_879),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_879),
.A2(n_890),
.B(n_880),
.Y(n_1044)
);

AO31x2_ASAP7_75t_L g1045 ( 
.A1(n_920),
.A2(n_899),
.A3(n_887),
.B(n_760),
.Y(n_1045)
);

NAND2x1p5_ASAP7_75t_L g1046 ( 
.A(n_857),
.B(n_873),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_811),
.A2(n_842),
.B(n_871),
.Y(n_1047)
);

OAI21x1_ASAP7_75t_L g1048 ( 
.A1(n_811),
.A2(n_842),
.B(n_871),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_811),
.A2(n_842),
.B(n_871),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_793),
.A2(n_880),
.B(n_879),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_885),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_793),
.A2(n_880),
.B(n_879),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_812),
.A2(n_913),
.B1(n_755),
.B2(n_852),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_811),
.A2(n_842),
.B(n_871),
.Y(n_1054)
);

AOI221xp5_ASAP7_75t_SL g1055 ( 
.A1(n_812),
.A2(n_828),
.B1(n_850),
.B2(n_904),
.C(n_899),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_879),
.A2(n_890),
.B(n_880),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_852),
.B(n_755),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_L g1058 ( 
.A1(n_811),
.A2(n_842),
.B(n_871),
.Y(n_1058)
);

AND2x2_ASAP7_75t_SL g1059 ( 
.A(n_912),
.B(n_867),
.Y(n_1059)
);

AO31x2_ASAP7_75t_L g1060 ( 
.A1(n_920),
.A2(n_899),
.A3(n_887),
.B(n_760),
.Y(n_1060)
);

AOI21xp33_ASAP7_75t_L g1061 ( 
.A1(n_755),
.A2(n_913),
.B(n_812),
.Y(n_1061)
);

AOI21xp33_ASAP7_75t_L g1062 ( 
.A1(n_755),
.A2(n_913),
.B(n_812),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_755),
.A2(n_913),
.B(n_850),
.C(n_867),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_879),
.A2(n_890),
.B(n_880),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_756),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_811),
.A2(n_842),
.B(n_871),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_820),
.B(n_821),
.Y(n_1067)
);

OR2x2_ASAP7_75t_L g1068 ( 
.A(n_860),
.B(n_737),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_1007),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_954),
.B(n_939),
.Y(n_1070)
);

OAI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_968),
.A2(n_967),
.B(n_1041),
.Y(n_1071)
);

OR2x6_ASAP7_75t_SL g1072 ( 
.A(n_965),
.B(n_1033),
.Y(n_1072)
);

O2A1O1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_1041),
.A2(n_1053),
.B(n_949),
.C(n_1061),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_1061),
.A2(n_1062),
.B(n_967),
.C(n_934),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_989),
.Y(n_1075)
);

INVx3_ASAP7_75t_L g1076 ( 
.A(n_985),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_1053),
.A2(n_1057),
.B1(n_934),
.B2(n_1059),
.Y(n_1077)
);

BUFx12f_ASAP7_75t_L g1078 ( 
.A(n_938),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_985),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_963),
.Y(n_1080)
);

NAND2x1p5_ASAP7_75t_L g1081 ( 
.A(n_985),
.B(n_982),
.Y(n_1081)
);

NAND2x1p5_ASAP7_75t_L g1082 ( 
.A(n_985),
.B(n_982),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_966),
.B(n_948),
.Y(n_1083)
);

AOI22xp33_ASAP7_75t_L g1084 ( 
.A1(n_1062),
.A2(n_1006),
.B1(n_940),
.B2(n_952),
.Y(n_1084)
);

INVx1_ASAP7_75t_SL g1085 ( 
.A(n_1023),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_977),
.B(n_1005),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_R g1087 ( 
.A(n_1030),
.B(n_988),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_938),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_950),
.B(n_961),
.Y(n_1089)
);

OAI21xp33_ASAP7_75t_L g1090 ( 
.A1(n_993),
.A2(n_978),
.B(n_970),
.Y(n_1090)
);

BUFx3_ASAP7_75t_L g1091 ( 
.A(n_979),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1025),
.A2(n_1026),
.B(n_1056),
.Y(n_1092)
);

AND2x4_ASAP7_75t_L g1093 ( 
.A(n_966),
.B(n_948),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1065),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_954),
.B(n_973),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_1067),
.B(n_1009),
.Y(n_1096)
);

BUFx2_ASAP7_75t_L g1097 ( 
.A(n_1051),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1029),
.A2(n_1044),
.B(n_1064),
.Y(n_1098)
);

INVx2_ASAP7_75t_SL g1099 ( 
.A(n_994),
.Y(n_1099)
);

BUFx4_ASAP7_75t_SL g1100 ( 
.A(n_1068),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_987),
.B(n_975),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1035),
.A2(n_1042),
.B(n_943),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1014),
.Y(n_1103)
);

BUFx3_ASAP7_75t_L g1104 ( 
.A(n_1017),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_956),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_SL g1106 ( 
.A(n_940),
.B(n_1020),
.Y(n_1106)
);

NOR3xp33_ASAP7_75t_L g1107 ( 
.A(n_997),
.B(n_983),
.C(n_1063),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_955),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1011),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_943),
.A2(n_1043),
.B(n_1050),
.Y(n_1110)
);

OR2x6_ASAP7_75t_L g1111 ( 
.A(n_956),
.B(n_1046),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_1067),
.B(n_974),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_978),
.B(n_944),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1043),
.A2(n_1052),
.B(n_1050),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1034),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_939),
.A2(n_1039),
.B1(n_1028),
.B2(n_1027),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_974),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_955),
.B(n_956),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1032),
.B(n_1027),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_969),
.B(n_972),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1052),
.A2(n_959),
.B(n_1018),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_1028),
.B(n_1039),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_998),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_936),
.B(n_1038),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_980),
.A2(n_984),
.B(n_991),
.C(n_998),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_981),
.B(n_1004),
.Y(n_1126)
);

O2A1O1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_991),
.A2(n_1004),
.B(n_981),
.C(n_964),
.Y(n_1127)
);

AOI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_1012),
.A2(n_937),
.B1(n_964),
.B2(n_990),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_996),
.Y(n_1129)
);

BUFx8_ASAP7_75t_SL g1130 ( 
.A(n_941),
.Y(n_1130)
);

BUFx2_ASAP7_75t_L g1131 ( 
.A(n_941),
.Y(n_1131)
);

OR2x6_ASAP7_75t_L g1132 ( 
.A(n_1046),
.B(n_1015),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_990),
.A2(n_1019),
.B(n_1013),
.C(n_995),
.Y(n_1133)
);

INVx1_ASAP7_75t_SL g1134 ( 
.A(n_1002),
.Y(n_1134)
);

AO21x2_ASAP7_75t_L g1135 ( 
.A1(n_1024),
.A2(n_958),
.B(n_951),
.Y(n_1135)
);

HB1xp67_ASAP7_75t_L g1136 ( 
.A(n_1010),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_1010),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_1016),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1031),
.B(n_1055),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1008),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_1016),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1008),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1055),
.B(n_986),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_996),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1008),
.B(n_947),
.Y(n_1145)
);

INVx3_ASAP7_75t_L g1146 ( 
.A(n_992),
.Y(n_1146)
);

AOI21xp33_ASAP7_75t_SL g1147 ( 
.A1(n_1000),
.A2(n_976),
.B(n_942),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_1003),
.B(n_957),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_962),
.B(n_1060),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_971),
.Y(n_1150)
);

OAI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_946),
.A2(n_1037),
.B1(n_1060),
.B2(n_1021),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_999),
.A2(n_1047),
.B(n_1058),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_1040),
.B(n_1048),
.Y(n_1153)
);

INVx8_ASAP7_75t_L g1154 ( 
.A(n_1021),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1022),
.B(n_1036),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1022),
.B(n_1036),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1049),
.A2(n_1054),
.B(n_1066),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_962),
.B(n_1060),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_SL g1159 ( 
.A1(n_1045),
.A2(n_1022),
.B(n_962),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1045),
.B(n_950),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1045),
.B(n_950),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_954),
.B(n_939),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_950),
.B(n_961),
.Y(n_1163)
);

A2O1A1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_968),
.A2(n_850),
.B(n_913),
.C(n_755),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_966),
.B(n_948),
.Y(n_1165)
);

BUFx3_ASAP7_75t_L g1166 ( 
.A(n_1030),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_953),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_1007),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_1007),
.Y(n_1169)
);

INVx5_ASAP7_75t_L g1170 ( 
.A(n_956),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_968),
.A2(n_850),
.B(n_913),
.C(n_755),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_953),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_966),
.B(n_948),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_953),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_945),
.A2(n_960),
.B(n_935),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_977),
.B(n_594),
.Y(n_1176)
);

NAND3xp33_ASAP7_75t_L g1177 ( 
.A(n_968),
.B(n_913),
.C(n_755),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_966),
.B(n_948),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_966),
.B(n_948),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_953),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_954),
.B(n_939),
.Y(n_1181)
);

BUFx2_ASAP7_75t_L g1182 ( 
.A(n_963),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_977),
.B(n_594),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_977),
.B(n_594),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_954),
.B(n_939),
.Y(n_1185)
);

INVxp67_ASAP7_75t_SL g1186 ( 
.A(n_978),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_954),
.B(n_939),
.Y(n_1187)
);

INVx3_ASAP7_75t_SL g1188 ( 
.A(n_965),
.Y(n_1188)
);

OA21x2_ASAP7_75t_L g1189 ( 
.A1(n_964),
.A2(n_1043),
.B(n_943),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_945),
.A2(n_960),
.B(n_935),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_968),
.A2(n_755),
.B1(n_913),
.B2(n_812),
.Y(n_1191)
);

NOR2x1_ASAP7_75t_SL g1192 ( 
.A(n_985),
.B(n_956),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_963),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_965),
.Y(n_1194)
);

INVx1_ASAP7_75t_SL g1195 ( 
.A(n_1023),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_953),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_968),
.A2(n_755),
.B1(n_913),
.B2(n_812),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1094),
.Y(n_1198)
);

AO21x1_ASAP7_75t_L g1199 ( 
.A1(n_1191),
.A2(n_1197),
.B(n_1073),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_1130),
.Y(n_1200)
);

INVx6_ASAP7_75t_L g1201 ( 
.A(n_1069),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1075),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_SL g1203 ( 
.A1(n_1192),
.A2(n_1077),
.B(n_1127),
.Y(n_1203)
);

AOI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1191),
.A2(n_1197),
.B1(n_1107),
.B2(n_1177),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1167),
.Y(n_1205)
);

NAND2x1p5_ASAP7_75t_L g1206 ( 
.A(n_1170),
.B(n_1076),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1172),
.Y(n_1207)
);

AO21x1_ASAP7_75t_L g1208 ( 
.A1(n_1071),
.A2(n_1106),
.B(n_1151),
.Y(n_1208)
);

NAND2x1p5_ASAP7_75t_L g1209 ( 
.A(n_1170),
.B(n_1079),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1174),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1180),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1196),
.Y(n_1212)
);

INVx6_ASAP7_75t_L g1213 ( 
.A(n_1069),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1095),
.A2(n_1113),
.B1(n_1186),
.B2(n_1119),
.Y(n_1214)
);

BUFx12f_ASAP7_75t_L g1215 ( 
.A(n_1078),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1071),
.A2(n_1177),
.B1(n_1084),
.B2(n_1106),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_1085),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_SL g1218 ( 
.A1(n_1089),
.A2(n_1163),
.B1(n_1096),
.B2(n_1104),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1090),
.A2(n_1124),
.B1(n_1128),
.B2(n_1122),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1109),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_1112),
.Y(n_1221)
);

OAI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1070),
.A2(n_1185),
.B1(n_1162),
.B2(n_1181),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1157),
.A2(n_1152),
.B(n_1175),
.Y(n_1223)
);

AO21x2_ASAP7_75t_L g1224 ( 
.A1(n_1147),
.A2(n_1152),
.B(n_1121),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1150),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1150),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1103),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1115),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1070),
.B(n_1162),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1123),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1124),
.A2(n_1116),
.B1(n_1181),
.B2(n_1187),
.Y(n_1231)
);

BUFx4_ASAP7_75t_R g1232 ( 
.A(n_1166),
.Y(n_1232)
);

INVx3_ASAP7_75t_L g1233 ( 
.A(n_1111),
.Y(n_1233)
);

AO21x2_ASAP7_75t_L g1234 ( 
.A1(n_1110),
.A2(n_1114),
.B(n_1190),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1117),
.Y(n_1235)
);

AO21x2_ASAP7_75t_L g1236 ( 
.A1(n_1092),
.A2(n_1098),
.B(n_1102),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1138),
.Y(n_1237)
);

NAND3xp33_ASAP7_75t_L g1238 ( 
.A(n_1164),
.B(n_1171),
.C(n_1074),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1116),
.A2(n_1185),
.B1(n_1187),
.B2(n_1126),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1189),
.A2(n_1195),
.B1(n_1085),
.B2(n_1139),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1138),
.Y(n_1241)
);

OAI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1195),
.A2(n_1091),
.B1(n_1108),
.B2(n_1188),
.Y(n_1242)
);

INVx11_ASAP7_75t_L g1243 ( 
.A(n_1100),
.Y(n_1243)
);

OR2x2_ASAP7_75t_L g1244 ( 
.A(n_1086),
.B(n_1097),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1101),
.A2(n_1139),
.B1(n_1099),
.B2(n_1120),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1176),
.B(n_1183),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1149),
.B(n_1161),
.Y(n_1247)
);

OR2x6_ASAP7_75t_L g1248 ( 
.A(n_1125),
.B(n_1132),
.Y(n_1248)
);

OR2x6_ASAP7_75t_L g1249 ( 
.A(n_1132),
.B(n_1111),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1133),
.A2(n_1146),
.B(n_1151),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1184),
.B(n_1096),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1138),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_1168),
.Y(n_1253)
);

INVx2_ASAP7_75t_SL g1254 ( 
.A(n_1118),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_1087),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1141),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1141),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1141),
.Y(n_1258)
);

INVxp67_ASAP7_75t_L g1259 ( 
.A(n_1080),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1136),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_1182),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1135),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1118),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1140),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1160),
.B(n_1158),
.Y(n_1265)
);

AND2x4_ASAP7_75t_L g1266 ( 
.A(n_1083),
.B(n_1165),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1093),
.B(n_1179),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_1193),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1142),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1131),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1137),
.Y(n_1271)
);

INVx4_ASAP7_75t_SL g1272 ( 
.A(n_1111),
.Y(n_1272)
);

CKINVDCx14_ASAP7_75t_R g1273 ( 
.A(n_1194),
.Y(n_1273)
);

CKINVDCx6p67_ASAP7_75t_R g1274 ( 
.A(n_1072),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1137),
.Y(n_1275)
);

OAI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1144),
.A2(n_1168),
.B1(n_1169),
.B2(n_1105),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1154),
.A2(n_1179),
.B1(n_1178),
.B2(n_1173),
.Y(n_1277)
);

OR2x2_ASAP7_75t_L g1278 ( 
.A(n_1093),
.B(n_1178),
.Y(n_1278)
);

BUFx2_ASAP7_75t_L g1279 ( 
.A(n_1165),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1173),
.B(n_1169),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1105),
.B(n_1132),
.Y(n_1281)
);

INVx4_ASAP7_75t_L g1282 ( 
.A(n_1169),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1145),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1154),
.A2(n_1143),
.B1(n_1156),
.B2(n_1155),
.Y(n_1284)
);

AND2x4_ASAP7_75t_L g1285 ( 
.A(n_1143),
.B(n_1153),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1134),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1129),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1081),
.A2(n_1082),
.B1(n_1159),
.B2(n_1088),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1134),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1077),
.B(n_1126),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1191),
.A2(n_755),
.B1(n_913),
.B2(n_812),
.Y(n_1291)
);

BUFx3_ASAP7_75t_L g1292 ( 
.A(n_1130),
.Y(n_1292)
);

BUFx2_ASAP7_75t_L g1293 ( 
.A(n_1091),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_SL g1294 ( 
.A1(n_1192),
.A2(n_991),
.B(n_1013),
.Y(n_1294)
);

INVx4_ASAP7_75t_L g1295 ( 
.A(n_1170),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1077),
.B(n_1126),
.Y(n_1296)
);

INVxp33_ASAP7_75t_L g1297 ( 
.A(n_1086),
.Y(n_1297)
);

AND2x4_ASAP7_75t_L g1298 ( 
.A(n_1118),
.B(n_1112),
.Y(n_1298)
);

AOI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1148),
.A2(n_1001),
.B(n_1024),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1094),
.Y(n_1300)
);

OR2x2_ASAP7_75t_L g1301 ( 
.A(n_1085),
.B(n_1195),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1094),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_1130),
.Y(n_1303)
);

HB1xp67_ASAP7_75t_L g1304 ( 
.A(n_1085),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1247),
.B(n_1265),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1264),
.Y(n_1306)
);

BUFx2_ASAP7_75t_L g1307 ( 
.A(n_1248),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1247),
.B(n_1265),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1269),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1290),
.B(n_1296),
.Y(n_1310)
);

OR2x2_ASAP7_75t_L g1311 ( 
.A(n_1285),
.B(n_1289),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1283),
.Y(n_1312)
);

AO21x1_ASAP7_75t_SL g1313 ( 
.A1(n_1216),
.A2(n_1204),
.B(n_1291),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1217),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1229),
.B(n_1214),
.Y(n_1315)
);

AND2x2_ASAP7_75t_SL g1316 ( 
.A(n_1284),
.B(n_1239),
.Y(n_1316)
);

OR2x2_ASAP7_75t_L g1317 ( 
.A(n_1285),
.B(n_1286),
.Y(n_1317)
);

BUFx2_ASAP7_75t_L g1318 ( 
.A(n_1248),
.Y(n_1318)
);

NAND2x1_ASAP7_75t_L g1319 ( 
.A(n_1248),
.B(n_1249),
.Y(n_1319)
);

OR2x2_ASAP7_75t_L g1320 ( 
.A(n_1240),
.B(n_1284),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_L g1321 ( 
.A(n_1281),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1223),
.A2(n_1250),
.B(n_1299),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1222),
.B(n_1304),
.Y(n_1323)
);

OA21x2_ASAP7_75t_L g1324 ( 
.A1(n_1208),
.A2(n_1199),
.B(n_1262),
.Y(n_1324)
);

OR2x2_ASAP7_75t_L g1325 ( 
.A(n_1245),
.B(n_1238),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1199),
.B(n_1258),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1301),
.Y(n_1327)
);

OAI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1219),
.A2(n_1231),
.B(n_1246),
.Y(n_1328)
);

AO21x2_ASAP7_75t_L g1329 ( 
.A1(n_1294),
.A2(n_1203),
.B(n_1224),
.Y(n_1329)
);

CKINVDCx20_ASAP7_75t_R g1330 ( 
.A(n_1273),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_SL g1331 ( 
.A(n_1255),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1230),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1297),
.B(n_1202),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1270),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1297),
.B(n_1205),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1249),
.B(n_1233),
.Y(n_1336)
);

OA21x2_ASAP7_75t_L g1337 ( 
.A1(n_1225),
.A2(n_1226),
.B(n_1210),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1207),
.B(n_1211),
.Y(n_1338)
);

INVxp67_ASAP7_75t_L g1339 ( 
.A(n_1244),
.Y(n_1339)
);

OR2x6_ASAP7_75t_L g1340 ( 
.A(n_1295),
.B(n_1288),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1242),
.A2(n_1279),
.B1(n_1251),
.B2(n_1274),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1260),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1212),
.B(n_1234),
.Y(n_1343)
);

HB1xp67_ASAP7_75t_L g1344 ( 
.A(n_1237),
.Y(n_1344)
);

OA21x2_ASAP7_75t_L g1345 ( 
.A1(n_1226),
.A2(n_1220),
.B(n_1302),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1241),
.B(n_1256),
.Y(n_1346)
);

INVxp33_ASAP7_75t_L g1347 ( 
.A(n_1293),
.Y(n_1347)
);

OR2x2_ASAP7_75t_L g1348 ( 
.A(n_1236),
.B(n_1218),
.Y(n_1348)
);

HB1xp67_ASAP7_75t_L g1349 ( 
.A(n_1252),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1257),
.B(n_1235),
.Y(n_1350)
);

INVx4_ASAP7_75t_L g1351 ( 
.A(n_1272),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1228),
.B(n_1198),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1227),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1300),
.Y(n_1354)
);

AO31x2_ASAP7_75t_L g1355 ( 
.A1(n_1271),
.A2(n_1275),
.A3(n_1295),
.B(n_1267),
.Y(n_1355)
);

CKINVDCx20_ASAP7_75t_R g1356 ( 
.A(n_1273),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1306),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1305),
.B(n_1277),
.Y(n_1358)
);

AO21x1_ASAP7_75t_L g1359 ( 
.A1(n_1325),
.A2(n_1276),
.B(n_1206),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1343),
.B(n_1268),
.Y(n_1360)
);

AOI211xp5_ASAP7_75t_L g1361 ( 
.A1(n_1328),
.A2(n_1259),
.B(n_1278),
.C(n_1280),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_1355),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1305),
.B(n_1277),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1308),
.B(n_1263),
.Y(n_1364)
);

INVx1_ASAP7_75t_SL g1365 ( 
.A(n_1314),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1315),
.B(n_1261),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_SL g1367 ( 
.A1(n_1316),
.A2(n_1232),
.B1(n_1298),
.B2(n_1215),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1343),
.B(n_1254),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1306),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1309),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1345),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1337),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1345),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1347),
.B(n_1287),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1345),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1317),
.B(n_1274),
.Y(n_1376)
);

NAND2x1p5_ASAP7_75t_L g1377 ( 
.A(n_1319),
.B(n_1282),
.Y(n_1377)
);

AOI33xp33_ASAP7_75t_L g1378 ( 
.A1(n_1310),
.A2(n_1266),
.A3(n_1232),
.B1(n_1243),
.B2(n_1201),
.B3(n_1213),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1355),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1326),
.B(n_1206),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1326),
.B(n_1209),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1333),
.B(n_1266),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1333),
.B(n_1266),
.Y(n_1383)
);

NAND2x1_ASAP7_75t_L g1384 ( 
.A(n_1340),
.B(n_1221),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1312),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1312),
.Y(n_1386)
);

INVxp67_ASAP7_75t_SL g1387 ( 
.A(n_1324),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1361),
.A2(n_1316),
.B(n_1325),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1365),
.B(n_1327),
.Y(n_1389)
);

NOR3xp33_ASAP7_75t_L g1390 ( 
.A(n_1361),
.B(n_1323),
.C(n_1348),
.Y(n_1390)
);

OAI21xp33_ASAP7_75t_L g1391 ( 
.A1(n_1378),
.A2(n_1320),
.B(n_1341),
.Y(n_1391)
);

NOR3xp33_ASAP7_75t_L g1392 ( 
.A(n_1367),
.B(n_1348),
.C(n_1351),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1360),
.B(n_1307),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1368),
.B(n_1318),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1366),
.B(n_1335),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_SL g1396 ( 
.A(n_1359),
.B(n_1321),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1385),
.B(n_1324),
.Y(n_1397)
);

NAND4xp25_ASAP7_75t_L g1398 ( 
.A(n_1366),
.B(n_1339),
.C(n_1320),
.D(n_1311),
.Y(n_1398)
);

NAND3xp33_ASAP7_75t_L g1399 ( 
.A(n_1376),
.B(n_1332),
.C(n_1334),
.Y(n_1399)
);

OA21x2_ASAP7_75t_L g1400 ( 
.A1(n_1387),
.A2(n_1322),
.B(n_1371),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_SL g1401 ( 
.A(n_1359),
.B(n_1321),
.Y(n_1401)
);

NAND3xp33_ASAP7_75t_L g1402 ( 
.A(n_1376),
.B(n_1342),
.C(n_1353),
.Y(n_1402)
);

NAND3xp33_ASAP7_75t_L g1403 ( 
.A(n_1374),
.B(n_1344),
.C(n_1349),
.Y(n_1403)
);

NAND3xp33_ASAP7_75t_L g1404 ( 
.A(n_1379),
.B(n_1354),
.C(n_1350),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1382),
.B(n_1383),
.Y(n_1405)
);

NAND3xp33_ASAP7_75t_L g1406 ( 
.A(n_1379),
.B(n_1354),
.C(n_1350),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1357),
.Y(n_1407)
);

NAND3xp33_ASAP7_75t_L g1408 ( 
.A(n_1362),
.B(n_1352),
.C(n_1346),
.Y(n_1408)
);

AOI221xp5_ASAP7_75t_L g1409 ( 
.A1(n_1358),
.A2(n_1363),
.B1(n_1362),
.B2(n_1381),
.C(n_1380),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1385),
.B(n_1324),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1369),
.B(n_1324),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1358),
.A2(n_1313),
.B1(n_1356),
.B2(n_1330),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1369),
.B(n_1336),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_SL g1414 ( 
.A(n_1377),
.B(n_1321),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1370),
.B(n_1329),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1364),
.B(n_1338),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1370),
.B(n_1329),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1415),
.B(n_1372),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1407),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1411),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1411),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1407),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1399),
.Y(n_1423)
);

INVxp67_ASAP7_75t_SL g1424 ( 
.A(n_1397),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1417),
.B(n_1386),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_1393),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_1413),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_R g1428 ( 
.A(n_1389),
.B(n_1255),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1397),
.Y(n_1429)
);

CKINVDCx6p67_ASAP7_75t_R g1430 ( 
.A(n_1396),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1410),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1395),
.B(n_1331),
.Y(n_1432)
);

NAND2x1p5_ASAP7_75t_L g1433 ( 
.A(n_1401),
.B(n_1384),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1400),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1409),
.B(n_1386),
.Y(n_1435)
);

INVxp67_ASAP7_75t_SL g1436 ( 
.A(n_1404),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1408),
.B(n_1373),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1408),
.B(n_1375),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1419),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1434),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1420),
.B(n_1405),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1419),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1422),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1422),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1425),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1423),
.B(n_1431),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1423),
.B(n_1390),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1423),
.B(n_1416),
.Y(n_1448)
);

OAI32xp33_ASAP7_75t_L g1449 ( 
.A1(n_1435),
.A2(n_1388),
.A3(n_1412),
.B1(n_1398),
.B2(n_1392),
.Y(n_1449)
);

INVx4_ASAP7_75t_L g1450 ( 
.A(n_1430),
.Y(n_1450)
);

OAI33xp33_ASAP7_75t_L g1451 ( 
.A1(n_1435),
.A2(n_1412),
.A3(n_1403),
.B1(n_1398),
.B2(n_1391),
.B3(n_1399),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1421),
.B(n_1404),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1431),
.B(n_1424),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1437),
.B(n_1406),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1427),
.B(n_1394),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1446),
.B(n_1436),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1450),
.B(n_1430),
.Y(n_1457)
);

AOI21xp33_ASAP7_75t_L g1458 ( 
.A1(n_1449),
.A2(n_1436),
.B(n_1388),
.Y(n_1458)
);

AOI21xp33_ASAP7_75t_L g1459 ( 
.A1(n_1449),
.A2(n_1391),
.B(n_1403),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1447),
.B(n_1429),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1440),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1450),
.B(n_1430),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1439),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1439),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1450),
.B(n_1426),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1442),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_L g1467 ( 
.A(n_1451),
.B(n_1200),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1450),
.B(n_1441),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1440),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1440),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1441),
.B(n_1426),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1442),
.Y(n_1472)
);

INVx2_ASAP7_75t_SL g1473 ( 
.A(n_1452),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1446),
.B(n_1454),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1441),
.B(n_1433),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1455),
.B(n_1433),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1454),
.B(n_1437),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1454),
.B(n_1438),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1443),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1455),
.B(n_1433),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1447),
.B(n_1429),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1444),
.Y(n_1482)
);

NOR3xp33_ASAP7_75t_L g1483 ( 
.A(n_1451),
.B(n_1282),
.C(n_1402),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1453),
.B(n_1438),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1453),
.B(n_1418),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1448),
.B(n_1200),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1455),
.B(n_1433),
.Y(n_1487)
);

NAND2x1p5_ASAP7_75t_L g1488 ( 
.A(n_1452),
.B(n_1351),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1448),
.B(n_1418),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1461),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1460),
.B(n_1481),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1461),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1474),
.B(n_1445),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1457),
.B(n_1452),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1463),
.Y(n_1495)
);

INVx1_ASAP7_75t_SL g1496 ( 
.A(n_1465),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1457),
.B(n_1452),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1463),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1472),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1461),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1472),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_1462),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1482),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1482),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1469),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1462),
.B(n_1452),
.Y(n_1506)
);

INVx2_ASAP7_75t_SL g1507 ( 
.A(n_1473),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1469),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1460),
.B(n_1445),
.Y(n_1509)
);

NAND2xp33_ASAP7_75t_L g1510 ( 
.A(n_1483),
.B(n_1428),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1469),
.Y(n_1511)
);

INVx1_ASAP7_75t_SL g1512 ( 
.A(n_1465),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1464),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1470),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1473),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1464),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1466),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1470),
.Y(n_1518)
);

INVx1_ASAP7_75t_SL g1519 ( 
.A(n_1474),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1470),
.Y(n_1520)
);

NAND2x1p5_ASAP7_75t_L g1521 ( 
.A(n_1468),
.B(n_1414),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1466),
.Y(n_1522)
);

INVxp67_ASAP7_75t_L g1523 ( 
.A(n_1467),
.Y(n_1523)
);

NOR3xp33_ASAP7_75t_L g1524 ( 
.A(n_1458),
.B(n_1282),
.C(n_1402),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1479),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_L g1526 ( 
.A(n_1523),
.B(n_1486),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1498),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1523),
.B(n_1483),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1496),
.B(n_1459),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1510),
.A2(n_1458),
.B1(n_1459),
.B2(n_1468),
.Y(n_1530)
);

AOI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1524),
.A2(n_1481),
.B1(n_1480),
.B2(n_1487),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1513),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1502),
.B(n_1473),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1496),
.B(n_1456),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1512),
.B(n_1456),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1513),
.Y(n_1536)
);

OAI21xp33_ASAP7_75t_SL g1537 ( 
.A1(n_1507),
.A2(n_1478),
.B(n_1477),
.Y(n_1537)
);

INVx2_ASAP7_75t_SL g1538 ( 
.A(n_1507),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1512),
.B(n_1471),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1524),
.A2(n_1478),
.B1(n_1477),
.B2(n_1488),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1516),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1494),
.B(n_1475),
.Y(n_1542)
);

OAI221xp5_ASAP7_75t_L g1543 ( 
.A1(n_1491),
.A2(n_1488),
.B1(n_1484),
.B2(n_1485),
.C(n_1489),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1502),
.B(n_1292),
.Y(n_1544)
);

A2O1A1Ixp33_ASAP7_75t_L g1545 ( 
.A1(n_1491),
.A2(n_1484),
.B(n_1480),
.C(n_1476),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1519),
.B(n_1471),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1516),
.Y(n_1547)
);

OAI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1519),
.A2(n_1488),
.B(n_1432),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1517),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1517),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_1533),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1532),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1536),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1541),
.Y(n_1554)
);

NAND2xp33_ASAP7_75t_L g1555 ( 
.A(n_1530),
.B(n_1515),
.Y(n_1555)
);

NOR2x1_ASAP7_75t_L g1556 ( 
.A(n_1544),
.B(n_1502),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1547),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1528),
.B(n_1494),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1526),
.B(n_1497),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1549),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1527),
.B(n_1529),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1550),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1546),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1533),
.B(n_1497),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1537),
.B(n_1506),
.Y(n_1565)
);

INVx1_ASAP7_75t_SL g1566 ( 
.A(n_1539),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1542),
.B(n_1538),
.Y(n_1567)
);

NOR2x1_ASAP7_75t_SL g1568 ( 
.A(n_1540),
.B(n_1507),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1534),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1535),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1551),
.B(n_1545),
.Y(n_1571)
);

AOI211x1_ASAP7_75t_L g1572 ( 
.A1(n_1565),
.A2(n_1548),
.B(n_1543),
.C(n_1540),
.Y(n_1572)
);

OAI211xp5_ASAP7_75t_SL g1573 ( 
.A1(n_1555),
.A2(n_1548),
.B(n_1531),
.C(n_1499),
.Y(n_1573)
);

OAI21xp5_ASAP7_75t_SL g1574 ( 
.A1(n_1566),
.A2(n_1506),
.B(n_1521),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1568),
.Y(n_1575)
);

BUFx2_ASAP7_75t_L g1576 ( 
.A(n_1556),
.Y(n_1576)
);

AOI21xp33_ASAP7_75t_L g1577 ( 
.A1(n_1555),
.A2(n_1499),
.B(n_1495),
.Y(n_1577)
);

AOI21xp33_ASAP7_75t_L g1578 ( 
.A1(n_1559),
.A2(n_1501),
.B(n_1495),
.Y(n_1578)
);

AOI221xp5_ASAP7_75t_L g1579 ( 
.A1(n_1561),
.A2(n_1501),
.B1(n_1504),
.B2(n_1503),
.C(n_1509),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1569),
.B(n_1509),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_SL g1581 ( 
.A(n_1569),
.B(n_1564),
.Y(n_1581)
);

AOI22x1_ASAP7_75t_SL g1582 ( 
.A1(n_1575),
.A2(n_1563),
.B1(n_1570),
.B2(n_1553),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1576),
.Y(n_1583)
);

NOR3xp33_ASAP7_75t_L g1584 ( 
.A(n_1573),
.B(n_1558),
.C(n_1567),
.Y(n_1584)
);

NOR3xp33_ASAP7_75t_L g1585 ( 
.A(n_1577),
.B(n_1554),
.C(n_1552),
.Y(n_1585)
);

AOI211xp5_ASAP7_75t_L g1586 ( 
.A1(n_1578),
.A2(n_1560),
.B(n_1562),
.C(n_1557),
.Y(n_1586)
);

NOR3xp33_ASAP7_75t_L g1587 ( 
.A(n_1581),
.B(n_1504),
.C(n_1503),
.Y(n_1587)
);

AND5x1_ASAP7_75t_L g1588 ( 
.A(n_1579),
.B(n_1568),
.C(n_1521),
.D(n_1493),
.E(n_1490),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_SL g1589 ( 
.A(n_1572),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1571),
.B(n_1493),
.Y(n_1590)
);

NAND3xp33_ASAP7_75t_SL g1591 ( 
.A(n_1584),
.B(n_1574),
.C(n_1580),
.Y(n_1591)
);

NAND4xp25_ASAP7_75t_L g1592 ( 
.A(n_1587),
.B(n_1303),
.C(n_1292),
.D(n_1522),
.Y(n_1592)
);

NOR3xp33_ASAP7_75t_L g1593 ( 
.A(n_1583),
.B(n_1585),
.C(n_1590),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1582),
.Y(n_1594)
);

AOI211xp5_ASAP7_75t_L g1595 ( 
.A1(n_1586),
.A2(n_1303),
.B(n_1525),
.C(n_1522),
.Y(n_1595)
);

NOR2xp67_ASAP7_75t_L g1596 ( 
.A(n_1592),
.B(n_1525),
.Y(n_1596)
);

AND2x4_ASAP7_75t_SL g1597 ( 
.A(n_1593),
.B(n_1243),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1594),
.Y(n_1598)
);

INVxp67_ASAP7_75t_L g1599 ( 
.A(n_1591),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1595),
.Y(n_1600)
);

AOI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1594),
.A2(n_1589),
.B1(n_1521),
.B2(n_1588),
.Y(n_1601)
);

OAI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1599),
.A2(n_1488),
.B1(n_1518),
.B2(n_1514),
.Y(n_1602)
);

NOR3xp33_ASAP7_75t_L g1603 ( 
.A(n_1598),
.B(n_1492),
.C(n_1490),
.Y(n_1603)
);

NAND3x1_ASAP7_75t_L g1604 ( 
.A(n_1601),
.B(n_1487),
.C(n_1476),
.Y(n_1604)
);

NOR2x1_ASAP7_75t_L g1605 ( 
.A(n_1600),
.B(n_1490),
.Y(n_1605)
);

AOI211xp5_ASAP7_75t_L g1606 ( 
.A1(n_1596),
.A2(n_1520),
.B(n_1518),
.C(n_1514),
.Y(n_1606)
);

XOR2x2_ASAP7_75t_L g1607 ( 
.A(n_1604),
.B(n_1597),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1605),
.B(n_1475),
.Y(n_1608)
);

OA22x2_ASAP7_75t_L g1609 ( 
.A1(n_1602),
.A2(n_1520),
.B1(n_1518),
.B2(n_1514),
.Y(n_1609)
);

XOR2xp5_ASAP7_75t_L g1610 ( 
.A(n_1607),
.B(n_1603),
.Y(n_1610)
);

NAND3xp33_ASAP7_75t_L g1611 ( 
.A(n_1610),
.B(n_1606),
.C(n_1608),
.Y(n_1611)
);

OAI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1611),
.A2(n_1609),
.B1(n_1520),
.B2(n_1511),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1611),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1613),
.Y(n_1614)
);

OR2x6_ASAP7_75t_L g1615 ( 
.A(n_1612),
.B(n_1201),
.Y(n_1615)
);

AOI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1614),
.A2(n_1511),
.B1(n_1508),
.B2(n_1505),
.Y(n_1616)
);

AOI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1615),
.A2(n_1511),
.B1(n_1508),
.B2(n_1505),
.Y(n_1617)
);

OA21x2_ASAP7_75t_L g1618 ( 
.A1(n_1616),
.A2(n_1500),
.B(n_1492),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1618),
.Y(n_1619)
);

OAI221xp5_ASAP7_75t_R g1620 ( 
.A1(n_1619),
.A2(n_1617),
.B1(n_1508),
.B2(n_1505),
.C(n_1500),
.Y(n_1620)
);

AOI211xp5_ASAP7_75t_L g1621 ( 
.A1(n_1620),
.A2(n_1500),
.B(n_1492),
.C(n_1253),
.Y(n_1621)
);


endmodule