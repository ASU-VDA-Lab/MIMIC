module fake_jpeg_19787_n_328 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx11_ASAP7_75t_SL g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_34),
.B(n_38),
.Y(n_44)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_0),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_16),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_55),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_38),
.B(n_20),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_16),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_31),
.B1(n_17),
.B2(n_25),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_56),
.A2(n_58),
.B1(n_35),
.B2(n_18),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_31),
.B1(n_17),
.B2(n_29),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_54),
.A2(n_24),
.B1(n_23),
.B2(n_20),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_40),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_61),
.B(n_62),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_41),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_63),
.A2(n_68),
.B1(n_69),
.B2(n_85),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_39),
.B1(n_35),
.B2(n_31),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_64),
.A2(n_76),
.B1(n_50),
.B2(n_56),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_65),
.B(n_79),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_43),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_52),
.Y(n_92)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_54),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_54),
.A2(n_24),
.B1(n_23),
.B2(n_31),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_18),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_88),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_73),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_41),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_74),
.Y(n_121)
);

NAND3xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_19),
.C(n_26),
.Y(n_75)
);

NAND3xp33_ASAP7_75t_SL g112 ( 
.A(n_75),
.B(n_71),
.C(n_19),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_55),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_46),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_50),
.A2(n_19),
.B1(n_25),
.B2(n_22),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_43),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_50),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_46),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_87),
.B(n_79),
.Y(n_119)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_91),
.Y(n_98)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_90),
.Y(n_100)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_106),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_104),
.A2(n_63),
.B1(n_64),
.B2(n_62),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_59),
.B(n_48),
.Y(n_106)
);

AO22x1_ASAP7_75t_SL g109 ( 
.A1(n_59),
.A2(n_58),
.B1(n_36),
.B2(n_42),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_109),
.B(n_116),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_114),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_67),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_71),
.B(n_66),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_115),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_61),
.B(n_48),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_61),
.B(n_58),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_117),
.B(n_119),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_62),
.A2(n_29),
.B(n_26),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_118),
.A2(n_26),
.B(n_29),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_120),
.B(n_106),
.Y(n_135)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_123),
.A2(n_145),
.B1(n_97),
.B2(n_99),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_74),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_126),
.A2(n_140),
.B(n_141),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_74),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_126),
.Y(n_163)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g130 ( 
.A1(n_116),
.A2(n_87),
.B(n_65),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_130),
.B(n_118),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_110),
.A2(n_82),
.B1(n_45),
.B2(n_91),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_131),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_117),
.A2(n_86),
.B1(n_90),
.B2(n_76),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_132),
.A2(n_139),
.B1(n_144),
.B2(n_146),
.Y(n_155)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_137),
.Y(n_151)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_136),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_96),
.B(n_77),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_96),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_138),
.B(n_30),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_84),
.B1(n_80),
.B2(n_78),
.Y(n_139)
);

NAND2x1_ASAP7_75t_SL g140 ( 
.A(n_100),
.B(n_22),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_95),
.Y(n_142)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_119),
.B(n_41),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_16),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_109),
.A2(n_88),
.B1(n_81),
.B2(n_47),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_104),
.A2(n_47),
.B1(n_89),
.B2(n_45),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_103),
.A2(n_45),
.B1(n_42),
.B2(n_41),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_103),
.A2(n_92),
.B1(n_121),
.B2(n_94),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_147),
.A2(n_100),
.B1(n_93),
.B2(n_114),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_16),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_149),
.A2(n_16),
.B(n_33),
.Y(n_175)
);

AO21x1_ASAP7_75t_L g196 ( 
.A1(n_150),
.A2(n_175),
.B(n_33),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_94),
.C(n_120),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_153),
.B(n_174),
.C(n_133),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_156),
.A2(n_177),
.B1(n_181),
.B2(n_143),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_122),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_157),
.B(n_162),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_158),
.B(n_161),
.Y(n_210)
);

OA22x2_ASAP7_75t_L g160 ( 
.A1(n_138),
.A2(n_97),
.B1(n_99),
.B2(n_108),
.Y(n_160)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_163),
.B(n_180),
.Y(n_187)
);

OAI32xp33_ASAP7_75t_L g164 ( 
.A1(n_148),
.A2(n_27),
.A3(n_45),
.B1(n_18),
.B2(n_32),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_146),
.Y(n_190)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_107),
.B(n_83),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_149),
.B(n_141),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_124),
.B(n_108),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_168),
.B(n_171),
.Y(n_211)
);

MAJx2_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_27),
.C(n_32),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_173),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_124),
.B(n_101),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_107),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_172),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_128),
.B(n_72),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_128),
.B(n_102),
.C(n_101),
.Y(n_174)
);

OAI22x1_ASAP7_75t_L g177 ( 
.A1(n_140),
.A2(n_27),
.B1(n_33),
.B2(n_22),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_142),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_179),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_125),
.B(n_27),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_135),
.B(n_72),
.Y(n_181)
);

A2O1A1O1Ixp25_ASAP7_75t_L g185 ( 
.A1(n_150),
.A2(n_125),
.B(n_148),
.C(n_149),
.D(n_137),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_185),
.B(n_201),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_155),
.A2(n_123),
.B1(n_145),
.B2(n_132),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_186),
.A2(n_189),
.B1(n_183),
.B2(n_210),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_188),
.B(n_198),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_155),
.A2(n_139),
.B1(n_144),
.B2(n_133),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_190),
.B(n_194),
.Y(n_230)
);

AOI21x1_ASAP7_75t_SL g229 ( 
.A1(n_192),
.A2(n_196),
.B(n_200),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_193),
.B(n_195),
.Y(n_233)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_163),
.B(n_140),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_178),
.A2(n_0),
.B(n_1),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_197),
.A2(n_199),
.B1(n_205),
.B2(n_207),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_166),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_178),
.A2(n_159),
.B1(n_156),
.B2(n_167),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_170),
.A2(n_25),
.B(n_30),
.Y(n_200)
);

XNOR2x1_ASAP7_75t_L g201 ( 
.A(n_153),
.B(n_32),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_170),
.A2(n_30),
.B(n_33),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_208),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_177),
.A2(n_102),
.B1(n_113),
.B2(n_21),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_113),
.C(n_16),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_175),
.C(n_152),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_164),
.A2(n_158),
.B1(n_151),
.B2(n_181),
.Y(n_207)
);

OAI32xp33_ASAP7_75t_L g208 ( 
.A1(n_151),
.A2(n_32),
.A3(n_21),
.B1(n_16),
.B2(n_10),
.Y(n_208)
);

NAND2xp33_ASAP7_75t_SL g213 ( 
.A(n_160),
.B(n_113),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_165),
.Y(n_223)
);

OA21x2_ASAP7_75t_L g214 ( 
.A1(n_160),
.A2(n_0),
.B(n_1),
.Y(n_214)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_209),
.Y(n_215)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_203),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_223),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_233),
.Y(n_242)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_209),
.Y(n_219)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_219),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_222),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_194),
.A2(n_173),
.B1(n_176),
.B2(n_182),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_224),
.A2(n_225),
.B1(n_236),
.B2(n_237),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_214),
.A2(n_154),
.B1(n_161),
.B2(n_169),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_227),
.A2(n_231),
.B1(n_13),
.B2(n_11),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_186),
.A2(n_180),
.B1(n_2),
.B2(n_3),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_193),
.B(n_15),
.C(n_14),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_2),
.C(n_3),
.Y(n_260)
);

NAND3xp33_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_13),
.C(n_12),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_184),
.Y(n_251)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_211),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_235),
.Y(n_255)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_214),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_238),
.A2(n_239),
.B1(n_183),
.B2(n_197),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_1),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_254),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_187),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_245),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_187),
.Y(n_245)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_221),
.B(n_204),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_250),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_218),
.B(n_195),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_257),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_204),
.C(n_192),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_256),
.C(n_250),
.Y(n_269)
);

AOI221xp5_ASAP7_75t_L g253 ( 
.A1(n_226),
.A2(n_189),
.B1(n_185),
.B2(n_202),
.C(n_191),
.Y(n_253)
);

AOI21xp33_ASAP7_75t_L g261 ( 
.A1(n_253),
.A2(n_239),
.B(n_217),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_190),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_200),
.C(n_196),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_213),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_228),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_220),
.B(n_10),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_229),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_260),
.B(n_256),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_261),
.A2(n_223),
.B(n_248),
.Y(n_281)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_263),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_240),
.A2(n_227),
.B1(n_236),
.B2(n_228),
.Y(n_265)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_265),
.Y(n_290)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_267),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_238),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_268),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_269),
.B(n_272),
.Y(n_288)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_243),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_273),
.Y(n_284)
);

NOR2x1_ASAP7_75t_SL g272 ( 
.A(n_259),
.B(n_229),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_246),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_241),
.B(n_224),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_275),
.Y(n_286)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_276),
.Y(n_282)
);

A2O1A1Ixp33_ASAP7_75t_SL g277 ( 
.A1(n_254),
.A2(n_223),
.B(n_231),
.C(n_252),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_277),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_242),
.C(n_244),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_283),
.Y(n_304)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_245),
.C(n_260),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_266),
.A2(n_2),
.B(n_3),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_285),
.A2(n_5),
.B(n_6),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_287),
.B(n_6),
.Y(n_301)
);

A2O1A1Ixp33_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_291)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_291),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_264),
.B(n_5),
.C(n_6),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_293),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_288),
.A2(n_262),
.B(n_277),
.Y(n_295)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_295),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_281),
.A2(n_277),
.B(n_278),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_296),
.A2(n_292),
.B(n_291),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_302),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_279),
.A2(n_275),
.B1(n_265),
.B2(n_278),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_299),
.A2(n_301),
.B1(n_287),
.B2(n_289),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_270),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_280),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_290),
.A2(n_270),
.B1(n_7),
.B2(n_8),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_305),
.B(n_308),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_298),
.B(n_286),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_307),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_294),
.A2(n_290),
.B(n_286),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_304),
.B(n_284),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_293),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_310),
.B(n_312),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_282),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_311),
.B(n_282),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_314),
.B(n_315),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_284),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_309),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_321),
.A2(n_322),
.B(n_319),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_316),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_320),
.C(n_318),
.Y(n_324)
);

OAI321xp33_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_307),
.A3(n_292),
.B1(n_303),
.B2(n_300),
.C(n_285),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_301),
.C(n_297),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_8),
.B(n_319),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_327),
.B(n_8),
.Y(n_328)
);


endmodule