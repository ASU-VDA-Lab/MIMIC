module fake_jpeg_26820_n_174 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_174);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_5),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_24),
.B(n_28),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_6),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_21),
.Y(n_30)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_29),
.A2(n_22),
.B1(n_18),
.B2(n_15),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_34),
.A2(n_35),
.B1(n_36),
.B2(n_11),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_30),
.A2(n_22),
.B1(n_15),
.B2(n_11),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_29),
.A2(n_22),
.B1(n_15),
.B2(n_11),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_40),
.B(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_42),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_27),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_32),
.B1(n_26),
.B2(n_33),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_46),
.B1(n_55),
.B2(n_37),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_21),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_45),
.B1(n_53),
.B2(n_54),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_21),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_26),
.B1(n_29),
.B2(n_25),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_28),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_49),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_31),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_52),
.Y(n_65)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_26),
.B1(n_19),
.B2(n_21),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_32),
.B1(n_37),
.B2(n_38),
.Y(n_73)
);

O2A1O1Ixp33_ASAP7_75t_SL g55 ( 
.A1(n_35),
.A2(n_25),
.B(n_23),
.C(n_19),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_35),
.B1(n_34),
.B2(n_32),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_57),
.A2(n_72),
.B1(n_73),
.B2(n_37),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_33),
.C(n_31),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_70),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_55),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_64),
.Y(n_78)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_17),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_69),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_33),
.C(n_31),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_45),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_53),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_72)
);

OAI32xp33_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_45),
.A3(n_55),
.B1(n_52),
.B2(n_14),
.Y(n_76)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_77),
.A2(n_87),
.B(n_91),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_85),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_64),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_88),
.Y(n_103)
);

CKINVDCx10_ASAP7_75t_R g82 ( 
.A(n_56),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_82),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_93),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_84),
.Y(n_113)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_50),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_17),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_89),
.B(n_12),
.Y(n_98)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_57),
.A2(n_51),
.B(n_1),
.Y(n_91)
);

OAI32xp33_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_19),
.A3(n_16),
.B1(n_12),
.B2(n_20),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_59),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_69),
.A2(n_38),
.B1(n_37),
.B2(n_25),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_94),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_96),
.B(n_84),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_63),
.B(n_70),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_98),
.B(n_74),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_58),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_109),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_63),
.B(n_1),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_105),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_0),
.B(n_1),
.Y(n_105)
);

AOI21x1_ASAP7_75t_SL g106 ( 
.A1(n_76),
.A2(n_38),
.B(n_23),
.Y(n_106)
);

NOR2x1_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_111),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_79),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_80),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_38),
.Y(n_109)
);

AOI221xp5_ASAP7_75t_L g110 ( 
.A1(n_91),
.A2(n_12),
.B1(n_20),
.B2(n_13),
.C(n_4),
.Y(n_110)
);

AOI221xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_92),
.B1(n_93),
.B2(n_10),
.C(n_4),
.Y(n_124)
);

AOI21x1_ASAP7_75t_L g111 ( 
.A1(n_78),
.A2(n_31),
.B(n_13),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_116),
.B(n_118),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_107),
.B(n_88),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_117),
.B(n_123),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_81),
.C(n_77),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_77),
.C(n_94),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_120),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_90),
.C(n_74),
.Y(n_120)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_85),
.B1(n_82),
.B2(n_48),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_125),
.A2(n_114),
.B1(n_102),
.B2(n_104),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_112),
.B(n_8),
.Y(n_126)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_23),
.B1(n_13),
.B2(n_20),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_128),
.A2(n_114),
.B1(n_95),
.B2(n_102),
.Y(n_133)
);

OA21x2_ASAP7_75t_L g130 ( 
.A1(n_127),
.A2(n_100),
.B(n_101),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_134),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_133),
.A2(n_121),
.B1(n_118),
.B2(n_103),
.Y(n_142)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

OAI21x1_ASAP7_75t_L g139 ( 
.A1(n_120),
.A2(n_111),
.B(n_106),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_139),
.A2(n_108),
.B(n_105),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_140),
.B(n_104),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_136),
.B(n_119),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_144),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_142),
.A2(n_121),
.B1(n_134),
.B2(n_127),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_135),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_129),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_147),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_140),
.B(n_129),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_146),
.B(n_130),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_108),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_149),
.B(n_115),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_7),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_155),
.B(n_149),
.C(n_103),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_146),
.A2(n_131),
.B1(n_128),
.B2(n_130),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_156),
.A2(n_148),
.B(n_131),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_157),
.A2(n_6),
.B(n_10),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_158),
.B(n_7),
.Y(n_164)
);

AOI322xp5_ASAP7_75t_L g159 ( 
.A1(n_155),
.A2(n_141),
.A3(n_96),
.B1(n_133),
.B2(n_145),
.C1(n_137),
.C2(n_12),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_159),
.B(n_160),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_20),
.C(n_23),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_153),
.C(n_156),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_161),
.B(n_162),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_13),
.C(n_4),
.Y(n_168)
);

NOR2xp67_ASAP7_75t_SL g165 ( 
.A(n_161),
.B(n_6),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_165),
.A2(n_167),
.B(n_8),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_168),
.A2(n_169),
.B(n_170),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_166),
.A2(n_9),
.B1(n_8),
.B2(n_3),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_170),
.A2(n_163),
.B(n_2),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_171),
.A2(n_0),
.B(n_2),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_172),
.Y(n_174)
);


endmodule