module real_jpeg_24633_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_0),
.B(n_15),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_0),
.B(n_49),
.Y(n_137)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_4),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_4),
.B(n_31),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_4),
.B(n_57),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_4),
.B(n_24),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_4),
.B(n_28),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_5),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_5),
.B(n_49),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_5),
.B(n_31),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_6),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_6),
.B(n_24),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_6),
.B(n_49),
.Y(n_67)
);

NAND2x1_ASAP7_75t_SL g82 ( 
.A(n_6),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_6),
.B(n_28),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_6),
.B(n_38),
.Y(n_150)
);

INVx8_ASAP7_75t_SL g120 ( 
.A(n_7),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_8),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_8),
.B(n_49),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_8),
.B(n_31),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_8),
.B(n_24),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_10),
.B(n_149),
.Y(n_148)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_11),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_12),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_12),
.B(n_24),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_12),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_12),
.B(n_49),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_12),
.B(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_14),
.B(n_28),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_14),
.B(n_31),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_14),
.B(n_49),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_14),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_14),
.B(n_38),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_14),
.B(n_118),
.Y(n_138)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_15),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_127),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_99),
.C(n_100),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_60),
.C(n_71),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_41),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_21),
.B(n_33),
.C(n_41),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_26),
.C(n_29),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_22),
.A2(n_23),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_32),
.B(n_89),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_34),
.B(n_36),
.C(n_37),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_51),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_42),
.B(n_52),
.C(n_53),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_47),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_46),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_56),
.B2(n_59),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_54),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_55),
.B(n_59),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g83 ( 
.A(n_58),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.C(n_70),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_64),
.A2(n_65),
.B1(n_70),
.B2(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_66),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_75)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_95),
.C(n_96),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_80),
.C(n_86),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_78),
.C(n_79),
.Y(n_95)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_81),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.C(n_90),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_89),
.B(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_113),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_114),
.C(n_126),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_109),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_108),
.C(n_109),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_104),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_107),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx24_ASAP7_75t_SL g163 ( 
.A(n_109),
.Y(n_163)
);

FAx1_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_111),
.CI(n_112),
.CON(n_109),
.SN(n_109)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_111),
.C(n_112),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_126),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_124),
.B2(n_125),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_117),
.Y(n_123)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_123),
.C(n_125),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_144),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_139),
.Y(n_134)
);

BUFx24_ASAP7_75t_SL g164 ( 
.A(n_135),
.Y(n_164)
);

FAx1_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_137),
.CI(n_138),
.CON(n_135),
.SN(n_135)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_152),
.B1(n_160),
.B2(n_161),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_147),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_150),
.B(n_151),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_148),
.B(n_150),
.Y(n_151)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_157),
.Y(n_152)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx11_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);


endmodule