module fake_jpeg_1414_n_126 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_126);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_126;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_20),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx4f_ASAP7_75t_SL g43 ( 
.A(n_10),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_17),
.B(n_19),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_54),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_43),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_42),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_40),
.Y(n_59)
);

NOR2x1_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_47),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_62),
.B(n_64),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_46),
.B1(n_43),
.B2(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_37),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_74),
.Y(n_85)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_77),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_39),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_78),
.B(n_86),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_44),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_82),
.Y(n_91)
);

AO21x2_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_48),
.B(n_53),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_63),
.B1(n_46),
.B2(n_2),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_41),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_36),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_88),
.B(n_89),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_75),
.B(n_76),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_51),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_34),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_63),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_93),
.Y(n_111)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_95),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_0),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_15),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_101),
.C(n_102),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_99),
.A2(n_100),
.B(n_103),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_22),
.C(n_32),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_14),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_97),
.A2(n_83),
.B(n_79),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_108),
.B1(n_24),
.B2(n_27),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_23),
.C(n_30),
.Y(n_106)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_11),
.B(n_29),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_33),
.Y(n_110)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_112),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_117)
);

XOR2x1_ASAP7_75t_SL g115 ( 
.A(n_111),
.B(n_3),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_115),
.A2(n_112),
.B(n_109),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_116),
.A2(n_117),
.B1(n_104),
.B2(n_107),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_119),
.C(n_120),
.Y(n_121)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_114),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_28),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_123),
.Y(n_124)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_115),
.C(n_6),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_8),
.Y(n_126)
);


endmodule