module fake_ariane_550_n_1452 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_332, n_294, n_197, n_176, n_34, n_172, n_347, n_183, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_367, n_345, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_349, n_346, n_214, n_348, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_327, n_77, n_15, n_23, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_267, n_335, n_350, n_291, n_344, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_11, n_129, n_126, n_282, n_328, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_333, n_221, n_321, n_86, n_361, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_343, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_358, n_105, n_30, n_131, n_263, n_360, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_118, n_121, n_353, n_22, n_241, n_29, n_357, n_191, n_80, n_211, n_97, n_322, n_251, n_116, n_351, n_39, n_359, n_155, n_127, n_1452);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_347;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_327;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_333;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_343;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_360;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_118;
input n_121;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_191;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_351;
input n_39;
input n_359;
input n_155;
input n_127;

output n_1452;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_995;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_559;
wire n_495;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1314;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_611;
wire n_1295;
wire n_1013;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1396;
wire n_1230;
wire n_612;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1391;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1432;
wire n_1108;
wire n_851;
wire n_444;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_436;
wire n_669;
wire n_931;
wire n_619;
wire n_437;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_479;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1363;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_1401;
wire n_1419;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1414;
wire n_1134;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_529;
wire n_502;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1371;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1218;
wire n_861;
wire n_1431;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_551;
wire n_417;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_608;
wire n_1037;
wire n_1329;
wire n_1257;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_649;
wire n_374;
wire n_1352;
wire n_643;
wire n_1441;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_1450;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1438;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_368;
wire n_467;
wire n_1422;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1440;
wire n_1370;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1420;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1444;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_1427;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1407;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_1361;
wire n_1057;
wire n_978;
wire n_1011;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_679;
wire n_663;
wire n_443;
wire n_1412;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_671;
wire n_1409;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1129;
wire n_1252;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_1434;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_675;

INVx1_ASAP7_75t_SL g368 ( 
.A(n_54),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_305),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_46),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_58),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_52),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_95),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_303),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_290),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_142),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_330),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_360),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_198),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_129),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_137),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_227),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_11),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_225),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_26),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_185),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_343),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_27),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_161),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_221),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_106),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_364),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_20),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_294),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_120),
.Y(n_395)
);

CKINVDCx14_ASAP7_75t_R g396 ( 
.A(n_19),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_134),
.Y(n_397)
);

CKINVDCx14_ASAP7_75t_R g398 ( 
.A(n_93),
.Y(n_398)
);

BUFx5_ASAP7_75t_L g399 ( 
.A(n_53),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_158),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_130),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_262),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_32),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_317),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_28),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_121),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_332),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_180),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_264),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_283),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_25),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_362),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_7),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_291),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_57),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_23),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_361),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_103),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_63),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_281),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_145),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_127),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_293),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_337),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_320),
.Y(n_425)
);

BUFx10_ASAP7_75t_L g426 ( 
.A(n_85),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_252),
.Y(n_427)
);

CKINVDCx14_ASAP7_75t_R g428 ( 
.A(n_24),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_278),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_86),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_266),
.Y(n_431)
);

INVx2_ASAP7_75t_SL g432 ( 
.A(n_59),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_273),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_254),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_0),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_0),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_329),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_300),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_4),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_243),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_344),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_298),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_186),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_335),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_351),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_178),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g447 ( 
.A(n_196),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_182),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_119),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_324),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_355),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_213),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_88),
.Y(n_453)
);

CKINVDCx14_ASAP7_75t_R g454 ( 
.A(n_125),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_191),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_367),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_189),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_248),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_353),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g460 ( 
.A(n_150),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_122),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_321),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_265),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_18),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_201),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_328),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_25),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_171),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_212),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_199),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_358),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_301),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_61),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_246),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_215),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_167),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_23),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_98),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_157),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_338),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_255),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_309),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_286),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_341),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_275),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_231),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_21),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_152),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_272),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_147),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_24),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_187),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_192),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_331),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_339),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_9),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_280),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_101),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_288),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_253),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_91),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_325),
.Y(n_502)
);

BUFx2_ASAP7_75t_SL g503 ( 
.A(n_159),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_308),
.Y(n_504)
);

CKINVDCx16_ASAP7_75t_R g505 ( 
.A(n_163),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_7),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_336),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_289),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_241),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_245),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_74),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_334),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_107),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_342),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_110),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_76),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_311),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_366),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_285),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_194),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_80),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_172),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_168),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_118),
.Y(n_524)
);

CKINVDCx14_ASAP7_75t_R g525 ( 
.A(n_256),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_81),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_104),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_184),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_322),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_346),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_222),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_327),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_45),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_148),
.Y(n_534)
);

INVxp67_ASAP7_75t_SL g535 ( 
.A(n_333),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_356),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_234),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_149),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_44),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_230),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_4),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_314),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_116),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_40),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_15),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_33),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_68),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_268),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_173),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_117),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_295),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_220),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_3),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_349),
.Y(n_554)
);

BUFx10_ASAP7_75t_L g555 ( 
.A(n_357),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_165),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_138),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_123),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_345),
.Y(n_559)
);

BUFx2_ASAP7_75t_L g560 ( 
.A(n_229),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_77),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_340),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_49),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_115),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_354),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_144),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_143),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_270),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_70),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_6),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_219),
.Y(n_571)
);

INVxp67_ASAP7_75t_SL g572 ( 
.A(n_160),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_32),
.Y(n_573)
);

INVxp33_ASAP7_75t_R g574 ( 
.A(n_17),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_316),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_18),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_388),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_370),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_389),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_401),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_544),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_544),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_416),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_396),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_R g585 ( 
.A(n_398),
.B(n_43),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_428),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_402),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_467),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_438),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_506),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_553),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_436),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_576),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_436),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_541),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_560),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_426),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_426),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_555),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_386),
.B(n_1),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_480),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_383),
.Y(n_602)
);

INVxp33_ASAP7_75t_SL g603 ( 
.A(n_385),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_483),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_555),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_386),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_377),
.B(n_1),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_485),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_497),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_395),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_512),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_397),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_533),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_400),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_412),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_536),
.Y(n_616)
);

INVxp33_ASAP7_75t_L g617 ( 
.A(n_574),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_556),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_414),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_393),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_415),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_557),
.Y(n_622)
);

INVxp67_ASAP7_75t_L g623 ( 
.A(n_403),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_405),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_419),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_411),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_413),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_471),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_424),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_471),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_435),
.Y(n_631)
);

INVxp67_ASAP7_75t_SL g632 ( 
.A(n_372),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_439),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_546),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_434),
.Y(n_635)
);

CKINVDCx16_ASAP7_75t_R g636 ( 
.A(n_505),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_453),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_464),
.Y(n_638)
);

NOR2xp67_ASAP7_75t_L g639 ( 
.A(n_477),
.B(n_2),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_454),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_455),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_487),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_491),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_525),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_456),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_406),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_465),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_496),
.Y(n_648)
);

CKINVDCx16_ASAP7_75t_R g649 ( 
.A(n_503),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_473),
.Y(n_650)
);

INVxp67_ASAP7_75t_SL g651 ( 
.A(n_372),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_474),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_478),
.Y(n_653)
);

CKINVDCx16_ASAP7_75t_R g654 ( 
.A(n_406),
.Y(n_654)
);

INVxp67_ASAP7_75t_SL g655 ( 
.A(n_425),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_479),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_482),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_486),
.B(n_2),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_545),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_570),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_489),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_504),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_515),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_573),
.Y(n_664)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_575),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_519),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_529),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_530),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_369),
.Y(n_669)
);

CKINVDCx14_ASAP7_75t_R g670 ( 
.A(n_371),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_534),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_373),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_548),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_558),
.Y(n_674)
);

CKINVDCx20_ASAP7_75t_R g675 ( 
.A(n_374),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_559),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_567),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_375),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_569),
.B(n_3),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_646),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_583),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_588),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_590),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_649),
.B(n_425),
.Y(n_684)
);

NAND2xp33_ASAP7_75t_SL g685 ( 
.A(n_600),
.B(n_432),
.Y(n_685)
);

XOR2xp5_ASAP7_75t_L g686 ( 
.A(n_589),
.B(n_376),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_591),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_646),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_646),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_646),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_654),
.B(n_447),
.Y(n_691)
);

BUFx8_ASAP7_75t_L g692 ( 
.A(n_626),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_606),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_593),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_628),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_670),
.B(n_484),
.Y(n_696)
);

BUFx2_ASAP7_75t_L g697 ( 
.A(n_660),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_577),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_672),
.B(n_517),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_584),
.B(n_517),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_630),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_678),
.B(n_384),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_636),
.B(n_627),
.Y(n_703)
);

HB1xp67_ASAP7_75t_L g704 ( 
.A(n_584),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_581),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_631),
.B(n_468),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_582),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_592),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_592),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_641),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_671),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_610),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_594),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_620),
.B(n_500),
.Y(n_714)
);

BUFx8_ASAP7_75t_L g715 ( 
.A(n_597),
.Y(n_715)
);

INVxp67_ASAP7_75t_L g716 ( 
.A(n_602),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_612),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_598),
.B(n_368),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_595),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_658),
.Y(n_720)
);

BUFx2_ASAP7_75t_L g721 ( 
.A(n_642),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_614),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_615),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_619),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_643),
.B(n_648),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_621),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_SL g727 ( 
.A(n_640),
.B(n_431),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_625),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_629),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_635),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_637),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_623),
.B(n_460),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_645),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_659),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_620),
.Y(n_735)
);

CKINVDCx20_ASAP7_75t_R g736 ( 
.A(n_634),
.Y(n_736)
);

NAND2xp33_ASAP7_75t_SL g737 ( 
.A(n_585),
.B(n_406),
.Y(n_737)
);

NOR2x1_ASAP7_75t_L g738 ( 
.A(n_599),
.B(n_463),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_647),
.Y(n_739)
);

OAI21x1_ASAP7_75t_L g740 ( 
.A1(n_650),
.A2(n_572),
.B(n_535),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_652),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_665),
.Y(n_742)
);

INVxp67_ASAP7_75t_L g743 ( 
.A(n_602),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_653),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_605),
.B(n_520),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_632),
.B(n_378),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_656),
.Y(n_747)
);

INVxp67_ASAP7_75t_L g748 ( 
.A(n_633),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_596),
.B(n_406),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_651),
.B(n_379),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_657),
.Y(n_751)
);

AND2x6_ASAP7_75t_L g752 ( 
.A(n_661),
.B(n_470),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_662),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_655),
.B(n_380),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_663),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_673),
.B(n_381),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_667),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_668),
.Y(n_758)
);

NAND2xp33_ASAP7_75t_SL g759 ( 
.A(n_585),
.B(n_470),
.Y(n_759)
);

INVx1_ASAP7_75t_SL g760 ( 
.A(n_578),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_674),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_676),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_677),
.B(n_382),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_666),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_666),
.Y(n_765)
);

CKINVDCx8_ASAP7_75t_R g766 ( 
.A(n_579),
.Y(n_766)
);

OR2x2_ASAP7_75t_L g767 ( 
.A(n_764),
.B(n_580),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_718),
.B(n_633),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_721),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_695),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_720),
.B(n_607),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_720),
.B(n_607),
.Y(n_772)
);

AND2x6_ASAP7_75t_L g773 ( 
.A(n_738),
.B(n_470),
.Y(n_773)
);

HB1xp67_ASAP7_75t_SL g774 ( 
.A(n_766),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_695),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_705),
.Y(n_776)
);

OR2x2_ASAP7_75t_L g777 ( 
.A(n_765),
.B(n_587),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_728),
.Y(n_778)
);

CKINVDCx20_ASAP7_75t_R g779 ( 
.A(n_736),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_728),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_695),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_732),
.B(n_603),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_720),
.B(n_679),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_707),
.Y(n_784)
);

INVx1_ASAP7_75t_SL g785 ( 
.A(n_760),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_701),
.Y(n_786)
);

INVx2_ASAP7_75t_SL g787 ( 
.A(n_718),
.Y(n_787)
);

BUFx2_ASAP7_75t_L g788 ( 
.A(n_692),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_701),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_701),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_719),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_735),
.B(n_624),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_728),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_747),
.Y(n_794)
);

NAND2xp33_ASAP7_75t_L g795 ( 
.A(n_696),
.B(n_387),
.Y(n_795)
);

INVx5_ASAP7_75t_L g796 ( 
.A(n_752),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_719),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_761),
.B(n_679),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_693),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_719),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_747),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_691),
.B(n_669),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_745),
.B(n_638),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_747),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_710),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_711),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_681),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_746),
.B(n_638),
.Y(n_808)
);

INVx5_ASAP7_75t_L g809 ( 
.A(n_752),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_713),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_745),
.B(n_699),
.Y(n_811)
);

INVx3_ASAP7_75t_L g812 ( 
.A(n_761),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_680),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_712),
.B(n_399),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_716),
.B(n_664),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_688),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_750),
.B(n_664),
.Y(n_817)
);

AND2x2_ASAP7_75t_SL g818 ( 
.A(n_727),
.B(n_644),
.Y(n_818)
);

OR2x2_ASAP7_75t_L g819 ( 
.A(n_708),
.B(n_604),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_682),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_702),
.B(n_675),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_683),
.Y(n_822)
);

CKINVDCx16_ASAP7_75t_R g823 ( 
.A(n_686),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_704),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_717),
.B(n_399),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_743),
.B(n_586),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_687),
.Y(n_827)
);

OR2x2_ASAP7_75t_SL g828 ( 
.A(n_698),
.B(n_617),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_690),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_692),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_726),
.Y(n_831)
);

BUFx3_ASAP7_75t_L g832 ( 
.A(n_694),
.Y(n_832)
);

OR2x2_ASAP7_75t_L g833 ( 
.A(n_709),
.B(n_608),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_739),
.Y(n_834)
);

INVx1_ASAP7_75t_SL g835 ( 
.A(n_697),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_744),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_751),
.Y(n_837)
);

AND2x2_ASAP7_75t_SL g838 ( 
.A(n_742),
.B(n_601),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_722),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_723),
.Y(n_840)
);

OR2x2_ASAP7_75t_L g841 ( 
.A(n_748),
.B(n_609),
.Y(n_841)
);

AND2x4_ASAP7_75t_L g842 ( 
.A(n_700),
.B(n_639),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_689),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_754),
.B(n_611),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_724),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_689),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_734),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_729),
.A2(n_470),
.B1(n_399),
.B2(n_391),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_700),
.B(n_616),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_684),
.Y(n_850)
);

INVx4_ASAP7_75t_L g851 ( 
.A(n_752),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_730),
.A2(n_618),
.B1(n_622),
.B2(n_613),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_715),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_749),
.B(n_390),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_731),
.B(n_399),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_763),
.B(n_392),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_740),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_689),
.Y(n_858)
);

NOR2xp67_ASAP7_75t_L g859 ( 
.A(n_802),
.B(n_725),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_785),
.B(n_703),
.Y(n_860)
);

OAI221xp5_ASAP7_75t_L g861 ( 
.A1(n_808),
.A2(n_685),
.B1(n_741),
.B2(n_753),
.C(n_733),
.Y(n_861)
);

BUFx8_ASAP7_75t_L g862 ( 
.A(n_788),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_785),
.B(n_769),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_776),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_784),
.Y(n_865)
);

AOI22xp5_ASAP7_75t_L g866 ( 
.A1(n_808),
.A2(n_737),
.B1(n_759),
.B2(n_706),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_834),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_807),
.Y(n_868)
);

AO22x2_ASAP7_75t_L g869 ( 
.A1(n_852),
.A2(n_749),
.B1(n_757),
.B2(n_755),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_831),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_820),
.Y(n_871)
);

CKINVDCx11_ASAP7_75t_R g872 ( 
.A(n_779),
.Y(n_872)
);

AO22x2_ASAP7_75t_L g873 ( 
.A1(n_852),
.A2(n_758),
.B1(n_762),
.B2(n_714),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_835),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_822),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_827),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_831),
.Y(n_877)
);

AND2x4_ASAP7_75t_L g878 ( 
.A(n_830),
.B(n_756),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_839),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_840),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_845),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_817),
.B(n_752),
.Y(n_882)
);

CKINVDCx20_ASAP7_75t_R g883 ( 
.A(n_823),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_787),
.A2(n_715),
.B1(n_399),
.B2(n_404),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_791),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_799),
.Y(n_886)
);

INVxp67_ASAP7_75t_L g887 ( 
.A(n_835),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_768),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_836),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_837),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_810),
.Y(n_891)
);

OR2x2_ASAP7_75t_SL g892 ( 
.A(n_841),
.B(n_5),
.Y(n_892)
);

AO22x2_ASAP7_75t_L g893 ( 
.A1(n_768),
.A2(n_8),
.B1(n_5),
.B2(n_6),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_805),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_817),
.B(n_394),
.Y(n_895)
);

NAND3xp33_ASAP7_75t_SL g896 ( 
.A(n_847),
.B(n_571),
.C(n_408),
.Y(n_896)
);

AO22x2_ASAP7_75t_L g897 ( 
.A1(n_803),
.A2(n_777),
.B1(n_767),
.B2(n_819),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_806),
.Y(n_898)
);

INVxp67_ASAP7_75t_L g899 ( 
.A(n_849),
.Y(n_899)
);

AO22x2_ASAP7_75t_L g900 ( 
.A1(n_803),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_900)
);

AO22x2_ASAP7_75t_L g901 ( 
.A1(n_833),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_824),
.B(n_407),
.Y(n_902)
);

INVxp67_ASAP7_75t_L g903 ( 
.A(n_774),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_812),
.B(n_409),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_812),
.B(n_410),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_856),
.B(n_417),
.Y(n_906)
);

BUFx8_ASAP7_75t_L g907 ( 
.A(n_826),
.Y(n_907)
);

OAI221xp5_ASAP7_75t_L g908 ( 
.A1(n_771),
.A2(n_421),
.B1(n_422),
.B2(n_420),
.C(n_418),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_856),
.B(n_423),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_832),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_813),
.Y(n_911)
);

AO22x2_ASAP7_75t_L g912 ( 
.A1(n_811),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_814),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_844),
.A2(n_427),
.B1(n_430),
.B2(n_429),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_814),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_816),
.Y(n_916)
);

OR2x6_ASAP7_75t_SL g917 ( 
.A(n_853),
.B(n_433),
.Y(n_917)
);

OAI221xp5_ASAP7_75t_L g918 ( 
.A1(n_771),
.A2(n_568),
.B1(n_566),
.B2(n_565),
.C(n_564),
.Y(n_918)
);

OAI221xp5_ASAP7_75t_L g919 ( 
.A1(n_772),
.A2(n_563),
.B1(n_562),
.B2(n_561),
.C(n_554),
.Y(n_919)
);

INVxp67_ASAP7_75t_L g920 ( 
.A(n_774),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_782),
.B(n_437),
.Y(n_921)
);

AO22x2_ASAP7_75t_L g922 ( 
.A1(n_850),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_825),
.Y(n_923)
);

INVxp67_ASAP7_75t_L g924 ( 
.A(n_792),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_829),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_772),
.B(n_440),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_825),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_855),
.Y(n_928)
);

OAI22xp33_ASAP7_75t_SL g929 ( 
.A1(n_821),
.A2(n_442),
.B1(n_443),
.B2(n_441),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_786),
.Y(n_930)
);

AO22x2_ASAP7_75t_L g931 ( 
.A1(n_842),
.A2(n_19),
.B1(n_16),
.B2(n_17),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_778),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_855),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_778),
.Y(n_934)
);

BUFx8_ASAP7_75t_L g935 ( 
.A(n_815),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_801),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_780),
.Y(n_937)
);

AO22x2_ASAP7_75t_L g938 ( 
.A1(n_842),
.A2(n_21),
.B1(n_16),
.B2(n_20),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_783),
.B(n_798),
.Y(n_939)
);

BUFx10_ASAP7_75t_L g940 ( 
.A(n_838),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_804),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_780),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_783),
.B(n_444),
.Y(n_943)
);

NAND2x1p5_ASAP7_75t_L g944 ( 
.A(n_793),
.B(n_22),
.Y(n_944)
);

AO22x2_ASAP7_75t_L g945 ( 
.A1(n_818),
.A2(n_27),
.B1(n_22),
.B2(n_26),
.Y(n_945)
);

OAI221xp5_ASAP7_75t_L g946 ( 
.A1(n_798),
.A2(n_552),
.B1(n_551),
.B2(n_550),
.C(n_549),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_800),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_794),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_770),
.Y(n_949)
);

AO22x2_ASAP7_75t_L g950 ( 
.A1(n_854),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_775),
.Y(n_951)
);

OR2x2_ASAP7_75t_SL g952 ( 
.A(n_828),
.B(n_29),
.Y(n_952)
);

AO22x2_ASAP7_75t_L g953 ( 
.A1(n_781),
.A2(n_33),
.B1(n_30),
.B2(n_31),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_791),
.Y(n_954)
);

OA22x2_ASAP7_75t_L g955 ( 
.A1(n_790),
.A2(n_792),
.B1(n_857),
.B2(n_773),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_924),
.B(n_791),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_859),
.B(n_797),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_863),
.B(n_797),
.Y(n_958)
);

NAND2xp33_ASAP7_75t_SL g959 ( 
.A(n_939),
.B(n_797),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_866),
.B(n_902),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_887),
.B(n_789),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_860),
.B(n_789),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_895),
.B(n_773),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_926),
.B(n_789),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_943),
.B(n_848),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_899),
.B(n_848),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_874),
.B(n_851),
.Y(n_967)
);

NAND2xp33_ASAP7_75t_SL g968 ( 
.A(n_906),
.B(n_851),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_888),
.B(n_857),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_897),
.B(n_773),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_929),
.B(n_796),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_935),
.B(n_796),
.Y(n_972)
);

NAND2xp33_ASAP7_75t_SL g973 ( 
.A(n_909),
.B(n_795),
.Y(n_973)
);

NAND2xp33_ASAP7_75t_SL g974 ( 
.A(n_864),
.B(n_843),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_910),
.B(n_796),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_878),
.B(n_809),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_882),
.B(n_809),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_903),
.B(n_809),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_914),
.B(n_858),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_904),
.B(n_846),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_905),
.B(n_445),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_921),
.B(n_446),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_865),
.B(n_448),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_868),
.B(n_449),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_871),
.B(n_773),
.Y(n_985)
);

XNOR2xp5_ASAP7_75t_L g986 ( 
.A(n_883),
.B(n_450),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_875),
.B(n_451),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_876),
.B(n_452),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_879),
.B(n_457),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_880),
.B(n_458),
.Y(n_990)
);

NAND2xp33_ASAP7_75t_SL g991 ( 
.A(n_881),
.B(n_547),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_885),
.B(n_459),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_897),
.B(n_940),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_894),
.B(n_461),
.Y(n_994)
);

NAND2xp33_ASAP7_75t_SL g995 ( 
.A(n_898),
.B(n_462),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_920),
.B(n_913),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_915),
.B(n_466),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_923),
.B(n_469),
.Y(n_998)
);

NAND2xp33_ASAP7_75t_SL g999 ( 
.A(n_927),
.B(n_543),
.Y(n_999)
);

NAND2xp33_ASAP7_75t_SL g1000 ( 
.A(n_928),
.B(n_472),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_933),
.B(n_475),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_867),
.B(n_476),
.Y(n_1002)
);

NAND2xp33_ASAP7_75t_SL g1003 ( 
.A(n_932),
.B(n_542),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_870),
.B(n_481),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_873),
.B(n_488),
.Y(n_1005)
);

NAND2xp33_ASAP7_75t_SL g1006 ( 
.A(n_934),
.B(n_490),
.Y(n_1006)
);

NAND2xp33_ASAP7_75t_SL g1007 ( 
.A(n_937),
.B(n_540),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_877),
.B(n_492),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_930),
.B(n_907),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_884),
.B(n_493),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_948),
.B(n_494),
.Y(n_1011)
);

NAND2xp33_ASAP7_75t_SL g1012 ( 
.A(n_942),
.B(n_539),
.Y(n_1012)
);

NAND2xp33_ASAP7_75t_SL g1013 ( 
.A(n_936),
.B(n_941),
.Y(n_1013)
);

NAND2xp33_ASAP7_75t_SL g1014 ( 
.A(n_886),
.B(n_495),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_944),
.B(n_498),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_954),
.B(n_499),
.Y(n_1016)
);

NAND2xp33_ASAP7_75t_SL g1017 ( 
.A(n_890),
.B(n_538),
.Y(n_1017)
);

NAND2xp33_ASAP7_75t_SL g1018 ( 
.A(n_891),
.B(n_501),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_955),
.B(n_502),
.Y(n_1019)
);

NAND2xp33_ASAP7_75t_SL g1020 ( 
.A(n_892),
.B(n_507),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_889),
.B(n_508),
.Y(n_1021)
);

NAND2xp33_ASAP7_75t_SL g1022 ( 
.A(n_896),
.B(n_509),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_873),
.B(n_510),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_947),
.B(n_511),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_949),
.B(n_513),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_951),
.B(n_514),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_962),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_L g1028 ( 
.A1(n_977),
.A2(n_916),
.B(n_911),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_986),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_958),
.Y(n_1030)
);

CKINVDCx20_ASAP7_75t_R g1031 ( 
.A(n_972),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_L g1032 ( 
.A1(n_964),
.A2(n_925),
.B(n_869),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_973),
.A2(n_861),
.B(n_946),
.Y(n_1033)
);

INVxp67_ASAP7_75t_SL g1034 ( 
.A(n_960),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_966),
.B(n_869),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_956),
.Y(n_1036)
);

AOI21x1_ASAP7_75t_L g1037 ( 
.A1(n_965),
.A2(n_912),
.B(n_953),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_985),
.Y(n_1038)
);

AOI21x1_ASAP7_75t_L g1039 ( 
.A1(n_963),
.A2(n_912),
.B(n_953),
.Y(n_1039)
);

O2A1O1Ixp5_ASAP7_75t_SL g1040 ( 
.A1(n_1019),
.A2(n_950),
.B(n_901),
.C(n_945),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_980),
.A2(n_399),
.B(n_922),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_978),
.B(n_872),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_1013),
.A2(n_908),
.B(n_919),
.C(n_918),
.Y(n_1043)
);

NOR2xp67_ASAP7_75t_L g1044 ( 
.A(n_978),
.B(n_982),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_998),
.A2(n_518),
.B(n_516),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_997),
.A2(n_901),
.B(n_950),
.C(n_900),
.Y(n_1046)
);

AO31x2_ASAP7_75t_L g1047 ( 
.A1(n_1005),
.A2(n_1023),
.A3(n_987),
.B(n_959),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_968),
.A2(n_922),
.B(n_931),
.Y(n_1048)
);

AO21x2_ASAP7_75t_L g1049 ( 
.A1(n_969),
.A2(n_945),
.B(n_938),
.Y(n_1049)
);

BUFx12f_ASAP7_75t_L g1050 ( 
.A(n_978),
.Y(n_1050)
);

BUFx10_ASAP7_75t_L g1051 ( 
.A(n_1022),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_961),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_993),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_981),
.A2(n_938),
.B(n_931),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_970),
.B(n_893),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_SL g1056 ( 
.A1(n_999),
.A2(n_917),
.B(n_952),
.C(n_900),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_979),
.A2(n_957),
.B(n_971),
.Y(n_1057)
);

INVx1_ASAP7_75t_SL g1058 ( 
.A(n_1009),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_975),
.A2(n_48),
.B(n_47),
.Y(n_1059)
);

AO31x2_ASAP7_75t_L g1060 ( 
.A1(n_974),
.A2(n_893),
.A3(n_209),
.B(n_210),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_996),
.Y(n_1061)
);

INVxp67_ASAP7_75t_SL g1062 ( 
.A(n_967),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_1020),
.A2(n_862),
.B1(n_537),
.B2(n_532),
.Y(n_1063)
);

AO31x2_ASAP7_75t_L g1064 ( 
.A1(n_1001),
.A2(n_206),
.A3(n_365),
.B(n_363),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_1000),
.A2(n_531),
.B(n_528),
.C(n_527),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_976),
.B(n_31),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_991),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1024),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_995),
.A2(n_526),
.B(n_524),
.C(n_523),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_983),
.A2(n_522),
.B(n_521),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_1015),
.B(n_1002),
.Y(n_1071)
);

NAND2x1_ASAP7_75t_L g1072 ( 
.A(n_1017),
.B(n_50),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_984),
.A2(n_34),
.B(n_35),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1014),
.B(n_34),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1025),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_988),
.B(n_35),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_1016),
.A2(n_55),
.B(n_51),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_989),
.B(n_36),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_990),
.A2(n_60),
.B(n_56),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_994),
.A2(n_64),
.B(n_62),
.Y(n_1080)
);

AO31x2_ASAP7_75t_L g1081 ( 
.A1(n_1018),
.A2(n_205),
.A3(n_352),
.B(n_350),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_1026),
.A2(n_66),
.B(n_65),
.Y(n_1082)
);

CKINVDCx11_ASAP7_75t_R g1083 ( 
.A(n_1003),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1011),
.B(n_36),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_1006),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1004),
.B(n_37),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1008),
.A2(n_69),
.B(n_67),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1021),
.Y(n_1088)
);

INVx1_ASAP7_75t_SL g1089 ( 
.A(n_1058),
.Y(n_1089)
);

HB1xp67_ASAP7_75t_L g1090 ( 
.A(n_1035),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_1057),
.A2(n_992),
.B(n_1010),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1061),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_1050),
.Y(n_1093)
);

OR2x2_ASAP7_75t_L g1094 ( 
.A(n_1029),
.B(n_1007),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1034),
.B(n_1012),
.Y(n_1095)
);

NOR2x1_ASAP7_75t_SL g1096 ( 
.A(n_1036),
.B(n_37),
.Y(n_1096)
);

AO21x2_ASAP7_75t_L g1097 ( 
.A1(n_1032),
.A2(n_72),
.B(n_71),
.Y(n_1097)
);

OAI221xp5_ASAP7_75t_SL g1098 ( 
.A1(n_1046),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.C(n_41),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_1042),
.B(n_359),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_1028),
.A2(n_75),
.B(n_73),
.Y(n_1100)
);

NOR2xp67_ASAP7_75t_L g1101 ( 
.A(n_1067),
.B(n_78),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_1055),
.B(n_38),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1041),
.A2(n_82),
.B(n_79),
.Y(n_1103)
);

HB1xp67_ASAP7_75t_L g1104 ( 
.A(n_1038),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_1042),
.Y(n_1105)
);

INVx2_ASAP7_75t_SL g1106 ( 
.A(n_1051),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_1053),
.B(n_39),
.Y(n_1107)
);

OAI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1033),
.A2(n_1043),
.B(n_1048),
.Y(n_1108)
);

NAND3xp33_ASAP7_75t_L g1109 ( 
.A(n_1073),
.B(n_41),
.C(n_42),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1027),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1030),
.Y(n_1111)
);

AO21x2_ASAP7_75t_L g1112 ( 
.A1(n_1037),
.A2(n_84),
.B(n_83),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_1054),
.A2(n_42),
.B1(n_87),
.B2(n_89),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1052),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1066),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1088),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1049),
.B(n_90),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_1059),
.A2(n_92),
.B(n_94),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1078),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_1031),
.Y(n_1120)
);

AOI22xp33_ASAP7_75t_L g1121 ( 
.A1(n_1068),
.A2(n_96),
.B1(n_97),
.B2(n_99),
.Y(n_1121)
);

OA21x2_ASAP7_75t_L g1122 ( 
.A1(n_1082),
.A2(n_100),
.B(n_102),
.Y(n_1122)
);

AOI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_1074),
.A2(n_105),
.B1(n_108),
.B2(n_109),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_1077),
.A2(n_1039),
.B(n_1079),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_1080),
.A2(n_111),
.B(n_112),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_1047),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_1045),
.A2(n_113),
.B(n_114),
.C(n_124),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1086),
.Y(n_1128)
);

A2O1A1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_1044),
.A2(n_126),
.B(n_128),
.C(n_131),
.Y(n_1129)
);

INVx6_ASAP7_75t_L g1130 ( 
.A(n_1051),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_1083),
.Y(n_1131)
);

OAI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1087),
.A2(n_132),
.B(n_133),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1075),
.A2(n_135),
.B1(n_136),
.B2(n_139),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_1085),
.Y(n_1134)
);

HB1xp67_ASAP7_75t_L g1135 ( 
.A(n_1047),
.Y(n_1135)
);

BUFx12f_ASAP7_75t_L g1136 ( 
.A(n_1071),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_1071),
.B(n_348),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_1072),
.A2(n_140),
.B(n_141),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1040),
.A2(n_1062),
.B(n_1084),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1076),
.B(n_146),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1070),
.A2(n_151),
.B(n_153),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1063),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1126),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_1116),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1104),
.Y(n_1145)
);

OA21x2_ASAP7_75t_L g1146 ( 
.A1(n_1108),
.A2(n_1065),
.B(n_1047),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1104),
.Y(n_1147)
);

HB1xp67_ASAP7_75t_L g1148 ( 
.A(n_1114),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1110),
.Y(n_1149)
);

NAND2x1p5_ASAP7_75t_L g1150 ( 
.A(n_1091),
.B(n_1060),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1102),
.B(n_1060),
.Y(n_1151)
);

OR2x2_ASAP7_75t_L g1152 ( 
.A(n_1090),
.B(n_1060),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1126),
.Y(n_1153)
);

AND2x4_ASAP7_75t_L g1154 ( 
.A(n_1137),
.B(n_1081),
.Y(n_1154)
);

INVx4_ASAP7_75t_L g1155 ( 
.A(n_1105),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1111),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_1130),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1124),
.A2(n_1108),
.B(n_1100),
.Y(n_1158)
);

OA21x2_ASAP7_75t_L g1159 ( 
.A1(n_1135),
.A2(n_1069),
.B(n_1081),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1135),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1090),
.B(n_1081),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1117),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1117),
.Y(n_1163)
);

BUFx3_ASAP7_75t_L g1164 ( 
.A(n_1130),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1137),
.B(n_1064),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1092),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_1103),
.A2(n_1064),
.B(n_1056),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1140),
.B(n_1064),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1097),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1097),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1112),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1107),
.B(n_162),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_1095),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1112),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1139),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_1095),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1122),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1128),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1122),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1119),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1115),
.Y(n_1181)
);

INVx2_ASAP7_75t_SL g1182 ( 
.A(n_1130),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1118),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1141),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1099),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_1131),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_1089),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1089),
.B(n_1134),
.Y(n_1188)
);

INVxp67_ASAP7_75t_SL g1189 ( 
.A(n_1105),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1125),
.A2(n_164),
.B(n_166),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1138),
.Y(n_1191)
);

INVxp67_ASAP7_75t_L g1192 ( 
.A(n_1120),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1096),
.Y(n_1193)
);

BUFx3_ASAP7_75t_L g1194 ( 
.A(n_1105),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1099),
.B(n_169),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1123),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1109),
.Y(n_1197)
);

INVx2_ASAP7_75t_SL g1198 ( 
.A(n_1136),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1101),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_1093),
.Y(n_1200)
);

XNOR2xp5_ASAP7_75t_L g1201 ( 
.A(n_1188),
.B(n_1094),
.Y(n_1201)
);

XNOR2xp5_ASAP7_75t_L g1202 ( 
.A(n_1187),
.B(n_1106),
.Y(n_1202)
);

CKINVDCx12_ASAP7_75t_R g1203 ( 
.A(n_1195),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1149),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_1194),
.B(n_1129),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_R g1206 ( 
.A(n_1186),
.B(n_1113),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_R g1207 ( 
.A(n_1186),
.B(n_1121),
.Y(n_1207)
);

OR2x6_ASAP7_75t_L g1208 ( 
.A(n_1198),
.B(n_1132),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_R g1209 ( 
.A(n_1157),
.B(n_1133),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1194),
.B(n_1127),
.Y(n_1210)
);

INVxp67_ASAP7_75t_L g1211 ( 
.A(n_1145),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1149),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_1189),
.B(n_1132),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_R g1214 ( 
.A(n_1157),
.B(n_1142),
.Y(n_1214)
);

NAND2xp33_ASAP7_75t_SL g1215 ( 
.A(n_1195),
.B(n_1098),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_1200),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1164),
.B(n_170),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1173),
.B(n_1098),
.Y(n_1218)
);

INVxp67_ASAP7_75t_L g1219 ( 
.A(n_1147),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_1164),
.B(n_174),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1200),
.B(n_175),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1144),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1173),
.B(n_176),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1176),
.B(n_177),
.Y(n_1224)
);

NAND2xp33_ASAP7_75t_R g1225 ( 
.A(n_1176),
.B(n_179),
.Y(n_1225)
);

INVxp67_ASAP7_75t_L g1226 ( 
.A(n_1148),
.Y(n_1226)
);

OR2x6_ASAP7_75t_L g1227 ( 
.A(n_1198),
.B(n_181),
.Y(n_1227)
);

BUFx2_ASAP7_75t_SL g1228 ( 
.A(n_1182),
.Y(n_1228)
);

XNOR2xp5_ASAP7_75t_L g1229 ( 
.A(n_1192),
.B(n_183),
.Y(n_1229)
);

INVxp67_ASAP7_75t_L g1230 ( 
.A(n_1178),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1180),
.B(n_188),
.Y(n_1231)
);

NAND2xp33_ASAP7_75t_R g1232 ( 
.A(n_1172),
.B(n_190),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_R g1233 ( 
.A(n_1182),
.B(n_1185),
.Y(n_1233)
);

BUFx4f_ASAP7_75t_L g1234 ( 
.A(n_1172),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_1155),
.B(n_193),
.Y(n_1235)
);

NAND2xp33_ASAP7_75t_R g1236 ( 
.A(n_1154),
.B(n_195),
.Y(n_1236)
);

XNOR2xp5_ASAP7_75t_L g1237 ( 
.A(n_1151),
.B(n_197),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_R g1238 ( 
.A(n_1155),
.B(n_200),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1156),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1181),
.B(n_202),
.Y(n_1240)
);

INVx2_ASAP7_75t_SL g1241 ( 
.A(n_1155),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1193),
.B(n_203),
.Y(n_1242)
);

INVxp67_ASAP7_75t_L g1243 ( 
.A(n_1181),
.Y(n_1243)
);

INVxp67_ASAP7_75t_L g1244 ( 
.A(n_1166),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1156),
.B(n_204),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1162),
.B(n_207),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_R g1247 ( 
.A(n_1199),
.B(n_208),
.Y(n_1247)
);

INVxp67_ASAP7_75t_L g1248 ( 
.A(n_1197),
.Y(n_1248)
);

NAND2xp33_ASAP7_75t_R g1249 ( 
.A(n_1154),
.B(n_1165),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1151),
.B(n_211),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1193),
.B(n_1199),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1168),
.B(n_214),
.Y(n_1252)
);

CKINVDCx16_ASAP7_75t_R g1253 ( 
.A(n_1154),
.Y(n_1253)
);

AND2x4_ASAP7_75t_L g1254 ( 
.A(n_1165),
.B(n_216),
.Y(n_1254)
);

NAND2xp33_ASAP7_75t_R g1255 ( 
.A(n_1146),
.B(n_217),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1222),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1239),
.Y(n_1257)
);

BUFx2_ASAP7_75t_L g1258 ( 
.A(n_1216),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1226),
.B(n_1168),
.Y(n_1259)
);

NAND2x1p5_ASAP7_75t_SL g1260 ( 
.A(n_1241),
.B(n_1196),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1253),
.B(n_1161),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1215),
.A2(n_1196),
.B1(n_1163),
.B2(n_1162),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1204),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_1234),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1230),
.B(n_1161),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1248),
.B(n_1163),
.Y(n_1266)
);

OR2x2_ASAP7_75t_L g1267 ( 
.A(n_1211),
.B(n_1219),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1237),
.A2(n_1197),
.B1(n_1152),
.B2(n_1146),
.Y(n_1268)
);

BUFx6f_ASAP7_75t_L g1269 ( 
.A(n_1217),
.Y(n_1269)
);

AND2x6_ASAP7_75t_L g1270 ( 
.A(n_1254),
.B(n_1143),
.Y(n_1270)
);

OR2x2_ASAP7_75t_L g1271 ( 
.A(n_1244),
.B(n_1152),
.Y(n_1271)
);

INVx4_ASAP7_75t_L g1272 ( 
.A(n_1208),
.Y(n_1272)
);

OR2x2_ASAP7_75t_L g1273 ( 
.A(n_1212),
.B(n_1143),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1243),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1251),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1202),
.B(n_1146),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_SL g1277 ( 
.A1(n_1218),
.A2(n_1146),
.B1(n_1159),
.B2(n_1174),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1213),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1202),
.B(n_1175),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1224),
.Y(n_1280)
);

INVx5_ASAP7_75t_L g1281 ( 
.A(n_1208),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1228),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1250),
.A2(n_1174),
.B1(n_1171),
.B2(n_1169),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1223),
.B(n_1153),
.Y(n_1284)
);

INVx4_ASAP7_75t_L g1285 ( 
.A(n_1210),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1245),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1201),
.B(n_1175),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1201),
.B(n_1153),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1252),
.B(n_1160),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1246),
.B(n_1160),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1227),
.A2(n_1150),
.B1(n_1159),
.B2(n_1191),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1233),
.B(n_1159),
.Y(n_1292)
);

INVx4_ASAP7_75t_R g1293 ( 
.A(n_1203),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1240),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1221),
.B(n_1169),
.Y(n_1295)
);

INVxp67_ASAP7_75t_SL g1296 ( 
.A(n_1255),
.Y(n_1296)
);

HB1xp67_ASAP7_75t_L g1297 ( 
.A(n_1231),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1242),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1205),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1227),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1229),
.B(n_1159),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1247),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_1258),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1280),
.B(n_1150),
.Y(n_1304)
);

AO21x2_ASAP7_75t_L g1305 ( 
.A1(n_1291),
.A2(n_1171),
.B(n_1170),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1276),
.B(n_1150),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1267),
.Y(n_1307)
);

OAI221xp5_ASAP7_75t_L g1308 ( 
.A1(n_1296),
.A2(n_1232),
.B1(n_1225),
.B2(n_1236),
.C(n_1249),
.Y(n_1308)
);

OAI221xp5_ASAP7_75t_L g1309 ( 
.A1(n_1296),
.A2(n_1206),
.B1(n_1184),
.B2(n_1191),
.C(n_1170),
.Y(n_1309)
);

INVxp67_ASAP7_75t_SL g1310 ( 
.A(n_1292),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1256),
.Y(n_1311)
);

NAND4xp25_ASAP7_75t_L g1312 ( 
.A(n_1282),
.B(n_1220),
.C(n_1183),
.D(n_1184),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1266),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1297),
.B(n_1177),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1266),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1259),
.B(n_1158),
.Y(n_1316)
);

OR2x2_ASAP7_75t_L g1317 ( 
.A(n_1271),
.B(n_1177),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1287),
.B(n_1158),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1268),
.A2(n_1214),
.B1(n_1209),
.B2(n_1207),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1257),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1281),
.B(n_1179),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_1302),
.Y(n_1322)
);

OAI31xp33_ASAP7_75t_L g1323 ( 
.A1(n_1291),
.A2(n_1235),
.A3(n_1238),
.B(n_1179),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1273),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1274),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1263),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1279),
.B(n_1183),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1278),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1315),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1313),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1320),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1319),
.A2(n_1301),
.B1(n_1262),
.B2(n_1277),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1303),
.B(n_1272),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1324),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1303),
.B(n_1307),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1327),
.B(n_1272),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1322),
.B(n_1300),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1327),
.B(n_1265),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_SL g1339 ( 
.A(n_1323),
.B(n_1281),
.Y(n_1339)
);

INVx3_ASAP7_75t_L g1340 ( 
.A(n_1316),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1317),
.Y(n_1341)
);

AOI21xp33_ASAP7_75t_L g1342 ( 
.A1(n_1309),
.A2(n_1286),
.B(n_1294),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1317),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1314),
.B(n_1288),
.Y(n_1344)
);

OR2x2_ASAP7_75t_L g1345 ( 
.A(n_1324),
.B(n_1284),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1318),
.B(n_1289),
.Y(n_1346)
);

CKINVDCx20_ASAP7_75t_R g1347 ( 
.A(n_1335),
.Y(n_1347)
);

OAI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1339),
.A2(n_1308),
.B1(n_1312),
.B2(n_1281),
.Y(n_1348)
);

INVx4_ASAP7_75t_L g1349 ( 
.A(n_1333),
.Y(n_1349)
);

AO221x2_ASAP7_75t_L g1350 ( 
.A1(n_1329),
.A2(n_1311),
.B1(n_1293),
.B2(n_1292),
.C(n_1299),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1330),
.B(n_1310),
.Y(n_1351)
);

NOR2x1_ASAP7_75t_L g1352 ( 
.A(n_1337),
.B(n_1264),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_1337),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_1344),
.Y(n_1354)
);

NAND2xp33_ASAP7_75t_SL g1355 ( 
.A(n_1346),
.B(n_1264),
.Y(n_1355)
);

NOR2x1_ASAP7_75t_L g1356 ( 
.A(n_1331),
.B(n_1264),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1334),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1357),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1354),
.Y(n_1359)
);

INVx8_ASAP7_75t_L g1360 ( 
.A(n_1347),
.Y(n_1360)
);

INVx2_ASAP7_75t_SL g1361 ( 
.A(n_1349),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1351),
.B(n_1338),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1353),
.B(n_1345),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1350),
.B(n_1342),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1349),
.B(n_1340),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1350),
.B(n_1352),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1356),
.Y(n_1367)
);

INVx1_ASAP7_75t_SL g1368 ( 
.A(n_1355),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1348),
.B(n_1340),
.Y(n_1369)
);

INVx1_ASAP7_75t_SL g1370 ( 
.A(n_1347),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1349),
.B(n_1340),
.Y(n_1371)
);

OR2x2_ASAP7_75t_L g1372 ( 
.A(n_1351),
.B(n_1284),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1363),
.B(n_1318),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1358),
.Y(n_1374)
);

OAI32xp33_ASAP7_75t_L g1375 ( 
.A1(n_1364),
.A2(n_1332),
.A3(n_1339),
.B1(n_1285),
.B2(n_1336),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1368),
.A2(n_1332),
.B1(n_1285),
.B2(n_1316),
.Y(n_1376)
);

OAI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1370),
.A2(n_1277),
.B(n_1290),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1361),
.B(n_1341),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1358),
.Y(n_1379)
);

NAND2x1p5_ASAP7_75t_L g1380 ( 
.A(n_1359),
.B(n_1269),
.Y(n_1380)
);

AOI322xp5_ASAP7_75t_L g1381 ( 
.A1(n_1360),
.A2(n_1306),
.A3(n_1341),
.B1(n_1343),
.B2(n_1290),
.C1(n_1261),
.C2(n_1283),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1360),
.Y(n_1382)
);

OR2x2_ASAP7_75t_L g1383 ( 
.A(n_1373),
.B(n_1372),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1382),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1374),
.B(n_1362),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1379),
.B(n_1367),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1378),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1380),
.B(n_1365),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1376),
.Y(n_1389)
);

INVxp67_ASAP7_75t_L g1390 ( 
.A(n_1384),
.Y(n_1390)
);

INVx1_ASAP7_75t_SL g1391 ( 
.A(n_1386),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1385),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1387),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1383),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1388),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1389),
.B(n_1375),
.Y(n_1396)
);

NOR3xp33_ASAP7_75t_L g1397 ( 
.A(n_1396),
.B(n_1390),
.C(n_1391),
.Y(n_1397)
);

NOR3xp33_ASAP7_75t_L g1398 ( 
.A(n_1391),
.B(n_1377),
.C(n_1366),
.Y(n_1398)
);

NOR3x1_ASAP7_75t_L g1399 ( 
.A(n_1394),
.B(n_1367),
.C(n_1369),
.Y(n_1399)
);

OAI21xp5_ASAP7_75t_SL g1400 ( 
.A1(n_1395),
.A2(n_1371),
.B(n_1381),
.Y(n_1400)
);

NAND4xp25_ASAP7_75t_SL g1401 ( 
.A(n_1392),
.B(n_1381),
.C(n_1293),
.D(n_1304),
.Y(n_1401)
);

OAI211xp5_ASAP7_75t_SL g1402 ( 
.A1(n_1393),
.A2(n_1325),
.B(n_1343),
.C(n_1298),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1395),
.B(n_1269),
.Y(n_1403)
);

OAI221xp5_ASAP7_75t_L g1404 ( 
.A1(n_1396),
.A2(n_1269),
.B1(n_1306),
.B2(n_1328),
.C(n_1326),
.Y(n_1404)
);

OAI221xp5_ASAP7_75t_L g1405 ( 
.A1(n_1400),
.A2(n_1326),
.B1(n_1328),
.B2(n_1275),
.C(n_1260),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1403),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1397),
.Y(n_1407)
);

A2O1A1Ixp33_ASAP7_75t_SL g1408 ( 
.A1(n_1398),
.A2(n_1401),
.B(n_1399),
.C(n_1404),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1402),
.A2(n_1305),
.B1(n_1270),
.B2(n_1295),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1397),
.Y(n_1410)
);

OAI31xp33_ASAP7_75t_L g1411 ( 
.A1(n_1400),
.A2(n_1321),
.A3(n_1295),
.B(n_1305),
.Y(n_1411)
);

NOR2x1_ASAP7_75t_L g1412 ( 
.A(n_1407),
.B(n_1305),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1406),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1410),
.Y(n_1414)
);

INVx2_ASAP7_75t_SL g1415 ( 
.A(n_1408),
.Y(n_1415)
);

OAI21xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1411),
.A2(n_1167),
.B(n_1190),
.Y(n_1416)
);

OAI211xp5_ASAP7_75t_SL g1417 ( 
.A1(n_1405),
.A2(n_1409),
.B(n_1270),
.C(n_224),
.Y(n_1417)
);

XOR2x2_ASAP7_75t_L g1418 ( 
.A(n_1407),
.B(n_1321),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1406),
.B(n_1270),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1406),
.B(n_1270),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1415),
.B(n_1321),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_R g1422 ( 
.A(n_1413),
.B(n_218),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_SL g1423 ( 
.A(n_1414),
.B(n_1167),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_R g1424 ( 
.A(n_1420),
.B(n_223),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1418),
.B(n_1190),
.Y(n_1425)
);

NAND2xp33_ASAP7_75t_SL g1426 ( 
.A(n_1419),
.B(n_226),
.Y(n_1426)
);

NAND3xp33_ASAP7_75t_SL g1427 ( 
.A(n_1417),
.B(n_347),
.C(n_232),
.Y(n_1427)
);

NAND2xp33_ASAP7_75t_SL g1428 ( 
.A(n_1416),
.B(n_228),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_R g1429 ( 
.A(n_1412),
.B(n_233),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1421),
.Y(n_1430)
);

AOI211xp5_ASAP7_75t_L g1431 ( 
.A1(n_1428),
.A2(n_235),
.B(n_236),
.C(n_237),
.Y(n_1431)
);

AOI211xp5_ASAP7_75t_L g1432 ( 
.A1(n_1426),
.A2(n_238),
.B(n_239),
.C(n_240),
.Y(n_1432)
);

NOR3xp33_ASAP7_75t_L g1433 ( 
.A(n_1427),
.B(n_242),
.C(n_244),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1425),
.A2(n_1423),
.B(n_1424),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1422),
.B(n_247),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_SL g1436 ( 
.A1(n_1429),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1430),
.B(n_257),
.Y(n_1437)
);

OAI221xp5_ASAP7_75t_L g1438 ( 
.A1(n_1434),
.A2(n_258),
.B1(n_259),
.B2(n_260),
.C(n_261),
.Y(n_1438)
);

OA22x2_ASAP7_75t_L g1439 ( 
.A1(n_1436),
.A2(n_263),
.B1(n_267),
.B2(n_269),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1438),
.A2(n_1431),
.B1(n_1432),
.B2(n_1435),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_SL g1441 ( 
.A1(n_1439),
.A2(n_1433),
.B1(n_274),
.B2(n_276),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1437),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1442),
.A2(n_271),
.B1(n_277),
.B2(n_279),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1441),
.A2(n_282),
.B1(n_284),
.B2(n_287),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1444),
.B(n_1440),
.Y(n_1445)
);

O2A1O1Ixp33_ASAP7_75t_L g1446 ( 
.A1(n_1443),
.A2(n_292),
.B(n_296),
.C(n_297),
.Y(n_1446)
);

OAI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1446),
.A2(n_299),
.B(n_302),
.Y(n_1447)
);

AOI222xp33_ASAP7_75t_L g1448 ( 
.A1(n_1445),
.A2(n_304),
.B1(n_306),
.B2(n_307),
.C1(n_310),
.C2(n_312),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1447),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1448),
.Y(n_1450)
);

AOI221xp5_ASAP7_75t_L g1451 ( 
.A1(n_1450),
.A2(n_313),
.B1(n_315),
.B2(n_318),
.C(n_319),
.Y(n_1451)
);

AOI211xp5_ASAP7_75t_L g1452 ( 
.A1(n_1451),
.A2(n_1449),
.B(n_323),
.C(n_326),
.Y(n_1452)
);


endmodule