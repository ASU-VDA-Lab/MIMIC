module fake_jpeg_22623_n_105 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_105);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g26 ( 
.A(n_23),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_27),
.Y(n_36)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_0),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_0),
.Y(n_41)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_12),
.B(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_30),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_22),
.B1(n_23),
.B2(n_13),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_37),
.B1(n_40),
.B2(n_21),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_26),
.A2(n_22),
.B1(n_21),
.B2(n_19),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_16),
.B1(n_14),
.B2(n_13),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_28),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_47),
.B(n_55),
.Y(n_68)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_51),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_24),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_46),
.B(n_49),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_25),
.B(n_27),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_52),
.B1(n_59),
.B2(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_19),
.B1(n_18),
.B2(n_12),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_32),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_54),
.B(n_56),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_15),
.C(n_30),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_35),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_24),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_15),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_58),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_1),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_67),
.B1(n_43),
.B2(n_39),
.Y(n_78)
);

OR2x2_ASAP7_75t_SL g62 ( 
.A(n_46),
.B(n_34),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_55),
.Y(n_74)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_42),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_39),
.B1(n_33),
.B2(n_43),
.Y(n_67)
);

AND2x6_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_5),
.Y(n_69)
);

NAND3xp33_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_51),
.C(n_6),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_65),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_75),
.Y(n_86)
);

AND2x4_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_49),
.Y(n_73)
);

NOR4xp25_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_74),
.C(n_77),
.D(n_79),
.Y(n_88)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_78),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_44),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_39),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_80),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_53),
.C(n_16),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_68),
.C(n_67),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_87),
.C(n_73),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_66),
.C(n_60),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_90),
.C(n_84),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_74),
.C(n_66),
.Y(n_90)
);

BUFx24_ASAP7_75t_SL g91 ( 
.A(n_86),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_69),
.B(n_60),
.Y(n_92)
);

OAI21x1_ASAP7_75t_SL g96 ( 
.A1(n_92),
.A2(n_87),
.B(n_83),
.Y(n_96)
);

BUFx24_ASAP7_75t_SL g93 ( 
.A(n_85),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

AO21x1_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_76),
.B(n_64),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_97),
.B(n_10),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_100),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_95),
.C(n_10),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_94),
.A2(n_16),
.B1(n_14),
.B2(n_20),
.Y(n_100)
);

AOI322xp5_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_6),
.A3(n_9),
.B1(n_2),
.B2(n_3),
.C1(n_14),
.C2(n_20),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_102),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_9),
.Y(n_105)
);


endmodule