module fake_aes_4725_n_492 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_492);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_492;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_217;
wire n_388;
wire n_139;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_2), .Y(n_77) );
BUFx3_ASAP7_75t_L g78 ( .A(n_48), .Y(n_78) );
CKINVDCx16_ASAP7_75t_R g79 ( .A(n_70), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_61), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_24), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_65), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_19), .Y(n_83) );
CKINVDCx16_ASAP7_75t_R g84 ( .A(n_34), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_6), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_0), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_14), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_0), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_52), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_76), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_63), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_58), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_10), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_12), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_33), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_22), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_51), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_23), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_72), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_44), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_39), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_29), .Y(n_102) );
BUFx3_ASAP7_75t_L g103 ( .A(n_42), .Y(n_103) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_55), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_17), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_32), .Y(n_106) );
INVxp67_ASAP7_75t_SL g107 ( .A(n_40), .Y(n_107) );
INVxp33_ASAP7_75t_SL g108 ( .A(n_71), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_8), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_69), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_11), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_10), .Y(n_112) );
BUFx3_ASAP7_75t_L g113 ( .A(n_8), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_36), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_27), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_77), .B(n_1), .Y(n_116) );
INVx3_ASAP7_75t_L g117 ( .A(n_113), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_104), .Y(n_118) );
INVx3_ASAP7_75t_L g119 ( .A(n_113), .Y(n_119) );
AND2x2_ASAP7_75t_L g120 ( .A(n_79), .B(n_1), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_105), .Y(n_121) );
NOR2xp33_ASAP7_75t_L g122 ( .A(n_95), .B(n_2), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_82), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_82), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_104), .Y(n_125) );
INVx6_ASAP7_75t_L g126 ( .A(n_104), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_84), .B(n_3), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_83), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_105), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_80), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_83), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_104), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_89), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_104), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_87), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_89), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_90), .Y(n_137) );
BUFx3_ASAP7_75t_L g138 ( .A(n_117), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_118), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_118), .Y(n_140) );
BUFx3_ASAP7_75t_L g141 ( .A(n_117), .Y(n_141) );
INVx2_ASAP7_75t_SL g142 ( .A(n_123), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_130), .B(n_108), .Y(n_143) );
BUFx3_ASAP7_75t_L g144 ( .A(n_117), .Y(n_144) );
INVxp67_ASAP7_75t_L g145 ( .A(n_120), .Y(n_145) );
AOI22xp33_ASAP7_75t_L g146 ( .A1(n_123), .A2(n_86), .B1(n_93), .B2(n_112), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_118), .Y(n_147) );
NAND3xp33_ASAP7_75t_L g148 ( .A(n_124), .B(n_115), .C(n_114), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_118), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_118), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_136), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_124), .B(n_96), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_125), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_117), .Y(n_154) );
OAI21xp5_ASAP7_75t_L g155 ( .A1(n_128), .A2(n_114), .B(n_90), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_119), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_119), .B(n_87), .Y(n_157) );
AOI22xp33_ASAP7_75t_L g158 ( .A1(n_128), .A2(n_88), .B1(n_112), .B2(n_86), .Y(n_158) );
OR2x2_ASAP7_75t_L g159 ( .A(n_120), .B(n_85), .Y(n_159) );
XNOR2xp5_ASAP7_75t_L g160 ( .A(n_127), .B(n_108), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_133), .B(n_137), .Y(n_161) );
HB1xp67_ASAP7_75t_SL g162 ( .A(n_160), .Y(n_162) );
INVx2_ASAP7_75t_SL g163 ( .A(n_142), .Y(n_163) );
BUFx3_ASAP7_75t_L g164 ( .A(n_138), .Y(n_164) );
INVx2_ASAP7_75t_SL g165 ( .A(n_142), .Y(n_165) );
OAI22xp5_ASAP7_75t_SL g166 ( .A1(n_160), .A2(n_116), .B1(n_109), .B2(n_93), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_151), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_142), .B(n_127), .Y(n_168) );
INVx5_ASAP7_75t_L g169 ( .A(n_154), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_154), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_151), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_154), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_145), .B(n_133), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_161), .B(n_137), .Y(n_174) );
AND2x4_ASAP7_75t_L g175 ( .A(n_155), .B(n_131), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_155), .B(n_136), .Y(n_176) );
OR2x4_ASAP7_75t_L g177 ( .A(n_143), .B(n_122), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_154), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_156), .Y(n_179) );
OAI22xp5_ASAP7_75t_L g180 ( .A1(n_146), .A2(n_136), .B1(n_131), .B2(n_88), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_152), .B(n_119), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_156), .Y(n_182) );
BUFx2_ASAP7_75t_L g183 ( .A(n_145), .Y(n_183) );
AO22x1_ASAP7_75t_L g184 ( .A1(n_157), .A2(n_107), .B1(n_80), .B2(n_81), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_159), .B(n_81), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_156), .Y(n_186) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_138), .Y(n_187) );
INVx3_ASAP7_75t_L g188 ( .A(n_156), .Y(n_188) );
OAI21xp5_ASAP7_75t_L g189 ( .A1(n_148), .A2(n_119), .B(n_115), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_138), .Y(n_190) );
BUFx3_ASAP7_75t_L g191 ( .A(n_141), .Y(n_191) );
BUFx3_ASAP7_75t_L g192 ( .A(n_141), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_159), .B(n_135), .Y(n_193) );
INVx3_ASAP7_75t_L g194 ( .A(n_141), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_173), .B(n_157), .Y(n_195) );
BUFx2_ASAP7_75t_L g196 ( .A(n_183), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_170), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_170), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_163), .A2(n_152), .B(n_144), .Y(n_199) );
BUFx2_ASAP7_75t_L g200 ( .A(n_183), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_170), .Y(n_201) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_187), .Y(n_202) );
INVx3_ASAP7_75t_L g203 ( .A(n_164), .Y(n_203) );
NOR2xp67_ASAP7_75t_L g204 ( .A(n_169), .B(n_148), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_167), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_173), .B(n_146), .Y(n_206) );
INVx5_ASAP7_75t_L g207 ( .A(n_187), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_185), .B(n_158), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_166), .A2(n_157), .B1(n_144), .B2(n_158), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_167), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_171), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_171), .Y(n_212) );
OR2x2_ASAP7_75t_L g213 ( .A(n_166), .B(n_157), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_178), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_193), .B(n_157), .Y(n_215) );
INVx2_ASAP7_75t_SL g216 ( .A(n_169), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_172), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_163), .A2(n_144), .B(n_92), .Y(n_218) );
BUFx2_ASAP7_75t_L g219 ( .A(n_164), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_175), .A2(n_102), .B1(n_91), .B2(n_85), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_187), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_172), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_172), .Y(n_223) );
INVx2_ASAP7_75t_SL g224 ( .A(n_169), .Y(n_224) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_175), .A2(n_111), .B1(n_94), .B2(n_129), .Y(n_225) );
OAI22xp33_ASAP7_75t_L g226 ( .A1(n_177), .A2(n_94), .B1(n_111), .B2(n_91), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_196), .A2(n_175), .B1(n_168), .B2(n_193), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g228 ( .A1(n_211), .A2(n_175), .B1(n_176), .B2(n_181), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_196), .A2(n_188), .B1(n_179), .B2(n_178), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g230 ( .A1(n_200), .A2(n_179), .B1(n_188), .B2(n_186), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g231 ( .A1(n_200), .A2(n_179), .B1(n_188), .B2(n_186), .Y(n_231) );
OAI22xp5_ASAP7_75t_L g232 ( .A1(n_211), .A2(n_176), .B1(n_181), .B2(n_177), .Y(n_232) );
INVx1_ASAP7_75t_SL g233 ( .A(n_215), .Y(n_233) );
OR2x2_ASAP7_75t_L g234 ( .A(n_213), .B(n_184), .Y(n_234) );
BUFx4f_ASAP7_75t_SL g235 ( .A(n_215), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_206), .Y(n_236) );
NAND3xp33_ASAP7_75t_L g237 ( .A(n_225), .B(n_184), .C(n_180), .Y(n_237) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_215), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_206), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_195), .A2(n_179), .B1(n_188), .B2(n_186), .Y(n_240) );
AND2x4_ASAP7_75t_L g241 ( .A(n_195), .B(n_169), .Y(n_241) );
OAI22xp5_ASAP7_75t_L g242 ( .A1(n_211), .A2(n_177), .B1(n_165), .B2(n_163), .Y(n_242) );
CKINVDCx11_ASAP7_75t_R g243 ( .A(n_195), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_215), .Y(n_244) );
NAND2x1_ASAP7_75t_L g245 ( .A(n_216), .B(n_194), .Y(n_245) );
OAI22xp5_ASAP7_75t_L g246 ( .A1(n_208), .A2(n_177), .B1(n_165), .B2(n_191), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_202), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_195), .A2(n_182), .B1(n_192), .B2(n_191), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_213), .A2(n_182), .B1(n_192), .B2(n_191), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_205), .B(n_169), .Y(n_250) );
AOI221xp5_ASAP7_75t_L g251 ( .A1(n_226), .A2(n_180), .B1(n_174), .B2(n_189), .C(n_135), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_205), .B(n_169), .Y(n_252) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_220), .A2(n_162), .B1(n_174), .B2(n_165), .Y(n_253) );
INVxp67_ASAP7_75t_SL g254 ( .A(n_228), .Y(n_254) );
AOI22x1_ASAP7_75t_L g255 ( .A1(n_250), .A2(n_210), .B1(n_212), .B2(n_199), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g256 ( .A1(n_236), .A2(n_210), .B1(n_212), .B2(n_209), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_236), .A2(n_214), .B1(n_219), .B2(n_204), .Y(n_257) );
OAI221xp5_ASAP7_75t_L g258 ( .A1(n_253), .A2(n_189), .B1(n_218), .B2(n_214), .C(n_204), .Y(n_258) );
OAI21xp33_ASAP7_75t_L g259 ( .A1(n_239), .A2(n_121), .B(n_129), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g260 ( .A1(n_239), .A2(n_162), .B1(n_219), .B2(n_224), .Y(n_260) );
AO31x2_ASAP7_75t_L g261 ( .A1(n_246), .A2(n_217), .A3(n_223), .B(n_222), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_234), .A2(n_203), .B1(n_182), .B2(n_192), .Y(n_262) );
AOI221xp5_ASAP7_75t_L g263 ( .A1(n_232), .A2(n_135), .B1(n_121), .B2(n_92), .C(n_110), .Y(n_263) );
OR2x2_ASAP7_75t_L g264 ( .A(n_233), .B(n_197), .Y(n_264) );
AOI221xp5_ASAP7_75t_L g265 ( .A1(n_227), .A2(n_135), .B1(n_106), .B2(n_101), .C(n_97), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_244), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_238), .B(n_197), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_237), .A2(n_203), .B1(n_164), .B2(n_194), .Y(n_268) );
OAI22xp5_ASAP7_75t_L g269 ( .A1(n_249), .A2(n_207), .B1(n_223), .B2(n_222), .Y(n_269) );
OAI21x1_ASAP7_75t_L g270 ( .A1(n_245), .A2(n_217), .B(n_198), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_243), .A2(n_203), .B1(n_194), .B2(n_201), .Y(n_271) );
OR2x6_ASAP7_75t_L g272 ( .A(n_241), .B(n_216), .Y(n_272) );
INVx3_ASAP7_75t_L g273 ( .A(n_241), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_250), .Y(n_274) );
AOI22xp33_ASAP7_75t_SL g275 ( .A1(n_235), .A2(n_203), .B1(n_207), .B2(n_103), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_251), .B(n_198), .Y(n_276) );
OA222x2_ASAP7_75t_L g277 ( .A1(n_256), .A2(n_243), .B1(n_242), .B2(n_78), .C1(n_103), .C2(n_99), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_264), .Y(n_278) );
NOR2x1_ASAP7_75t_SL g279 ( .A(n_269), .B(n_247), .Y(n_279) );
OAI221xp5_ASAP7_75t_L g280 ( .A1(n_259), .A2(n_229), .B1(n_230), .B2(n_231), .C(n_240), .Y(n_280) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_272), .Y(n_281) );
INVx4_ASAP7_75t_L g282 ( .A(n_272), .Y(n_282) );
OR2x2_ASAP7_75t_L g283 ( .A(n_256), .B(n_241), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_274), .B(n_252), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_266), .B(n_252), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_273), .B(n_201), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_255), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g288 ( .A1(n_254), .A2(n_248), .B1(n_78), .B2(n_224), .Y(n_288) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_270), .Y(n_289) );
AOI221xp5_ASAP7_75t_L g290 ( .A1(n_265), .A2(n_98), .B1(n_100), .B2(n_102), .C(n_134), .Y(n_290) );
AOI22xp5_ASAP7_75t_L g291 ( .A1(n_260), .A2(n_194), .B1(n_169), .B2(n_190), .Y(n_291) );
AND2x4_ASAP7_75t_L g292 ( .A(n_273), .B(n_247), .Y(n_292) );
AO21x2_ASAP7_75t_L g293 ( .A1(n_269), .A2(n_134), .B(n_190), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_261), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_267), .B(n_247), .Y(n_295) );
INVxp67_ASAP7_75t_SL g296 ( .A(n_257), .Y(n_296) );
OAI211xp5_ASAP7_75t_L g297 ( .A1(n_263), .A2(n_134), .B(n_132), .C(n_125), .Y(n_297) );
NAND3xp33_ASAP7_75t_L g298 ( .A(n_275), .B(n_125), .C(n_132), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_294), .Y(n_299) );
INVxp67_ASAP7_75t_SL g300 ( .A(n_278), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_294), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_289), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_289), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_282), .B(n_272), .Y(n_304) );
NAND3xp33_ASAP7_75t_L g305 ( .A(n_288), .B(n_258), .C(n_268), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_283), .B(n_261), .Y(n_306) );
AND2x4_ASAP7_75t_L g307 ( .A(n_279), .B(n_261), .Y(n_307) );
AND3x1_ASAP7_75t_L g308 ( .A(n_277), .B(n_271), .C(n_262), .Y(n_308) );
OAI221xp5_ASAP7_75t_SL g309 ( .A1(n_283), .A2(n_276), .B1(n_4), .B2(n_5), .C(n_6), .Y(n_309) );
AOI211xp5_ASAP7_75t_L g310 ( .A1(n_277), .A2(n_125), .B(n_132), .C(n_5), .Y(n_310) );
AND2x4_ASAP7_75t_L g311 ( .A(n_279), .B(n_247), .Y(n_311) );
BUFx3_ASAP7_75t_L g312 ( .A(n_282), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_296), .A2(n_207), .B1(n_221), .B2(n_202), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_282), .Y(n_314) );
AOI33xp33_ASAP7_75t_L g315 ( .A1(n_284), .A2(n_3), .A3(n_4), .B1(n_7), .B2(n_9), .B3(n_11), .Y(n_315) );
OAI21xp33_ASAP7_75t_SL g316 ( .A1(n_295), .A2(n_190), .B(n_9), .Y(n_316) );
OAI31xp33_ASAP7_75t_L g317 ( .A1(n_281), .A2(n_7), .A3(n_12), .B(n_13), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_287), .Y(n_318) );
OAI31xp33_ASAP7_75t_L g319 ( .A1(n_280), .A2(n_13), .A3(n_14), .B(n_150), .Y(n_319) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_295), .Y(n_320) );
OR2x2_ASAP7_75t_L g321 ( .A(n_285), .B(n_221), .Y(n_321) );
OAI221xp5_ASAP7_75t_L g322 ( .A1(n_291), .A2(n_126), .B1(n_207), .B2(n_125), .C(n_132), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_289), .Y(n_323) );
INVx2_ASAP7_75t_SL g324 ( .A(n_292), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_289), .Y(n_325) );
INVx5_ASAP7_75t_L g326 ( .A(n_289), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_320), .B(n_293), .Y(n_327) );
INVx1_ASAP7_75t_SL g328 ( .A(n_314), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_299), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_300), .B(n_293), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_299), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_301), .B(n_284), .Y(n_332) );
INVx3_ASAP7_75t_L g333 ( .A(n_326), .Y(n_333) );
NAND4xp25_ASAP7_75t_L g334 ( .A(n_310), .B(n_290), .C(n_284), .D(n_286), .Y(n_334) );
NOR3xp33_ASAP7_75t_SL g335 ( .A(n_309), .B(n_297), .C(n_298), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_321), .B(n_286), .Y(n_336) );
AOI211x1_ASAP7_75t_L g337 ( .A1(n_308), .A2(n_15), .B(n_16), .C(n_18), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_321), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_306), .B(n_292), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_306), .B(n_293), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_307), .B(n_292), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_314), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_307), .B(n_132), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_324), .B(n_132), .Y(n_344) );
INVx4_ASAP7_75t_L g345 ( .A(n_312), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_315), .B(n_125), .Y(n_346) );
INVx3_ASAP7_75t_L g347 ( .A(n_326), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_324), .B(n_126), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_318), .B(n_221), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_318), .B(n_221), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_307), .B(n_126), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_303), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_310), .B(n_207), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_307), .B(n_20), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_312), .B(n_221), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_312), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_304), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_316), .Y(n_358) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_311), .Y(n_359) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_311), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_308), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_302), .B(n_21), .Y(n_362) );
AND2x2_ASAP7_75t_SL g363 ( .A(n_311), .B(n_202), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_317), .A2(n_202), .B1(n_207), .B2(n_187), .Y(n_364) );
AOI221xp5_ASAP7_75t_L g365 ( .A1(n_319), .A2(n_305), .B1(n_322), .B2(n_313), .C(n_302), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_331), .Y(n_366) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_328), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_361), .B(n_305), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_338), .B(n_311), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_357), .B(n_302), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_340), .B(n_302), .Y(n_371) );
XOR2xp5_ASAP7_75t_L g372 ( .A(n_336), .B(n_325), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_332), .B(n_326), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_329), .Y(n_374) );
OAI21xp33_ASAP7_75t_L g375 ( .A1(n_358), .A2(n_303), .B(n_323), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_342), .Y(n_376) );
OAI21xp5_ASAP7_75t_SL g377 ( .A1(n_334), .A2(n_326), .B(n_202), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_330), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_340), .B(n_326), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_345), .Y(n_380) );
AOI31xp33_ASAP7_75t_L g381 ( .A1(n_354), .A2(n_326), .A3(n_26), .B(n_28), .Y(n_381) );
NAND3xp33_ASAP7_75t_SL g382 ( .A(n_353), .B(n_345), .C(n_365), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_345), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_339), .B(n_25), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_330), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_341), .B(n_30), .Y(n_386) );
INVx2_ASAP7_75t_SL g387 ( .A(n_333), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_341), .B(n_31), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_356), .B(n_35), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_343), .B(n_37), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_327), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_343), .B(n_359), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_360), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_351), .Y(n_394) );
NAND2x1_ASAP7_75t_L g395 ( .A(n_333), .B(n_153), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_352), .B(n_38), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_351), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_344), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_333), .B(n_41), .Y(n_399) );
INVxp33_ASAP7_75t_SL g400 ( .A(n_354), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_363), .B(n_43), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_363), .B(n_45), .Y(n_402) );
NOR3xp33_ASAP7_75t_L g403 ( .A(n_346), .B(n_150), .C(n_147), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_348), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_362), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_347), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_368), .B(n_347), .Y(n_407) );
INVx1_ASAP7_75t_SL g408 ( .A(n_383), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_367), .B(n_355), .Y(n_409) );
INVx3_ASAP7_75t_L g410 ( .A(n_387), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_366), .Y(n_411) );
OAI32xp33_ASAP7_75t_L g412 ( .A1(n_400), .A2(n_337), .A3(n_364), .B1(n_349), .B2(n_350), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_368), .B(n_350), .Y(n_413) );
O2A1O1Ixp33_ASAP7_75t_L g414 ( .A1(n_381), .A2(n_377), .B(n_382), .C(n_404), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_376), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_378), .B(n_335), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_393), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_374), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_385), .B(n_46), .Y(n_419) );
OAI222xp33_ASAP7_75t_L g420 ( .A1(n_372), .A2(n_47), .B1(n_49), .B2(n_50), .C1(n_53), .C2(n_54), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_391), .B(n_56), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_400), .A2(n_187), .B1(n_147), .B2(n_140), .Y(n_422) );
INVx1_ASAP7_75t_SL g423 ( .A(n_372), .Y(n_423) );
INVx1_ASAP7_75t_SL g424 ( .A(n_392), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_398), .B(n_57), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_370), .B(n_59), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_371), .B(n_60), .Y(n_427) );
XNOR2xp5_ASAP7_75t_L g428 ( .A(n_386), .B(n_62), .Y(n_428) );
NOR2xp67_ASAP7_75t_L g429 ( .A(n_387), .B(n_64), .Y(n_429) );
INVx1_ASAP7_75t_SL g430 ( .A(n_386), .Y(n_430) );
INVxp67_ASAP7_75t_L g431 ( .A(n_406), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_369), .B(n_66), .Y(n_432) );
INVx2_ASAP7_75t_SL g433 ( .A(n_395), .Y(n_433) );
AOI21xp33_ASAP7_75t_L g434 ( .A1(n_394), .A2(n_67), .B(n_68), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_397), .B(n_73), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_406), .B(n_74), .Y(n_436) );
XOR2x2_ASAP7_75t_L g437 ( .A(n_388), .B(n_75), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g438 ( .A(n_375), .B(n_139), .Y(n_438) );
INVxp33_ASAP7_75t_L g439 ( .A(n_399), .Y(n_439) );
XNOR2xp5_ASAP7_75t_L g440 ( .A(n_379), .B(n_140), .Y(n_440) );
XOR2x2_ASAP7_75t_L g441 ( .A(n_390), .B(n_187), .Y(n_441) );
O2A1O1Ixp33_ASAP7_75t_L g442 ( .A1(n_384), .A2(n_399), .B(n_389), .C(n_403), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g443 ( .A1(n_405), .A2(n_139), .B1(n_149), .B2(n_153), .C(n_373), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_396), .Y(n_444) );
O2A1O1Ixp33_ASAP7_75t_L g445 ( .A1(n_401), .A2(n_149), .B(n_153), .C(n_402), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_366), .Y(n_446) );
OAI211xp5_ASAP7_75t_SL g447 ( .A1(n_368), .A2(n_149), .B(n_153), .C(n_361), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_380), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_378), .B(n_149), .Y(n_449) );
OAI33xp33_ASAP7_75t_L g450 ( .A1(n_404), .A2(n_149), .A3(n_153), .B1(n_361), .B2(n_385), .B3(n_378), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_377), .A2(n_153), .B(n_381), .Y(n_451) );
O2A1O1Ixp33_ASAP7_75t_SL g452 ( .A1(n_377), .A2(n_380), .B(n_383), .C(n_400), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_L g453 ( .A1(n_382), .A2(n_361), .B(n_368), .C(n_381), .Y(n_453) );
NOR2x1p5_ASAP7_75t_L g454 ( .A(n_382), .B(n_361), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_380), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_400), .A2(n_377), .B1(n_308), .B2(n_310), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_456), .A2(n_454), .B1(n_416), .B2(n_423), .Y(n_457) );
INVxp67_ASAP7_75t_L g458 ( .A(n_417), .Y(n_458) );
AOI221xp5_ASAP7_75t_L g459 ( .A1(n_453), .A2(n_456), .B1(n_412), .B2(n_414), .C(n_450), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_452), .A2(n_433), .B(n_451), .Y(n_460) );
NOR2x1_ASAP7_75t_SL g461 ( .A(n_448), .B(n_455), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_446), .Y(n_462) );
NOR3xp33_ASAP7_75t_L g463 ( .A(n_420), .B(n_447), .C(n_445), .Y(n_463) );
AOI221xp5_ASAP7_75t_L g464 ( .A1(n_411), .A2(n_424), .B1(n_415), .B2(n_407), .C(n_408), .Y(n_464) );
NOR3xp33_ASAP7_75t_L g465 ( .A(n_420), .B(n_425), .C(n_419), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_409), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_L g467 ( .A1(n_438), .A2(n_442), .B(n_422), .C(n_421), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_410), .B(n_413), .Y(n_468) );
XOR2x2_ASAP7_75t_L g469 ( .A(n_437), .B(n_428), .Y(n_469) );
AOI211xp5_ASAP7_75t_SL g470 ( .A1(n_459), .A2(n_429), .B(n_434), .C(n_427), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_461), .Y(n_471) );
INVx2_ASAP7_75t_SL g472 ( .A(n_466), .Y(n_472) );
AOI221xp5_ASAP7_75t_L g473 ( .A1(n_457), .A2(n_430), .B1(n_439), .B2(n_431), .C(n_418), .Y(n_473) );
NOR2x2_ASAP7_75t_L g474 ( .A(n_469), .B(n_444), .Y(n_474) );
OAI211xp5_ASAP7_75t_L g475 ( .A1(n_460), .A2(n_443), .B(n_432), .C(n_435), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_462), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_463), .A2(n_441), .B1(n_440), .B2(n_439), .Y(n_477) );
NAND5xp2_ASAP7_75t_L g478 ( .A(n_470), .B(n_465), .C(n_467), .D(n_464), .E(n_436), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_472), .B(n_471), .Y(n_479) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_476), .Y(n_480) );
NAND3xp33_ASAP7_75t_SL g481 ( .A(n_470), .B(n_458), .C(n_468), .Y(n_481) );
NOR3xp33_ASAP7_75t_L g482 ( .A(n_475), .B(n_426), .C(n_449), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_480), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_479), .Y(n_484) );
XNOR2xp5_ASAP7_75t_L g485 ( .A(n_481), .B(n_477), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_485), .A2(n_482), .B1(n_473), .B2(n_478), .Y(n_486) );
XNOR2x1_ASAP7_75t_L g487 ( .A(n_484), .B(n_474), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_487), .Y(n_488) );
INVx2_ASAP7_75t_SL g489 ( .A(n_486), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_489), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_490), .B(n_483), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_491), .A2(n_488), .B(n_483), .Y(n_492) );
endmodule