module fake_jpeg_7997_n_303 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_303);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_303;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_152;
wire n_73;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_228;
wire n_178;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx3_ASAP7_75t_SL g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_7),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_0),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_52),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_23),
.Y(n_49)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_57),
.Y(n_70)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_34),
.A2(n_17),
.B1(n_33),
.B2(n_22),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_58),
.A2(n_32),
.B1(n_19),
.B2(n_16),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_59),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_33),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_42),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_35),
.A2(n_18),
.B1(n_27),
.B2(n_17),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_18),
.B1(n_27),
.B2(n_33),
.Y(n_68)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_63),
.B(n_65),
.Y(n_114)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_45),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_68),
.A2(n_81),
.B1(n_87),
.B2(n_28),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_45),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_69),
.B(n_76),
.Y(n_99)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_72),
.A2(n_20),
.B1(n_31),
.B2(n_30),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_59),
.Y(n_76)
);

AO22x1_ASAP7_75t_L g77 ( 
.A1(n_44),
.A2(n_42),
.B1(n_35),
.B2(n_39),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_77),
.A2(n_80),
.B1(n_55),
.B2(n_24),
.Y(n_112)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_44),
.A2(n_42),
.B1(n_35),
.B2(n_39),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_48),
.A2(n_23),
.B1(n_29),
.B2(n_22),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_52),
.A2(n_29),
.B1(n_28),
.B2(n_32),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_24),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_50),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_89),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_60),
.A2(n_42),
.B1(n_35),
.B2(n_20),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_90),
.A2(n_47),
.B1(n_25),
.B2(n_19),
.Y(n_106)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_43),
.C(n_60),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_70),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_104),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_56),
.C(n_53),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_51),
.C(n_47),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_103),
.B(n_118),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_46),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_106),
.A2(n_117),
.B1(n_120),
.B2(n_20),
.Y(n_150)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_115),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_85),
.A2(n_47),
.B1(n_46),
.B2(n_55),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_74),
.B1(n_91),
.B2(n_79),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_92),
.B1(n_63),
.B2(n_78),
.Y(n_137)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_30),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_90),
.A2(n_25),
.B1(n_21),
.B2(n_16),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_119),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_104),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_141),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_124),
.B(n_125),
.Y(n_158)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_126),
.B(n_127),
.Y(n_161)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_133),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_102),
.B(n_79),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_131),
.B(n_9),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_96),
.A2(n_75),
.B(n_24),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_132),
.A2(n_143),
.B(n_146),
.Y(n_171)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

AO21x1_ASAP7_75t_L g178 ( 
.A1(n_135),
.A2(n_138),
.B(n_147),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

INVxp33_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

AO22x1_ASAP7_75t_L g180 ( 
.A1(n_137),
.A2(n_113),
.B1(n_24),
.B2(n_20),
.Y(n_180)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_96),
.A2(n_92),
.B1(n_84),
.B2(n_74),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_140),
.A2(n_142),
.B1(n_145),
.B2(n_150),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_80),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_82),
.B1(n_83),
.B2(n_77),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_107),
.A2(n_24),
.B(n_30),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_93),
.B(n_77),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_100),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_71),
.B1(n_64),
.B2(n_55),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_24),
.B(n_31),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_149),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_127),
.A2(n_118),
.B1(n_102),
.B2(n_109),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_152),
.A2(n_164),
.B1(n_176),
.B2(n_30),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

AND2x6_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_97),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_154),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_155),
.B(n_143),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_100),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_162),
.Y(n_186)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_73),
.B(n_11),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_159),
.A2(n_170),
.B(n_9),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_123),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_128),
.A2(n_108),
.B1(n_94),
.B2(n_111),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_131),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_166),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_108),
.Y(n_169)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_132),
.A2(n_105),
.B(n_94),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_129),
.Y(n_172)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_172),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_122),
.B(n_31),
.Y(n_173)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

CKINVDCx12_ASAP7_75t_R g174 ( 
.A(n_133),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_174),
.B(n_182),
.Y(n_187)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_137),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_135),
.A2(n_138),
.B1(n_147),
.B2(n_130),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_122),
.B(n_31),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_146),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_124),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_179),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_180),
.A2(n_181),
.B1(n_105),
.B2(n_125),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_134),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_183),
.A2(n_189),
.B(n_199),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_190),
.C(n_195),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_157),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_171),
.A2(n_156),
.B(n_169),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_148),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_194),
.A2(n_196),
.B1(n_198),
.B2(n_200),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_148),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_175),
.A2(n_130),
.B1(n_150),
.B2(n_137),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_151),
.B(n_126),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_204),
.C(n_205),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_163),
.B1(n_165),
.B2(n_158),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_171),
.A2(n_137),
.B(n_113),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_176),
.A2(n_30),
.B1(n_1),
.B2(n_2),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_201),
.A2(n_203),
.B1(n_165),
.B2(n_168),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_155),
.A2(n_0),
.B(n_1),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_151),
.B(n_7),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_162),
.B(n_0),
.C(n_2),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_209),
.B(n_182),
.Y(n_225)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_212),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_186),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_207),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_214),
.A2(n_226),
.B1(n_230),
.B2(n_231),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_187),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_224),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_188),
.Y(n_233)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_203),
.Y(n_217)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_218),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_192),
.A2(n_152),
.B1(n_158),
.B2(n_164),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_219),
.A2(n_183),
.B1(n_165),
.B2(n_168),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_172),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_220),
.A2(n_222),
.B(n_180),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_184),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_160),
.C(n_154),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_209),
.C(n_195),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_202),
.B(n_166),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_225),
.Y(n_242)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_189),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_161),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_227),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_228),
.A2(n_180),
.B1(n_167),
.B2(n_178),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_194),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_183),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_174),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_232),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_233),
.B(n_216),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_235),
.C(n_243),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_185),
.C(n_208),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_238),
.A2(n_249),
.B1(n_227),
.B2(n_219),
.Y(n_254)
);

FAx1_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_200),
.CI(n_199),
.CON(n_240),
.SN(n_240)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_240),
.A2(n_226),
.B(n_213),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_170),
.C(n_204),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_205),
.C(n_167),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_221),
.C(n_220),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_246),
.A2(n_218),
.B1(n_217),
.B2(n_229),
.Y(n_253)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_247),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_231),
.A2(n_178),
.B1(n_10),
.B2(n_11),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_242),
.B(n_220),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_259),
.Y(n_268)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_253),
.Y(n_265)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_254),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_214),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_255),
.Y(n_270)
);

OAI321xp33_ASAP7_75t_L g269 ( 
.A1(n_256),
.A2(n_240),
.A3(n_222),
.B1(n_245),
.B2(n_234),
.C(n_243),
.Y(n_269)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_241),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_260),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_239),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_249),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_261),
.A2(n_250),
.B1(n_233),
.B2(n_237),
.Y(n_266)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_238),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_263),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_248),
.A2(n_222),
.B1(n_178),
.B2(n_221),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_264),
.A2(n_240),
.B1(n_235),
.B2(n_11),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_272),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_256),
.A2(n_246),
.B1(n_244),
.B2(n_247),
.Y(n_267)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_267),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_269),
.A2(n_258),
.B(n_6),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_251),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_273),
.B(n_264),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_257),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_261),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_277),
.B(n_278),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_268),
.Y(n_278)
);

OA21x2_ASAP7_75t_SL g280 ( 
.A1(n_272),
.A2(n_263),
.B(n_258),
.Y(n_280)
);

AOI322xp5_ASAP7_75t_L g288 ( 
.A1(n_280),
.A2(n_265),
.A3(n_275),
.B1(n_274),
.B2(n_266),
.C1(n_271),
.C2(n_273),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_271),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_282),
.A2(n_13),
.B(n_15),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_6),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_283),
.B(n_284),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_6),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_2),
.C(n_3),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_4),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_292),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_288),
.B(n_289),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_15),
.C(n_12),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_286),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_294),
.A2(n_296),
.B(n_295),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_290),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_298),
.A2(n_299),
.B(n_285),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_279),
.C(n_290),
.Y(n_299)
);

O2A1O1Ixp33_ASAP7_75t_L g301 ( 
.A1(n_300),
.A2(n_281),
.B(n_286),
.C(n_291),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_301),
.A2(n_13),
.B1(n_4),
.B2(n_5),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_302),
.A2(n_4),
.B1(n_5),
.B2(n_260),
.Y(n_303)
);


endmodule