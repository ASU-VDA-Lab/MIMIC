module real_jpeg_13479_n_17 (n_5, n_4, n_8, n_0, n_12, n_337, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_337;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_5),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_5),
.A2(n_63),
.B1(n_64),
.B2(n_79),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_5),
.A2(n_53),
.B1(n_54),
.B2(n_79),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_79),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_6),
.A2(n_63),
.B1(n_64),
.B2(n_160),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_6),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_6),
.B(n_54),
.C(n_67),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_6),
.B(n_88),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_6),
.A2(n_123),
.B(n_176),
.Y(n_192)
);

O2A1O1Ixp33_ASAP7_75t_L g202 ( 
.A1(n_6),
.A2(n_23),
.B(n_87),
.C(n_203),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_160),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_6),
.B(n_21),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_6),
.B(n_30),
.Y(n_247)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_7),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_8),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_8),
.A2(n_30),
.B1(n_31),
.B2(n_90),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_8),
.A2(n_63),
.B1(n_64),
.B2(n_90),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_8),
.A2(n_53),
.B1(n_54),
.B2(n_90),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_9),
.A2(n_30),
.B1(n_31),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_9),
.A2(n_38),
.B1(n_63),
.B2(n_64),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_38),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_9),
.A2(n_38),
.B1(n_53),
.B2(n_54),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_22)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_10),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

NAND2xp33_ASAP7_75t_SL g260 ( 
.A(n_10),
.B(n_24),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_11),
.A2(n_63),
.B1(n_64),
.B2(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_11),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_11),
.A2(n_53),
.B1(n_54),
.B2(n_172),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_11),
.A2(n_23),
.B1(n_24),
.B2(n_172),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_172),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_12),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_12),
.A2(n_23),
.B1(n_24),
.B2(n_62),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_12),
.A2(n_30),
.B1(n_31),
.B2(n_62),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_12),
.A2(n_53),
.B1(n_54),
.B2(n_62),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_13),
.A2(n_34),
.B1(n_53),
.B2(n_54),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_13),
.A2(n_34),
.B1(n_63),
.B2(n_64),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_13),
.A2(n_23),
.B1(n_24),
.B2(n_34),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_14),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_14),
.A2(n_23),
.B1(n_24),
.B2(n_75),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_14),
.A2(n_53),
.B1(n_54),
.B2(n_75),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_14),
.A2(n_63),
.B1(n_64),
.B2(n_75),
.Y(n_253)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_16),
.A2(n_30),
.B1(n_31),
.B2(n_132),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_16),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_16),
.A2(n_53),
.B1(n_54),
.B2(n_132),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_16),
.A2(n_63),
.B1(n_64),
.B2(n_132),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_16),
.A2(n_23),
.B1(n_24),
.B2(n_132),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_41),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_39),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_35),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_27),
.B(n_33),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_21),
.A2(n_27),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_21),
.A2(n_27),
.B1(n_37),
.B2(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_22),
.B(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_22),
.A2(n_74),
.B(n_76),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_22),
.A2(n_28),
.B1(n_74),
.B2(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_22),
.B(n_78),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_22),
.A2(n_28),
.B1(n_108),
.B2(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_22),
.A2(n_76),
.B(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_22),
.A2(n_28),
.B1(n_131),
.B2(n_274),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_23),
.A2(n_24),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

AOI32xp33_ASAP7_75t_L g259 ( 
.A1(n_23),
.A2(n_26),
.A3(n_31),
.B1(n_247),
.B2(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_27),
.B(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_28),
.A2(n_131),
.B(n_133),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g245 ( 
.A1(n_28),
.A2(n_31),
.B(n_160),
.C(n_246),
.Y(n_245)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_35),
.B(n_335),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_36),
.B(n_332),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_331),
.B(n_333),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_319),
.B(n_330),
.Y(n_42)
);

AO21x1_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_148),
.B(n_316),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_135),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_110),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_46),
.B(n_110),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_80),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_47),
.B(n_81),
.C(n_96),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_51),
.B(n_73),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_48),
.A2(n_49),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_59),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_50),
.A2(n_51),
.B1(n_73),
.B2(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_50),
.A2(n_51),
.B1(n_59),
.B2(n_60),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_56),
.B(n_57),
.Y(n_51)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_52),
.A2(n_56),
.B1(n_181),
.B2(n_183),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_52),
.B(n_177),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_52),
.A2(n_56),
.B1(n_122),
.B2(n_264),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_54),
.B1(n_67),
.B2(n_68),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_53),
.B(n_194),
.Y(n_193)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_56),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_56),
.B(n_177),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_58),
.A2(n_121),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_65),
.B1(n_70),
.B2(n_72),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_61),
.A2(n_65),
.B1(n_72),
.B2(n_127),
.Y(n_126)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_64),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

AO22x1_ASAP7_75t_SL g88 ( 
.A1(n_63),
.A2(n_64),
.B1(n_86),
.B2(n_87),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_63),
.B(n_164),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g203 ( 
.A1(n_64),
.A2(n_86),
.B(n_160),
.Y(n_203)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_65),
.A2(n_72),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_65),
.B(n_162),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_65),
.A2(n_72),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_65),
.A2(n_72),
.B1(n_127),
.B2(n_253),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_69),
.A2(n_71),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_69),
.A2(n_171),
.B(n_173),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_69),
.B(n_160),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_69),
.A2(n_173),
.B(n_252),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_72),
.B(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_96),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_81),
.A2(n_82),
.B(n_93),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_93),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_89),
.B1(n_91),
.B2(n_92),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_83),
.A2(n_89),
.B1(n_91),
.B2(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_83),
.A2(n_91),
.B1(n_101),
.B2(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_83),
.A2(n_208),
.B(n_209),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_83),
.A2(n_91),
.B1(n_223),
.B2(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_83),
.A2(n_209),
.B(n_250),
.Y(n_272)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_88),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_84),
.B(n_210),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_84),
.A2(n_88),
.B(n_323),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_88),
.B(n_210),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_91),
.A2(n_223),
.B(n_224),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_91),
.A2(n_129),
.B(n_224),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_94),
.A2(n_159),
.B(n_161),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_94),
.A2(n_161),
.B(n_235),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_106),
.B1(n_107),
.B2(n_109),
.Y(n_96)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_98),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_SL g146 ( 
.A(n_98),
.B(n_103),
.C(n_107),
.Y(n_146)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_102),
.A2(n_103),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_103),
.B(n_140),
.C(n_144),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_107),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_107),
.B(n_139),
.C(n_146),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_116),
.C(n_117),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_111),
.A2(n_112),
.B1(n_116),
.B2(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_116),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_117),
.B(n_313),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_128),
.C(n_130),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_118),
.A2(n_119),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_125),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_120),
.A2(n_125),
.B1(n_126),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_120),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_123),
.A2(n_175),
.B(n_176),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_123),
.A2(n_124),
.B1(n_205),
.B2(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_123),
.A2(n_124),
.B1(n_230),
.B2(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_124),
.A2(n_182),
.B(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_124),
.B(n_160),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_124),
.A2(n_190),
.B(n_205),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_128),
.B(n_130),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_134),
.B(n_245),
.Y(n_244)
);

OAI21xp33_ASAP7_75t_L g316 ( 
.A1(n_135),
.A2(n_317),
.B(n_318),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_147),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_136),
.B(n_147),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_146),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_141),
.Y(n_325)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_145),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_310),
.B(n_315),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_298),
.B(n_309),
.Y(n_149)
);

OAI321xp33_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_266),
.A3(n_291),
.B1(n_296),
.B2(n_297),
.C(n_337),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_239),
.B(n_265),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_217),
.B(n_238),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_198),
.B(n_216),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_178),
.B(n_197),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_165),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_156),
.B(n_165),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_163),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_157),
.A2(n_158),
.B1(n_163),
.B2(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_163),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_174),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_170),
.C(n_174),
.Y(n_199)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_171),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_175),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_186),
.B(n_196),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_184),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_180),
.B(n_184),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_191),
.B(n_195),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_188),
.B(n_189),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_199),
.B(n_200),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_206),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_211),
.C(n_215),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_204),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_211),
.B1(n_214),
.B2(n_215),
.Y(n_206)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_207),
.Y(n_215)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_213),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_218),
.B(n_219),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_231),
.B2(n_232),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_234),
.C(n_236),
.Y(n_240)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_225),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_226),
.C(n_229),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_236),
.B2(n_237),
.Y(n_232)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_233),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_234),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_240),
.B(n_241),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_255),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_242),
.B(n_256),
.C(n_257),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_248),
.B2(n_254),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_243),
.B(n_249),
.C(n_251),
.Y(n_280)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_248),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_261),
.B2(n_262),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_262),
.Y(n_276)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_281),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_267),
.B(n_281),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_277),
.C(n_280),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_268),
.A2(n_269),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_276),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_273),
.B2(n_275),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_275),
.C(n_276),
.Y(n_290)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_273),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_277),
.B(n_280),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_279),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_290),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_285),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_283),
.B(n_285),
.C(n_290),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_289),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_288),
.C(n_289),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_292),
.B(n_293),
.Y(n_296)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_308),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_308),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_303),
.C(n_304),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_304),
.B2(n_305),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_312),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_329),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_329),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_328),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_324),
.B1(n_326),
.B2(n_327),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_322),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_324),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_326),
.C(n_328),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_332),
.Y(n_335)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);


endmodule