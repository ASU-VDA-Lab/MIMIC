module fake_jpeg_854_n_144 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_144);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_24),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_13),
.C(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_58),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_52),
.B(n_0),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_59),
.A2(n_50),
.B1(n_51),
.B2(n_45),
.Y(n_62)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_69),
.Y(n_72)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_63),
.Y(n_80)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_57),
.A2(n_43),
.B1(n_40),
.B2(n_45),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_57),
.B1(n_56),
.B2(n_43),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_64),
.B(n_58),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_73),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_51),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_50),
.C(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_59),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_78),
.A2(n_61),
.B1(n_42),
.B2(n_41),
.Y(n_85)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_42),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_82),
.B(n_0),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_41),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_1),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_85),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_SL g86 ( 
.A1(n_73),
.A2(n_46),
.B(n_44),
.C(n_39),
.Y(n_86)
);

AO22x1_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_96),
.B1(n_81),
.B2(n_75),
.Y(n_101)
);

NOR2x1_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_38),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_94),
.Y(n_113)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_49),
.B(n_34),
.C(n_33),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_4),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_82),
.A2(n_49),
.B1(n_2),
.B2(n_3),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_98),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_99),
.B(n_74),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_101),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_75),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_110),
.C(n_106),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_90),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_105),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_104),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_108),
.Y(n_127)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_109),
.B(n_111),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_14),
.C(n_28),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_86),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_115),
.Y(n_122)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_117),
.B(n_126),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_107),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_121),
.Y(n_130)
);

OAI32xp33_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_113),
.A3(n_101),
.B1(n_116),
.B2(n_110),
.Y(n_124)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

AOI22x1_ASAP7_75t_L g125 ( 
.A1(n_116),
.A2(n_17),
.B1(n_25),
.B2(n_23),
.Y(n_125)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_114),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_126)
);

OAI21x1_ASAP7_75t_L g131 ( 
.A1(n_118),
.A2(n_9),
.B(n_10),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_128),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_117),
.C(n_119),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_132),
.C(n_122),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_135),
.A2(n_136),
.B1(n_128),
.B2(n_123),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_130),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_138),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_133),
.B1(n_127),
.B2(n_122),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_125),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_20),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_29),
.C(n_10),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_11),
.Y(n_144)
);


endmodule