module fake_jpeg_17066_n_348 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_348);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_348;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_45),
.Y(n_51)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_0),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_33),
.Y(n_56)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_22),
.Y(n_62)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_25),
.B1(n_19),
.B2(n_29),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_52),
.A2(n_65),
.B1(n_35),
.B2(n_33),
.Y(n_97)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_35),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_56),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_29),
.B(n_2),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_59),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_72),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_16),
.B(n_26),
.Y(n_59)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_62),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_25),
.B1(n_19),
.B2(n_29),
.Y(n_65)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_32),
.Y(n_71)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_35),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_20),
.Y(n_101)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_80),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_25),
.B1(n_47),
.B2(n_45),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_82),
.A2(n_68),
.B1(n_53),
.B2(n_21),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_55),
.C(n_76),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_84),
.B(n_70),
.Y(n_136)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_56),
.A2(n_25),
.B1(n_46),
.B2(n_26),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_88),
.A2(n_91),
.B1(n_24),
.B2(n_53),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_56),
.A2(n_16),
.B1(n_26),
.B2(n_24),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_51),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_102),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_95),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_97),
.A2(n_109),
.B1(n_93),
.B2(n_18),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_75),
.A2(n_17),
.B1(n_18),
.B2(n_32),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_104),
.B1(n_21),
.B2(n_20),
.Y(n_121)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_101),
.B(n_110),
.Y(n_119)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_105),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_69),
.A2(n_17),
.B1(n_18),
.B2(n_32),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_106),
.B(n_107),
.Y(n_145)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_63),
.B(n_16),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_63),
.B(n_17),
.Y(n_111)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_112),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_74),
.A2(n_34),
.B1(n_30),
.B2(n_28),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_L g118 ( 
.A1(n_113),
.A2(n_74),
.B1(n_70),
.B2(n_68),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_114),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_118),
.A2(n_141),
.B1(n_89),
.B2(n_114),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_98),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_126),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_137),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_69),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_133),
.Y(n_147)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_78),
.Y(n_125)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_125),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_134),
.Y(n_164)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_90),
.B(n_23),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_78),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_45),
.C(n_64),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_139),
.A2(n_135),
.B1(n_133),
.B2(n_137),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_140),
.B(n_99),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_90),
.A2(n_68),
.B1(n_53),
.B2(n_21),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_87),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_142),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_146),
.A2(n_151),
.B1(n_154),
.B2(n_173),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_92),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_149),
.B(n_170),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_165),
.C(n_149),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_130),
.A2(n_89),
.B1(n_83),
.B2(n_86),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_152),
.A2(n_158),
.B1(n_30),
.B2(n_31),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_141),
.A2(n_83),
.B(n_112),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_156),
.A2(n_27),
.B(n_143),
.Y(n_212)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_157),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_130),
.A2(n_86),
.B1(n_79),
.B2(n_33),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_124),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_159),
.B(n_160),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_119),
.B(n_104),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_124),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_162),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_127),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_122),
.B(n_135),
.C(n_129),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_127),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_177),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_67),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_167),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_126),
.A2(n_82),
.B1(n_113),
.B2(n_54),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_168),
.A2(n_178),
.B1(n_142),
.B2(n_128),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_144),
.A2(n_82),
.B1(n_23),
.B2(n_27),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_169),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_120),
.B(n_82),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_121),
.A2(n_23),
.B1(n_54),
.B2(n_80),
.Y(n_173)
);

OAI22x1_ASAP7_75t_SL g174 ( 
.A1(n_115),
.A2(n_27),
.B1(n_22),
.B2(n_28),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_174),
.A2(n_175),
.B1(n_180),
.B2(n_27),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_116),
.A2(n_54),
.B1(n_95),
.B2(n_12),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_145),
.A2(n_22),
.B(n_31),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_176),
.A2(n_31),
.B(n_28),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_116),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_117),
.A2(n_30),
.B1(n_28),
.B2(n_64),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_117),
.A2(n_10),
.B1(n_14),
.B2(n_11),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_181),
.B(n_200),
.C(n_206),
.Y(n_226)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_170),
.A2(n_115),
.B(n_123),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_183),
.A2(n_197),
.B(n_203),
.Y(n_233)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_153),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_194),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_150),
.B(n_134),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_189),
.B(n_210),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_154),
.A2(n_156),
.B1(n_151),
.B2(n_169),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_190),
.A2(n_191),
.B1(n_207),
.B2(n_213),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_155),
.A2(n_146),
.B1(n_147),
.B2(n_168),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_192),
.A2(n_209),
.B1(n_196),
.B2(n_195),
.Y(n_220)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_193),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_153),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_155),
.A2(n_78),
.B(n_2),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_205),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_199),
.A2(n_159),
.B(n_161),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_147),
.B(n_165),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_155),
.A2(n_1),
.B(n_2),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_157),
.B(n_125),
.Y(n_204)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_204),
.Y(n_236)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_162),
.B(n_67),
.C(n_143),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_174),
.A2(n_132),
.B1(n_143),
.B2(n_10),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_172),
.Y(n_208)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_31),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_166),
.Y(n_211)
);

NOR3xp33_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_30),
.C(n_3),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_178),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_214),
.B(n_175),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_177),
.Y(n_216)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_218),
.A2(n_197),
.B1(n_199),
.B2(n_205),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_220),
.A2(n_224),
.B1(n_229),
.B2(n_237),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_184),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_223),
.B(n_8),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_192),
.A2(n_179),
.B1(n_173),
.B2(n_171),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_160),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_231),
.C(n_243),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_211),
.Y(n_228)
);

INVx3_ASAP7_75t_SL g263 ( 
.A(n_228),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_181),
.B(n_180),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_191),
.A2(n_179),
.B1(n_171),
.B2(n_30),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_232),
.A2(n_188),
.B1(n_186),
.B2(n_182),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_207),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_195),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_237)
);

MAJx2_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_8),
.C(n_11),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_238),
.B(n_206),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_190),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_239),
.A2(n_240),
.B1(n_237),
.B2(n_224),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_202),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_202),
.B(n_183),
.C(n_210),
.Y(n_243)
);

NAND2x1p5_ASAP7_75t_R g245 ( 
.A(n_233),
.B(n_203),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_245),
.B(n_14),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_201),
.Y(n_246)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_246),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_212),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_256),
.C(n_260),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_248),
.B(n_262),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_222),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_267),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_215),
.Y(n_251)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_251),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_252),
.A2(n_227),
.B1(n_220),
.B2(n_239),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_215),
.Y(n_253)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_253),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_255),
.B(n_225),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_208),
.C(n_193),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_230),
.Y(n_257)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_217),
.Y(n_258)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_258),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_259),
.B(n_261),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_185),
.C(n_198),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_8),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_268),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_5),
.C(n_6),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_266),
.C(n_14),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_5),
.C(n_6),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_7),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_218),
.B(n_7),
.Y(n_268)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_269),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_244),
.A2(n_227),
.B1(n_219),
.B2(n_243),
.Y(n_271)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_271),
.Y(n_298)
);

XNOR2x1_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_233),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_274),
.A2(n_278),
.B1(n_267),
.B2(n_265),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_254),
.C(n_260),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_244),
.A2(n_219),
.B1(n_232),
.B2(n_221),
.Y(n_277)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_277),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_268),
.A2(n_240),
.B1(n_238),
.B2(n_7),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_246),
.B(n_9),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_284),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_255),
.B(n_10),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_288),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_287),
.B(n_278),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_250),
.A2(n_257),
.B1(n_263),
.B2(n_249),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_289),
.A2(n_277),
.B(n_269),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_290),
.B(n_295),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_263),
.Y(n_291)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_291),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_256),
.C(n_254),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_279),
.C(n_275),
.Y(n_312)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_276),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_282),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_259),
.Y(n_296)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_296),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_274),
.A2(n_247),
.B(n_266),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_297),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_270),
.A2(n_273),
.B1(n_283),
.B2(n_289),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_299),
.Y(n_318)
);

NOR3xp33_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_281),
.C(n_287),
.Y(n_303)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_303),
.Y(n_314)
);

AO22x1_ASAP7_75t_L g316 ( 
.A1(n_304),
.A2(n_285),
.B1(n_294),
.B2(n_298),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_305),
.B(n_295),
.Y(n_317)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_306),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_286),
.Y(n_308)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_308),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_271),
.Y(n_310)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_310),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_290),
.C(n_297),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_301),
.B(n_288),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_315),
.B(n_302),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_319),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_304),
.C(n_300),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_299),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_314),
.A2(n_298),
.B(n_292),
.Y(n_320)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_320),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_321),
.B(n_308),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_323),
.B(n_324),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_312),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_302),
.C(n_310),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_329),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_322),
.B(n_318),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_327),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_333),
.A2(n_319),
.B(n_307),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_326),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_334),
.A2(n_336),
.B(n_328),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_326),
.A2(n_309),
.B(n_318),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_337),
.B(n_338),
.C(n_339),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_334),
.B(n_313),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_340),
.B(n_341),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_335),
.A2(n_325),
.B1(n_321),
.B2(n_316),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_343),
.Y(n_344)
);

BUFx24_ASAP7_75t_SL g345 ( 
.A(n_344),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_345),
.Y(n_346)
);

OAI211xp5_ASAP7_75t_L g347 ( 
.A1(n_346),
.A2(n_342),
.B(n_330),
.C(n_331),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_338),
.Y(n_348)
);


endmodule