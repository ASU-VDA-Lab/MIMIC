module fake_jpeg_13087_n_402 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_402);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_402;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_48),
.Y(n_128)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_49),
.Y(n_138)
);

INVx5_ASAP7_75t_SL g50 ( 
.A(n_42),
.Y(n_50)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_50),
.Y(n_130)
);

BUFx24_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx11_ASAP7_75t_L g139 ( 
.A(n_51),
.Y(n_139)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_42),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g143 ( 
.A(n_52),
.Y(n_143)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_55),
.Y(n_129)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_16),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_59),
.B(n_81),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

BUFx24_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_31),
.B(n_15),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_65),
.B(n_75),
.Y(n_116)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_67),
.Y(n_132)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_70),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_72),
.Y(n_147)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_73),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_74),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_31),
.B(n_14),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

BUFx4f_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_79),
.Y(n_145)
);

BUFx4f_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_80),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_93),
.Y(n_94)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_85),
.Y(n_101)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_84),
.A2(n_27),
.B1(n_33),
.B2(n_35),
.Y(n_110)
);

BUFx12f_ASAP7_75t_SL g85 ( 
.A(n_47),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_47),
.A2(n_38),
.B1(n_32),
.B2(n_28),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_27),
.B1(n_35),
.B2(n_33),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_18),
.B(n_14),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_89),
.Y(n_103)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_88),
.B(n_29),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_18),
.B(n_26),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_19),
.B(n_14),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_91),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_19),
.B(n_13),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_25),
.B(n_0),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_26),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_62),
.C(n_38),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_95),
.B(n_142),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_61),
.A2(n_38),
.B1(n_27),
.B2(n_44),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_97),
.A2(n_93),
.B1(n_77),
.B2(n_82),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_62),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_107),
.B(n_0),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_108),
.A2(n_121),
.B1(n_125),
.B2(n_60),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_110),
.A2(n_74),
.B1(n_80),
.B2(n_60),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_111),
.B(n_119),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_25),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_113),
.B(n_133),
.Y(n_160)
);

O2A1O1Ixp33_ASAP7_75t_SL g115 ( 
.A1(n_50),
.A2(n_46),
.B(n_43),
.C(n_40),
.Y(n_115)
);

AO22x1_ASAP7_75t_L g155 ( 
.A1(n_115),
.A2(n_59),
.B1(n_52),
.B2(n_36),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_71),
.B(n_46),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_57),
.A2(n_35),
.B1(n_33),
.B2(n_45),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_51),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_122),
.B(n_126),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_L g125 ( 
.A1(n_67),
.A2(n_21),
.B1(n_44),
.B2(n_41),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_88),
.B(n_43),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_55),
.B(n_34),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_51),
.A2(n_45),
.B1(n_41),
.B2(n_23),
.Y(n_135)
);

XNOR2x1_ASAP7_75t_SL g178 ( 
.A(n_135),
.B(n_0),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_66),
.B(n_36),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_136),
.B(n_141),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_73),
.B(n_34),
.Y(n_141)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_145),
.Y(n_148)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_143),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_149),
.B(n_175),
.Y(n_202)
);

OAI21xp33_ASAP7_75t_L g150 ( 
.A1(n_101),
.A2(n_30),
.B(n_40),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_L g211 ( 
.A1(n_150),
.A2(n_155),
.B(n_178),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_104),
.B(n_21),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_186),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_130),
.A2(n_23),
.B1(n_29),
.B2(n_76),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_154),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_156),
.A2(n_158),
.B1(n_181),
.B2(n_184),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_130),
.A2(n_84),
.B1(n_30),
.B2(n_143),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_157),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_95),
.A2(n_97),
.B1(n_94),
.B2(n_110),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_118),
.Y(n_164)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_164),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_165),
.A2(n_168),
.B1(n_139),
.B2(n_102),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_144),
.A2(n_140),
.B1(n_147),
.B2(n_127),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_115),
.A2(n_135),
.B1(n_125),
.B2(n_105),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_169),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_177),
.Y(n_203)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_140),
.A2(n_54),
.B1(n_1),
.B2(n_2),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_173),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_106),
.Y(n_174)
);

INVx11_ASAP7_75t_L g214 ( 
.A(n_174),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_134),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_176),
.Y(n_215)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_137),
.Y(n_177)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_114),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_179),
.Y(n_198)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_117),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_180),
.B(n_182),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_132),
.A2(n_105),
.B1(n_100),
.B2(n_103),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_117),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_100),
.A2(n_54),
.B1(n_2),
.B2(n_3),
.Y(n_184)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_114),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_185),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_134),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_187),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_149),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_138),
.C(n_123),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_189),
.B(n_193),
.C(n_222),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_158),
.A2(n_159),
.B1(n_186),
.B2(n_175),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_192),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_153),
.B(n_138),
.C(n_123),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_200),
.A2(n_210),
.B1(n_182),
.B2(n_180),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_209),
.B(n_164),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_155),
.A2(n_146),
.B1(n_147),
.B2(n_127),
.Y(n_210)
);

OAI32xp33_ASAP7_75t_L g212 ( 
.A1(n_160),
.A2(n_116),
.A3(n_139),
.B1(n_146),
.B2(n_96),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_129),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_99),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_218),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_99),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_153),
.B(n_120),
.C(n_124),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_160),
.B(n_120),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_223),
.B(n_3),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_178),
.A2(n_129),
.B1(n_124),
.B2(n_98),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_224),
.Y(n_253)
);

OAI32xp33_ASAP7_75t_L g225 ( 
.A1(n_205),
.A2(n_166),
.A3(n_155),
.B1(n_151),
.B2(n_162),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_225),
.B(n_242),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_213),
.A2(n_187),
.B1(n_174),
.B2(n_185),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_226),
.A2(n_229),
.B1(n_233),
.B2(n_252),
.Y(n_255)
);

OA21x2_ASAP7_75t_L g227 ( 
.A1(n_200),
.A2(n_203),
.B(n_170),
.Y(n_227)
);

OA21x2_ASAP7_75t_L g280 ( 
.A1(n_227),
.A2(n_214),
.B(n_204),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_228),
.B(n_236),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_203),
.A2(n_156),
.B1(n_181),
.B2(n_184),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_230),
.B(n_232),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_203),
.A2(n_148),
.B1(n_171),
.B2(n_169),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_197),
.A2(n_163),
.B1(n_154),
.B2(n_161),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_234),
.A2(n_238),
.B1(n_199),
.B2(n_201),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_177),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_219),
.Y(n_237)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

OAI22x1_ASAP7_75t_SL g238 ( 
.A1(n_197),
.A2(n_98),
.B1(n_179),
.B2(n_176),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_187),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_239),
.B(n_240),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_174),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_96),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_243),
.B(n_244),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_191),
.B(n_112),
.Y(n_244)
);

BUFx12_ASAP7_75t_L g245 ( 
.A(n_214),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_245),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_191),
.B(n_124),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_248),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_190),
.A2(n_117),
.B(n_5),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_247),
.A2(n_221),
.B(n_201),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_202),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_206),
.Y(n_249)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_249),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_112),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_207),
.Y(n_267)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_196),
.Y(n_251)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_251),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_205),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_196),
.Y(n_254)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_254),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_231),
.C(n_222),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_235),
.C(n_248),
.Y(n_286)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_249),
.Y(n_260)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_260),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_229),
.A2(n_224),
.B1(n_202),
.B2(n_194),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_267),
.Y(n_281)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_266),
.Y(n_292)
);

AND2x6_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_211),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_SL g293 ( 
.A(n_270),
.B(n_225),
.C(n_227),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_228),
.B(n_198),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_271),
.B(n_272),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_198),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_229),
.A2(n_189),
.B1(n_193),
.B2(n_212),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_276),
.Y(n_291)
);

AO22x1_ASAP7_75t_L g295 ( 
.A1(n_274),
.A2(n_247),
.B1(n_227),
.B2(n_254),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_241),
.A2(n_221),
.B1(n_220),
.B2(n_216),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_231),
.A2(n_221),
.B1(n_220),
.B2(n_207),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_242),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_227),
.A2(n_195),
.B1(n_216),
.B2(n_206),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_278),
.A2(n_240),
.B1(n_239),
.B2(n_233),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_280),
.A2(n_230),
.B(n_252),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_235),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_283),
.B(n_286),
.C(n_289),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_271),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_284),
.B(n_285),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_236),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_287),
.A2(n_300),
.B1(n_280),
.B2(n_274),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_267),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_294),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_244),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_253),
.C(n_243),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_290),
.B(n_298),
.C(n_301),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_293),
.B(n_280),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_277),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_302),
.B(n_279),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_261),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_264),
.B(n_237),
.C(n_251),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_257),
.Y(n_299)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_299),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_278),
.A2(n_238),
.B1(n_234),
.B2(n_247),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_238),
.C(n_250),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_226),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_303),
.B(n_262),
.Y(n_305)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_257),
.Y(n_304)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_304),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_305),
.B(n_320),
.Y(n_331)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_306),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_301),
.A2(n_279),
.B1(n_255),
.B2(n_276),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_307),
.A2(n_322),
.B(n_295),
.Y(n_333)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_282),
.Y(n_308)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_308),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_259),
.Y(n_313)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_313),
.Y(n_342)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_299),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_314),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_315),
.B(n_325),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_265),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_316),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_283),
.B(n_270),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_310),
.C(n_286),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_321),
.Y(n_329)
);

NOR4xp25_ASAP7_75t_L g320 ( 
.A(n_291),
.B(n_275),
.C(n_270),
.D(n_268),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_304),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_292),
.A2(n_255),
.B1(n_275),
.B2(n_280),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_323),
.A2(n_326),
.B1(n_281),
.B2(n_302),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_289),
.B(n_268),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_292),
.A2(n_263),
.B1(n_261),
.B2(n_266),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_327),
.B(n_333),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_328),
.A2(n_322),
.B1(n_315),
.B2(n_326),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_310),
.B(n_290),
.C(n_291),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_332),
.B(n_336),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_306),
.A2(n_281),
.B1(n_300),
.B2(n_287),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_334),
.A2(n_325),
.B1(n_312),
.B2(n_309),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_307),
.A2(n_295),
.B(n_293),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_319),
.B(n_263),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_337),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_323),
.A2(n_296),
.B1(n_303),
.B2(n_282),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_338),
.A2(n_256),
.B1(n_195),
.B2(n_208),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_317),
.B(n_324),
.C(n_305),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_339),
.B(n_341),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_324),
.B(n_269),
.C(n_215),
.Y(n_341)
);

XNOR2x1_ASAP7_75t_L g345 ( 
.A(n_335),
.B(n_338),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_345),
.B(n_351),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_340),
.B(n_318),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_346),
.B(n_341),
.Y(n_369)
);

BUFx24_ASAP7_75t_SL g348 ( 
.A(n_342),
.Y(n_348)
);

BUFx24_ASAP7_75t_SL g363 ( 
.A(n_348),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_350),
.A2(n_358),
.B1(n_343),
.B2(n_330),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_339),
.B(n_311),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_353),
.B(n_328),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_334),
.A2(n_308),
.B1(n_252),
.B2(n_269),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_354),
.B(n_355),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_337),
.A2(n_260),
.B1(n_256),
.B2(n_215),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_335),
.B(n_214),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_357),
.B(n_359),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_331),
.B(n_245),
.Y(n_359)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_352),
.Y(n_361)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_361),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_362),
.A2(n_365),
.B1(n_367),
.B2(n_357),
.Y(n_378)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_352),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_364),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_356),
.A2(n_329),
.B1(n_332),
.B2(n_343),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_359),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_366),
.B(n_331),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_369),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_351),
.A2(n_336),
.B(n_333),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_371),
.A2(n_345),
.B1(n_347),
.B2(n_344),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_360),
.B(n_349),
.C(n_327),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_373),
.B(n_376),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_367),
.A2(n_329),
.B(n_370),
.Y(n_374)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_374),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_375),
.B(n_370),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_360),
.B(n_347),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_378),
.A2(n_374),
.B1(n_381),
.B2(n_377),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_379),
.B(n_245),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_363),
.B(n_344),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_380),
.B(n_368),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_384),
.B(n_386),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_385),
.B(n_387),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_373),
.A2(n_195),
.B(n_245),
.Y(n_386)
);

AOI322xp5_ASAP7_75t_L g387 ( 
.A1(n_372),
.A2(n_245),
.A3(n_208),
.B1(n_10),
.B2(n_11),
.C1(n_8),
.C2(n_4),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_388),
.B(n_4),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_389),
.Y(n_392)
);

FAx1_ASAP7_75t_SL g393 ( 
.A(n_383),
.B(n_376),
.CI(n_208),
.CON(n_393),
.SN(n_393)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_393),
.B(n_394),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_391),
.A2(n_382),
.B(n_384),
.Y(n_395)
);

OAI21x1_ASAP7_75t_L g398 ( 
.A1(n_395),
.A2(n_397),
.B(n_396),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_390),
.B(n_385),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_398),
.B(n_399),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_395),
.A2(n_392),
.B(n_393),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_400),
.A2(n_11),
.B1(n_8),
.B2(n_10),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_401),
.B(n_10),
.Y(n_402)
);


endmodule