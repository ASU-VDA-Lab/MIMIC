module real_jpeg_935_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_286;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx2_ASAP7_75t_L g105 ( 
.A(n_0),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_1),
.B(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_1),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_1),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_1),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_1),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_1),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_1),
.B(n_26),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_2),
.Y(n_125)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_3),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_3),
.B(n_26),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_3),
.B(n_61),
.Y(n_258)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_4),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_4),
.B(n_38),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_4),
.B(n_31),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_4),
.B(n_49),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_5),
.B(n_26),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_5),
.B(n_38),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_5),
.B(n_31),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_5),
.B(n_61),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_5),
.B(n_49),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_5),
.B(n_103),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_5),
.B(n_81),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_5),
.B(n_125),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_6),
.B(n_26),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_6),
.B(n_38),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_6),
.B(n_31),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_6),
.B(n_49),
.Y(n_107)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_6),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_6),
.B(n_103),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_8),
.B(n_26),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_8),
.B(n_38),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_8),
.B(n_31),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_8),
.B(n_49),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_8),
.B(n_61),
.Y(n_289)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g81 ( 
.A(n_10),
.Y(n_81)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_13),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_13),
.B(n_38),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_13),
.B(n_31),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_26),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_14),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_14),
.B(n_31),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_14),
.B(n_49),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_14),
.B(n_81),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_14),
.B(n_61),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_14),
.B(n_103),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_14),
.B(n_125),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI31xp33_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_25),
.A3(n_163),
.B(n_323),
.Y(n_17)
);

OAI211xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_42),
.B(n_89),
.C(n_322),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_64),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_21),
.B(n_64),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_50),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_42),
.B2(n_43),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B1(n_29),
.B2(n_41),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_25),
.B(n_75),
.C(n_76),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_25),
.A2(n_41),
.B1(n_118),
.B2(n_120),
.Y(n_117)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_26),
.Y(n_197)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_34),
.B(n_40),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_34),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_44),
.C(n_47),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_30),
.A2(n_47),
.B1(n_48),
.B2(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_30),
.B(n_193),
.C(n_200),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_30),
.A2(n_54),
.B1(n_200),
.B2(n_234),
.Y(n_233)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_31),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_34),
.A2(n_35),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_35),
.B(n_102),
.C(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_37),
.B(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_37),
.B(n_167),
.Y(n_166)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_40),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_45),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_44),
.A2(n_45),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_45),
.B(n_114),
.C(n_116),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_47),
.A2(n_48),
.B1(n_59),
.B2(n_60),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_47),
.A2(n_48),
.B1(n_186),
.B2(n_265),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_57),
.C(n_59),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_48),
.B(n_115),
.C(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_SL g220 ( 
.A(n_49),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_55),
.C(n_56),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_56),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_57),
.A2(n_58),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_59),
.A2(n_60),
.B1(n_79),
.B2(n_80),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_59),
.A2(n_60),
.B1(n_108),
.B2(n_148),
.Y(n_278)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_79),
.C(n_82),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_60),
.B(n_108),
.C(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_61),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_86),
.C(n_87),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_65),
.A2(n_66),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_78),
.C(n_83),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_67),
.A2(n_68),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_74),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_73),
.C(n_74),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_70),
.A2(n_71),
.B1(n_126),
.B2(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_70),
.A2(n_71),
.B1(n_171),
.B2(n_172),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_71),
.B(n_122),
.C(n_126),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_71),
.B(n_165),
.C(n_171),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_75),
.A2(n_76),
.B1(n_77),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_75),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_75),
.B(n_166),
.C(n_168),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_75),
.A2(n_119),
.B1(n_166),
.B2(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_78),
.B(n_83),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_79),
.A2(n_80),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_SL g133 ( 
.A(n_79),
.B(n_97),
.C(n_101),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_79),
.A2(n_80),
.B1(n_257),
.B2(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_80),
.B(n_257),
.C(n_258),
.Y(n_256)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_81),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_82),
.B(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_86),
.B(n_87),
.Y(n_319)
);

A2O1A1O1Ixp25_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_201),
.B(n_313),
.C(n_316),
.D(n_321),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_173),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_91),
.A2(n_314),
.B(n_315),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_139),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_92),
.B(n_139),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_127),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_93),
.B(n_128),
.C(n_138),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_117),
.C(n_121),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_94),
.B(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_106),
.C(n_110),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_95),
.A2(n_96),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_101),
.A2(n_102),
.B1(n_124),
.B2(n_154),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_106),
.B(n_110),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.C(n_109),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_107),
.B(n_109),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_108),
.Y(n_148)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_113),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_114),
.A2(n_115),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_121),
.Y(n_141)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_118),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_122),
.A2(n_123),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_153),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_124),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_184)
);

INVx3_ASAP7_75t_SL g255 ( 
.A(n_125),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_126),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_134),
.B1(n_137),
.B2(n_138),
.Y(n_127)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_132),
.C(n_133),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_129),
.A2(n_130),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_132),
.B(n_133),
.Y(n_143)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_134),
.Y(n_138)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.C(n_145),
.Y(n_139)
);

FAx1_ASAP7_75t_SL g174 ( 
.A(n_140),
.B(n_142),
.CI(n_145),
.CON(n_174),
.SN(n_174)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_143),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_160),
.C(n_164),
.Y(n_145)
);

FAx1_ASAP7_75t_SL g176 ( 
.A(n_146),
.B(n_160),
.CI(n_164),
.CON(n_176),
.SN(n_176)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.C(n_157),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_147),
.B(n_151),
.Y(n_238)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_149),
.Y(n_150)
);

O2A1O1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_154),
.B(n_155),
.C(n_156),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_152),
.B(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_152),
.A2(n_153),
.B1(n_254),
.B2(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_155),
.B(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_156),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_157),
.B(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_158),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_191),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_167),
.B(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_167),
.B(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_170),
.B(n_228),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_170),
.B(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_174),
.B(n_175),
.Y(n_314)
);

BUFx24_ASAP7_75t_SL g325 ( 
.A(n_174),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.C(n_180),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_176),
.B(n_177),
.Y(n_311)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_176),
.Y(n_324)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_178),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_180),
.B(n_311),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_190),
.C(n_192),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_181),
.A2(n_182),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.C(n_187),
.Y(n_182)
);

FAx1_ASAP7_75t_SL g267 ( 
.A(n_183),
.B(n_185),
.CI(n_187),
.CON(n_267),
.SN(n_267)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_186),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_190),
.B(n_192),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_193),
.A2(n_194),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_198),
.C(n_199),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_198),
.A2(n_199),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_198),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_199),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_200),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_268),
.B(n_307),
.C(n_308),
.D(n_312),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_243),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_204),
.B(n_243),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_235),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_205),
.B(n_236),
.C(n_242),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_223),
.C(n_231),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_206),
.A2(n_207),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_212),
.C(n_216),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_208),
.B(n_299),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_212),
.A2(n_213),
.B1(n_216),
.B2(n_300),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_213),
.A2(n_214),
.B(n_215),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_216),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_219),
.C(n_221),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_217),
.A2(n_218),
.B1(n_221),
.B2(n_222),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_251),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_223),
.B(n_231),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_227),
.C(n_229),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_225),
.B(n_278),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_229),
.Y(n_260)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_239),
.B2(n_242),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_239),
.Y(n_242)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_240),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_247),
.C(n_266),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_244),
.A2(n_266),
.B1(n_267),
.B2(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_244),
.Y(n_304)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_247),
.B(n_303),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_259),
.C(n_261),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_248),
.B(n_295),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_252),
.C(n_256),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_249),
.A2(n_250),
.B1(n_280),
.B2(n_282),
.Y(n_279)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_252),
.A2(n_253),
.B1(n_256),
.B2(n_281),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_254),
.Y(n_292)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_256),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_257),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_259),
.A2(n_261),
.B1(n_262),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_259),
.Y(n_296)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_267),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_301),
.B(n_306),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_293),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_279),
.C(n_283),
.Y(n_270)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_271),
.Y(n_326)
);

FAx1_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_276),
.CI(n_277),
.CON(n_271),
.SN(n_271)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_276),
.C(n_277),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.C(n_275),
.Y(n_272)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_280),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_287),
.C(n_291),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.C(n_290),
.Y(n_287)
);

BUFx24_ASAP7_75t_SL g329 ( 
.A(n_293),
.Y(n_329)
);

FAx1_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_297),
.CI(n_298),
.CON(n_293),
.SN(n_293)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_297),
.C(n_298),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_305),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_305),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_309),
.B(n_310),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_318),
.Y(n_321)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_319),
.Y(n_320)
);


endmodule