module fake_aes_7779_n_1142 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_1142);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1142;
wire n_663;
wire n_791;
wire n_707;
wire n_361;
wire n_513;
wire n_963;
wire n_1092;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_252;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_1056;
wire n_802;
wire n_985;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_1122;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_1128;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_786;
wire n_724;
wire n_857;
wire n_345;
wire n_360;
wire n_1090;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1024;
wire n_1016;
wire n_1078;
wire n_572;
wire n_1017;
wire n_324;
wire n_1097;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_975;
wire n_279;
wire n_303;
wire n_968;
wire n_1042;
wire n_1060;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_1011;
wire n_1025;
wire n_1132;
wire n_880;
wire n_1101;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_818;
wire n_769;
wire n_844;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_293;
wire n_1138;
wire n_533;
wire n_506;
wire n_393;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_1091;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_950;
wire n_1046;
wire n_460;
wire n_935;
wire n_478;
wire n_415;
wire n_482;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_1140;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_990;
wire n_751;
wire n_800;
wire n_626;
wire n_941;
wire n_466;
wire n_302;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_703;
wire n_839;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_285;
wire n_446;
wire n_420;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_1089;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_1066;
wire n_539;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_1135;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_681;
wire n_1139;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_419;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_1125;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_955;
wire n_1133;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_1110;
wire n_325;
wire n_1131;
wire n_1102;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1123;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_912;
wire n_924;
wire n_841;
wire n_947;
wire n_1141;
wire n_378;
wire n_582;
wire n_1043;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_1096;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_1136;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1117;
wire n_1040;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_1112;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_901;
wire n_834;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_281;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_695;
wire n_650;
wire n_625;
wire n_469;
wire n_1104;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_1134;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_1137;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_257;
wire n_992;
wire n_1127;
wire n_269;
INVx1_ASAP7_75t_L g251 ( .A(n_8), .Y(n_251) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_232), .Y(n_252) );
BUFx2_ASAP7_75t_L g253 ( .A(n_110), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_133), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_97), .Y(n_255) );
CKINVDCx20_ASAP7_75t_R g256 ( .A(n_27), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_191), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_202), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_4), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_247), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_131), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_201), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_192), .Y(n_263) );
INVx4_ASAP7_75t_R g264 ( .A(n_25), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_64), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_132), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_2), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_222), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_90), .Y(n_269) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_37), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_25), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_194), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_106), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_185), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_34), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_119), .Y(n_276) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_76), .Y(n_277) );
INVxp67_ASAP7_75t_L g278 ( .A(n_183), .Y(n_278) );
INVx1_ASAP7_75t_SL g279 ( .A(n_76), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_149), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_49), .Y(n_281) );
CKINVDCx20_ASAP7_75t_R g282 ( .A(n_60), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_236), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_181), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_77), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_205), .Y(n_286) );
CKINVDCx16_ASAP7_75t_R g287 ( .A(n_176), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_86), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_197), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_128), .Y(n_290) );
INVxp33_ASAP7_75t_SL g291 ( .A(n_121), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_219), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_175), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_104), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_182), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_136), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_221), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_122), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_63), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_99), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_195), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_160), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_209), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_116), .Y(n_304) );
CKINVDCx16_ASAP7_75t_R g305 ( .A(n_212), .Y(n_305) );
CKINVDCx20_ASAP7_75t_R g306 ( .A(n_170), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_45), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_174), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_166), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_71), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_100), .Y(n_311) );
CKINVDCx20_ASAP7_75t_R g312 ( .A(n_51), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_240), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_89), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_187), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_96), .Y(n_316) );
CKINVDCx20_ASAP7_75t_R g317 ( .A(n_225), .Y(n_317) );
CKINVDCx16_ASAP7_75t_R g318 ( .A(n_203), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_91), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_24), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_40), .Y(n_321) );
CKINVDCx20_ASAP7_75t_R g322 ( .A(n_109), .Y(n_322) );
BUFx3_ASAP7_75t_L g323 ( .A(n_233), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_142), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_143), .Y(n_325) );
INVxp67_ASAP7_75t_L g326 ( .A(n_190), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_22), .Y(n_327) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_169), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_180), .Y(n_329) );
BUFx3_ASAP7_75t_L g330 ( .A(n_231), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_218), .Y(n_331) );
INVx1_ASAP7_75t_SL g332 ( .A(n_151), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_73), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_85), .Y(n_334) );
CKINVDCx14_ASAP7_75t_R g335 ( .A(n_112), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_164), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_177), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_102), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_27), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_238), .Y(n_340) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_227), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_188), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_65), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_208), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_178), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_3), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_193), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_38), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_125), .Y(n_349) );
BUFx10_ASAP7_75t_L g350 ( .A(n_150), .Y(n_350) );
INVxp67_ASAP7_75t_L g351 ( .A(n_83), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_118), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_145), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_235), .Y(n_354) );
BUFx10_ASAP7_75t_L g355 ( .A(n_153), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_89), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_101), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_173), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_52), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_171), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_8), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_126), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_250), .Y(n_363) );
CKINVDCx20_ASAP7_75t_R g364 ( .A(n_140), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_46), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_196), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_53), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_130), .Y(n_368) );
INVxp67_ASAP7_75t_L g369 ( .A(n_9), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_54), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_92), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_216), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_127), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_55), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_94), .Y(n_375) );
BUFx2_ASAP7_75t_L g376 ( .A(n_88), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_214), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_155), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_108), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_60), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_234), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_114), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_228), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_167), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_103), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_86), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_35), .Y(n_387) );
NOR2xp67_ASAP7_75t_L g388 ( .A(n_211), .B(n_159), .Y(n_388) );
INVxp67_ASAP7_75t_SL g389 ( .A(n_135), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_51), .Y(n_390) );
INVx1_ASAP7_75t_SL g391 ( .A(n_28), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_58), .Y(n_392) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_30), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_45), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_139), .Y(n_395) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_154), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_16), .Y(n_397) );
CKINVDCx5p33_ASAP7_75t_R g398 ( .A(n_83), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_50), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_287), .Y(n_400) );
INVx3_ASAP7_75t_L g401 ( .A(n_350), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_327), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_253), .B(n_0), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_327), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_387), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_387), .Y(n_406) );
AND2x4_ASAP7_75t_L g407 ( .A(n_254), .B(n_0), .Y(n_407) );
INVx3_ASAP7_75t_L g408 ( .A(n_350), .Y(n_408) );
AND2x4_ASAP7_75t_L g409 ( .A(n_254), .B(n_1), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_255), .Y(n_410) );
OAI22xp5_ASAP7_75t_SL g411 ( .A1(n_256), .A2(n_3), .B1(n_1), .B2(n_2), .Y(n_411) );
AND2x4_ASAP7_75t_L g412 ( .A(n_292), .B(n_4), .Y(n_412) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_252), .Y(n_413) );
CKINVDCx16_ASAP7_75t_R g414 ( .A(n_305), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_257), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_252), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_252), .Y(n_417) );
NOR2x1_ASAP7_75t_L g418 ( .A(n_258), .B(n_5), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_270), .Y(n_419) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_252), .Y(n_420) );
AND2x4_ASAP7_75t_L g421 ( .A(n_292), .B(n_5), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_341), .B(n_6), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_376), .B(n_7), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_306), .A2(n_10), .B1(n_7), .B2(n_9), .Y(n_424) );
OA21x2_ASAP7_75t_L g425 ( .A1(n_349), .A2(n_10), .B(n_11), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_328), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_328), .Y(n_427) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_328), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_261), .Y(n_429) );
AND2x4_ASAP7_75t_L g430 ( .A(n_349), .B(n_11), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_262), .Y(n_431) );
INVx3_ASAP7_75t_L g432 ( .A(n_350), .Y(n_432) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_328), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_396), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_306), .A2(n_12), .B1(n_13), .B2(n_14), .Y(n_435) );
INVx1_ASAP7_75t_SL g436 ( .A(n_419), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_425), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_414), .A2(n_322), .B1(n_364), .B2(n_317), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_425), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_425), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_401), .B(n_318), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_414), .Y(n_442) );
BUFx10_ASAP7_75t_L g443 ( .A(n_407), .Y(n_443) );
OAI22xp33_ASAP7_75t_L g444 ( .A1(n_419), .A2(n_269), .B1(n_275), .B2(n_265), .Y(n_444) );
INVx4_ASAP7_75t_L g445 ( .A(n_401), .Y(n_445) );
AO22x2_ASAP7_75t_L g446 ( .A1(n_424), .A2(n_259), .B1(n_267), .B2(n_251), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_401), .B(n_278), .Y(n_447) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_413), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_425), .Y(n_449) );
BUFx2_ASAP7_75t_L g450 ( .A(n_400), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_425), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_423), .B(n_277), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_407), .A2(n_281), .B1(n_285), .B2(n_271), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_416), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_401), .B(n_326), .Y(n_455) );
BUFx4f_ASAP7_75t_L g456 ( .A(n_407), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_408), .B(n_335), .Y(n_457) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_408), .B(n_355), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_408), .B(n_265), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_425), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_408), .B(n_355), .Y(n_461) );
BUFx4f_ASAP7_75t_L g462 ( .A(n_407), .Y(n_462) );
INVx3_ASAP7_75t_L g463 ( .A(n_407), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_416), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_408), .B(n_335), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_416), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_432), .B(n_355), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_417), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_409), .A2(n_299), .B1(n_310), .B2(n_288), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_423), .B(n_380), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_409), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_409), .A2(n_322), .B1(n_364), .B2(n_317), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_403), .B(n_269), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_409), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_409), .Y(n_475) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_413), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_412), .Y(n_477) );
INVx4_ASAP7_75t_L g478 ( .A(n_432), .Y(n_478) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_413), .Y(n_479) );
INVx4_ASAP7_75t_L g480 ( .A(n_432), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_403), .B(n_319), .Y(n_481) );
INVx3_ASAP7_75t_L g482 ( .A(n_412), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_412), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_412), .Y(n_484) );
AND2x6_ASAP7_75t_SL g485 ( .A(n_442), .B(n_422), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_456), .B(n_462), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_436), .A2(n_432), .B1(n_422), .B2(n_412), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_471), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_459), .B(n_410), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_471), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_473), .A2(n_421), .B1(n_430), .B2(n_424), .Y(n_491) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_438), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_437), .Y(n_493) );
NAND2x1_ASAP7_75t_L g494 ( .A(n_445), .B(n_421), .Y(n_494) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_473), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_437), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_456), .A2(n_430), .B1(n_421), .B2(n_410), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_456), .B(n_421), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_441), .B(n_415), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_452), .B(n_319), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_462), .A2(n_430), .B1(n_421), .B2(n_429), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_474), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_452), .B(n_435), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_439), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_462), .B(n_430), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_443), .B(n_430), .Y(n_506) );
AND2x6_ASAP7_75t_SL g507 ( .A(n_446), .B(n_411), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_439), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_457), .B(n_429), .Y(n_509) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_443), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g511 ( .A1(n_481), .A2(n_435), .B1(n_411), .B2(n_321), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_457), .B(n_431), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_465), .B(n_445), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_465), .B(n_431), .Y(n_514) );
INVx1_ASAP7_75t_SL g515 ( .A(n_470), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_475), .Y(n_516) );
O2A1O1Ixp5_ASAP7_75t_L g517 ( .A1(n_440), .A2(n_389), .B(n_266), .C(n_268), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_450), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_446), .A2(n_321), .B1(n_334), .B2(n_320), .Y(n_519) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_443), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_440), .Y(n_521) );
INVx2_ASAP7_75t_SL g522 ( .A(n_478), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_450), .B(n_334), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_475), .Y(n_524) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_444), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_458), .B(n_291), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_472), .A2(n_346), .B1(n_365), .B2(n_339), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_478), .B(n_260), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_461), .B(n_291), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_467), .B(n_260), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_480), .B(n_280), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_447), .B(n_296), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_449), .B(n_263), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_449), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_455), .B(n_296), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_451), .B(n_272), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_451), .B(n_273), .Y(n_537) );
OAI22x1_ASAP7_75t_SL g538 ( .A1(n_446), .A2(n_282), .B1(n_312), .B2(n_256), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_453), .B(n_297), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_477), .B(n_324), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_469), .B(n_324), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_477), .B(n_339), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_483), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_484), .A2(n_463), .B1(n_482), .B2(n_460), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_460), .B(n_274), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_484), .B(n_325), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_463), .A2(n_418), .B1(n_333), .B2(n_343), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_482), .B(n_336), .Y(n_548) );
NAND2x1p5_ASAP7_75t_L g549 ( .A(n_472), .B(n_418), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_446), .A2(n_348), .B1(n_356), .B2(n_314), .Y(n_550) );
AND3x1_ASAP7_75t_L g551 ( .A(n_454), .B(n_361), .C(n_359), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_454), .B(n_336), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_464), .B(n_276), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_464), .Y(n_554) );
O2A1O1Ixp33_ASAP7_75t_L g555 ( .A1(n_466), .A2(n_369), .B(n_351), .C(n_402), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_466), .A2(n_365), .B1(n_370), .B2(n_346), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_468), .B(n_342), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_468), .B(n_342), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_448), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_448), .Y(n_560) );
NAND2xp33_ASAP7_75t_L g561 ( .A(n_448), .B(n_347), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_448), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_448), .A2(n_386), .B1(n_390), .B2(n_367), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_476), .B(n_347), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_476), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_476), .B(n_358), .Y(n_566) );
INVx5_ASAP7_75t_L g567 ( .A(n_476), .Y(n_567) );
BUFx5_ASAP7_75t_L g568 ( .A(n_476), .Y(n_568) );
INVx3_ASAP7_75t_L g569 ( .A(n_479), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_479), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_479), .A2(n_392), .B1(n_397), .B2(n_394), .Y(n_571) );
INVx4_ASAP7_75t_L g572 ( .A(n_479), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_459), .B(n_358), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_456), .A2(n_399), .B1(n_393), .B2(n_402), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_515), .B(n_374), .Y(n_575) );
BUFx4f_ASAP7_75t_L g576 ( .A(n_503), .Y(n_576) );
NAND2x1p5_ASAP7_75t_L g577 ( .A(n_510), .B(n_404), .Y(n_577) );
BUFx3_ASAP7_75t_L g578 ( .A(n_518), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_491), .A2(n_312), .B1(n_282), .B2(n_404), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_495), .B(n_279), .Y(n_580) );
O2A1O1Ixp33_ASAP7_75t_L g581 ( .A1(n_525), .A2(n_391), .B(n_406), .C(n_405), .Y(n_581) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_510), .Y(n_582) );
NOR2xp67_ASAP7_75t_L g583 ( .A(n_511), .B(n_378), .Y(n_583) );
NOR3xp33_ASAP7_75t_L g584 ( .A(n_527), .B(n_398), .C(n_307), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_500), .B(n_378), .Y(n_585) );
A2O1A1Ixp33_ASAP7_75t_L g586 ( .A1(n_488), .A2(n_406), .B(n_405), .C(n_283), .Y(n_586) );
BUFx12f_ASAP7_75t_L g587 ( .A(n_485), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_490), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_533), .A2(n_290), .B(n_289), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_523), .B(n_383), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_510), .B(n_284), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_510), .B(n_286), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_497), .A2(n_393), .B1(n_295), .B2(n_300), .Y(n_593) );
A2O1A1Ixp33_ASAP7_75t_L g594 ( .A1(n_502), .A2(n_301), .B(n_302), .C(n_294), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_542), .B(n_332), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_501), .A2(n_393), .B1(n_304), .B2(n_308), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_542), .B(n_518), .Y(n_597) );
INVx3_ASAP7_75t_L g598 ( .A(n_520), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_549), .B(n_12), .Y(n_599) );
O2A1O1Ixp33_ASAP7_75t_L g600 ( .A1(n_498), .A2(n_303), .B(n_315), .C(n_313), .Y(n_600) );
A2O1A1Ixp33_ASAP7_75t_L g601 ( .A1(n_516), .A2(n_329), .B(n_337), .C(n_331), .Y(n_601) );
NOR2xp33_ASAP7_75t_SL g602 ( .A(n_520), .B(n_293), .Y(n_602) );
AOI21xp5_ASAP7_75t_L g603 ( .A1(n_536), .A2(n_340), .B(n_338), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_536), .A2(n_345), .B(n_344), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_499), .B(n_298), .Y(n_605) );
AO32x2_ASAP7_75t_L g606 ( .A1(n_572), .A2(n_413), .A3(n_433), .B1(n_428), .B2(n_420), .Y(n_606) );
INVxp67_ASAP7_75t_L g607 ( .A(n_551), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_509), .B(n_309), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_492), .B(n_13), .Y(n_609) );
NAND2xp5_ASAP7_75t_SL g610 ( .A(n_520), .B(n_311), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_512), .B(n_316), .Y(n_611) );
BUFx2_ASAP7_75t_R g612 ( .A(n_492), .Y(n_612) );
BUFx4f_ASAP7_75t_L g613 ( .A(n_520), .Y(n_613) );
AND2x6_ASAP7_75t_SL g614 ( .A(n_538), .B(n_264), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_524), .Y(n_615) );
BUFx2_ASAP7_75t_L g616 ( .A(n_519), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_543), .Y(n_617) );
O2A1O1Ixp33_ASAP7_75t_L g618 ( .A1(n_498), .A2(n_353), .B(n_354), .C(n_352), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_556), .B(n_14), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_496), .A2(n_360), .B1(n_363), .B2(n_362), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_514), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_504), .A2(n_366), .B1(n_371), .B2(n_368), .Y(n_622) );
AOI21x1_ASAP7_75t_L g623 ( .A1(n_537), .A2(n_388), .B(n_375), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_537), .A2(n_379), .B(n_372), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_489), .B(n_381), .Y(n_625) );
BUFx3_ASAP7_75t_L g626 ( .A(n_494), .Y(n_626) );
OA22x2_ASAP7_75t_L g627 ( .A1(n_507), .A2(n_384), .B1(n_385), .B2(n_382), .Y(n_627) );
AOI21xp5_ASAP7_75t_L g628 ( .A1(n_545), .A2(n_395), .B(n_373), .Y(n_628) );
O2A1O1Ixp33_ASAP7_75t_L g629 ( .A1(n_505), .A2(n_373), .B(n_377), .C(n_357), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_545), .A2(n_377), .B(n_357), .Y(n_630) );
BUFx6f_ASAP7_75t_L g631 ( .A(n_504), .Y(n_631) );
AND2x4_ASAP7_75t_L g632 ( .A(n_486), .B(n_323), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_550), .A2(n_330), .B1(n_434), .B2(n_427), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g634 ( .A1(n_513), .A2(n_434), .B(n_427), .Y(n_634) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_508), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_487), .B(n_15), .Y(n_636) );
A2O1A1Ixp33_ASAP7_75t_L g637 ( .A1(n_517), .A2(n_434), .B(n_427), .C(n_417), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_548), .Y(n_638) );
CKINVDCx5p33_ASAP7_75t_R g639 ( .A(n_526), .Y(n_639) );
XNOR2xp5_ASAP7_75t_L g640 ( .A(n_547), .B(n_16), .Y(n_640) );
INVx5_ASAP7_75t_L g641 ( .A(n_522), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_521), .A2(n_426), .B1(n_433), .B2(n_428), .Y(n_642) );
CKINVDCx5p33_ASAP7_75t_R g643 ( .A(n_529), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_546), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g645 ( .A1(n_534), .A2(n_426), .B(n_420), .Y(n_645) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_506), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_540), .B(n_532), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_544), .A2(n_426), .B1(n_433), .B2(n_428), .Y(n_648) );
NOR2x1p5_ASAP7_75t_L g649 ( .A(n_539), .B(n_17), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_574), .A2(n_433), .B1(n_428), .B2(n_420), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_541), .B(n_17), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_530), .B(n_18), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_535), .A2(n_433), .B1(n_428), .B2(n_420), .Y(n_653) );
O2A1O1Ixp33_ASAP7_75t_L g654 ( .A1(n_555), .A2(n_18), .B(n_19), .C(n_20), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_531), .B(n_19), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_553), .Y(n_656) );
A2O1A1Ixp33_ASAP7_75t_L g657 ( .A1(n_573), .A2(n_433), .B(n_428), .C(n_420), .Y(n_657) );
OA22x2_ASAP7_75t_L g658 ( .A1(n_553), .A2(n_21), .B1(n_23), .B2(n_24), .Y(n_658) );
A2O1A1Ixp33_ASAP7_75t_L g659 ( .A1(n_528), .A2(n_433), .B(n_428), .C(n_29), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_552), .B(n_26), .Y(n_660) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_557), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_558), .Y(n_662) );
BUFx3_ASAP7_75t_L g663 ( .A(n_554), .Y(n_663) );
NOR2x1_ASAP7_75t_R g664 ( .A(n_562), .B(n_29), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_563), .Y(n_665) );
NOR2xp67_ASAP7_75t_L g666 ( .A(n_571), .B(n_30), .Y(n_666) );
NOR3xp33_ASAP7_75t_SL g667 ( .A(n_562), .B(n_31), .C(n_32), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_564), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_566), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_561), .B(n_31), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_561), .B(n_32), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_572), .Y(n_672) );
OAI21xp5_ASAP7_75t_L g673 ( .A1(n_559), .A2(n_95), .B(n_93), .Y(n_673) );
AOI22x1_ASAP7_75t_L g674 ( .A1(n_560), .A2(n_163), .B1(n_248), .B2(n_246), .Y(n_674) );
NOR2xp33_ASAP7_75t_SL g675 ( .A(n_567), .B(n_98), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_568), .B(n_33), .Y(n_676) );
BUFx2_ASAP7_75t_L g677 ( .A(n_568), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_568), .Y(n_678) );
O2A1O1Ixp33_ASAP7_75t_SL g679 ( .A1(n_565), .A2(n_165), .B(n_245), .C(n_244), .Y(n_679) );
A2O1A1Ixp33_ASAP7_75t_L g680 ( .A1(n_569), .A2(n_34), .B(n_35), .C(n_36), .Y(n_680) );
OR2x6_ASAP7_75t_L g681 ( .A(n_569), .B(n_36), .Y(n_681) );
AOI21xp5_ASAP7_75t_L g682 ( .A1(n_565), .A2(n_107), .B(n_105), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_569), .A2(n_38), .B1(n_39), .B2(n_40), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_570), .A2(n_113), .B(n_111), .Y(n_684) );
INVx1_ASAP7_75t_SL g685 ( .A(n_567), .Y(n_685) );
A2O1A1Ixp33_ASAP7_75t_L g686 ( .A1(n_570), .A2(n_39), .B(n_41), .C(n_42), .Y(n_686) );
BUFx6f_ASAP7_75t_L g687 ( .A(n_567), .Y(n_687) );
A2O1A1Ixp33_ASAP7_75t_L g688 ( .A1(n_568), .A2(n_41), .B(n_42), .C(n_43), .Y(n_688) );
AND2x4_ASAP7_75t_SL g689 ( .A(n_568), .B(n_43), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g690 ( .A(n_568), .B(n_44), .Y(n_690) );
NOR2xp33_ASAP7_75t_SL g691 ( .A(n_510), .B(n_115), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g692 ( .A1(n_533), .A2(n_120), .B(n_117), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_515), .B(n_44), .Y(n_693) );
AND2x4_ASAP7_75t_L g694 ( .A(n_542), .B(n_46), .Y(n_694) );
CKINVDCx5p33_ASAP7_75t_R g695 ( .A(n_518), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g696 ( .A1(n_491), .A2(n_47), .B1(n_48), .B2(n_49), .Y(n_696) );
BUFx3_ASAP7_75t_L g697 ( .A(n_518), .Y(n_697) );
AO31x2_ASAP7_75t_L g698 ( .A1(n_659), .A2(n_47), .A3(n_48), .B(n_50), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_597), .B(n_616), .Y(n_699) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_647), .A2(n_124), .B(n_123), .Y(n_700) );
INVx3_ASAP7_75t_L g701 ( .A(n_613), .Y(n_701) );
INVx4_ASAP7_75t_L g702 ( .A(n_613), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_579), .A2(n_55), .B1(n_56), .B2(n_57), .C(n_58), .Y(n_703) );
BUFx3_ASAP7_75t_L g704 ( .A(n_578), .Y(n_704) );
O2A1O1Ixp33_ASAP7_75t_SL g705 ( .A1(n_637), .A2(n_189), .B(n_243), .C(n_242), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_576), .B(n_56), .Y(n_706) );
OAI21xp5_ASAP7_75t_L g707 ( .A1(n_668), .A2(n_186), .B(n_241), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_631), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_576), .B(n_57), .Y(n_709) );
BUFx3_ASAP7_75t_L g710 ( .A(n_697), .Y(n_710) );
CKINVDCx5p33_ASAP7_75t_R g711 ( .A(n_587), .Y(n_711) );
NAND2xp5_ASAP7_75t_SL g712 ( .A(n_602), .B(n_59), .Y(n_712) );
NOR2x1_ASAP7_75t_R g713 ( .A(n_695), .B(n_59), .Y(n_713) );
OAI22xp33_ASAP7_75t_L g714 ( .A1(n_607), .A2(n_681), .B1(n_575), .B2(n_619), .Y(n_714) );
OAI21xp5_ASAP7_75t_L g715 ( .A1(n_669), .A2(n_184), .B(n_239), .Y(n_715) );
OAI221xp5_ASAP7_75t_L g716 ( .A1(n_584), .A2(n_61), .B1(n_62), .B2(n_63), .C(n_64), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_694), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_631), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_621), .Y(n_719) );
INVx2_ASAP7_75t_SL g720 ( .A(n_681), .Y(n_720) );
OA21x2_ASAP7_75t_L g721 ( .A1(n_673), .A2(n_179), .B(n_237), .Y(n_721) );
A2O1A1Ixp33_ASAP7_75t_L g722 ( .A1(n_651), .A2(n_61), .B(n_62), .C(n_65), .Y(n_722) );
INVx2_ASAP7_75t_SL g723 ( .A(n_681), .Y(n_723) );
AND2x4_ASAP7_75t_L g724 ( .A(n_641), .B(n_66), .Y(n_724) );
OR2x2_ASAP7_75t_L g725 ( .A(n_580), .B(n_66), .Y(n_725) );
BUFx3_ASAP7_75t_L g726 ( .A(n_687), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_696), .Y(n_727) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_577), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_588), .B(n_67), .Y(n_729) );
O2A1O1Ixp33_ASAP7_75t_L g730 ( .A1(n_581), .A2(n_67), .B(n_68), .C(n_69), .Y(n_730) );
OAI21xp33_ASAP7_75t_L g731 ( .A1(n_585), .A2(n_68), .B(n_69), .Y(n_731) );
NAND2x1p5_ASAP7_75t_L g732 ( .A(n_582), .B(n_70), .Y(n_732) );
BUFx10_ASAP7_75t_L g733 ( .A(n_689), .Y(n_733) );
A2O1A1Ixp33_ASAP7_75t_L g734 ( .A1(n_662), .A2(n_70), .B(n_71), .C(n_72), .Y(n_734) );
AOI31xp67_ASAP7_75t_L g735 ( .A1(n_653), .A2(n_198), .A3(n_230), .B(n_229), .Y(n_735) );
BUFx2_ASAP7_75t_R g736 ( .A(n_639), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_635), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_590), .B(n_74), .Y(n_738) );
A2O1A1Ixp33_ASAP7_75t_L g739 ( .A1(n_660), .A2(n_75), .B(n_77), .C(n_78), .Y(n_739) );
AND2x4_ASAP7_75t_L g740 ( .A(n_641), .B(n_75), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_615), .B(n_78), .Y(n_741) );
O2A1O1Ixp33_ASAP7_75t_L g742 ( .A1(n_654), .A2(n_79), .B(n_80), .C(n_81), .Y(n_742) );
AO32x2_ASAP7_75t_L g743 ( .A1(n_696), .A2(n_79), .A3(n_80), .B1(n_81), .B2(n_82), .Y(n_743) );
AO31x2_ASAP7_75t_L g744 ( .A1(n_648), .A2(n_586), .A3(n_633), .B(n_594), .Y(n_744) );
BUFx12f_ASAP7_75t_L g745 ( .A(n_614), .Y(n_745) );
A2O1A1Ixp33_ASAP7_75t_L g746 ( .A1(n_652), .A2(n_82), .B(n_84), .C(n_85), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_617), .B(n_84), .Y(n_747) );
O2A1O1Ixp33_ASAP7_75t_L g748 ( .A1(n_601), .A2(n_596), .B(n_593), .C(n_636), .Y(n_748) );
AOI221xp5_ASAP7_75t_SL g749 ( .A1(n_600), .A2(n_87), .B1(n_91), .B2(n_129), .C(n_134), .Y(n_749) );
OAI22x1_ASAP7_75t_L g750 ( .A1(n_649), .A2(n_137), .B1(n_138), .B2(n_141), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_661), .B(n_144), .Y(n_751) );
AO31x2_ASAP7_75t_L g752 ( .A1(n_648), .A2(n_146), .A3(n_147), .B(n_148), .Y(n_752) );
A2O1A1Ixp33_ASAP7_75t_L g753 ( .A1(n_618), .A2(n_152), .B(n_156), .C(n_157), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_646), .Y(n_754) );
CKINVDCx5p33_ASAP7_75t_R g755 ( .A(n_612), .Y(n_755) );
A2O1A1Ixp33_ASAP7_75t_L g756 ( .A1(n_629), .A2(n_158), .B(n_161), .C(n_162), .Y(n_756) );
AO32x2_ASAP7_75t_L g757 ( .A1(n_633), .A2(n_168), .A3(n_172), .B1(n_199), .B2(n_200), .Y(n_757) );
O2A1O1Ixp33_ASAP7_75t_SL g758 ( .A1(n_676), .A2(n_204), .B(n_206), .C(n_207), .Y(n_758) );
INVxp67_ASAP7_75t_L g759 ( .A(n_664), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g760 ( .A(n_643), .B(n_210), .Y(n_760) );
INVxp67_ASAP7_75t_L g761 ( .A(n_693), .Y(n_761) );
CKINVDCx5p33_ASAP7_75t_R g762 ( .A(n_640), .Y(n_762) );
AND2x4_ASAP7_75t_L g763 ( .A(n_641), .B(n_213), .Y(n_763) );
OA21x2_ASAP7_75t_L g764 ( .A1(n_673), .A2(n_215), .B(n_217), .Y(n_764) );
INVx2_ASAP7_75t_L g765 ( .A(n_635), .Y(n_765) );
OR2x2_ASAP7_75t_L g766 ( .A(n_609), .B(n_220), .Y(n_766) );
OR2x2_ASAP7_75t_L g767 ( .A(n_595), .B(n_223), .Y(n_767) );
AOI21x1_ASAP7_75t_L g768 ( .A1(n_623), .A2(n_224), .B(n_226), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_627), .A2(n_249), .B1(n_583), .B2(n_599), .Y(n_769) );
O2A1O1Ixp33_ASAP7_75t_SL g770 ( .A1(n_690), .A2(n_671), .B(n_670), .C(n_685), .Y(n_770) );
AO31x2_ASAP7_75t_L g771 ( .A1(n_642), .A2(n_686), .A3(n_688), .B(n_650), .Y(n_771) );
A2O1A1Ixp33_ASAP7_75t_L g772 ( .A1(n_589), .A2(n_624), .B(n_604), .C(n_603), .Y(n_772) );
O2A1O1Ixp33_ASAP7_75t_L g773 ( .A1(n_625), .A2(n_680), .B(n_622), .C(n_620), .Y(n_773) );
AOI21xp5_ASAP7_75t_L g774 ( .A1(n_605), .A2(n_611), .B(n_608), .Y(n_774) );
OAI21xp5_ASAP7_75t_L g775 ( .A1(n_656), .A2(n_628), .B(n_630), .Y(n_775) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_577), .A2(n_665), .B1(n_663), .B2(n_641), .Y(n_776) );
AOI22xp5_ASAP7_75t_L g777 ( .A1(n_602), .A2(n_666), .B1(n_632), .B2(n_667), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_683), .Y(n_778) );
AOI21xp5_ASAP7_75t_L g779 ( .A1(n_678), .A2(n_634), .B(n_672), .Y(n_779) );
O2A1O1Ixp33_ASAP7_75t_L g780 ( .A1(n_591), .A2(n_592), .B(n_610), .C(n_650), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_626), .B(n_582), .Y(n_781) );
OAI21x1_ASAP7_75t_L g782 ( .A1(n_674), .A2(n_684), .B(n_682), .Y(n_782) );
O2A1O1Ixp33_ASAP7_75t_L g783 ( .A1(n_679), .A2(n_692), .B(n_598), .C(n_645), .Y(n_783) );
NOR2xp33_ASAP7_75t_L g784 ( .A(n_598), .B(n_677), .Y(n_784) );
A2O1A1Ixp33_ASAP7_75t_L g785 ( .A1(n_675), .A2(n_691), .B(n_687), .C(n_658), .Y(n_785) );
AOI21xp5_ASAP7_75t_SL g786 ( .A1(n_687), .A2(n_658), .B(n_675), .Y(n_786) );
INVx3_ASAP7_75t_L g787 ( .A(n_691), .Y(n_787) );
AOI21xp5_ASAP7_75t_L g788 ( .A1(n_606), .A2(n_496), .B(n_493), .Y(n_788) );
AO31x2_ASAP7_75t_L g789 ( .A1(n_606), .A2(n_659), .A3(n_657), .B(n_637), .Y(n_789) );
O2A1O1Ixp5_ASAP7_75t_L g790 ( .A1(n_606), .A2(n_652), .B(n_655), .C(n_660), .Y(n_790) );
A2O1A1Ixp33_ASAP7_75t_L g791 ( .A1(n_647), .A2(n_638), .B(n_651), .C(n_644), .Y(n_791) );
AND2x4_ASAP7_75t_L g792 ( .A(n_621), .B(n_694), .Y(n_792) );
AOI21xp5_ASAP7_75t_L g793 ( .A1(n_647), .A2(n_496), .B(n_493), .Y(n_793) );
AOI21xp5_ASAP7_75t_L g794 ( .A1(n_647), .A2(n_496), .B(n_493), .Y(n_794) );
OR2x2_ASAP7_75t_L g795 ( .A(n_579), .B(n_515), .Y(n_795) );
OR2x2_ASAP7_75t_L g796 ( .A(n_579), .B(n_515), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g797 ( .A1(n_621), .A2(n_491), .B1(n_456), .B2(n_462), .Y(n_797) );
NOR2xp67_ASAP7_75t_SL g798 ( .A(n_578), .B(n_518), .Y(n_798) );
NOR2xp33_ASAP7_75t_L g799 ( .A(n_597), .B(n_515), .Y(n_799) );
OAI22xp5_ASAP7_75t_L g800 ( .A1(n_621), .A2(n_491), .B1(n_456), .B2(n_462), .Y(n_800) );
BUFx4f_ASAP7_75t_SL g801 ( .A(n_587), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g802 ( .A1(n_621), .A2(n_491), .B1(n_456), .B2(n_462), .Y(n_802) );
INVx2_ASAP7_75t_L g803 ( .A(n_631), .Y(n_803) );
O2A1O1Ixp33_ASAP7_75t_L g804 ( .A1(n_581), .A2(n_654), .B(n_696), .C(n_647), .Y(n_804) );
O2A1O1Ixp33_ASAP7_75t_SL g805 ( .A1(n_659), .A2(n_657), .B(n_637), .C(n_655), .Y(n_805) );
AND2x4_ASAP7_75t_L g806 ( .A(n_621), .B(n_694), .Y(n_806) );
AO31x2_ASAP7_75t_L g807 ( .A1(n_659), .A2(n_657), .A3(n_637), .B(n_648), .Y(n_807) );
BUFx2_ASAP7_75t_L g808 ( .A(n_578), .Y(n_808) );
AOI21xp5_ASAP7_75t_L g809 ( .A1(n_647), .A2(n_496), .B(n_493), .Y(n_809) );
OR2x2_ASAP7_75t_L g810 ( .A(n_579), .B(n_515), .Y(n_810) );
AOI21xp5_ASAP7_75t_L g811 ( .A1(n_647), .A2(n_496), .B(n_493), .Y(n_811) );
OR2x2_ASAP7_75t_L g812 ( .A(n_579), .B(n_515), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_621), .B(n_515), .Y(n_813) );
INVx5_ASAP7_75t_L g814 ( .A(n_681), .Y(n_814) );
AOI22xp5_ASAP7_75t_L g815 ( .A1(n_579), .A2(n_515), .B1(n_438), .B2(n_518), .Y(n_815) );
A2O1A1Ixp33_ASAP7_75t_L g816 ( .A1(n_647), .A2(n_638), .B(n_651), .C(n_644), .Y(n_816) );
NAND3xp33_ASAP7_75t_L g817 ( .A(n_659), .B(n_667), .C(n_585), .Y(n_817) );
A2O1A1Ixp33_ASAP7_75t_L g818 ( .A1(n_647), .A2(n_638), .B(n_651), .C(n_644), .Y(n_818) );
O2A1O1Ixp33_ASAP7_75t_SL g819 ( .A1(n_659), .A2(n_657), .B(n_637), .C(n_655), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_694), .Y(n_820) );
INVx3_ASAP7_75t_L g821 ( .A(n_702), .Y(n_821) );
AO31x2_ASAP7_75t_L g822 ( .A1(n_785), .A2(n_788), .A3(n_816), .B(n_818), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_813), .B(n_719), .Y(n_823) );
AOI21xp5_ASAP7_75t_L g824 ( .A1(n_793), .A2(n_809), .B(n_794), .Y(n_824) );
OAI22xp5_ASAP7_75t_L g825 ( .A1(n_814), .A2(n_727), .B1(n_714), .B2(n_795), .Y(n_825) );
INVx3_ASAP7_75t_L g826 ( .A(n_702), .Y(n_826) );
NAND2xp5_ASAP7_75t_SL g827 ( .A(n_814), .B(n_815), .Y(n_827) );
CKINVDCx20_ASAP7_75t_R g828 ( .A(n_801), .Y(n_828) );
AO21x2_ASAP7_75t_L g829 ( .A1(n_786), .A2(n_770), .B(n_715), .Y(n_829) );
AND2x2_ASAP7_75t_L g830 ( .A(n_799), .B(n_796), .Y(n_830) );
CKINVDCx20_ASAP7_75t_R g831 ( .A(n_711), .Y(n_831) );
AOI21x1_ASAP7_75t_L g832 ( .A1(n_721), .A2(n_764), .B(n_768), .Y(n_832) );
AOI22xp33_ASAP7_75t_SL g833 ( .A1(n_814), .A2(n_699), .B1(n_812), .B2(n_810), .Y(n_833) );
OR2x6_ASAP7_75t_L g834 ( .A(n_720), .B(n_723), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_729), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_741), .Y(n_836) );
NOR2xp33_ASAP7_75t_L g837 ( .A(n_792), .B(n_806), .Y(n_837) );
AND2x2_ASAP7_75t_L g838 ( .A(n_725), .B(n_706), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_778), .B(n_717), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_747), .Y(n_840) );
INVx3_ASAP7_75t_L g841 ( .A(n_726), .Y(n_841) );
INVx8_ASAP7_75t_L g842 ( .A(n_724), .Y(n_842) );
AOI21xp5_ASAP7_75t_L g843 ( .A1(n_811), .A2(n_774), .B(n_791), .Y(n_843) );
AO21x2_ASAP7_75t_L g844 ( .A1(n_707), .A2(n_819), .B(n_805), .Y(n_844) );
OAI22xp5_ASAP7_75t_SL g845 ( .A1(n_755), .A2(n_762), .B1(n_745), .B2(n_759), .Y(n_845) );
OR2x6_ASAP7_75t_L g846 ( .A(n_724), .B(n_740), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_754), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_740), .Y(n_848) );
INVxp67_ASAP7_75t_L g849 ( .A(n_798), .Y(n_849) );
AND2x4_ASAP7_75t_SL g850 ( .A(n_733), .B(n_701), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_817), .A2(n_797), .B1(n_802), .B2(n_800), .Y(n_851) );
OAI21xp5_ASAP7_75t_L g852 ( .A1(n_790), .A2(n_804), .B(n_773), .Y(n_852) );
AOI21xp5_ASAP7_75t_L g853 ( .A1(n_783), .A2(n_775), .B(n_779), .Y(n_853) );
A2O1A1Ixp33_ASAP7_75t_L g854 ( .A1(n_748), .A2(n_742), .B(n_730), .C(n_731), .Y(n_854) );
INVx2_ASAP7_75t_L g855 ( .A(n_732), .Y(n_855) );
A2O1A1Ixp33_ASAP7_75t_L g856 ( .A1(n_722), .A2(n_746), .B(n_738), .C(n_777), .Y(n_856) );
A2O1A1Ixp33_ASAP7_75t_L g857 ( .A1(n_739), .A2(n_780), .B(n_709), .C(n_761), .Y(n_857) );
AOI21xp5_ASAP7_75t_L g858 ( .A1(n_787), .A2(n_772), .B(n_705), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_820), .B(n_769), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_743), .Y(n_860) );
AOI21xp5_ASAP7_75t_L g861 ( .A1(n_721), .A2(n_764), .B(n_776), .Y(n_861) );
INVx2_ASAP7_75t_L g862 ( .A(n_763), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_743), .Y(n_863) );
INVx6_ASAP7_75t_L g864 ( .A(n_704), .Y(n_864) );
CKINVDCx16_ASAP7_75t_R g865 ( .A(n_710), .Y(n_865) );
A2O1A1Ixp33_ASAP7_75t_L g866 ( .A1(n_703), .A2(n_767), .B(n_749), .C(n_734), .Y(n_866) );
AND2x4_ASAP7_75t_L g867 ( .A(n_763), .B(n_701), .Y(n_867) );
AOI22xp33_ASAP7_75t_SL g868 ( .A1(n_733), .A2(n_716), .B1(n_808), .B2(n_760), .Y(n_868) );
O2A1O1Ixp33_ASAP7_75t_L g869 ( .A1(n_766), .A2(n_712), .B(n_753), .C(n_751), .Y(n_869) );
OR2x2_ASAP7_75t_L g870 ( .A(n_728), .B(n_781), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_744), .B(n_784), .Y(n_871) );
INVx2_ASAP7_75t_L g872 ( .A(n_698), .Y(n_872) );
BUFx4_ASAP7_75t_R g873 ( .A(n_736), .Y(n_873) );
OAI332xp33_ASAP7_75t_L g874 ( .A1(n_713), .A2(n_743), .A3(n_698), .B1(n_750), .B2(n_708), .B3(n_765), .C1(n_803), .C2(n_718), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_744), .B(n_771), .Y(n_875) );
AOI21xp5_ASAP7_75t_L g876 ( .A1(n_758), .A2(n_756), .B(n_700), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_698), .Y(n_877) );
AOI21xp5_ASAP7_75t_L g878 ( .A1(n_737), .A2(n_735), .B(n_807), .Y(n_878) );
NOR2x1_ASAP7_75t_L g879 ( .A(n_757), .B(n_752), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_752), .Y(n_880) );
OAI221xp5_ASAP7_75t_L g881 ( .A1(n_807), .A2(n_511), .B1(n_815), .B2(n_799), .C(n_503), .Y(n_881) );
AOI21xp33_ASAP7_75t_L g882 ( .A1(n_789), .A2(n_804), .B(n_714), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_789), .B(n_757), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_813), .Y(n_884) );
AOI21xp5_ASAP7_75t_L g885 ( .A1(n_793), .A2(n_809), .B(n_794), .Y(n_885) );
AOI221xp5_ASAP7_75t_L g886 ( .A1(n_799), .A2(n_579), .B1(n_515), .B2(n_527), .C(n_446), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_813), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_719), .B(n_621), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_813), .Y(n_889) );
INVx11_ASAP7_75t_L g890 ( .A(n_745), .Y(n_890) );
AOI22xp33_ASAP7_75t_SL g891 ( .A1(n_727), .A2(n_438), .B1(n_579), .B2(n_492), .Y(n_891) );
INVx3_ASAP7_75t_L g892 ( .A(n_702), .Y(n_892) );
BUFx12f_ASAP7_75t_L g893 ( .A(n_711), .Y(n_893) );
AOI22xp33_ASAP7_75t_SL g894 ( .A1(n_727), .A2(n_438), .B1(n_579), .B2(n_492), .Y(n_894) );
A2O1A1Ixp33_ASAP7_75t_L g895 ( .A1(n_791), .A2(n_816), .B(n_818), .C(n_774), .Y(n_895) );
AOI221xp5_ASAP7_75t_L g896 ( .A1(n_799), .A2(n_579), .B1(n_515), .B2(n_527), .C(n_446), .Y(n_896) );
AOI21xp5_ASAP7_75t_L g897 ( .A1(n_793), .A2(n_809), .B(n_794), .Y(n_897) );
OAI22xp5_ASAP7_75t_L g898 ( .A1(n_814), .A2(n_727), .B1(n_491), .B2(n_681), .Y(n_898) );
AND2x2_ASAP7_75t_L g899 ( .A(n_813), .B(n_515), .Y(n_899) );
AOI21xp5_ASAP7_75t_L g900 ( .A1(n_793), .A2(n_809), .B(n_794), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_813), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_719), .B(n_621), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_719), .B(n_621), .Y(n_903) );
AO21x2_ASAP7_75t_L g904 ( .A1(n_785), .A2(n_788), .B(n_786), .Y(n_904) );
OA21x2_ASAP7_75t_L g905 ( .A1(n_790), .A2(n_782), .B(n_785), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_813), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_813), .Y(n_907) );
AOI221xp5_ASAP7_75t_L g908 ( .A1(n_799), .A2(n_579), .B1(n_515), .B2(n_527), .C(n_446), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_719), .B(n_621), .Y(n_909) );
AOI221xp5_ASAP7_75t_L g910 ( .A1(n_799), .A2(n_579), .B1(n_515), .B2(n_527), .C(n_446), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_719), .B(n_621), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_719), .B(n_621), .Y(n_912) );
BUFx6f_ASAP7_75t_SL g913 ( .A(n_704), .Y(n_913) );
CKINVDCx20_ASAP7_75t_R g914 ( .A(n_801), .Y(n_914) );
AOI21xp5_ASAP7_75t_L g915 ( .A1(n_793), .A2(n_809), .B(n_794), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_813), .Y(n_916) );
INVx3_ASAP7_75t_L g917 ( .A(n_702), .Y(n_917) );
INVx3_ASAP7_75t_L g918 ( .A(n_702), .Y(n_918) );
AOI21xp5_ASAP7_75t_L g919 ( .A1(n_793), .A2(n_809), .B(n_794), .Y(n_919) );
O2A1O1Ixp33_ASAP7_75t_L g920 ( .A1(n_791), .A2(n_818), .B(n_816), .C(n_714), .Y(n_920) );
AOI22xp5_ASAP7_75t_L g921 ( .A1(n_799), .A2(n_438), .B1(n_518), .B2(n_515), .Y(n_921) );
INVx2_ASAP7_75t_L g922 ( .A(n_719), .Y(n_922) );
INVxp67_ASAP7_75t_L g923 ( .A(n_813), .Y(n_923) );
NAND2xp5_ASAP7_75t_L g924 ( .A(n_719), .B(n_621), .Y(n_924) );
CKINVDCx5p33_ASAP7_75t_R g925 ( .A(n_801), .Y(n_925) );
OAI22xp5_ASAP7_75t_L g926 ( .A1(n_814), .A2(n_727), .B1(n_491), .B2(n_681), .Y(n_926) );
OAI22xp5_ASAP7_75t_L g927 ( .A1(n_814), .A2(n_727), .B1(n_491), .B2(n_681), .Y(n_927) );
AO21x2_ASAP7_75t_L g928 ( .A1(n_852), .A2(n_853), .B(n_882), .Y(n_928) );
OR2x6_ASAP7_75t_L g929 ( .A(n_846), .B(n_842), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_877), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_872), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_860), .Y(n_932) );
AO21x2_ASAP7_75t_L g933 ( .A1(n_852), .A2(n_882), .B(n_878), .Y(n_933) );
AND2x2_ASAP7_75t_L g934 ( .A(n_830), .B(n_884), .Y(n_934) );
INVx3_ASAP7_75t_L g935 ( .A(n_842), .Y(n_935) );
HB1xp67_ASAP7_75t_L g936 ( .A(n_923), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_825), .A2(n_927), .B1(n_926), .B2(n_898), .Y(n_937) );
OA21x2_ASAP7_75t_L g938 ( .A1(n_880), .A2(n_883), .B(n_875), .Y(n_938) );
AOI21xp5_ASAP7_75t_L g939 ( .A1(n_895), .A2(n_876), .B(n_843), .Y(n_939) );
BUFx3_ASAP7_75t_L g940 ( .A(n_842), .Y(n_940) );
INVx1_ASAP7_75t_SL g941 ( .A(n_864), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_863), .Y(n_942) );
OAI211xp5_ASAP7_75t_SL g943 ( .A1(n_921), .A2(n_894), .B(n_891), .C(n_910), .Y(n_943) );
AO21x2_ASAP7_75t_L g944 ( .A1(n_824), .A2(n_897), .B(n_919), .Y(n_944) );
INVx1_ASAP7_75t_L g945 ( .A(n_871), .Y(n_945) );
OAI21xp5_ASAP7_75t_L g946 ( .A1(n_866), .A2(n_857), .B(n_854), .Y(n_946) );
INVx3_ASAP7_75t_L g947 ( .A(n_846), .Y(n_947) );
OR2x2_ASAP7_75t_L g948 ( .A(n_887), .B(n_889), .Y(n_948) );
INVx2_ASAP7_75t_L g949 ( .A(n_905), .Y(n_949) );
AO21x2_ASAP7_75t_L g950 ( .A1(n_885), .A2(n_915), .B(n_900), .Y(n_950) );
OR2x6_ASAP7_75t_L g951 ( .A(n_898), .B(n_926), .Y(n_951) );
OR2x6_ASAP7_75t_L g952 ( .A(n_927), .B(n_862), .Y(n_952) );
OAI22xp33_ASAP7_75t_L g953 ( .A1(n_825), .A2(n_908), .B1(n_896), .B2(n_886), .Y(n_953) );
INVx2_ASAP7_75t_SL g954 ( .A(n_864), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_839), .Y(n_955) );
AND2x2_ASAP7_75t_L g956 ( .A(n_901), .B(n_906), .Y(n_956) );
HB1xp67_ASAP7_75t_L g957 ( .A(n_907), .Y(n_957) );
AO21x2_ASAP7_75t_L g958 ( .A1(n_844), .A2(n_829), .B(n_904), .Y(n_958) );
OAI33xp33_ASAP7_75t_L g959 ( .A1(n_920), .A2(n_847), .A3(n_916), .B1(n_849), .B2(n_823), .B3(n_836), .Y(n_959) );
INVx2_ASAP7_75t_L g960 ( .A(n_822), .Y(n_960) );
OAI211xp5_ASAP7_75t_L g961 ( .A1(n_868), .A2(n_833), .B(n_881), .C(n_827), .Y(n_961) );
OAI321xp33_ASAP7_75t_L g962 ( .A1(n_851), .A2(n_856), .A3(n_859), .B1(n_848), .B2(n_835), .C(n_840), .Y(n_962) );
INVx2_ASAP7_75t_L g963 ( .A(n_904), .Y(n_963) );
AOI221xp5_ASAP7_75t_L g964 ( .A1(n_888), .A2(n_912), .B1(n_909), .B2(n_924), .C(n_911), .Y(n_964) );
AND2x2_ASAP7_75t_L g965 ( .A(n_922), .B(n_909), .Y(n_965) );
INVx1_ASAP7_75t_L g966 ( .A(n_879), .Y(n_966) );
NOR2xp33_ASAP7_75t_L g967 ( .A(n_837), .B(n_838), .Y(n_967) );
INVx2_ASAP7_75t_L g968 ( .A(n_829), .Y(n_968) );
AND2x2_ASAP7_75t_L g969 ( .A(n_902), .B(n_903), .Y(n_969) );
OR2x2_ASAP7_75t_L g970 ( .A(n_902), .B(n_924), .Y(n_970) );
AND2x2_ASAP7_75t_L g971 ( .A(n_911), .B(n_912), .Y(n_971) );
AO21x2_ASAP7_75t_L g972 ( .A1(n_869), .A2(n_874), .B(n_855), .Y(n_972) );
AOI21xp5_ASAP7_75t_SL g973 ( .A1(n_867), .A2(n_874), .B(n_834), .Y(n_973) );
INVx1_ASAP7_75t_SL g974 ( .A(n_865), .Y(n_974) );
INVx2_ASAP7_75t_L g975 ( .A(n_870), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_841), .B(n_821), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_834), .Y(n_977) );
AND2x2_ASAP7_75t_L g978 ( .A(n_826), .B(n_892), .Y(n_978) );
CKINVDCx5p33_ASAP7_75t_R g979 ( .A(n_828), .Y(n_979) );
AND2x2_ASAP7_75t_L g980 ( .A(n_892), .B(n_918), .Y(n_980) );
INVx1_ASAP7_75t_SL g981 ( .A(n_914), .Y(n_981) );
OA21x2_ASAP7_75t_L g982 ( .A1(n_917), .A2(n_850), .B(n_913), .Y(n_982) );
OR2x2_ASAP7_75t_L g983 ( .A(n_845), .B(n_925), .Y(n_983) );
OR2x2_ASAP7_75t_L g984 ( .A(n_913), .B(n_873), .Y(n_984) );
AND2x2_ASAP7_75t_L g985 ( .A(n_893), .B(n_831), .Y(n_985) );
INVx2_ASAP7_75t_L g986 ( .A(n_890), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_877), .Y(n_987) );
BUFx2_ASAP7_75t_L g988 ( .A(n_846), .Y(n_988) );
AND2x2_ASAP7_75t_L g989 ( .A(n_830), .B(n_884), .Y(n_989) );
AOI21x1_ASAP7_75t_L g990 ( .A1(n_832), .A2(n_858), .B(n_861), .Y(n_990) );
OAI221xp5_ASAP7_75t_L g991 ( .A1(n_891), .A2(n_894), .B1(n_511), .B2(n_868), .C(n_815), .Y(n_991) );
INVxp67_ASAP7_75t_L g992 ( .A(n_899), .Y(n_992) );
INVx1_ASAP7_75t_L g993 ( .A(n_877), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_877), .Y(n_994) );
NAND2xp33_ASAP7_75t_SL g995 ( .A(n_937), .B(n_988), .Y(n_995) );
HB1xp67_ASAP7_75t_L g996 ( .A(n_931), .Y(n_996) );
AND2x2_ASAP7_75t_L g997 ( .A(n_951), .B(n_945), .Y(n_997) );
NOR2xp33_ASAP7_75t_L g998 ( .A(n_943), .B(n_991), .Y(n_998) );
OR2x2_ASAP7_75t_L g999 ( .A(n_951), .B(n_945), .Y(n_999) );
AO21x2_ASAP7_75t_L g1000 ( .A1(n_939), .A2(n_990), .B(n_946), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g1001 ( .A(n_969), .B(n_971), .Y(n_1001) );
NOR2xp67_ASAP7_75t_SL g1002 ( .A(n_973), .B(n_940), .Y(n_1002) );
INVx2_ASAP7_75t_SL g1003 ( .A(n_982), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_951), .B(n_928), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_951), .B(n_928), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_951), .B(n_928), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_928), .B(n_932), .Y(n_1007) );
AND2x2_ASAP7_75t_L g1008 ( .A(n_932), .B(n_942), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_930), .Y(n_1009) );
AND2x2_ASAP7_75t_L g1010 ( .A(n_942), .B(n_987), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1011 ( .A(n_993), .B(n_994), .Y(n_1011) );
INVx5_ASAP7_75t_L g1012 ( .A(n_929), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_966), .Y(n_1013) );
OR2x2_ASAP7_75t_L g1014 ( .A(n_975), .B(n_970), .Y(n_1014) );
NAND4xp25_ASAP7_75t_L g1015 ( .A(n_964), .B(n_973), .C(n_961), .D(n_967), .Y(n_1015) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_960), .B(n_938), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_960), .B(n_938), .Y(n_1017) );
OR2x2_ASAP7_75t_SL g1018 ( .A(n_982), .B(n_984), .Y(n_1018) );
BUFx2_ASAP7_75t_L g1019 ( .A(n_952), .Y(n_1019) );
INVxp67_ASAP7_75t_SL g1020 ( .A(n_970), .Y(n_1020) );
AND2x2_ASAP7_75t_L g1021 ( .A(n_933), .B(n_949), .Y(n_1021) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_953), .A2(n_959), .B1(n_952), .B2(n_989), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_933), .B(n_952), .Y(n_1023) );
HB1xp67_ASAP7_75t_L g1024 ( .A(n_957), .Y(n_1024) );
INVx2_ASAP7_75t_SL g1025 ( .A(n_982), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_933), .B(n_952), .Y(n_1026) );
HB1xp67_ASAP7_75t_L g1027 ( .A(n_975), .Y(n_1027) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_1004), .B(n_963), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_1001), .B(n_934), .Y(n_1029) );
OR2x2_ASAP7_75t_L g1030 ( .A(n_1020), .B(n_975), .Y(n_1030) );
OAI21xp5_ASAP7_75t_L g1031 ( .A1(n_998), .A2(n_962), .B(n_936), .Y(n_1031) );
NAND2xp5_ASAP7_75t_L g1032 ( .A(n_1001), .B(n_955), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_1004), .B(n_958), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_1005), .B(n_958), .Y(n_1034) );
NOR2x1p5_ASAP7_75t_L g1035 ( .A(n_1020), .B(n_947), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_1005), .B(n_958), .Y(n_1036) );
BUFx2_ASAP7_75t_SL g1037 ( .A(n_1003), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_1005), .B(n_958), .Y(n_1038) );
OR2x2_ASAP7_75t_L g1039 ( .A(n_999), .B(n_972), .Y(n_1039) );
NAND2x1p5_ASAP7_75t_L g1040 ( .A(n_1012), .B(n_982), .Y(n_1040) );
INVx1_ASAP7_75t_L g1041 ( .A(n_1009), .Y(n_1041) );
AND2x4_ASAP7_75t_L g1042 ( .A(n_1007), .B(n_968), .Y(n_1042) );
OR2x2_ASAP7_75t_L g1043 ( .A(n_999), .B(n_972), .Y(n_1043) );
NAND2xp33_ASAP7_75t_L g1044 ( .A(n_1012), .B(n_984), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_1024), .B(n_956), .Y(n_1045) );
AND2x2_ASAP7_75t_L g1046 ( .A(n_1006), .B(n_997), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_1006), .B(n_950), .Y(n_1047) );
AND2x2_ASAP7_75t_L g1048 ( .A(n_997), .B(n_950), .Y(n_1048) );
AOI22xp5_ASAP7_75t_L g1049 ( .A1(n_998), .A2(n_992), .B1(n_965), .B2(n_929), .Y(n_1049) );
INVxp67_ASAP7_75t_SL g1050 ( .A(n_996), .Y(n_1050) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_997), .B(n_950), .Y(n_1051) );
AND2x4_ASAP7_75t_SL g1052 ( .A(n_1003), .B(n_929), .Y(n_1052) );
OR2x2_ASAP7_75t_L g1053 ( .A(n_1027), .B(n_972), .Y(n_1053) );
HB1xp67_ASAP7_75t_L g1054 ( .A(n_996), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_1010), .B(n_944), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_1010), .B(n_944), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_1010), .B(n_944), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1058 ( .A(n_1011), .B(n_944), .Y(n_1058) );
INVx1_ASAP7_75t_L g1059 ( .A(n_1041), .Y(n_1059) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_1048), .B(n_1023), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1041), .Y(n_1061) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_1051), .B(n_1023), .Y(n_1062) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_1051), .B(n_1026), .Y(n_1063) );
INVx1_ASAP7_75t_SL g1064 ( .A(n_1037), .Y(n_1064) );
NOR2xp33_ASAP7_75t_L g1065 ( .A(n_1029), .B(n_974), .Y(n_1065) );
AND2x2_ASAP7_75t_L g1066 ( .A(n_1046), .B(n_1007), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_1047), .B(n_1007), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_1047), .B(n_1016), .Y(n_1068) );
OR2x2_ASAP7_75t_L g1069 ( .A(n_1045), .B(n_1014), .Y(n_1069) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_1055), .B(n_1016), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_1056), .B(n_1017), .Y(n_1071) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_1056), .B(n_1017), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_1057), .B(n_1017), .Y(n_1073) );
AND2x4_ASAP7_75t_L g1074 ( .A(n_1042), .B(n_1021), .Y(n_1074) );
INVxp67_ASAP7_75t_SL g1075 ( .A(n_1050), .Y(n_1075) );
OR2x6_ASAP7_75t_L g1076 ( .A(n_1037), .B(n_1019), .Y(n_1076) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_1058), .B(n_1008), .Y(n_1077) );
AOI21xp33_ASAP7_75t_L g1078 ( .A1(n_1031), .A2(n_1000), .B(n_1002), .Y(n_1078) );
NAND4xp25_ASAP7_75t_L g1079 ( .A(n_1049), .B(n_1015), .C(n_1022), .D(n_995), .Y(n_1079) );
NOR2xp67_ASAP7_75t_SL g1080 ( .A(n_1054), .B(n_1025), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_1033), .B(n_1019), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1059), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_1068), .B(n_1033), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1059), .Y(n_1084) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1061), .Y(n_1085) );
OAI22xp5_ASAP7_75t_L g1086 ( .A1(n_1064), .A2(n_1018), .B1(n_1049), .B2(n_1035), .Y(n_1086) );
NAND2xp5_ASAP7_75t_L g1087 ( .A(n_1077), .B(n_1032), .Y(n_1087) );
OAI21xp5_ASAP7_75t_SL g1088 ( .A1(n_1079), .A2(n_1040), .B(n_1052), .Y(n_1088) );
OR2x2_ASAP7_75t_L g1089 ( .A(n_1067), .B(n_1053), .Y(n_1089) );
NAND2x1p5_ASAP7_75t_L g1090 ( .A(n_1064), .B(n_1025), .Y(n_1090) );
OR2x2_ASAP7_75t_L g1091 ( .A(n_1067), .B(n_1053), .Y(n_1091) );
NOR2xp33_ASAP7_75t_L g1092 ( .A(n_1065), .B(n_983), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_1068), .B(n_1034), .Y(n_1093) );
AND2x4_ASAP7_75t_L g1094 ( .A(n_1074), .B(n_1035), .Y(n_1094) );
OR2x2_ASAP7_75t_L g1095 ( .A(n_1070), .B(n_1030), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1096 ( .A(n_1070), .B(n_1036), .Y(n_1096) );
INVxp67_ASAP7_75t_L g1097 ( .A(n_1075), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_1071), .B(n_1036), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_1071), .B(n_1038), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_1072), .B(n_1028), .Y(n_1100) );
OR2x2_ASAP7_75t_L g1101 ( .A(n_1095), .B(n_1073), .Y(n_1101) );
NOR2xp33_ASAP7_75t_L g1102 ( .A(n_1092), .B(n_1069), .Y(n_1102) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1082), .Y(n_1103) );
AND2x2_ASAP7_75t_L g1104 ( .A(n_1083), .B(n_1066), .Y(n_1104) );
AOI31xp33_ASAP7_75t_L g1105 ( .A1(n_1086), .A2(n_1040), .A3(n_983), .B(n_1078), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1084), .Y(n_1106) );
NAND2xp5_ASAP7_75t_SL g1107 ( .A(n_1094), .B(n_1040), .Y(n_1107) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1084), .Y(n_1108) );
NAND2xp5_ASAP7_75t_SL g1109 ( .A(n_1094), .B(n_1025), .Y(n_1109) );
OAI21xp33_ASAP7_75t_SL g1110 ( .A1(n_1097), .A2(n_1076), .B(n_1078), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1085), .Y(n_1111) );
AOI22xp5_ASAP7_75t_L g1112 ( .A1(n_1088), .A2(n_1002), .B1(n_1081), .B2(n_1074), .Y(n_1112) );
INVxp67_ASAP7_75t_SL g1113 ( .A(n_1090), .Y(n_1113) );
NOR2xp33_ASAP7_75t_L g1114 ( .A(n_1087), .B(n_1069), .Y(n_1114) );
OAI211xp5_ASAP7_75t_SL g1115 ( .A1(n_1110), .A2(n_981), .B(n_941), .C(n_1044), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1103), .Y(n_1116) );
O2A1O1Ixp5_ASAP7_75t_L g1117 ( .A1(n_1107), .A2(n_1080), .B(n_1002), .C(n_1013), .Y(n_1117) );
AOI22xp5_ASAP7_75t_L g1118 ( .A1(n_1102), .A2(n_1063), .B1(n_1062), .B2(n_1060), .Y(n_1118) );
NAND4xp25_ASAP7_75t_SL g1119 ( .A(n_1112), .B(n_1091), .C(n_1089), .D(n_1100), .Y(n_1119) );
NAND2xp5_ASAP7_75t_SL g1120 ( .A(n_1105), .B(n_1090), .Y(n_1120) );
NOR2xp33_ASAP7_75t_L g1121 ( .A(n_1114), .B(n_1093), .Y(n_1121) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1106), .Y(n_1122) );
NOR2x1_ASAP7_75t_L g1123 ( .A(n_1115), .B(n_1107), .Y(n_1123) );
AOI21xp5_ASAP7_75t_L g1124 ( .A1(n_1120), .A2(n_1109), .B(n_1113), .Y(n_1124) );
AOI211xp5_ASAP7_75t_L g1125 ( .A1(n_1119), .A2(n_985), .B(n_986), .C(n_1114), .Y(n_1125) );
NAND4xp75_ASAP7_75t_L g1126 ( .A(n_1117), .B(n_986), .C(n_954), .D(n_1104), .Y(n_1126) );
O2A1O1Ixp33_ASAP7_75t_L g1127 ( .A1(n_1117), .A2(n_954), .B(n_977), .C(n_948), .Y(n_1127) );
OAI211xp5_ASAP7_75t_SL g1128 ( .A1(n_1118), .A2(n_1091), .B(n_1101), .C(n_947), .Y(n_1128) );
NOR2x1_ASAP7_75t_L g1129 ( .A(n_1126), .B(n_940), .Y(n_1129) );
NAND5xp2_ASAP7_75t_L g1130 ( .A(n_1125), .B(n_1121), .C(n_1090), .D(n_988), .E(n_977), .Y(n_1130) );
OAI22xp5_ASAP7_75t_SL g1131 ( .A1(n_1123), .A2(n_979), .B1(n_929), .B2(n_1012), .Y(n_1131) );
NAND4xp25_ASAP7_75t_SL g1132 ( .A(n_1124), .B(n_1096), .C(n_1098), .D(n_1099), .Y(n_1132) );
NOR3xp33_ASAP7_75t_SL g1133 ( .A(n_1131), .B(n_1128), .C(n_1127), .Y(n_1133) );
OR2x2_ASAP7_75t_L g1134 ( .A(n_1132), .B(n_1116), .Y(n_1134) );
AND2x4_ASAP7_75t_L g1135 ( .A(n_1129), .B(n_1122), .Y(n_1135) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1134), .Y(n_1136) );
AOI22xp5_ASAP7_75t_L g1137 ( .A1(n_1136), .A2(n_1133), .B1(n_1135), .B2(n_1130), .Y(n_1137) );
CKINVDCx20_ASAP7_75t_R g1138 ( .A(n_1137), .Y(n_1138) );
OAI22xp5_ASAP7_75t_L g1139 ( .A1(n_1138), .A2(n_1012), .B1(n_1111), .B2(n_1108), .Y(n_1139) );
OAI21xp5_ASAP7_75t_L g1140 ( .A1(n_1139), .A2(n_935), .B(n_978), .Y(n_1140) );
AO21x2_ASAP7_75t_L g1141 ( .A1(n_1140), .A2(n_980), .B(n_976), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g1142 ( .A1(n_1141), .A2(n_1074), .B1(n_1043), .B2(n_1039), .Y(n_1142) );
endmodule