module real_aes_16112_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_571;
wire n_549;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1441;
wire n_875;
wire n_951;
wire n_1199;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1600;
wire n_805;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1583;
wire n_360;
wire n_1250;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1648;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_1606;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1620;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_334;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1580;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1175;
wire n_1170;
wire n_778;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_1268;
wire n_852;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1603;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1619;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1654;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1252;
wire n_1647;
wire n_430;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
OAI22xp5_ASAP7_75t_L g889 ( .A1(n_0), .A2(n_51), .B1(n_603), .B2(n_890), .Y(n_889) );
INVxp67_ASAP7_75t_SL g917 ( .A(n_0), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g1327 ( .A1(n_1), .A2(n_82), .B1(n_1302), .B2(n_1305), .Y(n_1327) );
OAI22xp33_ASAP7_75t_L g1155 ( .A1(n_2), .A2(n_279), .B1(n_449), .B2(n_458), .Y(n_1155) );
OAI22xp33_ASAP7_75t_SL g1165 ( .A1(n_2), .A2(n_279), .B1(n_468), .B2(n_951), .Y(n_1165) );
INVx1_ASAP7_75t_L g322 ( .A(n_3), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_3), .B(n_332), .Y(n_402) );
AND2x2_ASAP7_75t_L g1518 ( .A(n_3), .B(n_219), .Y(n_1518) );
AND2x2_ASAP7_75t_L g1541 ( .A(n_3), .B(n_457), .Y(n_1541) );
AOI22xp33_ASAP7_75t_L g1204 ( .A1(n_4), .A2(n_224), .B1(n_996), .B2(n_1205), .Y(n_1204) );
AOI22xp33_ASAP7_75t_L g1223 ( .A1(n_4), .A2(n_174), .B1(n_1224), .B2(n_1225), .Y(n_1223) );
INVx1_ASAP7_75t_L g727 ( .A(n_5), .Y(n_727) );
INVx1_ASAP7_75t_L g1031 ( .A(n_6), .Y(n_1031) );
INVx1_ASAP7_75t_L g970 ( .A(n_7), .Y(n_970) );
INVx1_ASAP7_75t_L g1195 ( .A(n_8), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g1230 ( .A1(n_8), .A2(n_224), .B1(n_1225), .B2(n_1231), .Y(n_1230) );
OAI22xp5_ASAP7_75t_L g1032 ( .A1(n_9), .A2(n_137), .B1(n_324), .B2(n_458), .Y(n_1032) );
OAI22xp5_ASAP7_75t_L g1034 ( .A1(n_9), .A2(n_137), .B1(n_469), .B2(n_1035), .Y(n_1034) );
CKINVDCx5p33_ASAP7_75t_R g793 ( .A(n_10), .Y(n_793) );
INVx1_ASAP7_75t_L g866 ( .A(n_11), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_12), .A2(n_40), .B1(n_615), .B2(n_640), .Y(n_639) );
OAI22xp33_ASAP7_75t_L g659 ( .A1(n_12), .A2(n_40), .B1(n_324), .B2(n_458), .Y(n_659) );
CKINVDCx5p33_ASAP7_75t_R g1049 ( .A(n_13), .Y(n_1049) );
OAI22xp33_ASAP7_75t_L g1162 ( .A1(n_14), .A2(n_261), .B1(n_532), .B2(n_1163), .Y(n_1162) );
OAI22xp33_ASAP7_75t_L g1169 ( .A1(n_14), .A2(n_261), .B1(n_489), .B2(n_490), .Y(n_1169) );
OAI22xp5_ASAP7_75t_L g766 ( .A1(n_15), .A2(n_275), .B1(n_656), .B2(n_706), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_15), .A2(n_275), .B1(n_630), .B2(n_631), .Y(n_769) );
INVx2_ASAP7_75t_L g350 ( .A(n_16), .Y(n_350) );
INVx1_ASAP7_75t_L g1630 ( .A(n_17), .Y(n_1630) );
INVx1_ASAP7_75t_L g1631 ( .A(n_18), .Y(n_1631) );
XNOR2xp5_ASAP7_75t_L g856 ( .A(n_19), .B(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g556 ( .A(n_20), .Y(n_556) );
INVx1_ASAP7_75t_L g1113 ( .A(n_21), .Y(n_1113) );
INVx1_ASAP7_75t_L g964 ( .A(n_22), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g1253 ( .A1(n_23), .A2(n_163), .B1(n_1254), .B2(n_1256), .Y(n_1253) );
AOI22xp33_ASAP7_75t_SL g1277 ( .A1(n_23), .A2(n_121), .B1(n_1278), .B2(n_1279), .Y(n_1277) );
AOI221xp5_ASAP7_75t_L g1612 ( .A1(n_24), .A2(n_78), .B1(n_802), .B2(n_1262), .C(n_1613), .Y(n_1612) );
AOI22xp33_ASAP7_75t_L g1652 ( .A1(n_24), .A2(n_39), .B1(n_1279), .B2(n_1653), .Y(n_1652) );
AOI22xp33_ASAP7_75t_SL g1000 ( .A1(n_25), .A2(n_150), .B1(n_914), .B2(n_996), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_25), .A2(n_181), .B1(n_521), .B2(n_1020), .Y(n_1019) );
INVx1_ASAP7_75t_L g548 ( .A(n_26), .Y(n_548) );
OAI211xp5_ASAP7_75t_L g594 ( .A1(n_27), .A2(n_595), .B(n_598), .C(n_605), .Y(n_594) );
INVx1_ASAP7_75t_L g628 ( .A(n_27), .Y(n_628) );
INVx1_ASAP7_75t_L g339 ( .A(n_28), .Y(n_339) );
OAI22xp5_ASAP7_75t_L g946 ( .A1(n_29), .A2(n_278), .B1(n_532), .B2(n_947), .Y(n_946) );
OAI22xp33_ASAP7_75t_L g957 ( .A1(n_29), .A2(n_278), .B1(n_489), .B2(n_490), .Y(n_957) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_30), .Y(n_318) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_30), .B(n_316), .Y(n_1296) );
OAI22xp33_ASAP7_75t_SL g705 ( .A1(n_31), .A2(n_155), .B1(n_656), .B2(n_706), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_31), .A2(n_155), .B1(n_630), .B2(n_710), .Y(n_709) );
OAI222xp33_ASAP7_75t_L g1244 ( .A1(n_32), .A2(n_178), .B1(n_301), .B2(n_920), .C1(n_921), .C2(n_1245), .Y(n_1244) );
OAI222xp33_ASAP7_75t_L g1285 ( .A1(n_32), .A2(n_178), .B1(n_301), .B2(n_603), .C1(n_735), .C2(n_890), .Y(n_1285) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_33), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g1326 ( .A1(n_34), .A2(n_57), .B1(n_1295), .B2(n_1312), .Y(n_1326) );
INVx1_ASAP7_75t_L g1543 ( .A(n_35), .Y(n_1543) );
AOI22xp5_ASAP7_75t_L g1508 ( .A1(n_36), .A2(n_42), .B1(n_1509), .B2(n_1510), .Y(n_1508) );
AOI22xp33_ASAP7_75t_L g1561 ( .A1(n_36), .A2(n_146), .B1(n_1020), .B2(n_1562), .Y(n_1561) );
INVx1_ASAP7_75t_L g829 ( .A(n_37), .Y(n_829) );
INVxp67_ASAP7_75t_SL g888 ( .A(n_38), .Y(n_888) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_38), .A2(n_51), .B1(n_920), .B2(n_921), .Y(n_919) );
AOI221xp5_ASAP7_75t_L g1614 ( .A1(n_39), .A2(n_64), .B1(n_802), .B2(n_1262), .C(n_1615), .Y(n_1614) );
OAI22xp33_ASAP7_75t_L g948 ( .A1(n_41), .A2(n_234), .B1(n_449), .B2(n_593), .Y(n_948) );
OAI22xp33_ASAP7_75t_SL g950 ( .A1(n_41), .A2(n_234), .B1(n_468), .B2(n_951), .Y(n_950) );
AOI22xp33_ASAP7_75t_SL g1556 ( .A1(n_42), .A2(n_156), .B1(n_1227), .B2(n_1261), .Y(n_1556) );
INVx1_ASAP7_75t_L g664 ( .A(n_43), .Y(n_664) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_44), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g1192 ( .A(n_45), .Y(n_1192) );
INVx1_ASAP7_75t_L g1142 ( .A(n_46), .Y(n_1142) );
AOI22xp33_ASAP7_75t_SL g988 ( .A1(n_47), .A2(n_181), .B1(n_989), .B2(n_992), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_47), .A2(n_150), .B1(n_1004), .B2(n_1005), .Y(n_1003) );
INVx1_ASAP7_75t_L g1618 ( .A(n_48), .Y(n_1618) );
AOI22xp33_ASAP7_75t_SL g1647 ( .A1(n_48), .A2(n_227), .B1(n_996), .B2(n_1648), .Y(n_1647) );
AOI22xp5_ASAP7_75t_L g1311 ( .A1(n_49), .A2(n_102), .B1(n_1295), .B2(n_1312), .Y(n_1311) );
AOI22xp5_ASAP7_75t_L g1332 ( .A1(n_50), .A2(n_226), .B1(n_1295), .B2(n_1312), .Y(n_1332) );
INVx1_ASAP7_75t_L g1120 ( .A(n_52), .Y(n_1120) );
OAI211xp5_ASAP7_75t_SL g641 ( .A1(n_53), .A2(n_620), .B(n_622), .C(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g654 ( .A(n_53), .Y(n_654) );
OAI22xp33_ASAP7_75t_L g645 ( .A1(n_54), .A2(n_159), .B1(n_630), .B2(n_631), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_54), .A2(n_159), .B1(n_656), .B2(n_657), .Y(n_655) );
INVx1_ASAP7_75t_L g892 ( .A(n_55), .Y(n_892) );
OAI222xp33_ASAP7_75t_L g1181 ( .A1(n_56), .A2(n_165), .B1(n_443), .B2(n_450), .C1(n_1182), .C2(n_1183), .Y(n_1181) );
OAI222xp33_ASAP7_75t_L g1211 ( .A1(n_56), .A2(n_165), .B1(n_192), .B2(n_1212), .C1(n_1213), .C2(n_1214), .Y(n_1211) );
INVx1_ASAP7_75t_L g969 ( .A(n_58), .Y(n_969) );
OAI22xp33_ASAP7_75t_L g847 ( .A1(n_59), .A2(n_263), .B1(n_324), .B2(n_458), .Y(n_847) );
OAI22xp33_ASAP7_75t_L g849 ( .A1(n_59), .A2(n_263), .B1(n_640), .B2(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g604 ( .A(n_60), .Y(n_604) );
OAI211xp5_ASAP7_75t_L g619 ( .A1(n_60), .A2(n_620), .B(n_622), .C(n_623), .Y(n_619) );
INVx1_ASAP7_75t_L g1141 ( .A(n_61), .Y(n_1141) );
AOI221xp5_ASAP7_75t_L g1512 ( .A1(n_62), .A2(n_291), .B1(n_912), .B2(n_980), .C(n_1513), .Y(n_1512) );
AOI221xp5_ASAP7_75t_L g1559 ( .A1(n_62), .A2(n_258), .B1(n_674), .B2(n_1252), .C(n_1560), .Y(n_1559) );
INVx1_ASAP7_75t_L g1026 ( .A(n_63), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g1649 ( .A1(n_64), .A2(n_78), .B1(n_1200), .B2(n_1650), .Y(n_1649) );
CKINVDCx5p33_ASAP7_75t_R g1059 ( .A(n_65), .Y(n_1059) );
INVx1_ASAP7_75t_L g897 ( .A(n_66), .Y(n_897) );
INVx1_ASAP7_75t_L g677 ( .A(n_67), .Y(n_677) );
INVxp67_ASAP7_75t_SL g1548 ( .A(n_68), .Y(n_1548) );
OAI22xp5_ASAP7_75t_L g1563 ( .A1(n_68), .A2(n_300), .B1(n_1564), .B2(n_1568), .Y(n_1563) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_69), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g1339 ( .A1(n_70), .A2(n_208), .B1(n_1295), .B2(n_1312), .Y(n_1339) );
OAI211xp5_ASAP7_75t_L g941 ( .A1(n_71), .A2(n_432), .B(n_942), .C(n_943), .Y(n_941) );
INVx1_ASAP7_75t_L g954 ( .A(n_71), .Y(n_954) );
INVx1_ASAP7_75t_L g883 ( .A(n_72), .Y(n_883) );
AOI22xp5_ASAP7_75t_L g1320 ( .A1(n_73), .A2(n_217), .B1(n_1302), .B2(n_1305), .Y(n_1320) );
INVx1_ASAP7_75t_L g747 ( .A(n_74), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g1321 ( .A1(n_75), .A2(n_93), .B1(n_1295), .B2(n_1322), .Y(n_1321) );
AO22x1_ASAP7_75t_L g1301 ( .A1(n_76), .A2(n_228), .B1(n_1302), .B2(n_1305), .Y(n_1301) );
XNOR2xp5_ASAP7_75t_L g496 ( .A(n_77), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g1623 ( .A(n_79), .Y(n_1623) );
OAI22xp5_ASAP7_75t_L g1639 ( .A1(n_79), .A2(n_173), .B1(n_468), .B2(n_489), .Y(n_1639) );
INVx1_ASAP7_75t_L g561 ( .A(n_80), .Y(n_561) );
INVx1_ASAP7_75t_L g447 ( .A(n_81), .Y(n_447) );
OAI211xp5_ASAP7_75t_L g472 ( .A1(n_81), .A2(n_473), .B(n_476), .C(n_480), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g1069 ( .A1(n_83), .A2(n_232), .B1(n_449), .B2(n_947), .Y(n_1069) );
OAI22xp5_ASAP7_75t_SL g1078 ( .A1(n_83), .A2(n_115), .B1(n_468), .B2(n_490), .Y(n_1078) );
INVx1_ASAP7_75t_L g676 ( .A(n_84), .Y(n_676) );
CKINVDCx5p33_ASAP7_75t_R g1073 ( .A(n_85), .Y(n_1073) );
INVx1_ASAP7_75t_L g973 ( .A(n_86), .Y(n_973) );
CKINVDCx5p33_ASAP7_75t_R g1048 ( .A(n_87), .Y(n_1048) );
OAI22xp33_ASAP7_75t_L g592 ( .A1(n_88), .A2(n_148), .B1(n_324), .B2(n_593), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_88), .A2(n_148), .B1(n_615), .B2(n_617), .Y(n_614) );
INVx1_ASAP7_75t_L g1633 ( .A(n_89), .Y(n_1633) );
AOI22xp33_ASAP7_75t_SL g1001 ( .A1(n_90), .A2(n_309), .B1(n_989), .B2(n_992), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_90), .A2(n_91), .B1(n_1011), .B2(n_1016), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_91), .A2(n_281), .B1(n_994), .B2(n_996), .Y(n_993) );
INVx1_ASAP7_75t_L g1134 ( .A(n_92), .Y(n_1134) );
CKINVDCx5p33_ASAP7_75t_R g513 ( .A(n_94), .Y(n_513) );
INVx1_ASAP7_75t_L g868 ( .A(n_95), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_95), .A2(n_254), .B1(n_907), .B2(n_914), .Y(n_913) );
CKINVDCx5p33_ASAP7_75t_R g1055 ( .A(n_96), .Y(n_1055) );
INVx1_ASAP7_75t_L g945 ( .A(n_97), .Y(n_945) );
INVx1_ASAP7_75t_L g835 ( .A(n_98), .Y(n_835) );
OAI211xp5_ASAP7_75t_L g430 ( .A1(n_99), .A2(n_431), .B(n_432), .C(n_438), .Y(n_430) );
INVx1_ASAP7_75t_L g487 ( .A(n_99), .Y(n_487) );
INVx1_ASAP7_75t_L g316 ( .A(n_100), .Y(n_316) );
INVx1_ASAP7_75t_L g879 ( .A(n_101), .Y(n_879) );
AO221x2_ASAP7_75t_L g1393 ( .A1(n_103), .A2(n_292), .B1(n_1302), .B2(n_1305), .C(n_1394), .Y(n_1393) );
OAI22xp33_ASAP7_75t_L g454 ( .A1(n_104), .A2(n_259), .B1(n_455), .B2(n_458), .Y(n_454) );
OAI22xp33_ASAP7_75t_L g488 ( .A1(n_104), .A2(n_143), .B1(n_489), .B2(n_490), .Y(n_488) );
XOR2xp5_ASAP7_75t_L g1174 ( .A(n_105), .B(n_1175), .Y(n_1174) );
INVx1_ASAP7_75t_L g703 ( .A(n_106), .Y(n_703) );
INVx1_ASAP7_75t_L g823 ( .A(n_107), .Y(n_823) );
OAI22xp33_ASAP7_75t_L g1584 ( .A1(n_108), .A2(n_153), .B1(n_1585), .B2(n_1588), .Y(n_1584) );
INVxp67_ASAP7_75t_SL g1593 ( .A(n_108), .Y(n_1593) );
INVx1_ASAP7_75t_L g864 ( .A(n_109), .Y(n_864) );
INVx1_ASAP7_75t_L g732 ( .A(n_110), .Y(n_732) );
INVx1_ASAP7_75t_L g1145 ( .A(n_111), .Y(n_1145) );
OAI22xp5_ASAP7_75t_L g1241 ( .A1(n_112), .A2(n_222), .B1(n_1242), .B2(n_1243), .Y(n_1241) );
OAI22xp5_ASAP7_75t_L g1284 ( .A1(n_112), .A2(n_222), .B1(n_609), .B2(n_899), .Y(n_1284) );
INVx1_ASAP7_75t_L g1116 ( .A(n_113), .Y(n_1116) );
OAI22xp33_ASAP7_75t_SL g1075 ( .A1(n_114), .A2(n_115), .B1(n_532), .B2(n_593), .Y(n_1075) );
OAI22xp5_ASAP7_75t_L g1082 ( .A1(n_114), .A2(n_120), .B1(n_1083), .B2(n_1084), .Y(n_1082) );
INVx1_ASAP7_75t_L g681 ( .A(n_116), .Y(n_681) );
INVx1_ASAP7_75t_L g1119 ( .A(n_117), .Y(n_1119) );
INVx1_ASAP7_75t_L g1158 ( .A(n_118), .Y(n_1158) );
CKINVDCx5p33_ASAP7_75t_R g789 ( .A(n_119), .Y(n_789) );
INVx1_ASAP7_75t_L g1074 ( .A(n_120), .Y(n_1074) );
AOI22xp33_ASAP7_75t_L g1260 ( .A1(n_121), .A2(n_252), .B1(n_1261), .B2(n_1262), .Y(n_1260) );
INVx1_ASAP7_75t_L g1117 ( .A(n_122), .Y(n_1117) );
AO22x1_ASAP7_75t_L g1317 ( .A1(n_123), .A2(n_297), .B1(n_1302), .B2(n_1305), .Y(n_1317) );
INVx1_ASAP7_75t_L g550 ( .A(n_124), .Y(n_550) );
OAI22xp33_ASAP7_75t_L g531 ( .A1(n_125), .A2(n_169), .B1(n_458), .B2(n_532), .Y(n_531) );
OAI22xp33_ASAP7_75t_L g538 ( .A1(n_125), .A2(n_162), .B1(n_489), .B2(n_490), .Y(n_538) );
CKINVDCx5p33_ASAP7_75t_R g511 ( .A(n_126), .Y(n_511) );
CKINVDCx5p33_ASAP7_75t_R g792 ( .A(n_127), .Y(n_792) );
CKINVDCx5p33_ASAP7_75t_R g502 ( .A(n_128), .Y(n_502) );
CKINVDCx5p33_ASAP7_75t_R g1052 ( .A(n_129), .Y(n_1052) );
OAI211xp5_ASAP7_75t_L g701 ( .A1(n_130), .A2(n_648), .B(n_651), .C(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g717 ( .A(n_130), .Y(n_717) );
INVx1_ASAP7_75t_L g704 ( .A(n_131), .Y(n_704) );
OAI211xp5_ASAP7_75t_L g712 ( .A1(n_131), .A2(n_476), .B(n_713), .C(n_715), .Y(n_712) );
INVx1_ASAP7_75t_L g669 ( .A(n_132), .Y(n_669) );
INVx1_ASAP7_75t_L g1136 ( .A(n_133), .Y(n_1136) );
AOI221xp5_ASAP7_75t_L g1525 ( .A1(n_134), .A2(n_146), .B1(n_1510), .B2(n_1526), .C(n_1528), .Y(n_1525) );
AOI221xp5_ASAP7_75t_L g1557 ( .A1(n_134), .A2(n_291), .B1(n_396), .B2(n_918), .C(n_1558), .Y(n_1557) );
INVx1_ASAP7_75t_L g643 ( .A(n_135), .Y(n_643) );
INVx1_ASAP7_75t_L g563 ( .A(n_136), .Y(n_563) );
INVx1_ASAP7_75t_L g729 ( .A(n_138), .Y(n_729) );
OAI211xp5_ASAP7_75t_L g842 ( .A1(n_139), .A2(n_650), .B(n_651), .C(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g854 ( .A(n_139), .Y(n_854) );
XNOR2xp5_ASAP7_75t_L g1607 ( .A(n_140), .B(n_1608), .Y(n_1607) );
INVx1_ASAP7_75t_L g844 ( .A(n_141), .Y(n_844) );
INVx1_ASAP7_75t_L g1030 ( .A(n_142), .Y(n_1030) );
OAI22xp33_ASAP7_75t_L g448 ( .A1(n_143), .A2(n_236), .B1(n_449), .B2(n_451), .Y(n_448) );
INVx1_ASAP7_75t_L g529 ( .A(n_144), .Y(n_529) );
OAI211xp5_ASAP7_75t_L g535 ( .A1(n_144), .A2(n_473), .B(n_476), .C(n_536), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_145), .Y(n_352) );
AO22x1_ASAP7_75t_L g1294 ( .A1(n_147), .A2(n_298), .B1(n_1295), .B2(n_1299), .Y(n_1294) );
CKINVDCx16_ASAP7_75t_R g1395 ( .A(n_149), .Y(n_1395) );
INVx1_ASAP7_75t_L g1114 ( .A(n_151), .Y(n_1114) );
OAI22xp5_ASAP7_75t_L g846 ( .A1(n_152), .A2(n_251), .B1(n_656), .B2(n_706), .Y(n_846) );
OAI22xp33_ASAP7_75t_L g855 ( .A1(n_152), .A2(n_251), .B1(n_630), .B2(n_710), .Y(n_855) );
INVxp67_ASAP7_75t_SL g1537 ( .A(n_153), .Y(n_1537) );
OAI211xp5_ASAP7_75t_L g525 ( .A1(n_154), .A2(n_431), .B(n_432), .C(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g537 ( .A(n_154), .Y(n_537) );
INVx1_ASAP7_75t_L g1529 ( .A(n_156), .Y(n_1529) );
INVx1_ASAP7_75t_L g746 ( .A(n_157), .Y(n_746) );
INVx1_ASAP7_75t_L g834 ( .A(n_158), .Y(n_834) );
OAI22xp33_ASAP7_75t_L g530 ( .A1(n_160), .A2(n_162), .B1(n_449), .B2(n_451), .Y(n_530) );
OAI22xp33_ASAP7_75t_L g534 ( .A1(n_160), .A2(n_169), .B1(n_468), .B2(n_469), .Y(n_534) );
INVx1_ASAP7_75t_L g644 ( .A(n_161), .Y(n_644) );
OAI211xp5_ASAP7_75t_L g647 ( .A1(n_161), .A2(n_648), .B(n_651), .C(n_652), .Y(n_647) );
AOI22xp33_ASAP7_75t_SL g1269 ( .A1(n_163), .A2(n_252), .B1(n_1270), .B2(n_1274), .Y(n_1269) );
INVx1_ASAP7_75t_L g818 ( .A(n_164), .Y(n_818) );
INVx1_ASAP7_75t_L g1110 ( .A(n_166), .Y(n_1110) );
INVx2_ASAP7_75t_L g1298 ( .A(n_167), .Y(n_1298) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_167), .B(n_260), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_167), .B(n_1304), .Y(n_1306) );
AO22x2_ASAP7_75t_L g1128 ( .A1(n_168), .A2(n_1129), .B1(n_1170), .B2(n_1171), .Y(n_1128) );
INVx1_ASAP7_75t_L g1170 ( .A(n_168), .Y(n_1170) );
CKINVDCx5p33_ASAP7_75t_R g507 ( .A(n_170), .Y(n_507) );
CKINVDCx5p33_ASAP7_75t_R g1054 ( .A(n_171), .Y(n_1054) );
INVx1_ASAP7_75t_L g666 ( .A(n_172), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g1627 ( .A1(n_173), .A2(n_243), .B1(n_532), .B2(n_947), .Y(n_1627) );
INVx1_ASAP7_75t_L g1196 ( .A(n_174), .Y(n_1196) );
AOI22xp33_ASAP7_75t_L g1258 ( .A1(n_175), .A2(n_286), .B1(n_1249), .B2(n_1259), .Y(n_1258) );
AOI22xp33_ASAP7_75t_L g1276 ( .A1(n_175), .A2(n_213), .B1(n_1270), .B2(n_1274), .Y(n_1276) );
XNOR2x2_ASAP7_75t_L g542 ( .A(n_176), .B(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g1096 ( .A(n_177), .Y(n_1096) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_179), .Y(n_379) );
INVx1_ASAP7_75t_L g944 ( .A(n_180), .Y(n_944) );
XOR2x2_ASAP7_75t_L g938 ( .A(n_182), .B(n_939), .Y(n_938) );
CKINVDCx5p33_ASAP7_75t_R g763 ( .A(n_183), .Y(n_763) );
OAI211xp5_ASAP7_75t_L g1177 ( .A1(n_184), .A2(n_1178), .B(n_1179), .C(n_1187), .Y(n_1177) );
INVx1_ASAP7_75t_L g1217 ( .A(n_184), .Y(n_1217) );
INVx1_ASAP7_75t_L g824 ( .A(n_185), .Y(n_824) );
OAI22xp33_ASAP7_75t_L g700 ( .A1(n_186), .A2(n_253), .B1(n_324), .B2(n_458), .Y(n_700) );
OAI22xp33_ASAP7_75t_L g718 ( .A1(n_186), .A2(n_253), .B1(n_719), .B2(n_721), .Y(n_718) );
INVx2_ASAP7_75t_L g349 ( .A(n_187), .Y(n_349) );
INVx1_ASAP7_75t_L g397 ( .A(n_187), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g1567 ( .A(n_187), .B(n_350), .Y(n_1567) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_188), .Y(n_358) );
OAI22xp33_ASAP7_75t_L g1092 ( .A1(n_189), .A2(n_240), .B1(n_532), .B2(n_947), .Y(n_1092) );
OAI22xp5_ASAP7_75t_SL g1099 ( .A1(n_189), .A2(n_211), .B1(n_468), .B2(n_489), .Y(n_1099) );
XOR2xp5_ASAP7_75t_L g1234 ( .A(n_190), .B(n_1235), .Y(n_1234) );
INVx1_ASAP7_75t_L g1186 ( .A(n_191), .Y(n_1186) );
OAI22xp5_ASAP7_75t_L g1215 ( .A1(n_191), .A2(n_218), .B1(n_489), .B2(n_490), .Y(n_1215) );
INVx1_ASAP7_75t_L g1180 ( .A(n_192), .Y(n_1180) );
BUFx3_ASAP7_75t_L g355 ( .A(n_193), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_194), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g514 ( .A(n_195), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g790 ( .A(n_196), .Y(n_790) );
XOR2xp5_ASAP7_75t_L g813 ( .A(n_197), .B(n_814), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g1340 ( .A1(n_197), .A2(n_199), .B1(n_1302), .B2(n_1305), .Y(n_1340) );
AOI22xp33_ASAP7_75t_L g1248 ( .A1(n_198), .A2(n_213), .B1(n_1249), .B2(n_1252), .Y(n_1248) );
AOI22xp33_ASAP7_75t_L g1266 ( .A1(n_198), .A2(n_286), .B1(n_1267), .B2(n_1268), .Y(n_1266) );
INVx1_ASAP7_75t_L g872 ( .A(n_200), .Y(n_872) );
INVx1_ASAP7_75t_L g765 ( .A(n_201), .Y(n_765) );
OAI211xp5_ASAP7_75t_L g770 ( .A1(n_201), .A2(n_476), .B(n_771), .C(n_773), .Y(n_770) );
INVx1_ASAP7_75t_L g1029 ( .A(n_202), .Y(n_1029) );
INVx1_ASAP7_75t_L g1191 ( .A(n_203), .Y(n_1191) );
NAND2xp5_ASAP7_75t_L g1226 ( .A(n_203), .B(n_1227), .Y(n_1226) );
INVx1_ASAP7_75t_L g1159 ( .A(n_204), .Y(n_1159) );
INVx1_ASAP7_75t_L g819 ( .A(n_205), .Y(n_819) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_206), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_207), .Y(n_367) );
INVx1_ASAP7_75t_L g734 ( .A(n_209), .Y(n_734) );
INVx1_ASAP7_75t_L g1095 ( .A(n_210), .Y(n_1095) );
OAI22xp33_ASAP7_75t_L g1097 ( .A1(n_211), .A2(n_245), .B1(n_449), .B2(n_593), .Y(n_1097) );
CKINVDCx5p33_ASAP7_75t_R g787 ( .A(n_212), .Y(n_787) );
INVx1_ASAP7_75t_L g877 ( .A(n_214), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_214), .A2(n_262), .B1(n_905), .B2(n_907), .Y(n_904) );
INVx1_ASAP7_75t_L g1133 ( .A(n_215), .Y(n_1133) );
INVx1_ASAP7_75t_L g966 ( .A(n_216), .Y(n_966) );
XOR2xp5_ASAP7_75t_L g1043 ( .A(n_217), .B(n_1044), .Y(n_1043) );
INVx1_ASAP7_75t_L g1188 ( .A(n_218), .Y(n_1188) );
BUFx3_ASAP7_75t_L g332 ( .A(n_219), .Y(n_332) );
INVx1_ASAP7_75t_L g457 ( .A(n_219), .Y(n_457) );
INVx1_ASAP7_75t_L g601 ( .A(n_220), .Y(n_601) );
CKINVDCx20_ASAP7_75t_R g1397 ( .A(n_221), .Y(n_1397) );
XOR2x2_ASAP7_75t_L g636 ( .A(n_223), .B(n_637), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g1331 ( .A1(n_223), .A2(n_233), .B1(n_1302), .B2(n_1305), .Y(n_1331) );
INVx1_ASAP7_75t_L g961 ( .A(n_225), .Y(n_961) );
AOI22xp5_ASAP7_75t_L g1611 ( .A1(n_227), .A2(n_249), .B1(n_1038), .B2(n_1231), .Y(n_1611) );
INVx1_ASAP7_75t_L g571 ( .A(n_229), .Y(n_571) );
INVx1_ASAP7_75t_L g1239 ( .A(n_230), .Y(n_1239) );
OAI211xp5_ASAP7_75t_L g1093 ( .A1(n_231), .A2(n_432), .B(n_735), .C(n_1094), .Y(n_1093) );
INVx1_ASAP7_75t_L g1104 ( .A(n_231), .Y(n_1104) );
NOR2xp33_ASAP7_75t_L g1077 ( .A(n_232), .B(n_489), .Y(n_1077) );
CKINVDCx5p33_ASAP7_75t_R g1058 ( .A(n_235), .Y(n_1058) );
OAI22xp33_ASAP7_75t_L g467 ( .A1(n_236), .A2(n_259), .B1(n_468), .B2(n_469), .Y(n_467) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_237), .Y(n_504) );
XOR2x2_ASAP7_75t_L g697 ( .A(n_238), .B(n_698), .Y(n_697) );
XOR2x2_ASAP7_75t_L g984 ( .A(n_239), .B(n_985), .Y(n_984) );
AOI22xp5_ASAP7_75t_L g1310 ( .A1(n_239), .A2(n_305), .B1(n_1302), .B2(n_1305), .Y(n_1310) );
OAI22xp33_ASAP7_75t_L g1105 ( .A1(n_240), .A2(n_245), .B1(n_469), .B2(n_490), .Y(n_1105) );
AO22x1_ASAP7_75t_L g1316 ( .A1(n_241), .A2(n_248), .B1(n_1295), .B2(n_1312), .Y(n_1316) );
INVx1_ASAP7_75t_L g1596 ( .A(n_241), .Y(n_1596) );
AOI22xp33_ASAP7_75t_L g1602 ( .A1(n_241), .A2(n_1603), .B1(n_1606), .B2(n_1654), .Y(n_1602) );
INVx1_ASAP7_75t_L g1027 ( .A(n_242), .Y(n_1027) );
OAI22xp5_ASAP7_75t_L g1643 ( .A1(n_243), .A2(n_280), .B1(n_469), .B2(n_490), .Y(n_1643) );
INVx1_ASAP7_75t_L g357 ( .A(n_244), .Y(n_357) );
INVx1_ASAP7_75t_L g364 ( .A(n_244), .Y(n_364) );
INVx1_ASAP7_75t_L g570 ( .A(n_246), .Y(n_570) );
INVx1_ASAP7_75t_L g554 ( .A(n_247), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g1651 ( .A1(n_249), .A2(n_283), .B1(n_1200), .B2(n_1650), .Y(n_1651) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_250), .A2(n_296), .B1(n_609), .B2(n_610), .Y(n_608) );
OAI22xp33_ASAP7_75t_L g629 ( .A1(n_250), .A2(n_296), .B1(n_630), .B2(n_631), .Y(n_629) );
INVx1_ASAP7_75t_L g875 ( .A(n_254), .Y(n_875) );
OAI22xp33_ASAP7_75t_L g767 ( .A1(n_255), .A2(n_257), .B1(n_324), .B2(n_458), .Y(n_767) );
OAI22xp33_ASAP7_75t_L g775 ( .A1(n_255), .A2(n_257), .B1(n_640), .B2(n_719), .Y(n_775) );
INVx1_ASAP7_75t_L g671 ( .A(n_256), .Y(n_671) );
INVx1_ASAP7_75t_L g1530 ( .A(n_258), .Y(n_1530) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_260), .B(n_1298), .Y(n_1297) );
INVx1_ASAP7_75t_L g1304 ( .A(n_260), .Y(n_1304) );
INVx1_ASAP7_75t_L g861 ( .A(n_262), .Y(n_861) );
INVx1_ASAP7_75t_L g962 ( .A(n_264), .Y(n_962) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_265), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g779 ( .A(n_266), .Y(n_779) );
INVx1_ASAP7_75t_L g1238 ( .A(n_267), .Y(n_1238) );
INVx1_ASAP7_75t_L g972 ( .A(n_268), .Y(n_972) );
INVx1_ASAP7_75t_L g882 ( .A(n_269), .Y(n_882) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_270), .Y(n_527) );
INVx1_ASAP7_75t_L g1144 ( .A(n_271), .Y(n_1144) );
CKINVDCx5p33_ASAP7_75t_R g1198 ( .A(n_272), .Y(n_1198) );
OAI211xp5_ASAP7_75t_SL g1070 ( .A1(n_273), .A2(n_432), .B(n_1071), .C(n_1072), .Y(n_1070) );
OAI211xp5_ASAP7_75t_SL g1079 ( .A1(n_273), .A2(n_622), .B(n_1080), .C(n_1081), .Y(n_1079) );
INVx1_ASAP7_75t_L g1111 ( .A(n_274), .Y(n_1111) );
XOR2x2_ASAP7_75t_L g1089 ( .A(n_276), .B(n_1090), .Y(n_1089) );
OAI211xp5_ASAP7_75t_L g760 ( .A1(n_277), .A2(n_650), .B(n_761), .C(n_762), .Y(n_760) );
INVx1_ASAP7_75t_L g774 ( .A(n_277), .Y(n_774) );
INVxp67_ASAP7_75t_SL g1625 ( .A(n_280), .Y(n_1625) );
AOI22xp33_ASAP7_75t_SL g1010 ( .A1(n_281), .A2(n_309), .B1(n_1011), .B2(n_1016), .Y(n_1010) );
INVx1_ASAP7_75t_L g845 ( .A(n_282), .Y(n_845) );
OAI211xp5_ASAP7_75t_L g852 ( .A1(n_282), .A2(n_476), .B(n_714), .C(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g1617 ( .A(n_283), .Y(n_1617) );
CKINVDCx5p33_ASAP7_75t_R g781 ( .A(n_284), .Y(n_781) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_285), .Y(n_328) );
INVx1_ASAP7_75t_L g740 ( .A(n_287), .Y(n_740) );
INVx1_ASAP7_75t_L g1137 ( .A(n_288), .Y(n_1137) );
INVx1_ASAP7_75t_L g828 ( .A(n_289), .Y(n_828) );
CKINVDCx5p33_ASAP7_75t_R g784 ( .A(n_290), .Y(n_784) );
INVxp67_ASAP7_75t_SL g1546 ( .A(n_293), .Y(n_1546) );
OAI221xp5_ASAP7_75t_L g1577 ( .A1(n_293), .A2(n_294), .B1(n_1578), .B2(n_1580), .C(n_1582), .Y(n_1577) );
OAI221xp5_ASAP7_75t_L g1514 ( .A1(n_294), .A2(n_300), .B1(n_1515), .B2(n_1521), .C(n_1523), .Y(n_1514) );
CKINVDCx5p33_ASAP7_75t_R g441 ( .A(n_295), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g1051 ( .A(n_299), .Y(n_1051) );
INVx1_ASAP7_75t_L g1161 ( .A(n_302), .Y(n_1161) );
XOR2x2_ASAP7_75t_L g757 ( .A(n_303), .B(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g347 ( .A(n_304), .Y(n_347) );
INVx2_ASAP7_75t_L g395 ( .A(n_304), .Y(n_395) );
INVx1_ASAP7_75t_L g589 ( .A(n_304), .Y(n_589) );
INVx1_ASAP7_75t_L g742 ( .A(n_306), .Y(n_742) );
AOI21xp33_ASAP7_75t_L g1199 ( .A1(n_307), .A2(n_1200), .B(n_1202), .Y(n_1199) );
INVx1_ASAP7_75t_L g1220 ( .A(n_307), .Y(n_1220) );
INVx1_ASAP7_75t_L g680 ( .A(n_308), .Y(n_680) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_310), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g1184 ( .A(n_311), .Y(n_1184) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_333), .B(n_1289), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_319), .Y(n_313) );
INVx1_ASAP7_75t_L g1601 ( .A(n_314), .Y(n_1601) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g1605 ( .A(n_315), .B(n_318), .Y(n_1605) );
INVx1_ASAP7_75t_L g1655 ( .A(n_315), .Y(n_1655) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g1657 ( .A(n_318), .B(n_1655), .Y(n_1657) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_323), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g463 ( .A(n_321), .B(n_464), .Y(n_463) );
AOI21xp5_ASAP7_75t_SL g1176 ( .A1(n_321), .A2(n_1177), .B(n_1189), .Y(n_1176) );
NOR2xp33_ASAP7_75t_L g1600 ( .A(n_321), .B(n_1601), .Y(n_1600) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x4_ASAP7_75t_L g428 ( .A(n_322), .B(n_332), .Y(n_428) );
AND2x4_ASAP7_75t_L g1203 ( .A(n_322), .B(n_331), .Y(n_1203) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_323), .A2(n_459), .B1(n_882), .B2(n_883), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g1282 ( .A1(n_323), .A2(n_459), .B1(n_1238), .B2(n_1239), .Y(n_1282) );
AND2x4_ASAP7_75t_SL g1599 ( .A(n_323), .B(n_1600), .Y(n_1599) );
INVx3_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OR2x6_ASAP7_75t_L g324 ( .A(n_325), .B(n_330), .Y(n_324) );
OR2x6_ASAP7_75t_L g455 ( .A(n_325), .B(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g532 ( .A(n_325), .B(n_456), .Y(n_532) );
BUFx4f_ASAP7_75t_L g728 ( .A(n_325), .Y(n_728) );
INVx1_ASAP7_75t_L g983 ( .A(n_325), .Y(n_983) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx4f_ASAP7_75t_L g405 ( .A(n_326), .Y(n_405) );
INVx3_ASAP7_75t_L g450 ( .A(n_326), .Y(n_450) );
INVx3_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx2_ASAP7_75t_L g411 ( .A(n_328), .Y(n_411) );
INVx2_ASAP7_75t_L g416 ( .A(n_328), .Y(n_416) );
NAND2x1_ASAP7_75t_L g420 ( .A(n_328), .B(n_329), .Y(n_420) );
AND2x2_ASAP7_75t_L g437 ( .A(n_328), .B(n_329), .Y(n_437) );
INVx1_ASAP7_75t_L g446 ( .A(n_328), .Y(n_446) );
AND2x2_ASAP7_75t_L g460 ( .A(n_328), .B(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_329), .B(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g415 ( .A(n_329), .B(n_416), .Y(n_415) );
BUFx2_ASAP7_75t_L g440 ( .A(n_329), .Y(n_440) );
INVx2_ASAP7_75t_L g461 ( .A(n_329), .Y(n_461) );
INVx1_ASAP7_75t_L g896 ( .A(n_329), .Y(n_896) );
AND2x2_ASAP7_75t_L g909 ( .A(n_329), .B(n_411), .Y(n_909) );
OR2x6_ASAP7_75t_L g449 ( .A(n_330), .B(n_450), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g1183 ( .A1(n_330), .A2(n_1184), .B1(n_1185), .B2(n_1186), .Y(n_1183) );
INVxp67_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g434 ( .A(n_331), .Y(n_434) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x4_ASAP7_75t_L g444 ( .A(n_332), .B(n_445), .Y(n_444) );
BUFx2_ASAP7_75t_L g453 ( .A(n_332), .Y(n_453) );
XNOR2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_933), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_336), .B1(n_539), .B2(n_932), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
XNOR2x1_ASAP7_75t_L g337 ( .A(n_338), .B(n_496), .Y(n_337) );
XNOR2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
AND3x1_ASAP7_75t_L g340 ( .A(n_341), .B(n_429), .C(n_466), .Y(n_340) );
NOR2xp33_ASAP7_75t_SL g341 ( .A(n_342), .B(n_399), .Y(n_341) );
OAI33xp33_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_351), .A3(n_366), .B1(n_378), .B2(n_387), .B3(n_393), .Y(n_342) );
OAI33xp33_ASAP7_75t_L g515 ( .A1(n_343), .A2(n_393), .A3(n_516), .B1(n_518), .B2(n_519), .B3(n_523), .Y(n_515) );
BUFx3_ASAP7_75t_L g859 ( .A(n_343), .Y(n_859) );
OAI33xp33_ASAP7_75t_L g959 ( .A1(n_343), .A2(n_393), .A3(n_960), .B1(n_963), .B2(n_967), .B3(n_971), .Y(n_959) );
OAI33xp33_ASAP7_75t_L g1046 ( .A1(n_343), .A2(n_393), .A3(n_1047), .B1(n_1050), .B2(n_1053), .B3(n_1057), .Y(n_1046) );
OAI33xp33_ASAP7_75t_L g1121 ( .A1(n_343), .A2(n_393), .A3(n_1122), .B1(n_1123), .B2(n_1124), .B3(n_1125), .Y(n_1121) );
BUFx4f_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx4f_ASAP7_75t_L g573 ( .A(n_344), .Y(n_573) );
BUFx2_ASAP7_75t_L g662 ( .A(n_344), .Y(n_662) );
BUFx8_ASAP7_75t_L g795 ( .A(n_344), .Y(n_795) );
OR2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_348), .Y(n_344) );
AND2x2_ASAP7_75t_SL g427 ( .A(n_345), .B(n_428), .Y(n_427) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_345), .Y(n_495) );
INVx1_ASAP7_75t_L g567 ( .A(n_345), .Y(n_567) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx2_ASAP7_75t_L g465 ( .A(n_346), .Y(n_465) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx2_ASAP7_75t_L g1560 ( .A(n_348), .Y(n_1560) );
NAND2xp33_ASAP7_75t_SL g348 ( .A(n_349), .B(n_350), .Y(n_348) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_349), .Y(n_493) );
AND3x4_ASAP7_75t_L g1008 ( .A(n_349), .B(n_483), .C(n_1009), .Y(n_1008) );
INVx1_ASAP7_75t_L g1576 ( .A(n_349), .Y(n_1576) );
INVx3_ASAP7_75t_L g398 ( .A(n_350), .Y(n_398) );
BUFx3_ASAP7_75t_L g483 ( .A(n_350), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_353), .B1(n_358), .B2(n_359), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_352), .A2(n_390), .B1(n_404), .B2(n_406), .Y(n_403) );
OAI22xp33_ASAP7_75t_L g960 ( .A1(n_353), .A2(n_517), .B1(n_961), .B2(n_962), .Y(n_960) );
OAI22xp33_ASAP7_75t_L g971 ( .A1(n_353), .A2(n_391), .B1(n_972), .B2(n_973), .Y(n_971) );
OAI22xp5_ASAP7_75t_L g1047 ( .A1(n_353), .A2(n_359), .B1(n_1048), .B2(n_1049), .Y(n_1047) );
OAI22xp5_ASAP7_75t_L g1057 ( .A1(n_353), .A2(n_391), .B1(n_1058), .B2(n_1059), .Y(n_1057) );
OAI22xp33_ASAP7_75t_L g1125 ( .A1(n_353), .A2(n_1111), .B1(n_1117), .B2(n_1126), .Y(n_1125) );
OAI22xp33_ASAP7_75t_L g1147 ( .A1(n_353), .A2(n_359), .B1(n_1136), .B2(n_1144), .Y(n_1147) );
OAI22xp33_ASAP7_75t_L g1153 ( .A1(n_353), .A2(n_391), .B1(n_1137), .B2(n_1145), .Y(n_1153) );
BUFx4f_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g389 ( .A(n_354), .Y(n_389) );
OR2x4_ASAP7_75t_L g468 ( .A(n_354), .B(n_398), .Y(n_468) );
OR2x4_ASAP7_75t_L g489 ( .A(n_354), .B(n_471), .Y(n_489) );
BUFx3_ASAP7_75t_L g577 ( .A(n_354), .Y(n_577) );
BUFx3_ASAP7_75t_L g665 ( .A(n_354), .Y(n_665) );
OR2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_355), .Y(n_365) );
INVx2_ASAP7_75t_L g372 ( .A(n_355), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_355), .B(n_364), .Y(n_377) );
AND2x4_ASAP7_75t_L g478 ( .A(n_355), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g1015 ( .A(n_356), .Y(n_1015) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVxp67_ASAP7_75t_L g371 ( .A(n_357), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_358), .A2(n_392), .B1(n_422), .B2(n_423), .Y(n_421) );
INVx3_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g667 ( .A(n_360), .Y(n_667) );
INVx2_ASAP7_75t_L g799 ( .A(n_360), .Y(n_799) );
INVx3_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx6f_ASAP7_75t_L g517 ( .A(n_361), .Y(n_517) );
INVx4_ASAP7_75t_L g621 ( .A(n_361), .Y(n_621) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx3_ASAP7_75t_L g391 ( .A(n_362), .Y(n_391) );
BUFx2_ASAP7_75t_L g475 ( .A(n_362), .Y(n_475) );
NAND2x1p5_ASAP7_75t_L g362 ( .A(n_363), .B(n_365), .Y(n_362) );
BUFx2_ASAP7_75t_L g486 ( .A(n_363), .Y(n_486) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g479 ( .A(n_364), .Y(n_479) );
BUFx2_ASAP7_75t_L g484 ( .A(n_365), .Y(n_484) );
AND2x4_ASAP7_75t_L g1006 ( .A(n_365), .B(n_1007), .Y(n_1006) );
INVx2_ASAP7_75t_L g1084 ( .A(n_365), .Y(n_1084) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .B1(n_373), .B2(n_374), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_367), .A2(n_379), .B1(n_413), .B2(n_417), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_368), .A2(n_374), .B1(n_506), .B2(n_513), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g1050 ( .A1(n_368), .A2(n_374), .B1(n_1051), .B2(n_1052), .Y(n_1050) );
OAI22xp5_ASAP7_75t_L g1124 ( .A1(n_368), .A2(n_1056), .B1(n_1114), .B2(n_1120), .Y(n_1124) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g470 ( .A(n_369), .B(n_471), .Y(n_470) );
AND2x4_ASAP7_75t_L g618 ( .A(n_369), .B(n_471), .Y(n_618) );
BUFx6f_ASAP7_75t_L g802 ( .A(n_369), .Y(n_802) );
INVx2_ASAP7_75t_L g804 ( .A(n_369), .Y(n_804) );
BUFx6f_ASAP7_75t_L g1222 ( .A(n_369), .Y(n_1222) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g382 ( .A(n_370), .Y(n_382) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_370), .Y(n_521) );
BUFx8_ASAP7_75t_L g871 ( .A(n_370), .Y(n_871) );
AND2x4_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
AND2x4_ASAP7_75t_L g1014 ( .A(n_372), .B(n_1015), .Y(n_1014) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_373), .A2(n_383), .B1(n_404), .B2(n_425), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g1123 ( .A1(n_374), .A2(n_675), .B1(n_1113), .B2(n_1119), .Y(n_1123) );
INVx3_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx3_ASAP7_75t_L g522 ( .A(n_375), .Y(n_522) );
CKINVDCx8_ASAP7_75t_R g582 ( .A(n_375), .Y(n_582) );
INVx3_ASAP7_75t_L g1056 ( .A(n_375), .Y(n_1056) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g874 ( .A(n_376), .Y(n_874) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx2_ASAP7_75t_L g386 ( .A(n_377), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .B1(n_383), .B2(n_384), .Y(n_378) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx3_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx2_ASAP7_75t_L g1229 ( .A(n_382), .Y(n_1229) );
BUFx2_ASAP7_75t_L g1255 ( .A(n_382), .Y(n_1255) );
INVx1_ASAP7_75t_L g1261 ( .A(n_382), .Y(n_1261) );
OR2x6_ASAP7_75t_SL g1585 ( .A(n_382), .B(n_1586), .Y(n_1585) );
OAI22xp5_ASAP7_75t_L g963 ( .A1(n_384), .A2(n_964), .B1(n_965), .B2(n_966), .Y(n_963) );
OAI22xp33_ASAP7_75t_SL g1148 ( .A1(n_384), .A2(n_581), .B1(n_1133), .B2(n_1141), .Y(n_1148) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx2_ASAP7_75t_L g754 ( .A(n_385), .Y(n_754) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
OR2x6_ASAP7_75t_L g490 ( .A(n_386), .B(n_398), .Y(n_490) );
BUFx3_ASAP7_75t_L g584 ( .A(n_386), .Y(n_584) );
OAI22xp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_390), .B1(n_391), .B2(n_392), .Y(n_387) );
OAI22xp33_ASAP7_75t_L g516 ( .A1(n_388), .A2(n_502), .B1(n_509), .B2(n_517), .Y(n_516) );
OAI22xp33_ASAP7_75t_L g523 ( .A1(n_388), .A2(n_391), .B1(n_504), .B2(n_511), .Y(n_523) );
INVx2_ASAP7_75t_SL g863 ( .A(n_388), .Y(n_863) );
OAI22xp33_ASAP7_75t_L g876 ( .A1(n_388), .A2(n_877), .B1(n_878), .B2(n_879), .Y(n_876) );
OAI22xp33_ASAP7_75t_L g1122 ( .A1(n_388), .A2(n_391), .B1(n_1110), .B2(n_1116), .Y(n_1122) );
INVx2_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
INVx3_ASAP7_75t_L g751 ( .A(n_389), .Y(n_751) );
INVx2_ASAP7_75t_L g579 ( .A(n_391), .Y(n_579) );
BUFx6f_ASAP7_75t_L g878 ( .A(n_391), .Y(n_878) );
OR2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_396), .Y(n_393) );
AND2x4_ASAP7_75t_L g401 ( .A(n_394), .B(n_402), .Y(n_401) );
OR2x6_ASAP7_75t_L g1152 ( .A(n_394), .B(n_396), .Y(n_1152) );
INVx1_ASAP7_75t_L g1207 ( .A(n_394), .Y(n_1207) );
BUFx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g1009 ( .A(n_395), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1517 ( .A(n_395), .B(n_1518), .Y(n_1517) );
NAND2x1p5_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
NAND3x1_ASAP7_75t_L g587 ( .A(n_397), .B(n_398), .C(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g471 ( .A(n_398), .Y(n_471) );
AND2x4_ASAP7_75t_L g477 ( .A(n_398), .B(n_478), .Y(n_477) );
AND2x4_ASAP7_75t_L g1575 ( .A(n_398), .B(n_1576), .Y(n_1575) );
OAI33xp33_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_403), .A3(n_412), .B1(n_421), .B2(n_424), .B3(n_426), .Y(n_399) );
OAI22xp5_ASAP7_75t_SL g902 ( .A1(n_400), .A2(n_691), .B1(n_903), .B2(n_910), .Y(n_902) );
OAI33xp33_ASAP7_75t_L g974 ( .A1(n_400), .A2(n_975), .A3(n_977), .B1(n_979), .B2(n_980), .B3(n_981), .Y(n_974) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g500 ( .A(n_401), .Y(n_500) );
INVx2_ASAP7_75t_L g546 ( .A(n_401), .Y(n_546) );
INVx1_ASAP7_75t_L g782 ( .A(n_401), .Y(n_782) );
INVx4_ASAP7_75t_L g998 ( .A(n_401), .Y(n_998) );
OAI221xp5_ASAP7_75t_L g1528 ( .A1(n_401), .A2(n_739), .B1(n_1071), .B2(n_1529), .C(n_1530), .Y(n_1528) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_404), .A2(n_502), .B1(n_503), .B2(n_504), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_404), .A2(n_406), .B1(n_513), .B2(n_514), .Y(n_512) );
OAI22xp33_ASAP7_75t_L g975 ( .A1(n_404), .A2(n_961), .B1(n_972), .B2(n_976), .Y(n_975) );
OAI22xp5_ASAP7_75t_L g1109 ( .A1(n_404), .A2(n_406), .B1(n_1110), .B2(n_1111), .Y(n_1109) );
OAI22xp5_ASAP7_75t_L g1118 ( .A1(n_404), .A2(n_503), .B1(n_1119), .B2(n_1120), .Y(n_1118) );
OAI22xp33_ASAP7_75t_L g1135 ( .A1(n_404), .A2(n_1136), .B1(n_1137), .B2(n_1138), .Y(n_1135) );
INVx4_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx3_ASAP7_75t_L g549 ( .A(n_405), .Y(n_549) );
BUFx6f_ASAP7_75t_L g745 ( .A(n_405), .Y(n_745) );
OAI22xp5_ASAP7_75t_L g1061 ( .A1(n_406), .A2(n_1048), .B1(n_1058), .B2(n_1062), .Y(n_1061) );
OAI22xp5_ASAP7_75t_L g1140 ( .A1(n_406), .A2(n_1062), .B1(n_1141), .B2(n_1142), .Y(n_1140) );
INVx1_ASAP7_75t_L g1509 ( .A(n_406), .Y(n_1509) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx4_ASAP7_75t_L g425 ( .A(n_408), .Y(n_425) );
INVx2_ASAP7_75t_SL g503 ( .A(n_408), .Y(n_503) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_408), .Y(n_552) );
INVx1_ASAP7_75t_L g976 ( .A(n_408), .Y(n_976) );
INVx1_ASAP7_75t_L g1138 ( .A(n_408), .Y(n_1138) );
INVx8_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g452 ( .A(n_409), .B(n_453), .Y(n_452) );
OR2x2_ASAP7_75t_L g947 ( .A(n_409), .B(n_434), .Y(n_947) );
BUFx2_ASAP7_75t_L g1527 ( .A(n_409), .Y(n_1527) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g505 ( .A1(n_413), .A2(n_423), .B1(n_506), .B2(n_507), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_413), .A2(n_509), .B1(n_510), .B2(n_511), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g1112 ( .A1(n_413), .A2(n_510), .B1(n_1113), .B2(n_1114), .Y(n_1112) );
OAI22xp5_ASAP7_75t_L g1115 ( .A1(n_413), .A2(n_1064), .B1(n_1116), .B2(n_1117), .Y(n_1115) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g555 ( .A(n_414), .Y(n_555) );
BUFx2_ASAP7_75t_L g688 ( .A(n_414), .Y(n_688) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx2_ASAP7_75t_L g422 ( .A(n_415), .Y(n_422) );
BUFx2_ASAP7_75t_L g560 ( .A(n_415), .Y(n_560) );
BUFx3_ASAP7_75t_L g739 ( .A(n_415), .Y(n_739) );
INVx1_ASAP7_75t_L g786 ( .A(n_415), .Y(n_786) );
AND2x2_ASAP7_75t_L g895 ( .A(n_416), .B(n_896), .Y(n_895) );
OAI22xp5_ASAP7_75t_L g977 ( .A1(n_417), .A2(n_964), .B1(n_969), .B2(n_978), .Y(n_977) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g431 ( .A(n_418), .Y(n_431) );
INVx2_ASAP7_75t_L g689 ( .A(n_418), .Y(n_689) );
INVx2_ASAP7_75t_L g1066 ( .A(n_418), .Y(n_1066) );
INVx1_ASAP7_75t_L g1194 ( .A(n_418), .Y(n_1194) );
INVx4_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_419), .Y(n_510) );
BUFx4f_ASAP7_75t_L g597 ( .A(n_419), .Y(n_597) );
BUFx4f_ASAP7_75t_L g741 ( .A(n_419), .Y(n_741) );
BUFx4f_ASAP7_75t_L g1064 ( .A(n_419), .Y(n_1064) );
BUFx4f_ASAP7_75t_L g1071 ( .A(n_419), .Y(n_1071) );
OR2x6_ASAP7_75t_L g1523 ( .A(n_419), .B(n_1524), .Y(n_1523) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx3_ASAP7_75t_L g423 ( .A(n_420), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_423), .A2(n_554), .B1(n_555), .B2(n_556), .Y(n_553) );
BUFx2_ASAP7_75t_SL g562 ( .A(n_423), .Y(n_562) );
BUFx3_ASAP7_75t_L g650 ( .A(n_423), .Y(n_650) );
INVx2_ASAP7_75t_SL g736 ( .A(n_423), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g979 ( .A1(n_423), .A2(n_962), .B1(n_973), .B2(n_978), .Y(n_979) );
OR2x2_ASAP7_75t_L g1545 ( .A(n_423), .B(n_1540), .Y(n_1545) );
OAI22xp5_ASAP7_75t_L g981 ( .A1(n_425), .A2(n_966), .B1(n_970), .B2(n_982), .Y(n_981) );
OAI22xp5_ASAP7_75t_L g1067 ( .A1(n_425), .A2(n_1052), .B1(n_1055), .B2(n_1062), .Y(n_1067) );
OAI33xp33_ASAP7_75t_L g499 ( .A1(n_426), .A2(n_500), .A3(n_501), .B1(n_505), .B2(n_508), .B3(n_512), .Y(n_499) );
OAI33xp33_ASAP7_75t_L g1108 ( .A1(n_426), .A2(n_500), .A3(n_1109), .B1(n_1112), .B2(n_1115), .B3(n_1118), .Y(n_1108) );
OAI33xp33_ASAP7_75t_L g1131 ( .A1(n_426), .A2(n_1132), .A3(n_1135), .B1(n_1139), .B2(n_1140), .B3(n_1143), .Y(n_1131) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g980 ( .A(n_427), .Y(n_980) );
NAND3xp33_ASAP7_75t_L g999 ( .A(n_427), .B(n_1000), .C(n_1001), .Y(n_999) );
AOI33xp33_ASAP7_75t_L g1645 ( .A1(n_427), .A2(n_1646), .A3(n_1647), .B1(n_1649), .B2(n_1651), .B3(n_1652), .Y(n_1645) );
AND2x4_ASAP7_75t_L g565 ( .A(n_428), .B(n_566), .Y(n_565) );
OAI221xp5_ASAP7_75t_L g1193 ( .A1(n_428), .A2(n_687), .B1(n_1194), .B2(n_1195), .C(n_1196), .Y(n_1193) );
OAI31xp33_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_448), .A3(n_454), .B(n_462), .Y(n_429) );
OAI22xp5_ASAP7_75t_L g690 ( .A1(n_431), .A2(n_666), .B1(n_681), .B2(n_687), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g783 ( .A1(n_431), .A2(n_784), .B1(n_785), .B2(n_787), .Y(n_783) );
OAI22xp33_ASAP7_75t_L g838 ( .A1(n_431), .A2(n_733), .B1(n_823), .B2(n_828), .Y(n_838) );
NAND3xp33_ASAP7_75t_L g1024 ( .A(n_432), .B(n_1025), .C(n_1028), .Y(n_1024) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g1636 ( .A(n_433), .Y(n_1636) );
AND2x2_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
AND2x2_ASAP7_75t_L g439 ( .A(n_434), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g606 ( .A(n_434), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g1635 ( .A(n_435), .Y(n_1635) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx2_ASAP7_75t_L g1275 ( .A(n_436), .Y(n_1275) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx6f_ASAP7_75t_L g607 ( .A(n_437), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_441), .B1(n_442), .B2(n_447), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_439), .A2(n_527), .B1(n_528), .B2(n_529), .Y(n_526) );
INVx1_ASAP7_75t_L g1182 ( .A(n_439), .Y(n_1182) );
AOI22xp33_ASAP7_75t_L g1629 ( .A1(n_439), .A2(n_444), .B1(n_1630), .B2(n_1631), .Y(n_1629) );
AND2x4_ASAP7_75t_L g600 ( .A(n_440), .B(n_453), .Y(n_600) );
AND2x2_ASAP7_75t_L g653 ( .A(n_440), .B(n_453), .Y(n_653) );
INVx1_ASAP7_75t_L g1520 ( .A(n_440), .Y(n_1520) );
AOI22xp33_ASAP7_75t_SL g480 ( .A1(n_441), .A2(n_481), .B1(n_485), .B2(n_487), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_442), .A2(n_600), .B1(n_844), .B2(n_845), .Y(n_843) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
BUFx3_ASAP7_75t_L g528 ( .A(n_444), .Y(n_528) );
INVx2_ASAP7_75t_L g603 ( .A(n_444), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_444), .A2(n_600), .B1(n_703), .B2(n_704), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g1522 ( .A(n_445), .B(n_1518), .Y(n_1522) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g1624 ( .A(n_449), .Y(n_1624) );
BUFx3_ASAP7_75t_L g569 ( .A(n_450), .Y(n_569) );
BUFx3_ASAP7_75t_L g1062 ( .A(n_450), .Y(n_1062) );
BUFx6f_ASAP7_75t_L g1511 ( .A(n_450), .Y(n_1511) );
INVx2_ASAP7_75t_SL g658 ( .A(n_451), .Y(n_658) );
BUFx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g611 ( .A(n_452), .Y(n_611) );
INVx1_ASAP7_75t_L g900 ( .A(n_452), .Y(n_900) );
AND2x2_ASAP7_75t_L g893 ( .A(n_453), .B(n_894), .Y(n_893) );
O2A1O1Ixp33_ASAP7_75t_L g1179 ( .A1(n_453), .A2(n_992), .B(n_1180), .C(n_1181), .Y(n_1179) );
INVx1_ASAP7_75t_L g1185 ( .A(n_453), .Y(n_1185) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_455), .Y(n_609) );
BUFx2_ASAP7_75t_L g656 ( .A(n_455), .Y(n_656) );
AND2x4_ASAP7_75t_L g459 ( .A(n_456), .B(n_460), .Y(n_459) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
CKINVDCx16_ASAP7_75t_R g458 ( .A(n_459), .Y(n_458) );
INVx4_ASAP7_75t_L g593 ( .A(n_459), .Y(n_593) );
INVx3_ASAP7_75t_SL g1178 ( .A(n_459), .Y(n_1178) );
AOI22xp5_ASAP7_75t_L g1622 ( .A1(n_459), .A2(n_1623), .B1(n_1624), .B2(n_1625), .Y(n_1622) );
BUFx3_ASAP7_75t_L g991 ( .A(n_460), .Y(n_991) );
BUFx6f_ASAP7_75t_L g1201 ( .A(n_460), .Y(n_1201) );
INVx2_ASAP7_75t_L g1273 ( .A(n_460), .Y(n_1273) );
OAI31xp33_ASAP7_75t_L g524 ( .A1(n_462), .A2(n_525), .A3(n_530), .B(n_531), .Y(n_524) );
OAI31xp33_ASAP7_75t_L g1154 ( .A1(n_462), .A2(n_1155), .A3(n_1156), .B(n_1162), .Y(n_1154) );
BUFx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx3_ASAP7_75t_L g612 ( .A(n_463), .Y(n_612) );
BUFx2_ASAP7_75t_SL g707 ( .A(n_463), .Y(n_707) );
INVx1_ASAP7_75t_L g901 ( .A(n_463), .Y(n_901) );
OAI31xp33_ASAP7_75t_L g1068 ( .A1(n_463), .A2(n_1069), .A3(n_1070), .B(n_1075), .Y(n_1068) );
OAI31xp33_ASAP7_75t_L g1091 ( .A1(n_463), .A2(n_1092), .A3(n_1093), .B(n_1097), .Y(n_1091) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
OR2x2_ASAP7_75t_L g1521 ( .A(n_465), .B(n_1522), .Y(n_1521) );
INVx1_ASAP7_75t_L g1552 ( .A(n_465), .Y(n_1552) );
OAI31xp33_ASAP7_75t_SL g466 ( .A1(n_467), .A2(n_472), .A3(n_488), .B(n_491), .Y(n_466) );
INVx2_ASAP7_75t_SL g616 ( .A(n_468), .Y(n_616) );
INVx1_ASAP7_75t_L g720 ( .A(n_468), .Y(n_720) );
INVx1_ASAP7_75t_L g851 ( .A(n_468), .Y(n_851) );
INVx2_ASAP7_75t_SL g923 ( .A(n_468), .Y(n_923) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AOI22xp33_ASAP7_75t_SL g1216 ( .A1(n_470), .A2(n_720), .B1(n_1184), .B2(n_1217), .Y(n_1216) );
OAI22xp33_ASAP7_75t_L g590 ( .A1(n_473), .A2(n_550), .B1(n_563), .B2(n_575), .Y(n_590) );
OAI22xp33_ASAP7_75t_L g679 ( .A1(n_473), .A2(n_665), .B1(n_680), .B2(n_681), .Y(n_679) );
OAI22xp33_ASAP7_75t_L g749 ( .A1(n_473), .A2(n_727), .B1(n_740), .B2(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g821 ( .A(n_475), .Y(n_821) );
OR2x6_ASAP7_75t_L g1582 ( .A(n_475), .B(n_1583), .Y(n_1582) );
NAND3xp33_ASAP7_75t_L g952 ( .A(n_476), .B(n_953), .C(n_955), .Y(n_952) );
NAND3xp33_ASAP7_75t_SL g1100 ( .A(n_476), .B(n_1101), .C(n_1103), .Y(n_1100) );
NAND3xp33_ASAP7_75t_SL g1640 ( .A(n_476), .B(n_1641), .C(n_1642), .Y(n_1640) );
CKINVDCx8_ASAP7_75t_R g476 ( .A(n_477), .Y(n_476) );
CKINVDCx8_ASAP7_75t_R g622 ( .A(n_477), .Y(n_622) );
AOI211xp5_ASAP7_75t_L g916 ( .A1(n_477), .A2(n_917), .B(n_918), .C(n_919), .Y(n_916) );
NOR3xp33_ASAP7_75t_L g1210 ( .A(n_477), .B(n_1211), .C(n_1215), .Y(n_1210) );
NOR3xp33_ASAP7_75t_L g1240 ( .A(n_477), .B(n_1241), .C(n_1244), .Y(n_1240) );
BUFx3_ASAP7_75t_L g918 ( .A(n_478), .Y(n_918) );
INVx2_ASAP7_75t_L g1017 ( .A(n_478), .Y(n_1017) );
BUFx2_ASAP7_75t_L g1038 ( .A(n_478), .Y(n_1038) );
BUFx2_ASAP7_75t_L g1102 ( .A(n_478), .Y(n_1102) );
BUFx2_ASAP7_75t_L g1225 ( .A(n_478), .Y(n_1225) );
AND2x2_ASAP7_75t_L g1569 ( .A(n_478), .B(n_1566), .Y(n_1569) );
INVx1_ASAP7_75t_L g1007 ( .A(n_479), .Y(n_1007) );
AOI22xp33_ASAP7_75t_SL g536 ( .A1(n_481), .A2(n_485), .B1(n_527), .B2(n_537), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g1081 ( .A1(n_481), .A2(n_1073), .B1(n_1082), .B2(n_1085), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_481), .A2(n_485), .B1(n_1095), .B2(n_1104), .Y(n_1103) );
INVx1_ASAP7_75t_L g1213 ( .A(n_481), .Y(n_1213) );
AOI22xp33_ASAP7_75t_L g1642 ( .A1(n_481), .A2(n_485), .B1(n_1630), .B2(n_1633), .Y(n_1642) );
AND2x4_ASAP7_75t_L g481 ( .A(n_482), .B(n_484), .Y(n_481) );
AND2x2_ASAP7_75t_L g485 ( .A(n_482), .B(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g625 ( .A(n_482), .B(n_484), .Y(n_625) );
AND2x4_ASAP7_75t_L g627 ( .A(n_482), .B(n_486), .Y(n_627) );
AND2x4_ASAP7_75t_L g716 ( .A(n_482), .B(n_484), .Y(n_716) );
INVx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_483), .B(n_1086), .Y(n_1085) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_485), .A2(n_716), .B1(n_944), .B2(n_954), .Y(n_953) );
INVxp67_ASAP7_75t_L g1080 ( .A(n_485), .Y(n_1080) );
INVxp67_ASAP7_75t_L g1214 ( .A(n_485), .Y(n_1214) );
BUFx3_ASAP7_75t_L g630 ( .A(n_489), .Y(n_630) );
INVx2_ASAP7_75t_SL g925 ( .A(n_489), .Y(n_925) );
BUFx2_ASAP7_75t_L g1242 ( .A(n_489), .Y(n_1242) );
INVx1_ASAP7_75t_L g632 ( .A(n_490), .Y(n_632) );
INVx1_ASAP7_75t_L g711 ( .A(n_490), .Y(n_711) );
INVx2_ASAP7_75t_L g926 ( .A(n_490), .Y(n_926) );
OAI31xp33_ASAP7_75t_SL g533 ( .A1(n_491), .A2(n_534), .A3(n_535), .B(n_538), .Y(n_533) );
OAI31xp33_ASAP7_75t_L g949 ( .A1(n_491), .A2(n_950), .A3(n_952), .B(n_957), .Y(n_949) );
OAI21xp5_ASAP7_75t_L g1033 ( .A1(n_491), .A2(n_1034), .B(n_1036), .Y(n_1033) );
OAI31xp33_ASAP7_75t_SL g1076 ( .A1(n_491), .A2(n_1077), .A3(n_1078), .B(n_1079), .Y(n_1076) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_494), .Y(n_491) );
AND2x2_ASAP7_75t_SL g634 ( .A(n_492), .B(n_494), .Y(n_634) );
AND2x2_ASAP7_75t_L g722 ( .A(n_492), .B(n_494), .Y(n_722) );
AND2x4_ASAP7_75t_L g928 ( .A(n_492), .B(n_494), .Y(n_928) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_492), .B(n_494), .Y(n_1106) );
INVx1_ASAP7_75t_SL g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND3x1_ASAP7_75t_L g497 ( .A(n_498), .B(n_524), .C(n_533), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_499), .B(n_515), .Y(n_498) );
BUFx6f_ASAP7_75t_L g725 ( .A(n_500), .Y(n_725) );
OAI33xp33_ASAP7_75t_L g1060 ( .A1(n_500), .A2(n_980), .A3(n_1061), .B1(n_1063), .B2(n_1065), .B3(n_1067), .Y(n_1060) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_507), .A2(n_514), .B1(n_520), .B2(n_522), .Y(n_519) );
HB1xp67_ASAP7_75t_L g942 ( .A(n_510), .Y(n_942) );
OAI22xp5_ASAP7_75t_L g1132 ( .A1(n_510), .A2(n_978), .B1(n_1133), .B2(n_1134), .Y(n_1132) );
INVx1_ASAP7_75t_L g772 ( .A(n_517), .Y(n_772) );
OAI22xp33_ASAP7_75t_L g860 ( .A1(n_517), .A2(n_861), .B1(n_862), .B2(n_864), .Y(n_860) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_520), .A2(n_556), .B1(n_571), .B2(n_584), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_520), .A2(n_732), .B1(n_746), .B2(n_753), .Y(n_752) );
OAI22xp5_ASAP7_75t_L g1053 ( .A1(n_520), .A2(n_1054), .B1(n_1055), .B2(n_1056), .Y(n_1053) );
INVx2_ASAP7_75t_SL g520 ( .A(n_521), .Y(n_520) );
INVx5_ASAP7_75t_L g581 ( .A(n_521), .Y(n_581) );
INVx3_ASAP7_75t_L g675 ( .A(n_521), .Y(n_675) );
INVx2_ASAP7_75t_SL g867 ( .A(n_521), .Y(n_867) );
HB1xp67_ASAP7_75t_L g1004 ( .A(n_521), .Y(n_1004) );
OAI22xp5_ASAP7_75t_L g865 ( .A1(n_522), .A2(n_866), .B1(n_867), .B2(n_868), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_528), .A2(n_600), .B1(n_944), .B2(n_945), .Y(n_943) );
AOI222xp33_ASAP7_75t_L g1028 ( .A1(n_528), .A2(n_600), .B1(n_992), .B2(n_1029), .C1(n_1030), .C2(n_1031), .Y(n_1028) );
AOI22xp5_ASAP7_75t_L g1072 ( .A1(n_528), .A2(n_600), .B1(n_1073), .B2(n_1074), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g1094 ( .A1(n_528), .A2(n_600), .B1(n_1095), .B2(n_1096), .Y(n_1094) );
AOI22xp33_ASAP7_75t_L g1157 ( .A1(n_528), .A2(n_653), .B1(n_1158), .B2(n_1159), .Y(n_1157) );
INVx2_ASAP7_75t_SL g932 ( .A(n_539), .Y(n_932) );
XOR2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_694), .Y(n_539) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_635), .B(n_693), .Y(n_540) );
INVx2_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
OR2x2_ASAP7_75t_L g693 ( .A(n_542), .B(n_636), .Y(n_693) );
NAND3xp33_ASAP7_75t_L g543 ( .A(n_544), .B(n_591), .C(n_613), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_545), .B(n_572), .Y(n_544) );
OAI33xp33_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_547), .A3(n_553), .B1(n_557), .B2(n_564), .B3(n_568), .Y(n_545) );
OAI33xp33_ASAP7_75t_L g682 ( .A1(n_546), .A2(n_683), .A3(n_686), .B1(n_690), .B2(n_691), .B3(n_692), .Y(n_682) );
OAI22xp5_ASAP7_75t_SL g547 ( .A1(n_548), .A2(n_549), .B1(n_550), .B2(n_551), .Y(n_547) );
OAI22xp33_ASAP7_75t_L g574 ( .A1(n_548), .A2(n_561), .B1(n_575), .B2(n_578), .Y(n_574) );
INVx2_ASAP7_75t_SL g685 ( .A(n_549), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_551), .A2(n_569), .B1(n_570), .B2(n_571), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_551), .A2(n_664), .B1(n_680), .B2(n_684), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_551), .A2(n_671), .B1(n_677), .B2(n_684), .Y(n_692) );
OAI22xp33_ASAP7_75t_L g778 ( .A1(n_551), .A2(n_779), .B1(n_780), .B2(n_781), .Y(n_778) );
OAI22xp33_ASAP7_75t_L g791 ( .A1(n_551), .A2(n_780), .B1(n_792), .B2(n_793), .Y(n_791) );
INVx6_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx5_ASAP7_75t_L g730 ( .A(n_552), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_554), .A2(n_570), .B1(n_581), .B2(n_582), .Y(n_580) );
OAI221xp5_ASAP7_75t_L g903 ( .A1(n_555), .A2(n_650), .B1(n_866), .B2(n_872), .C(n_904), .Y(n_903) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_561), .B1(n_562), .B2(n_563), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx4_ASAP7_75t_L g733 ( .A(n_559), .Y(n_733) );
INVx4_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OAI33xp33_ASAP7_75t_L g836 ( .A1(n_564), .A2(n_725), .A3(n_837), .B1(n_838), .B2(n_839), .B3(n_840), .Y(n_836) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
CKINVDCx5p33_ASAP7_75t_R g691 ( .A(n_565), .Y(n_691) );
AOI33xp33_ASAP7_75t_L g1264 ( .A1(n_565), .A2(n_1265), .A3(n_1266), .B1(n_1269), .B2(n_1276), .B3(n_1277), .Y(n_1264) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OAI33xp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_574), .A3(n_580), .B1(n_583), .B2(n_585), .B3(n_590), .Y(n_572) );
OAI33xp33_ASAP7_75t_L g748 ( .A1(n_573), .A2(n_678), .A3(n_749), .B1(n_752), .B2(n_755), .B3(n_756), .Y(n_748) );
OAI33xp33_ASAP7_75t_L g816 ( .A1(n_573), .A2(n_817), .A3(n_822), .B1(n_825), .B2(n_830), .B3(n_833), .Y(n_816) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVxp67_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g798 ( .A(n_577), .Y(n_798) );
INVx1_ASAP7_75t_L g808 ( .A(n_577), .Y(n_808) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
BUFx3_ASAP7_75t_L g670 ( .A(n_581), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_581), .A2(n_582), .B1(n_734), .B2(n_747), .Y(n_755) );
INVx8_ASAP7_75t_L g827 ( .A(n_581), .Y(n_827) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_582), .A2(n_669), .B1(n_670), .B2(n_671), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g825 ( .A1(n_582), .A2(n_826), .B1(n_828), .B2(n_829), .Y(n_825) );
OAI221xp5_ASAP7_75t_L g1228 ( .A1(n_582), .A2(n_1192), .B1(n_1198), .B2(n_1229), .C(n_1230), .Y(n_1228) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_584), .A2(n_673), .B1(n_676), .B2(n_677), .Y(n_672) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
CKINVDCx5p33_ASAP7_75t_R g678 ( .A(n_586), .Y(n_678) );
INVx2_ASAP7_75t_L g805 ( .A(n_586), .Y(n_805) );
INVx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx3_ASAP7_75t_L g832 ( .A(n_587), .Y(n_832) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g1534 ( .A(n_589), .Y(n_1534) );
NAND2xp5_ASAP7_75t_L g1540 ( .A(n_589), .B(n_1541), .Y(n_1540) );
OAI31xp33_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_594), .A3(n_608), .B(n_612), .Y(n_591) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g788 ( .A1(n_597), .A2(n_785), .B1(n_789), .B2(n_790), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_601), .B1(n_602), .B2(n_604), .Y(n_598) );
BUFx3_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g890 ( .A(n_600), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_601), .A2(n_624), .B1(n_626), .B2(n_628), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_602), .A2(n_643), .B1(n_653), .B2(n_654), .Y(n_652) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g764 ( .A(n_603), .Y(n_764) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g651 ( .A(n_606), .Y(n_651) );
INVx3_ASAP7_75t_L g761 ( .A(n_606), .Y(n_761) );
AOI211xp5_ASAP7_75t_L g884 ( .A1(n_606), .A2(n_885), .B(n_888), .C(n_889), .Y(n_884) );
NOR3xp33_ASAP7_75t_L g1283 ( .A(n_606), .B(n_1284), .C(n_1285), .Y(n_1283) );
BUFx6f_ASAP7_75t_L g887 ( .A(n_607), .Y(n_887) );
BUFx3_ASAP7_75t_L g992 ( .A(n_607), .Y(n_992) );
BUFx3_ASAP7_75t_L g1650 ( .A(n_607), .Y(n_1650) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g706 ( .A(n_611), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_611), .A2(n_893), .B1(n_1026), .B2(n_1027), .Y(n_1025) );
INVx1_ASAP7_75t_L g1163 ( .A(n_611), .Y(n_1163) );
OAI31xp33_ASAP7_75t_L g646 ( .A1(n_612), .A2(n_647), .A3(n_655), .B(n_659), .Y(n_646) );
OAI31xp33_ASAP7_75t_SL g841 ( .A1(n_612), .A2(n_842), .A3(n_846), .B(n_847), .Y(n_841) );
OAI31xp33_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_619), .A3(n_629), .B(n_633), .Y(n_613) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g640 ( .A(n_618), .Y(n_640) );
INVx1_ASAP7_75t_L g721 ( .A(n_618), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_618), .A2(n_882), .B1(n_883), .B2(n_923), .Y(n_922) );
INVx1_ASAP7_75t_L g951 ( .A(n_618), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g1237 ( .A1(n_618), .A2(n_923), .B1(n_1238), .B2(n_1239), .Y(n_1237) );
OAI22xp33_ASAP7_75t_L g806 ( .A1(n_620), .A2(n_781), .B1(n_790), .B2(n_807), .Y(n_806) );
OAI22xp33_ASAP7_75t_L g833 ( .A1(n_620), .A2(n_750), .B1(n_834), .B2(n_835), .Y(n_833) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g714 ( .A(n_621), .Y(n_714) );
INVx1_ASAP7_75t_L g1126 ( .A(n_621), .Y(n_1126) );
INVx2_ASAP7_75t_L g1212 ( .A(n_621), .Y(n_1212) );
INVx1_ASAP7_75t_L g1245 ( .A(n_621), .Y(n_1245) );
NAND3xp33_ASAP7_75t_L g1036 ( .A(n_622), .B(n_1037), .C(n_1040), .Y(n_1036) );
NAND3xp33_ASAP7_75t_L g1166 ( .A(n_622), .B(n_1167), .C(n_1168), .Y(n_1166) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_624), .A2(n_626), .B1(n_643), .B2(n_644), .Y(n_642) );
BUFx3_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
BUFx3_ASAP7_75t_L g1039 ( .A(n_625), .Y(n_1039) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_627), .A2(n_703), .B1(n_716), .B2(n_717), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_627), .A2(n_716), .B1(n_763), .B2(n_774), .Y(n_773) );
AOI22xp33_ASAP7_75t_SL g853 ( .A1(n_627), .A2(n_716), .B1(n_844), .B2(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g921 ( .A(n_627), .Y(n_921) );
AOI222xp33_ASAP7_75t_L g1037 ( .A1(n_627), .A2(n_1029), .B1(n_1030), .B2(n_1031), .C1(n_1038), .C2(n_1039), .Y(n_1037) );
AOI22xp33_ASAP7_75t_L g1167 ( .A1(n_627), .A2(n_716), .B1(n_1158), .B2(n_1161), .Y(n_1167) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OAI31xp33_ASAP7_75t_L g638 ( .A1(n_633), .A2(n_639), .A3(n_641), .B(n_645), .Y(n_638) );
BUFx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g1208 ( .A1(n_634), .A2(n_1209), .B(n_1218), .Y(n_1208) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NAND3xp33_ASAP7_75t_L g637 ( .A(n_638), .B(n_646), .C(n_660), .Y(n_637) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OAI221xp5_ASAP7_75t_L g910 ( .A1(n_650), .A2(n_864), .B1(n_879), .B2(n_911), .C(n_913), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_653), .A2(n_763), .B1(n_764), .B2(n_765), .Y(n_762) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_661), .B(n_682), .Y(n_660) );
OAI33xp33_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_663), .A3(n_668), .B1(n_672), .B2(n_678), .B3(n_679), .Y(n_661) );
OAI33xp33_ASAP7_75t_L g1146 ( .A1(n_662), .A2(n_1147), .A3(n_1148), .B1(n_1149), .B2(n_1152), .B3(n_1153), .Y(n_1146) );
OAI22xp5_ASAP7_75t_L g1218 ( .A1(n_662), .A2(n_678), .B1(n_1219), .B2(n_1228), .Y(n_1218) );
OAI22xp33_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_665), .B1(n_666), .B2(n_667), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_669), .A2(n_676), .B1(n_687), .B2(n_689), .Y(n_686) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
OAI22xp33_ASAP7_75t_SL g822 ( .A1(n_675), .A2(n_753), .B1(n_823), .B2(n_824), .Y(n_822) );
INVx1_ASAP7_75t_L g1263 ( .A(n_678), .Y(n_1263) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx4_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
OAI33xp33_ASAP7_75t_L g724 ( .A1(n_691), .A2(n_725), .A3(n_726), .B1(n_731), .B2(n_737), .B3(n_743), .Y(n_724) );
OAI33xp33_ASAP7_75t_L g777 ( .A1(n_691), .A2(n_778), .A3(n_782), .B1(n_783), .B2(n_788), .B3(n_791), .Y(n_777) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_810), .B1(n_811), .B2(n_931), .Y(n_694) );
INVx1_ASAP7_75t_L g931 ( .A(n_695), .Y(n_931) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .B1(n_757), .B2(n_809), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NAND3xp33_ASAP7_75t_L g698 ( .A(n_699), .B(n_708), .C(n_723), .Y(n_698) );
OAI31xp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_701), .A3(n_705), .B(n_707), .Y(n_699) );
OAI31xp33_ASAP7_75t_L g759 ( .A1(n_707), .A2(n_760), .A3(n_766), .B(n_767), .Y(n_759) );
OAI31xp33_ASAP7_75t_SL g940 ( .A1(n_707), .A2(n_941), .A3(n_946), .B(n_948), .Y(n_940) );
OAI21xp5_ASAP7_75t_L g1023 ( .A1(n_707), .A2(n_1024), .B(n_1032), .Y(n_1023) );
OAI31xp33_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_712), .A3(n_718), .B(n_722), .Y(n_708) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
OAI22xp33_ASAP7_75t_L g756 ( .A1(n_714), .A2(n_729), .B1(n_742), .B2(n_750), .Y(n_756) );
INVx1_ASAP7_75t_L g920 ( .A(n_716), .Y(n_920) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
OAI31xp33_ASAP7_75t_L g768 ( .A1(n_722), .A2(n_769), .A3(n_770), .B(n_775), .Y(n_768) );
OAI31xp33_ASAP7_75t_L g848 ( .A1(n_722), .A2(n_849), .A3(n_852), .B(n_855), .Y(n_848) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_724), .B(n_748), .Y(n_723) );
INVx1_ASAP7_75t_L g1265 ( .A(n_725), .Y(n_1265) );
OAI22xp33_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_728), .B1(n_729), .B2(n_730), .Y(n_726) );
OAI22xp33_ASAP7_75t_L g837 ( .A1(n_728), .A2(n_730), .B1(n_818), .B2(n_834), .Y(n_837) );
OAI22xp5_ASAP7_75t_L g1190 ( .A1(n_728), .A2(n_730), .B1(n_1191), .B2(n_1192), .Y(n_1190) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_730), .A2(n_744), .B1(n_746), .B2(n_747), .Y(n_743) );
OAI22xp5_ASAP7_75t_L g840 ( .A1(n_730), .A2(n_744), .B1(n_824), .B2(n_829), .Y(n_840) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_733), .B1(n_734), .B2(n_735), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_733), .A2(n_741), .B1(n_819), .B2(n_835), .Y(n_839) );
INVx5_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
OAI22xp33_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_740), .B1(n_741), .B2(n_742), .Y(n_737) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g912 ( .A(n_739), .Y(n_912) );
OAI22xp5_ASAP7_75t_L g1065 ( .A1(n_739), .A2(n_1049), .B1(n_1059), .B2(n_1066), .Y(n_1065) );
OAI22xp5_ASAP7_75t_L g1143 ( .A1(n_739), .A2(n_1064), .B1(n_1144), .B2(n_1145), .Y(n_1143) );
OAI211xp5_ASAP7_75t_SL g1197 ( .A1(n_741), .A2(n_1198), .B(n_1199), .C(n_1204), .Y(n_1197) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx3_ASAP7_75t_L g780 ( .A(n_745), .Y(n_780) );
OAI22xp33_ASAP7_75t_L g817 ( .A1(n_750), .A2(n_818), .B1(n_819), .B2(n_820), .Y(n_817) );
BUFx4f_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
OAI22xp5_ASAP7_75t_L g800 ( .A1(n_753), .A2(n_784), .B1(n_792), .B2(n_801), .Y(n_800) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_753), .A2(n_787), .B1(n_793), .B2(n_804), .Y(n_803) );
INVx3_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g809 ( .A(n_757), .Y(n_809) );
NAND3xp33_ASAP7_75t_SL g758 ( .A(n_759), .B(n_768), .C(n_776), .Y(n_758) );
NAND3xp33_ASAP7_75t_L g1156 ( .A(n_761), .B(n_1157), .C(n_1160), .Y(n_1156) );
INVx2_ASAP7_75t_SL g771 ( .A(n_772), .Y(n_771) );
NOR2xp33_ASAP7_75t_SL g776 ( .A(n_777), .B(n_794), .Y(n_776) );
OAI22xp33_ASAP7_75t_L g796 ( .A1(n_779), .A2(n_789), .B1(n_797), .B2(n_799), .Y(n_796) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx2_ASAP7_75t_L g978 ( .A(n_786), .Y(n_978) );
OAI33xp33_ASAP7_75t_L g794 ( .A1(n_795), .A2(n_796), .A3(n_800), .B1(n_803), .B2(n_805), .B3(n_806), .Y(n_794) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
AOI22xp5_ASAP7_75t_L g811 ( .A1(n_812), .A2(n_856), .B1(n_929), .B2(n_930), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
HB1xp67_ASAP7_75t_L g929 ( .A(n_813), .Y(n_929) );
NAND3xp33_ASAP7_75t_L g814 ( .A(n_815), .B(n_841), .C(n_848), .Y(n_814) );
NOR2xp33_ASAP7_75t_L g815 ( .A(n_816), .B(n_836), .Y(n_815) );
INVxp67_ASAP7_75t_SL g820 ( .A(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
OAI33xp33_ASAP7_75t_L g858 ( .A1(n_830), .A2(n_859), .A3(n_860), .B1(n_865), .B2(n_869), .B3(n_876), .Y(n_858) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
BUFx2_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
BUFx2_ASAP7_75t_L g1021 ( .A(n_832), .Y(n_1021) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g930 ( .A(n_856), .Y(n_930) );
NOR4xp25_ASAP7_75t_L g857 ( .A(n_858), .B(n_880), .C(n_902), .D(n_915), .Y(n_857) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
OAI22xp5_ASAP7_75t_L g869 ( .A1(n_870), .A2(n_872), .B1(n_873), .B2(n_875), .Y(n_869) );
INVx2_ASAP7_75t_SL g870 ( .A(n_871), .Y(n_870) );
INVx3_ASAP7_75t_L g965 ( .A(n_871), .Y(n_965) );
INVx2_ASAP7_75t_SL g968 ( .A(n_871), .Y(n_968) );
OAI22xp5_ASAP7_75t_L g967 ( .A1(n_873), .A2(n_968), .B1(n_969), .B2(n_970), .Y(n_967) );
BUFx3_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g1151 ( .A(n_874), .Y(n_1151) );
AOI31xp33_ASAP7_75t_SL g880 ( .A1(n_881), .A2(n_884), .A3(n_891), .B(n_901), .Y(n_880) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_892), .A2(n_893), .B1(n_897), .B2(n_898), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_892), .A2(n_897), .B1(n_925), .B2(n_926), .Y(n_924) );
BUFx6f_ASAP7_75t_L g914 ( .A(n_894), .Y(n_914) );
INVx3_ASAP7_75t_L g995 ( .A(n_894), .Y(n_995) );
BUFx6f_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
INVx3_ASAP7_75t_L g906 ( .A(n_895), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g1536 ( .A(n_895), .B(n_1518), .Y(n_1536) );
AND2x2_ASAP7_75t_L g1553 ( .A(n_895), .B(n_1541), .Y(n_1553) );
INVx2_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx2_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
NAND2xp5_ASAP7_75t_SL g1187 ( .A(n_900), .B(n_1188), .Y(n_1187) );
AO21x1_ASAP7_75t_L g1281 ( .A1(n_901), .A2(n_1282), .B(n_1283), .Y(n_1281) );
AO21x1_ASAP7_75t_L g1621 ( .A1(n_901), .A2(n_1622), .B(n_1626), .Y(n_1621) );
INVx2_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx2_ASAP7_75t_L g1205 ( .A(n_906), .Y(n_1205) );
INVx1_ASAP7_75t_L g1267 ( .A(n_906), .Y(n_1267) );
INVx2_ASAP7_75t_SL g1278 ( .A(n_906), .Y(n_1278) );
INVx2_ASAP7_75t_L g1648 ( .A(n_906), .Y(n_1648) );
BUFx2_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
BUFx6f_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
BUFx3_ASAP7_75t_L g996 ( .A(n_909), .Y(n_996) );
INVx2_ASAP7_75t_L g1280 ( .A(n_909), .Y(n_1280) );
INVx3_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
AOI31xp33_ASAP7_75t_L g915 ( .A1(n_916), .A2(n_922), .A3(n_924), .B(n_927), .Y(n_915) );
HB1xp67_ASAP7_75t_L g956 ( .A(n_918), .Y(n_956) );
INVx1_ASAP7_75t_L g1616 ( .A(n_918), .Y(n_1616) );
INVx2_ASAP7_75t_SL g1035 ( .A(n_923), .Y(n_1035) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_925), .A2(n_926), .B1(n_1026), .B2(n_1027), .Y(n_1040) );
INVx2_ASAP7_75t_L g1243 ( .A(n_926), .Y(n_1243) );
AO21x1_ASAP7_75t_L g1236 ( .A1(n_927), .A2(n_1237), .B(n_1240), .Y(n_1236) );
CKINVDCx14_ASAP7_75t_R g927 ( .A(n_928), .Y(n_927) );
AOI22xp33_ASAP7_75t_SL g933 ( .A1(n_934), .A2(n_935), .B1(n_1172), .B2(n_1288), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
XNOR2xp5_ASAP7_75t_L g935 ( .A(n_936), .B(n_1041), .Y(n_935) );
INVx2_ASAP7_75t_SL g936 ( .A(n_937), .Y(n_936) );
XNOR2x1_ASAP7_75t_L g937 ( .A(n_938), .B(n_984), .Y(n_937) );
NAND3xp33_ASAP7_75t_L g939 ( .A(n_940), .B(n_949), .C(n_958), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g955 ( .A(n_945), .B(n_956), .Y(n_955) );
NOR2xp33_ASAP7_75t_L g958 ( .A(n_959), .B(n_974), .Y(n_958) );
OAI22xp5_ASAP7_75t_L g1149 ( .A1(n_965), .A2(n_1134), .B1(n_1142), .B2(n_1150), .Y(n_1149) );
OAI22xp5_ASAP7_75t_L g1063 ( .A1(n_978), .A2(n_1051), .B1(n_1054), .B2(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
NAND3xp33_ASAP7_75t_L g985 ( .A(n_986), .B(n_1023), .C(n_1033), .Y(n_985) );
AND4x1_ASAP7_75t_L g986 ( .A(n_987), .B(n_999), .C(n_1002), .D(n_1018), .Y(n_986) );
NAND3xp33_ASAP7_75t_L g987 ( .A(n_988), .B(n_993), .C(n_997), .Y(n_987) );
INVx1_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g1160 ( .A(n_992), .B(n_1161), .Y(n_1160) );
INVx2_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
INVx1_ASAP7_75t_L g1653 ( .A(n_995), .Y(n_1653) );
HB1xp67_ASAP7_75t_L g1268 ( .A(n_996), .Y(n_1268) );
INVx1_ASAP7_75t_L g1139 ( .A(n_997), .Y(n_1139) );
INVx2_ASAP7_75t_SL g997 ( .A(n_998), .Y(n_997) );
INVx2_ASAP7_75t_SL g1646 ( .A(n_998), .Y(n_1646) );
NAND3xp33_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1008), .C(n_1010), .Y(n_1002) );
BUFx3_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
BUFx12f_ASAP7_75t_L g1020 ( .A(n_1006), .Y(n_1020) );
BUFx2_ASAP7_75t_L g1227 ( .A(n_1006), .Y(n_1227) );
INVx5_ASAP7_75t_L g1257 ( .A(n_1006), .Y(n_1257) );
AND2x4_ASAP7_75t_L g1589 ( .A(n_1006), .B(n_1587), .Y(n_1589) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1007), .Y(n_1086) );
BUFx3_ASAP7_75t_L g1247 ( .A(n_1008), .Y(n_1247) );
INVx1_ASAP7_75t_L g1613 ( .A(n_1008), .Y(n_1613) );
INVx1_ASAP7_75t_L g1591 ( .A(n_1009), .Y(n_1591) );
INVx1_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
INVx1_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
BUFx2_ASAP7_75t_L g1562 ( .A(n_1013), .Y(n_1562) );
BUFx3_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
BUFx3_ASAP7_75t_L g1224 ( .A(n_1014), .Y(n_1224) );
INVx8_ASAP7_75t_L g1232 ( .A(n_1014), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1565 ( .A(n_1014), .B(n_1566), .Y(n_1565) );
NAND2x1p5_ASAP7_75t_L g1574 ( .A(n_1014), .B(n_1575), .Y(n_1574) );
INVx1_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
INVx2_ASAP7_75t_L g1252 ( .A(n_1017), .Y(n_1252) );
NAND3xp33_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1021), .C(n_1022), .Y(n_1018) );
XNOR2xp5_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1087), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
NAND3xp33_ASAP7_75t_L g1044 ( .A(n_1045), .B(n_1068), .C(n_1076), .Y(n_1044) );
NOR2xp33_ASAP7_75t_SL g1045 ( .A(n_1046), .B(n_1060), .Y(n_1045) );
INVxp67_ASAP7_75t_SL g1513 ( .A(n_1071), .Y(n_1513) );
AND2x6_ASAP7_75t_L g1579 ( .A(n_1083), .B(n_1575), .Y(n_1579) );
INVx3_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1581 ( .A(n_1086), .B(n_1575), .Y(n_1581) );
OAI22xp5_ASAP7_75t_L g1087 ( .A1(n_1088), .A2(n_1089), .B1(n_1127), .B2(n_1128), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1089), .Y(n_1088) );
NAND3xp33_ASAP7_75t_SL g1090 ( .A(n_1091), .B(n_1098), .C(n_1107), .Y(n_1090) );
NAND2xp5_ASAP7_75t_L g1101 ( .A(n_1096), .B(n_1102), .Y(n_1101) );
OAI31xp33_ASAP7_75t_SL g1098 ( .A1(n_1099), .A2(n_1100), .A3(n_1105), .B(n_1106), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g1168 ( .A(n_1102), .B(n_1159), .Y(n_1168) );
OAI31xp33_ASAP7_75t_L g1164 ( .A1(n_1106), .A2(n_1165), .A3(n_1166), .B(n_1169), .Y(n_1164) );
OAI31xp33_ASAP7_75t_SL g1638 ( .A1(n_1106), .A2(n_1639), .A3(n_1640), .B(n_1643), .Y(n_1638) );
NOR2xp33_ASAP7_75t_L g1107 ( .A(n_1108), .B(n_1121), .Y(n_1107) );
INVx3_ASAP7_75t_SL g1127 ( .A(n_1128), .Y(n_1127) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1129), .Y(n_1171) );
NAND3xp33_ASAP7_75t_L g1129 ( .A(n_1130), .B(n_1154), .C(n_1164), .Y(n_1129) );
NOR2xp33_ASAP7_75t_L g1130 ( .A(n_1131), .B(n_1146), .Y(n_1130) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
INVx1_ASAP7_75t_L g1619 ( .A(n_1152), .Y(n_1619) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1172), .Y(n_1288) );
OAI22xp5_ASAP7_75t_L g1172 ( .A1(n_1173), .A2(n_1233), .B1(n_1286), .B2(n_1287), .Y(n_1172) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1173), .Y(n_1286) );
HB1xp67_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
OAI21xp5_ASAP7_75t_L g1175 ( .A1(n_1176), .A2(n_1206), .B(n_1208), .Y(n_1175) );
OAI21xp5_ASAP7_75t_L g1189 ( .A1(n_1190), .A2(n_1193), .B(n_1197), .Y(n_1189) );
BUFx6f_ASAP7_75t_L g1200 ( .A(n_1201), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1595 ( .A(n_1201), .B(n_1541), .Y(n_1595) );
INVx2_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
BUFx2_ASAP7_75t_L g1206 ( .A(n_1207), .Y(n_1206) );
NAND2xp5_ASAP7_75t_SL g1209 ( .A(n_1210), .B(n_1216), .Y(n_1209) );
OAI211xp5_ASAP7_75t_L g1219 ( .A1(n_1220), .A2(n_1221), .B(n_1223), .C(n_1226), .Y(n_1219) );
INVx2_ASAP7_75t_SL g1221 ( .A(n_1222), .Y(n_1221) );
INVx2_ASAP7_75t_SL g1251 ( .A(n_1224), .Y(n_1251) );
BUFx2_ASAP7_75t_L g1259 ( .A(n_1225), .Y(n_1259) );
INVx2_ASAP7_75t_L g1231 ( .A(n_1232), .Y(n_1231) );
INVx8_ASAP7_75t_L g1558 ( .A(n_1232), .Y(n_1558) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1233), .Y(n_1287) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
NAND4xp25_ASAP7_75t_SL g1235 ( .A(n_1236), .B(n_1246), .C(n_1264), .D(n_1281), .Y(n_1235) );
AOI33xp33_ASAP7_75t_L g1246 ( .A1(n_1247), .A2(n_1248), .A3(n_1253), .B1(n_1258), .B2(n_1260), .B3(n_1263), .Y(n_1246) );
BUFx2_ASAP7_75t_SL g1249 ( .A(n_1250), .Y(n_1249) );
INVx2_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
OAI221xp5_ASAP7_75t_L g1615 ( .A1(n_1251), .A2(n_1616), .B1(n_1617), .B2(n_1618), .C(n_1619), .Y(n_1615) );
NAND2xp5_ASAP7_75t_L g1641 ( .A(n_1252), .B(n_1631), .Y(n_1641) );
INVx2_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1257), .Y(n_1256) );
INVx2_ASAP7_75t_L g1262 ( .A(n_1257), .Y(n_1262) );
INVx2_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
INVx2_ASAP7_75t_L g1271 ( .A(n_1272), .Y(n_1271) );
INVx2_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1280), .Y(n_1279) );
INVx3_ASAP7_75t_L g1542 ( .A(n_1280), .Y(n_1542) );
OAI221xp5_ASAP7_75t_L g1289 ( .A1(n_1290), .A2(n_1500), .B1(n_1502), .B2(n_1597), .C(n_1602), .Y(n_1289) );
AOI21xp5_ASAP7_75t_L g1290 ( .A1(n_1291), .A2(n_1413), .B(n_1457), .Y(n_1290) );
OAI211xp5_ASAP7_75t_L g1291 ( .A1(n_1292), .A2(n_1307), .B(n_1353), .C(n_1399), .Y(n_1291) );
AOI22xp5_ASAP7_75t_L g1482 ( .A1(n_1292), .A2(n_1405), .B1(n_1483), .B2(n_1489), .Y(n_1482) );
CKINVDCx5p33_ASAP7_75t_R g1292 ( .A(n_1293), .Y(n_1292) );
CKINVDCx6p67_ASAP7_75t_R g1365 ( .A(n_1293), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1466 ( .A(n_1293), .B(n_1325), .Y(n_1466) );
OR2x2_ASAP7_75t_L g1484 ( .A(n_1293), .B(n_1325), .Y(n_1484) );
OR2x2_ASAP7_75t_L g1499 ( .A(n_1293), .B(n_1389), .Y(n_1499) );
OR2x6_ASAP7_75t_L g1293 ( .A(n_1294), .B(n_1301), .Y(n_1293) );
OR2x2_ASAP7_75t_L g1386 ( .A(n_1294), .B(n_1301), .Y(n_1386) );
INVx2_ASAP7_75t_L g1396 ( .A(n_1295), .Y(n_1396) );
AND2x6_ASAP7_75t_L g1295 ( .A(n_1296), .B(n_1297), .Y(n_1295) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1296), .B(n_1300), .Y(n_1299) );
AND2x4_ASAP7_75t_L g1302 ( .A(n_1296), .B(n_1303), .Y(n_1302) );
AND2x6_ASAP7_75t_L g1305 ( .A(n_1296), .B(n_1306), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1296), .B(n_1300), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1322 ( .A(n_1296), .B(n_1300), .Y(n_1322) );
OAI21xp5_ASAP7_75t_L g1654 ( .A1(n_1297), .A2(n_1655), .B(n_1656), .Y(n_1654) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_1298), .B(n_1304), .Y(n_1303) );
O2A1O1Ixp33_ASAP7_75t_L g1307 ( .A1(n_1308), .A2(n_1323), .B(n_1328), .C(n_1342), .Y(n_1307) );
NOR2xp33_ASAP7_75t_L g1308 ( .A(n_1309), .B(n_1313), .Y(n_1308) );
INVx2_ASAP7_75t_L g1336 ( .A(n_1309), .Y(n_1336) );
NAND2xp5_ASAP7_75t_L g1343 ( .A(n_1309), .B(n_1344), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1350 ( .A(n_1309), .B(n_1318), .Y(n_1350) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1309), .Y(n_1358) );
AND2x2_ASAP7_75t_L g1380 ( .A(n_1309), .B(n_1381), .Y(n_1380) );
OR2x2_ASAP7_75t_L g1423 ( .A(n_1309), .B(n_1385), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1455 ( .A(n_1309), .B(n_1338), .Y(n_1455) );
OR2x2_ASAP7_75t_L g1472 ( .A(n_1309), .B(n_1338), .Y(n_1472) );
AND2x2_ASAP7_75t_L g1309 ( .A(n_1310), .B(n_1311), .Y(n_1309) );
INVxp67_ASAP7_75t_L g1398 ( .A(n_1312), .Y(n_1398) );
OR2x2_ASAP7_75t_L g1313 ( .A(n_1314), .B(n_1318), .Y(n_1313) );
AND2x2_ASAP7_75t_L g1352 ( .A(n_1314), .B(n_1347), .Y(n_1352) );
AND3x1_ASAP7_75t_L g1369 ( .A(n_1314), .B(n_1330), .C(n_1335), .Y(n_1369) );
AND2x2_ASAP7_75t_L g1376 ( .A(n_1314), .B(n_1330), .Y(n_1376) );
AND2x2_ASAP7_75t_L g1488 ( .A(n_1314), .B(n_1318), .Y(n_1488) );
INVx2_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_1315), .B(n_1330), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1360 ( .A(n_1315), .B(n_1347), .Y(n_1360) );
NAND2xp5_ASAP7_75t_L g1385 ( .A(n_1315), .B(n_1318), .Y(n_1385) );
OR2x2_ASAP7_75t_L g1315 ( .A(n_1316), .B(n_1317), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1318), .B(n_1347), .Y(n_1346) );
OR2x2_ASAP7_75t_L g1371 ( .A(n_1318), .B(n_1330), .Y(n_1371) );
AND2x2_ASAP7_75t_L g1438 ( .A(n_1318), .B(n_1376), .Y(n_1438) );
AND2x2_ASAP7_75t_L g1453 ( .A(n_1318), .B(n_1330), .Y(n_1453) );
BUFx2_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
INVx2_ASAP7_75t_L g1335 ( .A(n_1319), .Y(n_1335) );
AND2x2_ASAP7_75t_L g1367 ( .A(n_1319), .B(n_1329), .Y(n_1367) );
AND2x2_ASAP7_75t_L g1388 ( .A(n_1319), .B(n_1352), .Y(n_1388) );
AND2x2_ASAP7_75t_L g1420 ( .A(n_1319), .B(n_1360), .Y(n_1420) );
OR2x2_ASAP7_75t_L g1441 ( .A(n_1319), .B(n_1442), .Y(n_1441) );
AND2x2_ASAP7_75t_L g1319 ( .A(n_1320), .B(n_1321), .Y(n_1319) );
O2A1O1Ixp33_ASAP7_75t_L g1328 ( .A1(n_1323), .A2(n_1329), .B(n_1333), .C(n_1337), .Y(n_1328) );
CKINVDCx14_ASAP7_75t_R g1323 ( .A(n_1324), .Y(n_1323) );
OAI22xp5_ASAP7_75t_L g1406 ( .A1(n_1324), .A2(n_1404), .B1(n_1407), .B2(n_1410), .Y(n_1406) );
NAND2xp5_ASAP7_75t_L g1424 ( .A(n_1324), .B(n_1392), .Y(n_1424) );
AOI211xp5_ASAP7_75t_L g1448 ( .A1(n_1324), .A2(n_1449), .B(n_1450), .C(n_1451), .Y(n_1448) );
AOI221xp5_ASAP7_75t_L g1458 ( .A1(n_1324), .A2(n_1369), .B1(n_1459), .B2(n_1461), .C(n_1462), .Y(n_1458) );
INVx3_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1325), .Y(n_1341) );
OR2x2_ASAP7_75t_L g1355 ( .A(n_1325), .B(n_1338), .Y(n_1355) );
AOI22xp5_ASAP7_75t_L g1379 ( .A1(n_1325), .A2(n_1380), .B1(n_1383), .B2(n_1384), .Y(n_1379) );
AND2x2_ASAP7_75t_L g1383 ( .A(n_1325), .B(n_1338), .Y(n_1383) );
AND2x2_ASAP7_75t_L g1390 ( .A(n_1325), .B(n_1344), .Y(n_1390) );
OR2x2_ASAP7_75t_L g1436 ( .A(n_1325), .B(n_1365), .Y(n_1436) );
AND2x2_ASAP7_75t_L g1454 ( .A(n_1325), .B(n_1455), .Y(n_1454) );
AND2x2_ASAP7_75t_L g1481 ( .A(n_1325), .B(n_1365), .Y(n_1481) );
AND2x4_ASAP7_75t_L g1325 ( .A(n_1326), .B(n_1327), .Y(n_1325) );
NAND2xp5_ASAP7_75t_L g1403 ( .A(n_1329), .B(n_1336), .Y(n_1403) );
INVx1_ASAP7_75t_L g1442 ( .A(n_1329), .Y(n_1442) );
AND2x2_ASAP7_75t_L g1486 ( .A(n_1329), .B(n_1350), .Y(n_1486) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1330), .Y(n_1347) );
NAND2xp5_ASAP7_75t_L g1382 ( .A(n_1330), .B(n_1335), .Y(n_1382) );
AND2x2_ASAP7_75t_L g1330 ( .A(n_1331), .B(n_1332), .Y(n_1330) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
AND2x2_ASAP7_75t_L g1491 ( .A(n_1334), .B(n_1352), .Y(n_1491) );
AND2x2_ASAP7_75t_L g1334 ( .A(n_1335), .B(n_1336), .Y(n_1334) );
AND2x2_ASAP7_75t_L g1359 ( .A(n_1335), .B(n_1360), .Y(n_1359) );
OR2x2_ASAP7_75t_L g1402 ( .A(n_1335), .B(n_1403), .Y(n_1402) );
AND2x2_ASAP7_75t_L g1445 ( .A(n_1335), .B(n_1352), .Y(n_1445) );
OR2x2_ASAP7_75t_L g1494 ( .A(n_1335), .B(n_1412), .Y(n_1494) );
NAND2xp5_ASAP7_75t_SL g1496 ( .A(n_1335), .B(n_1497), .Y(n_1496) );
NOR2xp33_ASAP7_75t_L g1374 ( .A(n_1336), .B(n_1375), .Y(n_1374) );
NOR2xp33_ASAP7_75t_L g1409 ( .A(n_1336), .B(n_1371), .Y(n_1409) );
NAND2xp5_ASAP7_75t_L g1419 ( .A(n_1336), .B(n_1364), .Y(n_1419) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1336), .Y(n_1447) );
NAND2xp5_ASAP7_75t_L g1479 ( .A(n_1336), .B(n_1453), .Y(n_1479) );
AND2x2_ASAP7_75t_L g1372 ( .A(n_1337), .B(n_1365), .Y(n_1372) );
INVx1_ASAP7_75t_L g1430 ( .A(n_1337), .Y(n_1430) );
AND2x2_ASAP7_75t_L g1337 ( .A(n_1338), .B(n_1341), .Y(n_1337) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1338), .Y(n_1344) );
AND2x2_ASAP7_75t_L g1338 ( .A(n_1339), .B(n_1340), .Y(n_1338) );
OAI21xp33_ASAP7_75t_L g1342 ( .A1(n_1343), .A2(n_1345), .B(n_1348), .Y(n_1342) );
INVx2_ASAP7_75t_L g1364 ( .A(n_1344), .Y(n_1364) );
AND2x2_ASAP7_75t_L g1377 ( .A(n_1344), .B(n_1365), .Y(n_1377) );
OAI211xp5_ASAP7_75t_SL g1415 ( .A1(n_1345), .A2(n_1416), .B(n_1417), .C(n_1421), .Y(n_1415) );
NAND2xp5_ASAP7_75t_L g1440 ( .A(n_1345), .B(n_1441), .Y(n_1440) );
INVx1_ASAP7_75t_L g1345 ( .A(n_1346), .Y(n_1345) );
A2O1A1Ixp33_ASAP7_75t_L g1373 ( .A1(n_1346), .A2(n_1358), .B(n_1374), .C(n_1377), .Y(n_1373) );
AOI221xp5_ASAP7_75t_L g1399 ( .A1(n_1346), .A2(n_1400), .B1(n_1401), .B2(n_1404), .C(n_1406), .Y(n_1399) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1348), .Y(n_1449) );
OR2x2_ASAP7_75t_L g1476 ( .A(n_1348), .B(n_1364), .Y(n_1476) );
OR2x2_ASAP7_75t_L g1348 ( .A(n_1349), .B(n_1351), .Y(n_1348) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1350), .Y(n_1349) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1352), .Y(n_1351) );
NAND2xp5_ASAP7_75t_L g1412 ( .A(n_1352), .B(n_1358), .Y(n_1412) );
AOI211xp5_ASAP7_75t_L g1353 ( .A1(n_1354), .A2(n_1356), .B(n_1361), .C(n_1378), .Y(n_1353) );
AND2x2_ASAP7_75t_L g1400 ( .A(n_1354), .B(n_1358), .Y(n_1400) );
OAI322xp33_ASAP7_75t_L g1427 ( .A1(n_1354), .A2(n_1371), .A3(n_1386), .B1(n_1403), .B2(n_1428), .C1(n_1431), .C2(n_1433), .Y(n_1427) );
AND2x2_ASAP7_75t_SL g1450 ( .A(n_1354), .B(n_1369), .Y(n_1450) );
NAND2xp5_ASAP7_75t_L g1460 ( .A(n_1354), .B(n_1357), .Y(n_1460) );
INVx2_ASAP7_75t_L g1354 ( .A(n_1355), .Y(n_1354) );
AND2x2_ASAP7_75t_L g1356 ( .A(n_1357), .B(n_1359), .Y(n_1356) );
NOR2xp33_ASAP7_75t_L g1370 ( .A(n_1357), .B(n_1371), .Y(n_1370) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1357), .Y(n_1432) );
AOI31xp33_ASAP7_75t_L g1439 ( .A1(n_1357), .A2(n_1435), .A3(n_1440), .B(n_1443), .Y(n_1439) );
AND2x2_ASAP7_75t_L g1480 ( .A(n_1357), .B(n_1369), .Y(n_1480) );
INVx2_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
NAND2xp5_ASAP7_75t_SL g1416 ( .A(n_1358), .B(n_1383), .Y(n_1416) );
AND2x2_ASAP7_75t_L g1437 ( .A(n_1358), .B(n_1438), .Y(n_1437) );
NAND2xp5_ASAP7_75t_L g1431 ( .A(n_1359), .B(n_1432), .Y(n_1431) );
OR2x2_ASAP7_75t_L g1497 ( .A(n_1360), .B(n_1376), .Y(n_1497) );
OAI211xp5_ASAP7_75t_L g1361 ( .A1(n_1362), .A2(n_1366), .B(n_1368), .C(n_1373), .Y(n_1361) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1363), .Y(n_1362) );
AND2x2_ASAP7_75t_L g1363 ( .A(n_1364), .B(n_1365), .Y(n_1363) );
INVx2_ASAP7_75t_L g1405 ( .A(n_1364), .Y(n_1405) );
A2O1A1Ixp33_ASAP7_75t_L g1477 ( .A1(n_1364), .A2(n_1478), .B(n_1480), .C(n_1481), .Y(n_1477) );
NAND2xp5_ASAP7_75t_L g1425 ( .A(n_1365), .B(n_1426), .Y(n_1425) );
NOR2xp33_ASAP7_75t_SL g1429 ( .A(n_1365), .B(n_1430), .Y(n_1429) );
NOR2xp33_ASAP7_75t_L g1471 ( .A(n_1365), .B(n_1472), .Y(n_1471) );
O2A1O1Ixp33_ASAP7_75t_L g1462 ( .A1(n_1366), .A2(n_1463), .B(n_1464), .C(n_1465), .Y(n_1462) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1367), .Y(n_1366) );
OAI21xp33_ASAP7_75t_L g1368 ( .A1(n_1369), .A2(n_1370), .B(n_1372), .Y(n_1368) );
NAND2xp5_ASAP7_75t_L g1456 ( .A(n_1372), .B(n_1388), .Y(n_1456) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1376), .Y(n_1375) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1377), .Y(n_1433) );
OAI221xp5_ASAP7_75t_L g1378 ( .A1(n_1379), .A2(n_1386), .B1(n_1387), .B2(n_1389), .C(n_1391), .Y(n_1378) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1382), .Y(n_1381) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1385), .Y(n_1384) );
AOI22xp5_ASAP7_75t_L g1467 ( .A1(n_1386), .A2(n_1468), .B1(n_1473), .B2(n_1475), .Y(n_1467) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1388), .Y(n_1387) );
CKINVDCx6p67_ASAP7_75t_R g1389 ( .A(n_1390), .Y(n_1389) );
NAND2xp5_ASAP7_75t_L g1446 ( .A(n_1390), .B(n_1447), .Y(n_1446) );
INVx3_ASAP7_75t_L g1391 ( .A(n_1392), .Y(n_1391) );
INVx2_ASAP7_75t_SL g1392 ( .A(n_1393), .Y(n_1392) );
OAI21xp33_ASAP7_75t_L g1421 ( .A1(n_1393), .A2(n_1422), .B(n_1424), .Y(n_1421) );
INVx2_ASAP7_75t_SL g1426 ( .A(n_1393), .Y(n_1426) );
OAI22xp5_ASAP7_75t_SL g1394 ( .A1(n_1395), .A2(n_1396), .B1(n_1397), .B2(n_1398), .Y(n_1394) );
CKINVDCx20_ASAP7_75t_R g1501 ( .A(n_1396), .Y(n_1501) );
INVx1_ASAP7_75t_L g1469 ( .A(n_1400), .Y(n_1469) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1402), .Y(n_1401) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1404), .B(n_1409), .Y(n_1408) );
AND2x2_ASAP7_75t_L g1461 ( .A(n_1404), .B(n_1449), .Y(n_1461) );
NAND2xp5_ASAP7_75t_L g1490 ( .A(n_1404), .B(n_1491), .Y(n_1490) );
INVx2_ASAP7_75t_L g1404 ( .A(n_1405), .Y(n_1404) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
INVx1_ASAP7_75t_L g1410 ( .A(n_1411), .Y(n_1410) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1412), .Y(n_1411) );
NAND5xp2_ASAP7_75t_L g1413 ( .A(n_1414), .B(n_1434), .C(n_1439), .D(n_1448), .E(n_1456), .Y(n_1413) );
AOI21xp5_ASAP7_75t_L g1414 ( .A1(n_1415), .A2(n_1425), .B(n_1427), .Y(n_1414) );
NAND2xp5_ASAP7_75t_L g1417 ( .A(n_1418), .B(n_1420), .Y(n_1417) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1419), .Y(n_1418) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1423), .Y(n_1422) );
NAND3xp33_ASAP7_75t_L g1478 ( .A(n_1423), .B(n_1444), .C(n_1479), .Y(n_1478) );
INVx1_ASAP7_75t_L g1428 ( .A(n_1429), .Y(n_1428) );
NAND2xp5_ASAP7_75t_L g1434 ( .A(n_1435), .B(n_1437), .Y(n_1434) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
OAI22xp5_ASAP7_75t_L g1483 ( .A1(n_1436), .A2(n_1484), .B1(n_1485), .B2(n_1487), .Y(n_1483) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1438), .Y(n_1474) );
AOI21xp33_ASAP7_75t_L g1443 ( .A1(n_1442), .A2(n_1444), .B(n_1446), .Y(n_1443) );
NAND2xp5_ASAP7_75t_L g1473 ( .A(n_1444), .B(n_1474), .Y(n_1473) );
INVx1_ASAP7_75t_L g1444 ( .A(n_1445), .Y(n_1444) );
INVxp67_ASAP7_75t_SL g1451 ( .A(n_1452), .Y(n_1451) );
NAND2xp5_ASAP7_75t_L g1452 ( .A(n_1453), .B(n_1454), .Y(n_1452) );
INVx1_ASAP7_75t_L g1463 ( .A(n_1453), .Y(n_1463) );
CKINVDCx14_ASAP7_75t_R g1464 ( .A(n_1455), .Y(n_1464) );
NAND5xp2_ASAP7_75t_L g1457 ( .A(n_1458), .B(n_1467), .C(n_1477), .D(n_1482), .E(n_1492), .Y(n_1457) );
INVx1_ASAP7_75t_L g1459 ( .A(n_1460), .Y(n_1459) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1466), .Y(n_1465) );
NAND2xp5_ASAP7_75t_SL g1468 ( .A(n_1469), .B(n_1470), .Y(n_1468) );
INVxp67_ASAP7_75t_L g1470 ( .A(n_1471), .Y(n_1470) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1476), .Y(n_1475) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1486), .Y(n_1485) );
CKINVDCx14_ASAP7_75t_R g1487 ( .A(n_1488), .Y(n_1487) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1490), .Y(n_1489) );
OAI21xp5_ASAP7_75t_L g1492 ( .A1(n_1493), .A2(n_1495), .B(n_1498), .Y(n_1492) );
INVx1_ASAP7_75t_L g1493 ( .A(n_1494), .Y(n_1493) );
INVxp67_ASAP7_75t_SL g1495 ( .A(n_1496), .Y(n_1495) );
INVx1_ASAP7_75t_L g1498 ( .A(n_1499), .Y(n_1498) );
CKINVDCx20_ASAP7_75t_R g1500 ( .A(n_1501), .Y(n_1500) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1503), .Y(n_1502) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1504), .Y(n_1503) );
XNOR2x1_ASAP7_75t_L g1504 ( .A(n_1505), .B(n_1596), .Y(n_1504) );
OR2x2_ASAP7_75t_L g1505 ( .A(n_1506), .B(n_1554), .Y(n_1505) );
NAND3xp33_ASAP7_75t_SL g1506 ( .A(n_1507), .B(n_1531), .C(n_1547), .Y(n_1506) );
AOI211xp5_ASAP7_75t_SL g1507 ( .A1(n_1508), .A2(n_1512), .B(n_1514), .C(n_1525), .Y(n_1507) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1511), .Y(n_1510) );
NAND2x2_ASAP7_75t_L g1515 ( .A(n_1516), .B(n_1519), .Y(n_1515) );
INVx1_ASAP7_75t_L g1524 ( .A(n_1516), .Y(n_1524) );
INVx2_ASAP7_75t_L g1516 ( .A(n_1517), .Y(n_1516) );
INVx2_ASAP7_75t_SL g1519 ( .A(n_1520), .Y(n_1519) );
INVx1_ASAP7_75t_L g1526 ( .A(n_1527), .Y(n_1526) );
AOI222xp33_ASAP7_75t_L g1531 ( .A1(n_1532), .A2(n_1537), .B1(n_1538), .B2(n_1543), .C1(n_1544), .C2(n_1546), .Y(n_1531) );
AND2x4_ASAP7_75t_L g1532 ( .A(n_1533), .B(n_1535), .Y(n_1532) );
INVx1_ASAP7_75t_L g1533 ( .A(n_1534), .Y(n_1533) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1536), .Y(n_1535) );
AND2x4_ASAP7_75t_L g1538 ( .A(n_1539), .B(n_1542), .Y(n_1538) );
INVx1_ASAP7_75t_L g1539 ( .A(n_1540), .Y(n_1539) );
AOI211xp5_ASAP7_75t_L g1570 ( .A1(n_1543), .A2(n_1571), .B(n_1577), .C(n_1584), .Y(n_1570) );
INVx2_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
NAND2xp5_ASAP7_75t_L g1547 ( .A(n_1548), .B(n_1549), .Y(n_1547) );
INVx1_ASAP7_75t_L g1549 ( .A(n_1550), .Y(n_1549) );
INVx3_ASAP7_75t_L g1550 ( .A(n_1551), .Y(n_1550) );
AND2x4_ASAP7_75t_L g1551 ( .A(n_1552), .B(n_1553), .Y(n_1551) );
AND2x4_ASAP7_75t_L g1594 ( .A(n_1552), .B(n_1595), .Y(n_1594) );
A2O1A1Ixp33_ASAP7_75t_L g1554 ( .A1(n_1555), .A2(n_1570), .B(n_1590), .C(n_1592), .Y(n_1554) );
AOI221xp5_ASAP7_75t_L g1555 ( .A1(n_1556), .A2(n_1557), .B1(n_1559), .B2(n_1561), .C(n_1563), .Y(n_1555) );
INVx2_ASAP7_75t_L g1564 ( .A(n_1565), .Y(n_1564) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
INVx1_ASAP7_75t_L g1587 ( .A(n_1567), .Y(n_1587) );
INVx1_ASAP7_75t_L g1568 ( .A(n_1569), .Y(n_1568) );
INVx1_ASAP7_75t_L g1571 ( .A(n_1572), .Y(n_1571) );
INVx2_ASAP7_75t_L g1572 ( .A(n_1573), .Y(n_1572) );
INVx2_ASAP7_75t_L g1573 ( .A(n_1574), .Y(n_1573) );
INVx1_ASAP7_75t_L g1583 ( .A(n_1575), .Y(n_1583) );
INVx4_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
INVx2_ASAP7_75t_L g1580 ( .A(n_1581), .Y(n_1580) );
INVx2_ASAP7_75t_L g1586 ( .A(n_1587), .Y(n_1586) );
INVx3_ASAP7_75t_L g1588 ( .A(n_1589), .Y(n_1588) );
BUFx2_ASAP7_75t_L g1590 ( .A(n_1591), .Y(n_1590) );
NAND2xp5_ASAP7_75t_L g1592 ( .A(n_1593), .B(n_1594), .Y(n_1592) );
INVx2_ASAP7_75t_L g1597 ( .A(n_1598), .Y(n_1597) );
BUFx3_ASAP7_75t_L g1598 ( .A(n_1599), .Y(n_1598) );
BUFx3_ASAP7_75t_L g1603 ( .A(n_1604), .Y(n_1603) );
BUFx3_ASAP7_75t_L g1604 ( .A(n_1605), .Y(n_1604) );
INVxp33_ASAP7_75t_SL g1606 ( .A(n_1607), .Y(n_1606) );
NOR4xp25_ASAP7_75t_L g1608 ( .A(n_1609), .B(n_1620), .C(n_1637), .D(n_1644), .Y(n_1608) );
INVx1_ASAP7_75t_L g1609 ( .A(n_1610), .Y(n_1609) );
AOI21xp5_ASAP7_75t_L g1610 ( .A1(n_1611), .A2(n_1612), .B(n_1614), .Y(n_1610) );
INVxp67_ASAP7_75t_SL g1620 ( .A(n_1621), .Y(n_1620) );
NOR2xp33_ASAP7_75t_L g1626 ( .A(n_1627), .B(n_1628), .Y(n_1626) );
NAND3xp33_ASAP7_75t_L g1628 ( .A(n_1629), .B(n_1632), .C(n_1636), .Y(n_1628) );
NAND2xp5_ASAP7_75t_L g1632 ( .A(n_1633), .B(n_1634), .Y(n_1632) );
INVx2_ASAP7_75t_L g1634 ( .A(n_1635), .Y(n_1634) );
INVxp67_ASAP7_75t_SL g1637 ( .A(n_1638), .Y(n_1637) );
INVx1_ASAP7_75t_L g1644 ( .A(n_1645), .Y(n_1644) );
INVx1_ASAP7_75t_L g1656 ( .A(n_1657), .Y(n_1656) );
endmodule