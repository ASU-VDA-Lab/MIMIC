module real_jpeg_32497_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_681, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_681;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_669;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_553;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_678;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_611;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_673;
wire n_631;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_195;
wire n_110;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_579;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_670;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_638;
wire n_497;
wire n_633;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_572;
wire n_412;
wire n_405;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_613;
wire n_265;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_667;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g225 ( 
.A(n_0),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_0),
.Y(n_228)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_0),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_0),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_0),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_1),
.A2(n_345),
.B1(n_346),
.B2(n_348),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_1),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_1),
.A2(n_345),
.B1(n_439),
.B2(n_441),
.Y(n_438)
);

AOI22xp33_ASAP7_75t_SL g552 ( 
.A1(n_1),
.A2(n_345),
.B1(n_553),
.B2(n_557),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_SL g590 ( 
.A1(n_1),
.A2(n_345),
.B1(n_591),
.B2(n_593),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_2),
.A2(n_68),
.B1(n_74),
.B2(n_75),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_2),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_2),
.A2(n_74),
.B1(n_173),
.B2(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_2),
.A2(n_74),
.B1(n_280),
.B2(n_282),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g413 ( 
.A1(n_2),
.A2(n_74),
.B1(n_414),
.B2(n_417),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_3),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_5),
.A2(n_149),
.B1(n_150),
.B2(n_154),
.Y(n_148)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_5),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_5),
.A2(n_154),
.B1(n_181),
.B2(n_186),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_5),
.A2(n_154),
.B1(n_236),
.B2(n_239),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_5),
.A2(n_154),
.B1(n_329),
.B2(n_333),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_6),
.A2(n_187),
.B1(n_246),
.B2(n_249),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_6),
.Y(n_249)
);

OAI22x1_ASAP7_75t_SL g355 ( 
.A1(n_6),
.A2(n_249),
.B1(n_356),
.B2(n_359),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_6),
.A2(n_249),
.B1(n_458),
.B2(n_460),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_6),
.A2(n_249),
.B1(n_515),
.B2(n_517),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_7),
.Y(n_185)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_8),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_8),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_9),
.A2(n_57),
.B1(n_58),
.B2(n_62),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_9),
.A2(n_57),
.B1(n_305),
.B2(n_308),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_9),
.A2(n_57),
.B1(n_282),
.B2(n_340),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_9),
.A2(n_57),
.B1(n_483),
.B2(n_486),
.Y(n_482)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_10),
.Y(n_84)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_10),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_10),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_10),
.Y(n_232)
);

AO22x1_ASAP7_75t_L g156 ( 
.A1(n_11),
.A2(n_157),
.B1(n_161),
.B2(n_162),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_11),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_11),
.A2(n_161),
.B1(n_206),
.B2(n_210),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_11),
.A2(n_161),
.B1(n_269),
.B2(n_271),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_12),
.B(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_12),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_12),
.B(n_66),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_12),
.B(n_521),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_SL g543 ( 
.A1(n_12),
.A2(n_452),
.B1(n_544),
.B2(n_547),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_12),
.B(n_155),
.Y(n_569)
);

OAI21xp33_ASAP7_75t_L g599 ( 
.A1(n_12),
.A2(n_272),
.B(n_579),
.Y(n_599)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_13),
.Y(n_88)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_13),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_14),
.B(n_256),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_14),
.Y(n_679)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_15),
.A2(n_108),
.B1(n_114),
.B2(n_115),
.Y(n_107)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_15),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_15),
.A2(n_114),
.B1(n_172),
.B2(n_175),
.Y(n_171)
);

AO22x1_ASAP7_75t_SL g229 ( 
.A1(n_15),
.A2(n_114),
.B1(n_230),
.B2(n_233),
.Y(n_229)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_16),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_16),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_16),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_16),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_17),
.A2(n_294),
.B1(n_295),
.B2(n_298),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_17),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_17),
.A2(n_294),
.B1(n_383),
.B2(n_385),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_SL g503 ( 
.A1(n_17),
.A2(n_294),
.B1(n_504),
.B2(n_508),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_SL g571 ( 
.A1(n_17),
.A2(n_294),
.B1(n_572),
.B2(n_577),
.Y(n_571)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_18),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_18),
.Y(n_160)
);

NAND4xp25_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_669),
.C(n_673),
.D(n_676),
.Y(n_19)
);

NAND3xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_253),
.C(n_319),
.Y(n_20)
);

NAND3xp33_ASAP7_75t_L g669 ( 
.A(n_21),
.B(n_253),
.C(n_670),
.Y(n_669)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_21),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_251),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_193),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_24),
.B(n_193),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_166),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_77),
.C(n_118),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_26),
.A2(n_27),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_L g194 ( 
.A1(n_26),
.A2(n_27),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_R g314 ( 
.A(n_26),
.B(n_200),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_26),
.B(n_199),
.Y(n_317)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_27),
.B(n_200),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_27),
.B(n_199),
.Y(n_318)
);

AO22x2_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_56),
.B1(n_65),
.B2(n_67),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_28),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_28),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_28),
.B(n_293),
.Y(n_292)
);

AO22x1_ASAP7_75t_SL g343 ( 
.A1(n_28),
.A2(n_66),
.B1(n_293),
.B2(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_28),
.B(n_447),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_44),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_34),
.B1(n_38),
.B2(n_41),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_37),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_37),
.Y(n_407)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_39),
.Y(n_248)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_40),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_40),
.Y(n_349)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B1(n_51),
.B2(n_54),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_49),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g444 ( 
.A(n_49),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_50),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_50),
.Y(n_362)
);

BUFx5_ASAP7_75t_L g404 ( 
.A(n_50),
.Y(n_404)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_53),
.Y(n_546)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_56),
.B(n_66),
.Y(n_250)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_64),
.Y(n_395)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_65),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_66),
.B(n_245),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_66),
.B(n_344),
.Y(n_380)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_67),
.Y(n_190)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_77),
.B(n_170),
.Y(n_169)
);

XOR2x2_ASAP7_75t_L g196 ( 
.A(n_77),
.B(n_118),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_107),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_97),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_79),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_79),
.A2(n_97),
.B1(n_205),
.B2(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_79),
.A2(n_97),
.B1(n_235),
.B2(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_79),
.A2(n_97),
.B1(n_279),
.B2(n_339),
.Y(n_338)
);

OAI22xp33_ASAP7_75t_L g551 ( 
.A1(n_79),
.A2(n_97),
.B1(n_503),
.B2(n_552),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_L g566 ( 
.A1(n_79),
.A2(n_552),
.B(n_567),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_SL g588 ( 
.A(n_79),
.B(n_452),
.Y(n_588)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_80),
.A2(n_203),
.B1(n_456),
.B2(n_457),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_80),
.B(n_457),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_98),
.Y(n_97)
);

OAI22x1_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B1(n_89),
.B2(n_93),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_82),
.Y(n_271)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_83),
.Y(n_416)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_84),
.Y(n_332)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_84),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_84),
.Y(n_621)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx6_ASAP7_75t_L g626 ( 
.A(n_91),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_94),
.Y(n_518)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_97),
.Y(n_203)
);

OAI21xp33_ASAP7_75t_SL g502 ( 
.A1(n_97),
.A2(n_503),
.B(n_509),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_100),
.Y(n_281)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_101),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_105),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_106),
.Y(n_507)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_106),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_107),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_201)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_112),
.Y(n_240)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_112),
.Y(n_463)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_117),
.Y(n_529)
);

AO22x1_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_148),
.B1(n_155),
.B2(n_156),
.Y(n_118)
);

AO22x1_ASAP7_75t_L g170 ( 
.A1(n_119),
.A2(n_155),
.B1(n_156),
.B2(n_171),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_119),
.A2(n_148),
.B1(n_155),
.B2(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_119),
.A2(n_155),
.B1(n_213),
.B2(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g363 ( 
.A(n_119),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_119),
.A2(n_155),
.B1(n_437),
.B2(n_438),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_119),
.B(n_355),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_134),
.Y(n_119)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

AOI22x1_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_124),
.B1(n_127),
.B2(n_131),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_123),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_130),
.Y(n_535)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_140),
.B1(n_143),
.B2(n_146),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_139),
.Y(n_392)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_153),
.Y(n_440)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_153),
.Y(n_526)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_155),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_155),
.B(n_355),
.Y(n_387)
);

INVx3_ASAP7_75t_SL g157 ( 
.A(n_158),
.Y(n_157)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx5_ASAP7_75t_L g358 ( 
.A(n_159),
.Y(n_358)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_160),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_160),
.Y(n_384)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_165),
.Y(n_531)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_165),
.Y(n_549)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2x1_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_178),
.Y(n_168)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVxp67_ASAP7_75t_SL g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_177),
.Y(n_309)
);

OA22x2_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_190),
.B2(n_191),
.Y(n_178)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_182),
.Y(n_400)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_184),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_185),
.Y(n_297)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx11_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.C(n_217),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_195),
.A2(n_196),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_195),
.A2(n_196),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_196),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

OA21x2_ASAP7_75t_SL g261 ( 
.A1(n_200),
.A2(n_201),
.B(n_212),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_212),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_203),
.B(n_457),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_203),
.B(n_644),
.Y(n_643)
);

INVxp67_ASAP7_75t_SL g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx6f_ASAP7_75t_SL g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_208),
.Y(n_342)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_209),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_209),
.Y(n_641)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_217),
.B(n_312),
.Y(n_311)
);

OA21x2_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_241),
.B(n_242),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_218),
.B(n_264),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_234),
.Y(n_218)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_219),
.B(n_243),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_219),
.A2(n_234),
.B1(n_241),
.B2(n_366),
.Y(n_365)
);

OA21x2_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_226),
.B(n_229),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_220),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_220),
.A2(n_328),
.B1(n_409),
.B2(n_412),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_220),
.B(n_514),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_220),
.A2(n_611),
.B1(n_612),
.B2(n_613),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_224),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_221),
.Y(n_270)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_222),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_222),
.Y(n_334)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_222),
.Y(n_418)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_223),
.Y(n_487)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_223),
.Y(n_636)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx8_ASAP7_75t_L g581 ( 
.A(n_225),
.Y(n_581)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_227),
.A2(n_272),
.B1(n_413),
.B2(n_482),
.Y(n_481)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_228),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_229),
.B(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_232),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_232),
.Y(n_592)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_234),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_240),
.Y(n_459)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_240),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_250),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_244),
.B(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.Y(n_253)
);

NAND4xp25_ASAP7_75t_L g673 ( 
.A(n_254),
.B(n_671),
.C(n_674),
.D(n_675),
.Y(n_673)
);

AOI31xp33_ASAP7_75t_L g676 ( 
.A1(n_254),
.A2(n_258),
.A3(n_675),
.B(n_677),
.Y(n_676)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_255),
.B(n_678),
.Y(n_677)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_258),
.Y(n_257)
);

NOR2xp67_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_311),
.Y(n_258)
);

NAND2xp33_ASAP7_75t_L g672 ( 
.A(n_259),
.B(n_311),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_265),
.B(n_310),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp33_ASAP7_75t_R g310 ( 
.A(n_261),
.B(n_262),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_261),
.B(n_263),
.Y(n_371)
);

INVxp33_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2x1_ASAP7_75t_L g370 ( 
.A(n_265),
.B(n_371),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_288),
.C(n_301),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_266),
.B(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_278),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_267),
.B(n_421),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_272),
.B(n_273),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_268),
.A2(n_272),
.B1(n_327),
.B2(n_335),
.Y(n_326)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g570 ( 
.A1(n_272),
.A2(n_571),
.B(n_579),
.Y(n_570)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_274),
.Y(n_512)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_277),
.Y(n_411)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_277),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_278),
.Y(n_421)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_284),
.Y(n_508)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_286),
.Y(n_631)
);

INVx5_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_290),
.B(n_303),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_291),
.B(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_297),
.Y(n_300)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_297),
.Y(n_347)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVxp33_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_304),
.Y(n_353)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_316),
.Y(n_312)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_319),
.Y(n_674)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_490),
.B(n_660),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_426),
.Y(n_321)
);

AOI21x1_ASAP7_75t_L g660 ( 
.A1(n_322),
.A2(n_661),
.B(n_665),
.Y(n_660)
);

OA21x2_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_370),
.B(n_372),
.Y(n_322)
);

NOR2x1_ASAP7_75t_SL g666 ( 
.A(n_323),
.B(n_370),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_323),
.B(n_370),
.Y(n_668)
);

MAJx2_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_364),
.C(n_367),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_324),
.B(n_374),
.Y(n_373)
);

MAJx2_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_343),
.C(n_350),
.Y(n_324)
);

XNOR2x1_ASAP7_75t_L g423 ( 
.A(n_325),
.B(n_424),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_338),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_326),
.B(n_338),
.Y(n_464)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_329),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

BUFx12f_ASAP7_75t_L g516 ( 
.A(n_332),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

BUFx4f_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_339),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_341),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_343),
.B(n_351),
.Y(n_424)
);

INVx2_ASAP7_75t_SL g346 ( 
.A(n_347),
.Y(n_346)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_352),
.A2(n_353),
.B1(n_354),
.B2(n_363),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_352),
.A2(n_479),
.B(n_480),
.Y(n_478)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_360),
.Y(n_386)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

OA21x2_ASAP7_75t_L g381 ( 
.A1(n_363),
.A2(n_382),
.B(n_387),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g542 ( 
.A1(n_363),
.A2(n_387),
.B(n_543),
.Y(n_542)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_365),
.B(n_368),
.Y(n_374)
);

INVxp33_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_375),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g667 ( 
.A(n_373),
.B(n_375),
.Y(n_667)
);

OAI21x1_ASAP7_75t_L g375 ( 
.A1(n_376),
.A2(n_422),
.B(n_425),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_419),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_377),
.B(n_419),
.Y(n_425)
);

XOR2x1_ASAP7_75t_L g465 ( 
.A(n_377),
.B(n_466),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_381),
.C(n_388),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_378),
.A2(n_379),
.B1(n_381),
.B2(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_381),
.Y(n_432)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_382),
.Y(n_437)
);

INVx8_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_388),
.B(n_431),
.Y(n_430)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_408),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_389),
.B(n_408),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_390),
.A2(n_393),
.B1(n_399),
.B2(n_401),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_396),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_399),
.Y(n_453)
);

NAND2xp33_ASAP7_75t_SL g401 ( 
.A(n_402),
.B(n_405),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_SL g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx2_ASAP7_75t_SL g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_SL g414 ( 
.A(n_415),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_420),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

XNOR2x1_ASAP7_75t_L g466 ( 
.A(n_423),
.B(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_428),
.A2(n_465),
.B(n_468),
.Y(n_427)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_428),
.Y(n_663)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_433),
.C(n_464),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_429),
.A2(n_430),
.B1(n_470),
.B2(n_471),
.Y(n_469)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_434),
.B(n_464),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_445),
.C(n_454),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_436),
.B(n_455),
.Y(n_474)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_438),
.Y(n_479)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g473 ( 
.A(n_445),
.B(n_474),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_448),
.A2(n_452),
.B(n_453),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx2_ASAP7_75t_SL g449 ( 
.A(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_452),
.B(n_528),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_452),
.B(n_602),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_452),
.B(n_629),
.Y(n_628)
);

OAI21xp33_ASAP7_75t_SL g644 ( 
.A1(n_452),
.A2(n_628),
.B(n_645),
.Y(n_644)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_465),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_472),
.Y(n_468)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_469),
.B(n_472),
.Y(n_662)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_470),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_475),
.C(n_476),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_473),
.B(n_493),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_475),
.A2(n_476),
.B1(n_477),
.B2(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_475),
.Y(n_494)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_481),
.C(n_488),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_SL g498 ( 
.A(n_478),
.B(n_499),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_481),
.A2(n_488),
.B1(n_489),
.B2(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_481),
.Y(n_500)
);

OA21x2_ASAP7_75t_L g511 ( 
.A1(n_482),
.A2(n_512),
.B(n_513),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_485),
.Y(n_607)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

AOI21x1_ASAP7_75t_L g490 ( 
.A1(n_491),
.A2(n_536),
.B(n_658),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_495),
.Y(n_491)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_492),
.Y(n_659)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_496),
.B(n_659),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_501),
.C(n_510),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_498),
.B(n_539),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_501),
.A2(n_502),
.B1(n_510),
.B2(n_540),
.Y(n_539)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx3_ASAP7_75t_SL g504 ( 
.A(n_505),
.Y(n_504)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx4_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_509),
.B(n_643),
.Y(n_642)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_510),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_519),
.Y(n_510)
);

XNOR2x1_ASAP7_75t_L g561 ( 
.A(n_511),
.B(n_519),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_SL g589 ( 
.A1(n_513),
.A2(n_590),
.B(n_594),
.Y(n_589)
);

NAND2xp33_ASAP7_75t_SL g579 ( 
.A(n_514),
.B(n_580),
.Y(n_579)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_520),
.A2(n_524),
.B1(n_527),
.B2(n_530),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_529),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_532),
.Y(n_530)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

AO21x2_ASAP7_75t_L g536 ( 
.A1(n_537),
.A2(n_562),
.B(n_657),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_538),
.B(n_541),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_538),
.B(n_541),
.Y(n_657)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_542),
.B(n_550),
.C(n_560),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_542),
.B(n_551),
.Y(n_584)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx3_ASAP7_75t_SL g545 ( 
.A(n_546),
.Y(n_545)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_560),
.A2(n_561),
.B1(n_583),
.B2(n_584),
.Y(n_582)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

OAI321xp33_ASAP7_75t_L g562 ( 
.A1(n_563),
.A2(n_585),
.A3(n_649),
.B1(n_655),
.B2(n_656),
.C(n_681),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_564),
.B(n_582),
.Y(n_563)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_564),
.B(n_582),
.Y(n_656)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_565),
.B(n_568),
.C(n_570),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_566),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g653 ( 
.A1(n_566),
.A2(n_568),
.B1(n_569),
.B2(n_654),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_566),
.Y(n_654)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_570),
.Y(n_652)
);

INVxp33_ASAP7_75t_SL g611 ( 
.A(n_571),
.Y(n_611)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_573),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_574),
.Y(n_573)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_574),
.Y(n_593)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_578),
.Y(n_577)
);

INVx5_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

AOI21xp5_ASAP7_75t_L g585 ( 
.A1(n_586),
.A2(n_609),
.B(n_648),
.Y(n_585)
);

OAI21xp5_ASAP7_75t_SL g586 ( 
.A1(n_587),
.A2(n_598),
.B(n_608),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_588),
.B(n_589),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_588),
.B(n_589),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g613 ( 
.A(n_590),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_592),
.Y(n_591)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_595),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_597),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_599),
.B(n_600),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_SL g600 ( 
.A(n_601),
.B(n_606),
.Y(n_600)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_604),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

INVx5_ASAP7_75t_L g606 ( 
.A(n_607),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_610),
.B(n_614),
.Y(n_609)
);

NOR2xp67_ASAP7_75t_L g648 ( 
.A(n_610),
.B(n_614),
.Y(n_648)
);

XNOR2xp5_ASAP7_75t_L g614 ( 
.A(n_615),
.B(n_642),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_615),
.B(n_642),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_616),
.A2(n_627),
.B1(n_632),
.B2(n_637),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_617),
.B(n_622),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_618),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_620),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_621),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_622),
.B(n_638),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g622 ( 
.A(n_623),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_624),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_625),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_626),
.Y(n_625)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_628),
.Y(n_627)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_630),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_631),
.Y(n_630)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_633),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_634),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_635),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_636),
.Y(n_635)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_639),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_640),
.Y(n_639)
);

INVx4_ASAP7_75t_L g640 ( 
.A(n_641),
.Y(n_640)
);

BUFx4f_ASAP7_75t_SL g645 ( 
.A(n_646),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_647),
.Y(n_646)
);

NOR2xp67_ASAP7_75t_L g649 ( 
.A(n_650),
.B(n_651),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_650),
.B(n_651),
.Y(n_655)
);

XNOR2xp5_ASAP7_75t_L g651 ( 
.A(n_652),
.B(n_653),
.Y(n_651)
);

MAJIxp5_ASAP7_75t_L g661 ( 
.A(n_662),
.B(n_663),
.C(n_664),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_L g665 ( 
.A1(n_666),
.A2(n_667),
.B(n_668),
.Y(n_665)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_671),
.Y(n_670)
);

HB1xp67_ASAP7_75t_L g671 ( 
.A(n_672),
.Y(n_671)
);

INVx6_ASAP7_75t_L g678 ( 
.A(n_679),
.Y(n_678)
);


endmodule