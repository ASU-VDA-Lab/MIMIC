module fake_jpeg_6255_n_109 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_109);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_109;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_8;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g13 ( 
.A(n_3),
.B(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_4),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_20),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_24),
.A2(n_22),
.B1(n_18),
.B2(n_16),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_31),
.B1(n_18),
.B2(n_22),
.Y(n_32)
);

AO22x1_ASAP7_75t_SL g31 ( 
.A1(n_24),
.A2(n_15),
.B1(n_12),
.B2(n_8),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_32),
.A2(n_24),
.B1(n_29),
.B2(n_11),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_38),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_37),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_26),
.B(n_19),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_16),
.B1(n_22),
.B2(n_18),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_29),
.B1(n_28),
.B2(n_27),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_26),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_41),
.Y(n_44)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_41),
.B(n_37),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_53),
.C(n_19),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_29),
.B1(n_23),
.B2(n_28),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_46),
.B1(n_25),
.B2(n_21),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_29),
.B1(n_23),
.B2(n_28),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_14),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_17),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_24),
.B1(n_35),
.B2(n_15),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_35),
.B1(n_15),
.B2(n_2),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_26),
.B(n_10),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_62),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_53),
.B(n_20),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_55),
.B(n_57),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_25),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_56),
.A2(n_52),
.B(n_48),
.Y(n_70)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_59),
.B(n_35),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_45),
.B(n_17),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_60),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_49),
.A2(n_9),
.B1(n_11),
.B2(n_21),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_48),
.B(n_15),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_25),
.Y(n_62)
);

OAI21xp33_ASAP7_75t_SL g63 ( 
.A1(n_49),
.A2(n_52),
.B(n_47),
.Y(n_63)
);

AO21x1_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_15),
.B(n_5),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_24),
.B1(n_10),
.B2(n_9),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_64),
.A2(n_65),
.B1(n_66),
.B2(n_46),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_43),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_72),
.C(n_54),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_62),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_75),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_74),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_64),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_78),
.B(n_72),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_61),
.Y(n_81)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_68),
.C(n_70),
.Y(n_86)
);

BUFx12f_ASAP7_75t_SL g89 ( 
.A(n_84),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_58),
.B1(n_65),
.B2(n_0),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_67),
.Y(n_90)
);

AOI321xp33_ASAP7_75t_L g94 ( 
.A1(n_86),
.A2(n_91),
.A3(n_80),
.B1(n_73),
.B2(n_77),
.C(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_76),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_89),
.A2(n_78),
.B(n_83),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_93),
.C(n_94),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_91),
.B(n_79),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_87),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_1),
.C(n_6),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_96),
.A2(n_88),
.B1(n_71),
.B2(n_3),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_100),
.B(n_7),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_SL g101 ( 
.A1(n_98),
.A2(n_2),
.B(n_6),
.C(n_7),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_102),
.A2(n_103),
.B(n_98),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_99),
.B(n_1),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_104),
.C(n_1),
.Y(n_107)
);

BUFx24_ASAP7_75t_SL g108 ( 
.A(n_107),
.Y(n_108)
);

BUFx24_ASAP7_75t_SL g109 ( 
.A(n_108),
.Y(n_109)
);


endmodule