module fake_jpeg_24064_n_233 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_233);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_233;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_32),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_18),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_23),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_29),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_39),
.Y(n_52)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_21),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_50),
.Y(n_73)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_35),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_24),
.B1(n_30),
.B2(n_17),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_49),
.B1(n_33),
.B2(n_34),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_30),
.B1(n_29),
.B2(n_24),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_33),
.B1(n_34),
.B2(n_39),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_29),
.B1(n_20),
.B2(n_23),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_48),
.A2(n_38),
.B1(n_33),
.B2(n_35),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_53),
.A2(n_68),
.B1(n_22),
.B2(n_19),
.Y(n_103)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_55),
.B(n_56),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_32),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_35),
.B1(n_38),
.B2(n_37),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_58),
.A2(n_39),
.B1(n_43),
.B2(n_49),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_31),
.Y(n_59)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_61),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_31),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_15),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_63),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_34),
.C(n_37),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_21),
.B1(n_26),
.B2(n_28),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_69),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_28),
.B1(n_26),
.B2(n_25),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_66),
.A2(n_79),
.B1(n_23),
.B2(n_22),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_25),
.Y(n_67)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_47),
.B(n_20),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_27),
.Y(n_70)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

OAI21xp33_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_34),
.B(n_37),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_71),
.B(n_49),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_47),
.B(n_1),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_76),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_49),
.B1(n_51),
.B2(n_39),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_41),
.B(n_1),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_45),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_81),
.A2(n_97),
.B1(n_100),
.B2(n_103),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_56),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_59),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_101),
.B1(n_76),
.B2(n_72),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_80),
.B(n_93),
.Y(n_116)
);

AO22x1_ASAP7_75t_SL g91 ( 
.A1(n_68),
.A2(n_23),
.B1(n_22),
.B2(n_15),
.Y(n_91)
);

AO22x1_ASAP7_75t_SL g110 ( 
.A1(n_91),
.A2(n_53),
.B1(n_75),
.B2(n_60),
.Y(n_110)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_102),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_63),
.A2(n_62),
.B1(n_58),
.B2(n_61),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_99),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_22),
.B1(n_27),
.B2(n_19),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_65),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

BUFx2_ASAP7_75t_SL g128 ( 
.A(n_104),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_118),
.B1(n_112),
.B2(n_110),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_106),
.A2(n_121),
.B(n_126),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_107),
.Y(n_148)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_108),
.A2(n_110),
.B1(n_111),
.B2(n_114),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_69),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_82),
.B(n_67),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_113),
.Y(n_140)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_116),
.A2(n_119),
.B(n_97),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_87),
.B(n_73),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_118),
.Y(n_147)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_80),
.A2(n_73),
.B(n_54),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_77),
.Y(n_122)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_84),
.B(n_73),
.Y(n_123)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_78),
.Y(n_124)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_84),
.B(n_79),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_125),
.Y(n_134)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_127),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_112),
.A2(n_93),
.B1(n_91),
.B2(n_89),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_129),
.A2(n_130),
.B1(n_141),
.B2(n_142),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_144),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_110),
.A2(n_120),
.B1(n_106),
.B2(n_91),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_136),
.B1(n_143),
.B2(n_151),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_120),
.A2(n_91),
.B1(n_81),
.B2(n_103),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_114),
.A2(n_96),
.B1(n_95),
.B2(n_87),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_111),
.A2(n_96),
.B1(n_83),
.B2(n_92),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_83),
.B1(n_78),
.B2(n_74),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_27),
.B(n_19),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_105),
.C(n_108),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_16),
.C(n_3),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_27),
.B(n_19),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_7),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_126),
.A2(n_74),
.B1(n_57),
.B2(n_19),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_158),
.C(n_162),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_2),
.Y(n_154)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_154),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_127),
.B1(n_115),
.B2(n_57),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_164),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_57),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_157),
.Y(n_186)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_16),
.C(n_14),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_16),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_160),
.B(n_161),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_128),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_16),
.C(n_5),
.Y(n_162)
);

AO22x1_ASAP7_75t_SL g163 ( 
.A1(n_135),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_163),
.A2(n_139),
.B1(n_134),
.B2(n_140),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_152),
.B(n_4),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_166),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_151),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_167),
.B(n_168),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_4),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_132),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_169),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_144),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_8),
.C(n_9),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_139),
.C(n_150),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_175),
.A2(n_185),
.B1(n_159),
.B2(n_129),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_181),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_165),
.Y(n_179)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_179),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_132),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_182),
.A2(n_177),
.B(n_162),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_166),
.A2(n_163),
.B1(n_159),
.B2(n_158),
.Y(n_185)
);

NAND4xp25_ASAP7_75t_SL g187 ( 
.A(n_174),
.B(n_163),
.C(n_137),
.D(n_143),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_193),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_186),
.Y(n_189)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_180),
.A2(n_148),
.B1(n_183),
.B2(n_145),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_190),
.A2(n_133),
.B1(n_182),
.B2(n_153),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_145),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_192),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_181),
.A2(n_141),
.B(n_142),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_176),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_194),
.A2(n_177),
.B1(n_178),
.B2(n_171),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_133),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_196),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_179),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_185),
.A2(n_154),
.B(n_172),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_184),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_189),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_195),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_208),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_202),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_204),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_198),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_8),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_190),
.Y(n_211)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_211),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_212),
.B(n_215),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_214),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_8),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_205),
.Y(n_221)
);

MAJx2_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_200),
.C(n_205),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_216),
.B(n_9),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_207),
.Y(n_217)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_217),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_219),
.B(n_221),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_219),
.A2(n_210),
.B(n_10),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_11),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_223),
.B(n_220),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_225),
.Y(n_230)
);

A2O1A1Ixp33_ASAP7_75t_SL g227 ( 
.A1(n_224),
.A2(n_218),
.B(n_12),
.C(n_13),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_228),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_229),
.A2(n_230),
.B(n_11),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_12),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_12),
.Y(n_233)
);


endmodule