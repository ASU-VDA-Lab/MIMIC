module fake_netlist_1_12498_n_690 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_690);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_690;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_624;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_482;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_466;
wire n_302;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_493;
wire n_418;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_12), .Y(n_89) );
INVxp67_ASAP7_75t_L g90 ( .A(n_69), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_47), .Y(n_91) );
INVx1_ASAP7_75t_SL g92 ( .A(n_48), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_42), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_84), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_2), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_71), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_34), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_0), .Y(n_98) );
HB1xp67_ASAP7_75t_L g99 ( .A(n_2), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_53), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_81), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_63), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_55), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_79), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_68), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_87), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_66), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_1), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_15), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_13), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_10), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_61), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_19), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_83), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_36), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_82), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_58), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_67), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_60), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_56), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_52), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_23), .Y(n_122) );
CKINVDCx16_ASAP7_75t_R g123 ( .A(n_3), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_38), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_4), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_76), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_24), .Y(n_127) );
INVx1_ASAP7_75t_SL g128 ( .A(n_80), .Y(n_128) );
NOR2xp67_ASAP7_75t_L g129 ( .A(n_22), .B(n_31), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_101), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_101), .Y(n_131) );
AND2x2_ASAP7_75t_SL g132 ( .A(n_106), .B(n_21), .Y(n_132) );
BUFx3_ASAP7_75t_L g133 ( .A(n_93), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_96), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_97), .Y(n_135) );
OAI22xp5_ASAP7_75t_L g136 ( .A1(n_108), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g137 ( .A(n_90), .B(n_4), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_105), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_123), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_107), .Y(n_140) );
OAI21x1_ASAP7_75t_L g141 ( .A1(n_114), .A2(n_41), .B(n_86), .Y(n_141) );
BUFx2_ASAP7_75t_L g142 ( .A(n_99), .Y(n_142) );
OA21x2_ASAP7_75t_L g143 ( .A1(n_117), .A2(n_5), .B(n_6), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_118), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_95), .B(n_5), .Y(n_145) );
OA21x2_ASAP7_75t_L g146 ( .A1(n_119), .A2(n_6), .B(n_7), .Y(n_146) );
INVx4_ASAP7_75t_L g147 ( .A(n_91), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_120), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_147), .B(n_91), .Y(n_149) );
OR2x2_ASAP7_75t_L g150 ( .A(n_142), .B(n_89), .Y(n_150) );
OAI22xp33_ASAP7_75t_L g151 ( .A1(n_142), .A2(n_89), .B1(n_111), .B2(n_113), .Y(n_151) );
AOI22xp33_ASAP7_75t_L g152 ( .A1(n_132), .A2(n_110), .B1(n_125), .B2(n_98), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_147), .B(n_94), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_148), .Y(n_154) );
OR2x2_ASAP7_75t_L g155 ( .A(n_142), .B(n_111), .Y(n_155) );
INVx2_ASAP7_75t_SL g156 ( .A(n_147), .Y(n_156) );
BUFx10_ASAP7_75t_L g157 ( .A(n_132), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_148), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_147), .B(n_121), .Y(n_159) );
BUFx3_ASAP7_75t_L g160 ( .A(n_133), .Y(n_160) );
INVx2_ASAP7_75t_SL g161 ( .A(n_147), .Y(n_161) );
AND3x2_ASAP7_75t_L g162 ( .A(n_132), .B(n_122), .C(n_126), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_148), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_148), .Y(n_164) );
BUFx2_ASAP7_75t_L g165 ( .A(n_132), .Y(n_165) );
INVx3_ASAP7_75t_L g166 ( .A(n_148), .Y(n_166) );
BUFx4f_ASAP7_75t_L g167 ( .A(n_143), .Y(n_167) );
OAI22xp33_ASAP7_75t_SL g168 ( .A1(n_136), .A2(n_113), .B1(n_100), .B2(n_102), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_148), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_131), .B(n_94), .Y(n_170) );
NAND2xp33_ASAP7_75t_SL g171 ( .A(n_139), .B(n_103), .Y(n_171) );
AOI22xp33_ASAP7_75t_L g172 ( .A1(n_131), .A2(n_112), .B1(n_100), .B2(n_127), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_134), .B(n_102), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_134), .B(n_104), .Y(n_174) );
NAND2xp33_ASAP7_75t_L g175 ( .A(n_135), .B(n_104), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_148), .Y(n_176) );
NOR2x1_ASAP7_75t_L g177 ( .A(n_150), .B(n_137), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_174), .B(n_135), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_174), .B(n_144), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_170), .B(n_144), .Y(n_180) );
INVx1_ASAP7_75t_SL g181 ( .A(n_150), .Y(n_181) );
INVx1_ASAP7_75t_SL g182 ( .A(n_155), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_154), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_170), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_155), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_165), .A2(n_137), .B1(n_136), .B2(n_139), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_173), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_159), .B(n_133), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_167), .B(n_133), .Y(n_189) );
AO22x1_ASAP7_75t_L g190 ( .A1(n_165), .A2(n_127), .B1(n_124), .B2(n_112), .Y(n_190) );
NAND2x1_ASAP7_75t_L g191 ( .A(n_166), .B(n_143), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_160), .B(n_133), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_160), .B(n_138), .Y(n_193) );
OAI22xp5_ASAP7_75t_SL g194 ( .A1(n_152), .A2(n_109), .B1(n_146), .B2(n_143), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_162), .B(n_145), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_149), .B(n_138), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_154), .Y(n_197) );
NAND2x1_ASAP7_75t_L g198 ( .A(n_166), .B(n_143), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_167), .B(n_148), .Y(n_199) );
INVx5_ASAP7_75t_L g200 ( .A(n_166), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_160), .B(n_138), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_175), .B(n_140), .Y(n_202) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_157), .A2(n_146), .B1(n_143), .B2(n_140), .Y(n_203) );
OR2x2_ASAP7_75t_L g204 ( .A(n_151), .B(n_145), .Y(n_204) );
BUFx2_ASAP7_75t_L g205 ( .A(n_162), .Y(n_205) );
NOR2xp33_ASAP7_75t_SL g206 ( .A(n_157), .B(n_115), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_154), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_153), .B(n_140), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_172), .B(n_130), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_158), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_167), .B(n_130), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g212 ( .A1(n_157), .A2(n_168), .B1(n_167), .B2(n_171), .Y(n_212) );
INVx1_ASAP7_75t_SL g213 ( .A(n_157), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_156), .B(n_130), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_211), .A2(n_156), .B(n_161), .Y(n_215) );
NAND3xp33_ASAP7_75t_L g216 ( .A(n_212), .B(n_161), .C(n_143), .Y(n_216) );
INVxp67_ASAP7_75t_L g217 ( .A(n_181), .Y(n_217) );
OAI21x1_ASAP7_75t_L g218 ( .A1(n_191), .A2(n_141), .B(n_158), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_206), .B(n_115), .Y(n_219) );
AND2x2_ASAP7_75t_L g220 ( .A(n_182), .B(n_146), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_184), .B(n_168), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_185), .A2(n_146), .B(n_92), .C(n_128), .Y(n_222) );
BUFx3_ASAP7_75t_L g223 ( .A(n_205), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_178), .B(n_116), .Y(n_224) );
OAI21xp5_ASAP7_75t_L g225 ( .A1(n_199), .A2(n_141), .B(n_176), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_204), .B(n_116), .Y(n_226) );
NOR2xp33_ASAP7_75t_SL g227 ( .A(n_205), .B(n_124), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_193), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g229 ( .A1(n_204), .A2(n_213), .B1(n_180), .B2(n_187), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_211), .A2(n_141), .B(n_176), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_179), .B(n_146), .Y(n_231) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_209), .A2(n_146), .B(n_169), .C(n_166), .Y(n_232) );
AND2x2_ASAP7_75t_SL g233 ( .A(n_195), .B(n_169), .Y(n_233) );
OAI22xp5_ASAP7_75t_L g234 ( .A1(n_186), .A2(n_129), .B1(n_163), .B2(n_158), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g235 ( .A1(n_195), .A2(n_164), .B1(n_163), .B2(n_9), .Y(n_235) );
INVx2_ASAP7_75t_SL g236 ( .A(n_190), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_SL g237 ( .A1(n_199), .A2(n_164), .B(n_163), .C(n_44), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_201), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_177), .B(n_7), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_195), .B(n_164), .Y(n_240) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_194), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_196), .B(n_8), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_202), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_189), .A2(n_45), .B(n_85), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_214), .B(n_11), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_208), .Y(n_246) );
CKINVDCx5p33_ASAP7_75t_R g247 ( .A(n_217), .Y(n_247) );
INVx3_ASAP7_75t_L g248 ( .A(n_223), .Y(n_248) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_233), .A2(n_203), .B1(n_188), .B2(n_189), .Y(n_249) );
NAND3xp33_ASAP7_75t_L g250 ( .A(n_234), .B(n_191), .C(n_198), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_246), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_221), .B(n_198), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_246), .Y(n_253) );
OAI21xp5_ASAP7_75t_L g254 ( .A1(n_216), .A2(n_192), .B(n_207), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_232), .A2(n_231), .B(n_230), .Y(n_255) );
AO31x2_ASAP7_75t_L g256 ( .A1(n_241), .A2(n_210), .A3(n_207), .B(n_197), .Y(n_256) );
AO21x1_ASAP7_75t_L g257 ( .A1(n_222), .A2(n_210), .B(n_197), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_239), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_228), .Y(n_259) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_228), .A2(n_183), .B(n_200), .Y(n_260) );
AO32x2_ASAP7_75t_L g261 ( .A1(n_235), .A2(n_11), .A3(n_12), .B1(n_13), .B2(n_14), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_L g262 ( .A1(n_229), .A2(n_183), .B(n_15), .C(n_16), .Y(n_262) );
AO31x2_ASAP7_75t_L g263 ( .A1(n_244), .A2(n_14), .A3(n_16), .B(n_17), .Y(n_263) );
AO31x2_ASAP7_75t_L g264 ( .A1(n_242), .A2(n_17), .A3(n_18), .B(n_19), .Y(n_264) );
AO21x1_ASAP7_75t_L g265 ( .A1(n_225), .A2(n_54), .B(n_88), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_215), .A2(n_200), .B(n_51), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_226), .B(n_200), .Y(n_267) );
INVx3_ASAP7_75t_L g268 ( .A(n_223), .Y(n_268) );
AO31x2_ASAP7_75t_L g269 ( .A1(n_245), .A2(n_18), .A3(n_20), .B(n_25), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_251), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_253), .B(n_238), .Y(n_271) );
AO21x2_ASAP7_75t_L g272 ( .A1(n_255), .A2(n_218), .B(n_237), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_259), .Y(n_273) );
OAI22xp33_ASAP7_75t_L g274 ( .A1(n_258), .A2(n_236), .B1(n_227), .B2(n_243), .Y(n_274) );
AO21x2_ASAP7_75t_L g275 ( .A1(n_255), .A2(n_218), .B(n_240), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_260), .B(n_233), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_247), .B(n_236), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_248), .B(n_233), .Y(n_278) );
OAI21xp5_ASAP7_75t_L g279 ( .A1(n_252), .A2(n_220), .B(n_238), .Y(n_279) );
OR2x2_ASAP7_75t_L g280 ( .A(n_252), .B(n_220), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_263), .Y(n_281) );
OAI21xp5_ASAP7_75t_L g282 ( .A1(n_249), .A2(n_224), .B(n_243), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_263), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_263), .Y(n_284) );
NOR2xp33_ASAP7_75t_SL g285 ( .A(n_262), .B(n_219), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_263), .Y(n_286) );
INVx2_ASAP7_75t_SL g287 ( .A(n_248), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_264), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_264), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_269), .Y(n_290) );
OA21x2_ASAP7_75t_L g291 ( .A1(n_257), .A2(n_57), .B(n_26), .Y(n_291) );
BUFx3_ASAP7_75t_L g292 ( .A(n_278), .Y(n_292) );
AOI21x1_ASAP7_75t_L g293 ( .A1(n_290), .A2(n_289), .B(n_288), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_280), .B(n_268), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_275), .Y(n_295) );
AO21x2_ASAP7_75t_L g296 ( .A1(n_288), .A2(n_254), .B(n_265), .Y(n_296) );
AND2x4_ASAP7_75t_L g297 ( .A(n_280), .B(n_250), .Y(n_297) );
INVxp67_ASAP7_75t_L g298 ( .A(n_273), .Y(n_298) );
AOI21xp33_ASAP7_75t_L g299 ( .A1(n_274), .A2(n_262), .B(n_249), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_275), .Y(n_300) );
OAI21x1_ASAP7_75t_L g301 ( .A1(n_286), .A2(n_266), .B(n_268), .Y(n_301) );
AO21x2_ASAP7_75t_L g302 ( .A1(n_289), .A2(n_266), .B(n_267), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_276), .B(n_261), .Y(n_303) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_291), .Y(n_304) );
AND2x4_ASAP7_75t_L g305 ( .A(n_280), .B(n_256), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_276), .B(n_261), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_286), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_275), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_276), .B(n_261), .Y(n_309) );
NOR2x1_ASAP7_75t_SL g310 ( .A(n_278), .B(n_261), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_270), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_270), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_273), .Y(n_313) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_290), .Y(n_314) );
OA21x2_ASAP7_75t_L g315 ( .A1(n_290), .A2(n_269), .B(n_256), .Y(n_315) );
NAND4xp25_ASAP7_75t_L g316 ( .A(n_277), .B(n_20), .C(n_264), .D(n_269), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_281), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_275), .Y(n_318) );
INVx3_ASAP7_75t_L g319 ( .A(n_278), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_275), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_303), .B(n_284), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_303), .B(n_284), .Y(n_322) );
OR2x2_ASAP7_75t_L g323 ( .A(n_313), .B(n_283), .Y(n_323) );
INVx3_ASAP7_75t_L g324 ( .A(n_307), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_313), .Y(n_325) );
BUFx2_ASAP7_75t_L g326 ( .A(n_314), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_303), .B(n_281), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_317), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_307), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_307), .Y(n_330) );
BUFx3_ASAP7_75t_L g331 ( .A(n_314), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_306), .B(n_283), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_307), .B(n_286), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_317), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_306), .B(n_309), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_293), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_293), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_306), .B(n_279), .Y(n_338) );
INVxp67_ASAP7_75t_SL g339 ( .A(n_298), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_293), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_309), .B(n_279), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_311), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_295), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_311), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_312), .Y(n_345) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_304), .Y(n_346) );
INVx4_ASAP7_75t_R g347 ( .A(n_292), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_309), .B(n_291), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_312), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_295), .Y(n_350) );
BUFx2_ASAP7_75t_L g351 ( .A(n_298), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_305), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_305), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_295), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_305), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_319), .B(n_282), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_305), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_292), .B(n_271), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_305), .B(n_291), .Y(n_359) );
AND2x2_ASAP7_75t_SL g360 ( .A(n_297), .B(n_291), .Y(n_360) );
BUFx3_ASAP7_75t_L g361 ( .A(n_294), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_300), .B(n_291), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_300), .Y(n_363) );
AND2x4_ASAP7_75t_L g364 ( .A(n_300), .B(n_272), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_308), .Y(n_365) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_294), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_308), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_292), .B(n_271), .Y(n_368) );
AND2x4_ASAP7_75t_L g369 ( .A(n_320), .B(n_272), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_335), .B(n_297), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_335), .B(n_297), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_335), .B(n_297), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_329), .Y(n_373) );
NOR2xp67_ASAP7_75t_L g374 ( .A(n_325), .B(n_316), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_321), .B(n_297), .Y(n_375) );
AND2x4_ASAP7_75t_L g376 ( .A(n_352), .B(n_320), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_321), .B(n_319), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_328), .Y(n_378) );
AND2x4_ASAP7_75t_L g379 ( .A(n_352), .B(n_320), .Y(n_379) );
INVx3_ASAP7_75t_L g380 ( .A(n_324), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_321), .B(n_319), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_358), .B(n_277), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_322), .B(n_319), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_366), .B(n_319), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_328), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_322), .B(n_318), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_322), .B(n_318), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_334), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_342), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_342), .B(n_292), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_344), .B(n_294), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_344), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_327), .B(n_318), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_329), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_327), .B(n_308), .Y(n_395) );
BUFx2_ASAP7_75t_SL g396 ( .A(n_331), .Y(n_396) );
INVx3_ASAP7_75t_L g397 ( .A(n_324), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_329), .Y(n_398) );
INVx4_ASAP7_75t_L g399 ( .A(n_331), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_345), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_327), .B(n_332), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_345), .B(n_310), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_349), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_349), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_330), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_337), .Y(n_406) );
INVx4_ASAP7_75t_L g407 ( .A(n_331), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_337), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_332), .B(n_315), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_340), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_332), .B(n_315), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_325), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_368), .B(n_316), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_338), .B(n_315), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_340), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_343), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_343), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_330), .Y(n_418) );
BUFx2_ASAP7_75t_SL g419 ( .A(n_330), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_338), .B(n_315), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_343), .Y(n_421) );
INVxp67_ASAP7_75t_L g422 ( .A(n_351), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_338), .B(n_315), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_350), .Y(n_424) );
AND2x4_ASAP7_75t_L g425 ( .A(n_355), .B(n_301), .Y(n_425) );
INVx3_ASAP7_75t_L g426 ( .A(n_324), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_368), .B(n_274), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_350), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_341), .B(n_299), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_350), .Y(n_430) );
INVx2_ASAP7_75t_SL g431 ( .A(n_347), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_341), .B(n_315), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_355), .B(n_296), .Y(n_433) );
NOR2x1_ASAP7_75t_SL g434 ( .A(n_347), .B(n_287), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_351), .B(n_282), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_357), .B(n_296), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_357), .B(n_296), .Y(n_437) );
AND2x4_ASAP7_75t_L g438 ( .A(n_353), .B(n_301), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g439 ( .A(n_326), .B(n_285), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_406), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_406), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_408), .Y(n_442) );
BUFx3_ASAP7_75t_L g443 ( .A(n_399), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_401), .B(n_353), .Y(n_444) );
INVxp67_ASAP7_75t_L g445 ( .A(n_412), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_378), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_401), .B(n_359), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_370), .B(n_339), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_370), .B(n_339), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_371), .B(n_361), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_371), .B(n_326), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_409), .B(n_323), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_378), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_372), .B(n_361), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_385), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_372), .B(n_361), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_385), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_382), .A2(n_356), .B1(n_360), .B2(n_359), .Y(n_458) );
NAND4xp25_ASAP7_75t_SL g459 ( .A(n_413), .B(n_359), .C(n_356), .D(n_323), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_414), .B(n_348), .Y(n_460) );
NAND2xp67_ASAP7_75t_L g461 ( .A(n_402), .B(n_348), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_414), .B(n_348), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_420), .B(n_423), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_388), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_388), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_389), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_377), .B(n_324), .Y(n_467) );
NAND2x1p5_ASAP7_75t_L g468 ( .A(n_431), .B(n_333), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_377), .B(n_333), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_374), .A2(n_360), .B1(n_287), .B2(n_333), .Y(n_470) );
BUFx3_ASAP7_75t_L g471 ( .A(n_399), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_409), .B(n_333), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_381), .B(n_333), .Y(n_473) );
INVx2_ASAP7_75t_SL g474 ( .A(n_399), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_411), .B(n_367), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_422), .B(n_287), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_408), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_435), .B(n_360), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_389), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_411), .B(n_367), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_386), .B(n_363), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_392), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_392), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_400), .Y(n_484) );
AND2x2_ASAP7_75t_SL g485 ( .A(n_407), .B(n_336), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_420), .B(n_365), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_423), .B(n_365), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_432), .B(n_365), .Y(n_488) );
INVxp67_ASAP7_75t_SL g489 ( .A(n_373), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_432), .B(n_354), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_400), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_403), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_429), .B(n_354), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_386), .B(n_363), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_387), .B(n_363), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_403), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_427), .B(n_285), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_410), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_383), .B(n_369), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_383), .B(n_364), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_404), .Y(n_501) );
BUFx2_ASAP7_75t_L g502 ( .A(n_431), .Y(n_502) );
NAND2x1p5_ASAP7_75t_L g503 ( .A(n_407), .B(n_336), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_404), .Y(n_504) );
INVx1_ASAP7_75t_SL g505 ( .A(n_396), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_410), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_387), .B(n_364), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_415), .Y(n_508) );
INVxp67_ASAP7_75t_L g509 ( .A(n_396), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_415), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_416), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_375), .B(n_369), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_375), .B(n_369), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_416), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_393), .B(n_369), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_393), .B(n_364), .Y(n_516) );
NAND2x1p5_ASAP7_75t_L g517 ( .A(n_407), .B(n_336), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_390), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_395), .B(n_369), .Y(n_519) );
INVxp67_ASAP7_75t_L g520 ( .A(n_419), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_395), .B(n_364), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_384), .B(n_364), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_433), .B(n_362), .Y(n_523) );
NAND2x1_ASAP7_75t_L g524 ( .A(n_474), .B(n_438), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_446), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_453), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_485), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_452), .B(n_463), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_455), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_518), .B(n_433), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_475), .B(n_417), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_457), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_485), .A2(n_434), .B(n_439), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_445), .B(n_391), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_445), .B(n_436), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_480), .B(n_417), .Y(n_536) );
NAND2x1p5_ASAP7_75t_L g537 ( .A(n_443), .B(n_434), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_447), .B(n_419), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_443), .Y(n_539) );
INVxp33_ASAP7_75t_L g540 ( .A(n_468), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_464), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_460), .B(n_436), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_460), .B(n_437), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_471), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_471), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_497), .A2(n_437), .B1(n_376), .B2(n_379), .Y(n_546) );
AND3x2_ASAP7_75t_L g547 ( .A(n_502), .B(n_438), .C(n_430), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_465), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_466), .Y(n_549) );
NOR2x1_ASAP7_75t_L g550 ( .A(n_505), .B(n_380), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_479), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_486), .B(n_421), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_448), .B(n_380), .Y(n_553) );
OAI21xp5_ASAP7_75t_L g554 ( .A1(n_509), .A2(n_438), .B(n_430), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_474), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_482), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_497), .A2(n_376), .B1(n_379), .B2(n_438), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_487), .B(n_428), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_483), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_484), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_491), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_462), .B(n_376), .Y(n_562) );
NOR2x1_ASAP7_75t_L g563 ( .A(n_470), .B(n_380), .Y(n_563) );
INVxp67_ASAP7_75t_L g564 ( .A(n_493), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_503), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_492), .Y(n_566) );
AND2x4_ASAP7_75t_L g567 ( .A(n_509), .B(n_425), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_496), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_462), .B(n_376), .Y(n_569) );
INVx2_ASAP7_75t_SL g570 ( .A(n_468), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_501), .Y(n_571) );
AND2x4_ASAP7_75t_L g572 ( .A(n_444), .B(n_425), .Y(n_572) );
INVx2_ASAP7_75t_SL g573 ( .A(n_444), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_447), .B(n_426), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_488), .B(n_428), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_504), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_523), .B(n_379), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_490), .B(n_424), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_469), .B(n_426), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_523), .B(n_421), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_473), .B(n_426), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_472), .B(n_424), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_481), .B(n_418), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_506), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_510), .Y(n_585) );
INVx2_ASAP7_75t_SL g586 ( .A(n_450), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_449), .B(n_397), .Y(n_587) );
NAND4xp25_ASAP7_75t_SL g588 ( .A(n_458), .B(n_362), .C(n_418), .D(n_405), .Y(n_588) );
AOI21xp33_ASAP7_75t_L g589 ( .A1(n_476), .A2(n_425), .B(n_302), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_512), .B(n_397), .Y(n_590) );
AND2x4_ASAP7_75t_L g591 ( .A(n_520), .B(n_397), .Y(n_591) );
O2A1O1Ixp33_ASAP7_75t_L g592 ( .A1(n_520), .A2(n_405), .B(n_398), .C(n_394), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_522), .B(n_394), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_440), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_451), .B(n_398), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_564), .B(n_461), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_588), .A2(n_459), .B1(n_478), .B2(n_476), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_582), .Y(n_598) );
OAI321xp33_ASAP7_75t_L g599 ( .A1(n_554), .A2(n_478), .A3(n_503), .B1(n_517), .B2(n_500), .C(n_507), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_525), .Y(n_600) );
INVx1_ASAP7_75t_SL g601 ( .A(n_528), .Y(n_601) );
OAI21xp5_ASAP7_75t_L g602 ( .A1(n_533), .A2(n_517), .B(n_489), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_526), .Y(n_603) );
A2O1A1Ixp33_ASAP7_75t_L g604 ( .A1(n_524), .A2(n_456), .B(n_454), .C(n_513), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_529), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_534), .B(n_516), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_532), .Y(n_607) );
NAND2xp33_ASAP7_75t_SL g608 ( .A(n_540), .B(n_519), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_572), .B(n_499), .Y(n_609) );
NOR2xp67_ASAP7_75t_L g610 ( .A(n_554), .B(n_521), .Y(n_610) );
INVxp67_ASAP7_75t_L g611 ( .A(n_555), .Y(n_611) );
OAI222xp33_ASAP7_75t_L g612 ( .A1(n_563), .A2(n_494), .B1(n_495), .B2(n_467), .C1(n_515), .C2(n_489), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_586), .B(n_495), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_535), .B(n_494), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_546), .A2(n_477), .B1(n_441), .B2(n_508), .Y(n_615) );
NOR2xp33_ASAP7_75t_R g616 ( .A(n_570), .B(n_27), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_546), .A2(n_477), .B1(n_441), .B2(n_508), .Y(n_617) );
NOR2x1_ASAP7_75t_L g618 ( .A(n_550), .B(n_514), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_539), .Y(n_619) );
INVxp33_ASAP7_75t_L g620 ( .A(n_537), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_530), .B(n_440), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_557), .A2(n_514), .B1(n_511), .B2(n_498), .Y(n_622) );
A2O1A1Ixp33_ASAP7_75t_L g623 ( .A1(n_563), .A2(n_442), .B(n_511), .C(n_373), .Y(n_623) );
INVxp67_ASAP7_75t_SL g624 ( .A(n_592), .Y(n_624) );
INVxp67_ASAP7_75t_L g625 ( .A(n_544), .Y(n_625) );
OR2x2_ASAP7_75t_L g626 ( .A(n_542), .B(n_543), .Y(n_626) );
OAI31xp33_ASAP7_75t_L g627 ( .A1(n_589), .A2(n_362), .A3(n_256), .B(n_302), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_574), .B(n_346), .Y(n_628) );
CKINVDCx5p33_ASAP7_75t_R g629 ( .A(n_545), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_531), .Y(n_630) );
NAND4xp25_ASAP7_75t_SL g631 ( .A(n_550), .B(n_304), .C(n_302), .D(n_346), .Y(n_631) );
NAND4xp25_ASAP7_75t_L g632 ( .A(n_589), .B(n_28), .C(n_29), .D(n_30), .Y(n_632) );
A2O1A1Ixp33_ASAP7_75t_SL g633 ( .A1(n_565), .A2(n_302), .B(n_33), .C(n_35), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_541), .Y(n_634) );
NOR3xp33_ASAP7_75t_L g635 ( .A(n_527), .B(n_301), .C(n_302), .Y(n_635) );
INVxp67_ASAP7_75t_L g636 ( .A(n_553), .Y(n_636) );
NOR3xp33_ASAP7_75t_L g637 ( .A(n_624), .B(n_571), .C(n_548), .Y(n_637) );
OAI211xp5_ASAP7_75t_L g638 ( .A1(n_616), .A2(n_538), .B(n_587), .C(n_573), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_600), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_598), .B(n_595), .Y(n_640) );
OAI221xp5_ASAP7_75t_L g641 ( .A1(n_608), .A2(n_549), .B1(n_551), .B2(n_556), .C(n_559), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_597), .A2(n_567), .B1(n_591), .B2(n_581), .Y(n_642) );
OAI211xp5_ASAP7_75t_L g643 ( .A1(n_602), .A2(n_569), .B(n_562), .C(n_580), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_604), .A2(n_620), .B1(n_601), .B2(n_610), .Y(n_644) );
OAI221xp5_ASAP7_75t_L g645 ( .A1(n_596), .A2(n_617), .B1(n_615), .B2(n_627), .C(n_623), .Y(n_645) );
AOI221xp5_ASAP7_75t_SL g646 ( .A1(n_612), .A2(n_577), .B1(n_579), .B2(n_590), .C(n_560), .Y(n_646) );
AOI222xp33_ASAP7_75t_L g647 ( .A1(n_612), .A2(n_567), .B1(n_561), .B2(n_566), .C1(n_585), .C2(n_584), .Y(n_647) );
OAI32xp33_ASAP7_75t_L g648 ( .A1(n_611), .A2(n_558), .A3(n_575), .B1(n_536), .B2(n_552), .Y(n_648) );
A2O1A1Ixp33_ASAP7_75t_L g649 ( .A1(n_599), .A2(n_591), .B(n_578), .C(n_583), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_603), .Y(n_650) );
OAI32xp33_ASAP7_75t_L g651 ( .A1(n_611), .A2(n_593), .A3(n_547), .B1(n_576), .B2(n_568), .Y(n_651) );
NOR2xp67_ASAP7_75t_L g652 ( .A(n_631), .B(n_594), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_626), .B(n_630), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_605), .Y(n_654) );
OR2x2_ASAP7_75t_L g655 ( .A(n_621), .B(n_296), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_629), .A2(n_304), .B1(n_346), .B2(n_296), .Y(n_656) );
AOI221xp5_ASAP7_75t_L g657 ( .A1(n_622), .A2(n_606), .B1(n_636), .B2(n_634), .C(n_607), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_618), .A2(n_32), .B(n_37), .Y(n_658) );
NAND5xp2_ASAP7_75t_L g659 ( .A(n_635), .B(n_39), .C(n_40), .D(n_43), .E(n_46), .Y(n_659) );
O2A1O1Ixp33_ASAP7_75t_L g660 ( .A1(n_619), .A2(n_49), .B(n_50), .C(n_59), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_614), .Y(n_661) );
OAI22xp33_ASAP7_75t_L g662 ( .A1(n_632), .A2(n_62), .B1(n_64), .B2(n_65), .Y(n_662) );
OAI211xp5_ASAP7_75t_SL g663 ( .A1(n_625), .A2(n_70), .B(n_72), .C(n_73), .Y(n_663) );
OAI221xp5_ASAP7_75t_L g664 ( .A1(n_613), .A2(n_74), .B1(n_75), .B2(n_77), .C(n_78), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_609), .A2(n_200), .B1(n_628), .B2(n_633), .Y(n_665) );
NOR3xp33_ASAP7_75t_SL g666 ( .A(n_599), .B(n_200), .C(n_612), .Y(n_666) );
AOI222xp33_ASAP7_75t_L g667 ( .A1(n_624), .A2(n_612), .B1(n_608), .B2(n_601), .C1(n_610), .C2(n_622), .Y(n_667) );
NOR3xp33_ASAP7_75t_SL g668 ( .A(n_638), .B(n_644), .C(n_649), .Y(n_668) );
O2A1O1Ixp33_ASAP7_75t_SL g669 ( .A1(n_638), .A2(n_648), .B(n_651), .C(n_657), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_654), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_637), .B(n_642), .Y(n_671) );
NOR2x1_ASAP7_75t_L g672 ( .A(n_662), .B(n_659), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_646), .B(n_661), .Y(n_673) );
NOR2x1_ASAP7_75t_L g674 ( .A(n_663), .B(n_658), .Y(n_674) );
NOR3xp33_ASAP7_75t_L g675 ( .A(n_669), .B(n_664), .C(n_645), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_671), .B(n_643), .Y(n_676) );
NOR2xp67_ASAP7_75t_L g677 ( .A(n_673), .B(n_643), .Y(n_677) );
NOR4xp25_ASAP7_75t_L g678 ( .A(n_670), .B(n_641), .C(n_660), .D(n_639), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_676), .B(n_650), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_677), .Y(n_680) );
NOR3xp33_ASAP7_75t_L g681 ( .A(n_675), .B(n_672), .C(n_674), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_680), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_681), .B(n_678), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_682), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_683), .Y(n_685) );
AO22x2_ASAP7_75t_L g686 ( .A1(n_684), .A2(n_679), .B1(n_668), .B2(n_665), .Y(n_686) );
O2A1O1Ixp33_ASAP7_75t_L g687 ( .A1(n_686), .A2(n_685), .B(n_667), .C(n_666), .Y(n_687) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_687), .A2(n_653), .B(n_647), .Y(n_688) );
AND2x4_ASAP7_75t_L g689 ( .A(n_688), .B(n_640), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_689), .A2(n_652), .B1(n_655), .B2(n_656), .Y(n_690) );
endmodule