module fake_netlist_1_3338_n_611 (n_117, n_44, n_133, n_149, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_125, n_9, n_161, n_10, n_130, n_103, n_19, n_87, n_137, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_165, n_146, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_169, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_46, n_31, n_58, n_122, n_138, n_126, n_118, n_32, n_0, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_166, n_162, n_75, n_163, n_105, n_159, n_72, n_136, n_43, n_76, n_89, n_68, n_144, n_27, n_53, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_15, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_611);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_125;
input n_9;
input n_161;
input n_10;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_165;
input n_146;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_169;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_46;
input n_31;
input n_58;
input n_122;
input n_138;
input n_126;
input n_118;
input n_32;
input n_0;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_166;
input n_162;
input n_75;
input n_163;
input n_105;
input n_159;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_68;
input n_144;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_15;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_611;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_431;
wire n_484;
wire n_496;
wire n_177;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_202;
wire n_386;
wire n_432;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_205;
wire n_330;
wire n_587;
wire n_387;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_517;
wire n_560;
wire n_479;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_527;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_178;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_295;
wire n_263;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_524;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_602;
wire n_198;
wire n_424;
wire n_569;
wire n_297;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_187;
wire n_375;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_421;
wire n_175;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx14_ASAP7_75t_R g173 ( .A(n_54), .Y(n_173) );
INVxp67_ASAP7_75t_L g174 ( .A(n_149), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_17), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_3), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_150), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_16), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_0), .Y(n_179) );
BUFx2_ASAP7_75t_L g180 ( .A(n_58), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_66), .Y(n_181) );
CKINVDCx5p33_ASAP7_75t_R g182 ( .A(n_95), .Y(n_182) );
INVxp33_ASAP7_75t_L g183 ( .A(n_70), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_33), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_72), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_43), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_77), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_153), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_126), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_140), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_42), .Y(n_191) );
INVxp67_ASAP7_75t_SL g192 ( .A(n_73), .Y(n_192) );
INVx1_ASAP7_75t_SL g193 ( .A(n_19), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_122), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_97), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_152), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_64), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_71), .Y(n_198) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_151), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_146), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_82), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_59), .Y(n_202) );
CKINVDCx14_ASAP7_75t_R g203 ( .A(n_55), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_163), .Y(n_204) );
BUFx3_ASAP7_75t_L g205 ( .A(n_129), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_41), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_84), .Y(n_207) );
BUFx2_ASAP7_75t_SL g208 ( .A(n_37), .Y(n_208) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_134), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_90), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_108), .Y(n_211) );
BUFx3_ASAP7_75t_L g212 ( .A(n_68), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_137), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_15), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_158), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_13), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_148), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_161), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_39), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_133), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_124), .Y(n_221) );
INVx3_ASAP7_75t_L g222 ( .A(n_24), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_142), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_50), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_48), .Y(n_225) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_160), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_154), .Y(n_227) );
INVxp67_ASAP7_75t_SL g228 ( .A(n_26), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g229 ( .A(n_162), .Y(n_229) );
CKINVDCx16_ASAP7_75t_R g230 ( .A(n_38), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_143), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_93), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_128), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_159), .Y(n_234) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_114), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_164), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_141), .Y(n_237) );
INVxp67_ASAP7_75t_SL g238 ( .A(n_76), .Y(n_238) );
BUFx2_ASAP7_75t_L g239 ( .A(n_166), .Y(n_239) );
BUFx10_ASAP7_75t_L g240 ( .A(n_51), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_29), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_5), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_35), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g244 ( .A(n_9), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_79), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_136), .Y(n_246) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_125), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_75), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_135), .Y(n_249) );
INVxp33_ASAP7_75t_L g250 ( .A(n_144), .Y(n_250) );
HB1xp67_ASAP7_75t_L g251 ( .A(n_52), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_49), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_12), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_102), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_53), .Y(n_255) );
CKINVDCx20_ASAP7_75t_R g256 ( .A(n_40), .Y(n_256) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_98), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_156), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_32), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_118), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_104), .Y(n_261) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_155), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_147), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_78), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_139), .Y(n_265) );
CKINVDCx16_ASAP7_75t_R g266 ( .A(n_157), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_138), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_61), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_5), .Y(n_269) );
INVxp67_ASAP7_75t_SL g270 ( .A(n_88), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_28), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_165), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_145), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_47), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_119), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_209), .B(n_0), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_229), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_222), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_209), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_247), .Y(n_280) );
INVx4_ASAP7_75t_L g281 ( .A(n_222), .Y(n_281) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_210), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_251), .Y(n_283) );
BUFx2_ASAP7_75t_L g284 ( .A(n_242), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_180), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_239), .Y(n_286) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_210), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_179), .B(n_1), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_202), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_216), .B(n_1), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_253), .Y(n_291) );
OA21x2_ASAP7_75t_L g292 ( .A1(n_175), .A2(n_111), .B(n_171), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_269), .B(n_207), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_256), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_240), .Y(n_295) );
NAND3xp33_ASAP7_75t_L g296 ( .A(n_288), .B(n_275), .C(n_178), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_278), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_277), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_278), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_295), .B(n_279), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_285), .B(n_183), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_281), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_281), .Y(n_303) );
NAND2x1p5_ASAP7_75t_L g304 ( .A(n_290), .B(n_193), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_290), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_280), .B(n_192), .Y(n_306) );
INVx3_ASAP7_75t_L g307 ( .A(n_293), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_276), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_308), .B(n_283), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_304), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_302), .Y(n_311) );
AND2x6_ASAP7_75t_SL g312 ( .A(n_301), .B(n_276), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_303), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_297), .Y(n_314) );
BUFx12f_ASAP7_75t_L g315 ( .A(n_298), .Y(n_315) );
BUFx6f_ASAP7_75t_L g316 ( .A(n_299), .Y(n_316) );
NAND2x1p5_ASAP7_75t_L g317 ( .A(n_306), .B(n_293), .Y(n_317) );
NOR2xp33_ASAP7_75t_R g318 ( .A(n_307), .B(n_294), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_306), .B(n_286), .Y(n_319) );
AOI222xp33_ASAP7_75t_L g320 ( .A1(n_309), .A2(n_301), .B1(n_307), .B2(n_291), .C1(n_300), .C2(n_284), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_309), .B(n_305), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_312), .B(n_304), .Y(n_322) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_317), .A2(n_296), .B1(n_266), .B2(n_230), .Y(n_323) );
BUFx2_ASAP7_75t_L g324 ( .A(n_318), .Y(n_324) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_311), .A2(n_292), .B(n_296), .Y(n_325) );
A2O1A1Ixp33_ASAP7_75t_L g326 ( .A1(n_319), .A2(n_288), .B(n_228), .C(n_238), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_317), .B(n_289), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_316), .Y(n_328) );
OAI21xp33_ASAP7_75t_SL g329 ( .A1(n_319), .A2(n_228), .B(n_192), .Y(n_329) );
INVx5_ASAP7_75t_L g330 ( .A(n_316), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_313), .A2(n_292), .B(n_270), .Y(n_331) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_324), .Y(n_332) );
OAI21x1_ASAP7_75t_L g333 ( .A1(n_331), .A2(n_292), .B(n_314), .Y(n_333) );
OAI21x1_ASAP7_75t_L g334 ( .A1(n_325), .A2(n_181), .B(n_177), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_330), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_321), .B(n_310), .Y(n_336) );
AND2x4_ASAP7_75t_SL g337 ( .A(n_322), .B(n_244), .Y(n_337) );
OAI21x1_ASAP7_75t_L g338 ( .A1(n_328), .A2(n_185), .B(n_184), .Y(n_338) );
OAI22xp33_ASAP7_75t_L g339 ( .A1(n_323), .A2(n_315), .B1(n_250), .B2(n_316), .Y(n_339) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_330), .A2(n_238), .B1(n_270), .B2(n_174), .Y(n_340) );
OAI21xp5_ASAP7_75t_L g341 ( .A1(n_329), .A2(n_174), .B(n_190), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_320), .B(n_240), .Y(n_342) );
OA21x2_ASAP7_75t_L g343 ( .A1(n_326), .A2(n_195), .B(n_191), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_330), .A2(n_173), .B1(n_203), .B2(n_206), .Y(n_344) );
O2A1O1Ixp33_ASAP7_75t_L g345 ( .A1(n_327), .A2(n_259), .B(n_225), .C(n_196), .Y(n_345) );
OAI21x1_ASAP7_75t_L g346 ( .A1(n_331), .A2(n_198), .B(n_197), .Y(n_346) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_325), .A2(n_201), .B(n_200), .Y(n_347) );
A2O1A1Ixp33_ASAP7_75t_L g348 ( .A1(n_329), .A2(n_233), .B(n_204), .C(n_221), .Y(n_348) );
OAI21x1_ASAP7_75t_L g349 ( .A1(n_331), .A2(n_214), .B(n_213), .Y(n_349) );
OAI21xp33_ASAP7_75t_L g350 ( .A1(n_342), .A2(n_212), .B(n_205), .Y(n_350) );
BUFx12f_ASAP7_75t_L g351 ( .A(n_332), .Y(n_351) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_337), .A2(n_236), .B1(n_218), .B2(n_219), .Y(n_352) );
AOI22xp33_ASAP7_75t_SL g353 ( .A1(n_344), .A2(n_208), .B1(n_176), .B2(n_193), .Y(n_353) );
OAI211xp5_ASAP7_75t_L g354 ( .A1(n_341), .A2(n_176), .B(n_227), .C(n_255), .Y(n_354) );
AOI22xp5_ASAP7_75t_L g355 ( .A1(n_336), .A2(n_252), .B1(n_220), .B2(n_223), .Y(n_355) );
NAND2xp5_ASAP7_75t_SL g356 ( .A(n_339), .B(n_182), .Y(n_356) );
OA21x2_ASAP7_75t_L g357 ( .A1(n_334), .A2(n_232), .B(n_224), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_341), .A2(n_176), .B1(n_246), .B2(n_245), .Y(n_358) );
AOI21xp5_ASAP7_75t_L g359 ( .A1(n_347), .A2(n_241), .B(n_234), .Y(n_359) );
OAI21x1_ASAP7_75t_L g360 ( .A1(n_333), .A2(n_237), .B(n_215), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_340), .Y(n_361) );
A2O1A1Ixp33_ASAP7_75t_L g362 ( .A1(n_345), .A2(n_348), .B(n_347), .C(n_336), .Y(n_362) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_335), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_344), .A2(n_254), .B1(n_258), .B2(n_260), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_343), .B(n_2), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_340), .A2(n_249), .B1(n_263), .B2(n_265), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_343), .A2(n_271), .B1(n_267), .B2(n_248), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_346), .A2(n_273), .B(n_268), .Y(n_368) );
AOI21xp5_ASAP7_75t_L g369 ( .A1(n_349), .A2(n_264), .B(n_261), .Y(n_369) );
OAI21xp5_ASAP7_75t_L g370 ( .A1(n_338), .A2(n_186), .B(n_187), .Y(n_370) );
OAI21x1_ASAP7_75t_L g371 ( .A1(n_334), .A2(n_257), .B(n_235), .Y(n_371) );
INVx2_ASAP7_75t_SL g372 ( .A(n_337), .Y(n_372) );
AO21x2_ASAP7_75t_L g373 ( .A1(n_347), .A2(n_287), .B(n_282), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_336), .B(n_2), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_336), .Y(n_375) );
AND2x4_ASAP7_75t_L g376 ( .A(n_336), .B(n_3), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_336), .Y(n_377) );
AOI222xp33_ASAP7_75t_L g378 ( .A1(n_342), .A2(n_257), .B1(n_210), .B2(n_235), .C1(n_188), .C2(n_189), .Y(n_378) );
OAI22xp33_ASAP7_75t_L g379 ( .A1(n_336), .A2(n_272), .B1(n_199), .B2(n_211), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_336), .B(n_4), .Y(n_380) );
OAI221xp5_ASAP7_75t_L g381 ( .A1(n_342), .A2(n_235), .B1(n_257), .B2(n_274), .C(n_262), .Y(n_381) );
BUFx3_ASAP7_75t_L g382 ( .A(n_332), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_342), .A2(n_243), .B1(n_231), .B2(n_226), .Y(n_383) );
CKINVDCx14_ASAP7_75t_R g384 ( .A(n_332), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_375), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_377), .B(n_376), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_376), .B(n_4), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_374), .B(n_6), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_380), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_360), .Y(n_390) );
OR2x2_ASAP7_75t_L g391 ( .A(n_363), .B(n_6), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_373), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_361), .B(n_372), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_373), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_366), .B(n_7), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_365), .Y(n_396) );
INVx3_ASAP7_75t_L g397 ( .A(n_357), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_357), .Y(n_398) );
INVxp67_ASAP7_75t_L g399 ( .A(n_382), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_369), .Y(n_400) );
BUFx2_ASAP7_75t_L g401 ( .A(n_351), .Y(n_401) );
OA21x2_ASAP7_75t_L g402 ( .A1(n_371), .A2(n_217), .B(n_194), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_355), .B(n_7), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_367), .B(n_8), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_354), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_362), .B(n_8), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_359), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_370), .Y(n_408) );
AOI21xp33_ASAP7_75t_L g409 ( .A1(n_350), .A2(n_287), .B(n_282), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_384), .Y(n_410) );
BUFx2_ASAP7_75t_L g411 ( .A(n_352), .Y(n_411) );
NOR3xp33_ASAP7_75t_L g412 ( .A(n_381), .B(n_9), .C(n_10), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_358), .B(n_10), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_370), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_364), .B(n_11), .Y(n_415) );
AND2x4_ASAP7_75t_L g416 ( .A(n_368), .B(n_14), .Y(n_416) );
OAI221xp5_ASAP7_75t_L g417 ( .A1(n_353), .A2(n_287), .B1(n_282), .B2(n_13), .C(n_12), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_378), .B(n_11), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_364), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_378), .A2(n_287), .B1(n_282), .B2(n_21), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_356), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_383), .B(n_18), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_379), .Y(n_423) );
INVxp67_ASAP7_75t_SL g424 ( .A(n_375), .Y(n_424) );
INVx3_ASAP7_75t_L g425 ( .A(n_376), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_375), .B(n_20), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_375), .B(n_22), .Y(n_427) );
INVx4_ASAP7_75t_L g428 ( .A(n_376), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_375), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_375), .B(n_23), .Y(n_430) );
INVx4_ASAP7_75t_L g431 ( .A(n_376), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_375), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_375), .B(n_25), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_375), .B(n_27), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_375), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_375), .B(n_172), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_375), .B(n_30), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_375), .Y(n_438) );
BUFx2_ASAP7_75t_L g439 ( .A(n_351), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_375), .B(n_31), .Y(n_440) );
NAND2xp33_ASAP7_75t_R g441 ( .A(n_357), .B(n_34), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_435), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g443 ( .A1(n_411), .A2(n_36), .B1(n_44), .B2(n_45), .C(n_46), .Y(n_443) );
INVx3_ASAP7_75t_L g444 ( .A(n_428), .Y(n_444) );
AOI322xp5_ASAP7_75t_L g445 ( .A1(n_415), .A2(n_56), .A3(n_57), .B1(n_60), .B2(n_62), .C1(n_63), .C2(n_65), .Y(n_445) );
BUFx3_ASAP7_75t_L g446 ( .A(n_401), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_419), .B(n_67), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_387), .B(n_69), .Y(n_448) );
NOR2x1_ASAP7_75t_L g449 ( .A(n_428), .B(n_431), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_415), .B(n_74), .Y(n_450) );
NAND2x1p5_ASAP7_75t_SL g451 ( .A(n_406), .B(n_80), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_424), .B(n_170), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_439), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_388), .B(n_81), .Y(n_454) );
INVx3_ASAP7_75t_L g455 ( .A(n_428), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_393), .B(n_169), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_391), .B(n_83), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_386), .B(n_85), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_385), .Y(n_459) );
INVx2_ASAP7_75t_SL g460 ( .A(n_410), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_429), .Y(n_461) );
NAND4xp75_ASAP7_75t_L g462 ( .A(n_418), .B(n_86), .C(n_87), .D(n_89), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_386), .B(n_168), .Y(n_463) );
AO21x2_ASAP7_75t_L g464 ( .A1(n_392), .A2(n_91), .B(n_92), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_432), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_396), .B(n_438), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_389), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_431), .B(n_425), .Y(n_468) );
INVx2_ASAP7_75t_SL g469 ( .A(n_431), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_398), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_404), .B(n_94), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_425), .B(n_167), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_406), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_404), .B(n_96), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_398), .Y(n_475) );
AND2x4_ASAP7_75t_L g476 ( .A(n_425), .B(n_99), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_408), .B(n_100), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_430), .Y(n_478) );
BUFx2_ASAP7_75t_L g479 ( .A(n_399), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_430), .B(n_101), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_433), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_397), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_397), .Y(n_483) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_421), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_433), .Y(n_485) );
AOI31xp33_ASAP7_75t_L g486 ( .A1(n_441), .A2(n_103), .A3(n_105), .B(n_106), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_397), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_434), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_434), .B(n_107), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_437), .Y(n_490) );
AOI31xp33_ASAP7_75t_SL g491 ( .A1(n_420), .A2(n_109), .A3(n_110), .B(n_112), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_437), .Y(n_492) );
AOI221xp5_ASAP7_75t_L g493 ( .A1(n_412), .A2(n_113), .B1(n_115), .B2(n_116), .C(n_117), .Y(n_493) );
CKINVDCx8_ASAP7_75t_R g494 ( .A(n_416), .Y(n_494) );
NAND2x1_ASAP7_75t_L g495 ( .A(n_416), .B(n_120), .Y(n_495) );
OAI21xp5_ASAP7_75t_L g496 ( .A1(n_420), .A2(n_121), .B(n_123), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_442), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_473), .B(n_408), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_461), .B(n_414), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_459), .Y(n_500) );
OAI21xp33_ASAP7_75t_L g501 ( .A1(n_445), .A2(n_421), .B(n_423), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_465), .Y(n_502) );
INVxp67_ASAP7_75t_SL g503 ( .A(n_470), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_467), .B(n_440), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_466), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_494), .B(n_440), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_466), .B(n_414), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_479), .B(n_427), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_446), .B(n_392), .Y(n_509) );
INVx1_ASAP7_75t_SL g510 ( .A(n_444), .Y(n_510) );
AND2x4_ASAP7_75t_L g511 ( .A(n_449), .B(n_394), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_447), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_475), .Y(n_513) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_482), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_484), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_490), .B(n_413), .Y(n_516) );
NOR2xp67_ASAP7_75t_L g517 ( .A(n_453), .B(n_416), .Y(n_517) );
AND2x4_ASAP7_75t_L g518 ( .A(n_444), .B(n_394), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_478), .B(n_407), .Y(n_519) );
NAND3xp33_ASAP7_75t_SL g520 ( .A(n_443), .B(n_445), .C(n_453), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_447), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_481), .B(n_413), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_446), .B(n_395), .Y(n_523) );
BUFx2_ASAP7_75t_L g524 ( .A(n_455), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_485), .B(n_400), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_460), .B(n_403), .Y(n_526) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_456), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_448), .B(n_422), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_488), .B(n_405), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_484), .Y(n_530) );
AND2x4_ASAP7_75t_L g531 ( .A(n_455), .B(n_469), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_492), .B(n_484), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_450), .B(n_436), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_468), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_458), .B(n_426), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_520), .A2(n_443), .B1(n_441), .B2(n_471), .Y(n_536) );
INVxp67_ASAP7_75t_L g537 ( .A(n_524), .Y(n_537) );
INVx1_ASAP7_75t_SL g538 ( .A(n_510), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_497), .B(n_483), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_534), .B(n_487), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_517), .B(n_486), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_500), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_505), .B(n_451), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_502), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_499), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_509), .B(n_452), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_513), .Y(n_547) );
BUFx2_ASAP7_75t_L g548 ( .A(n_531), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_529), .B(n_451), .Y(n_549) );
INVx2_ASAP7_75t_SL g550 ( .A(n_531), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_499), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_527), .B(n_454), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_522), .B(n_474), .Y(n_553) );
OAI22xp33_ASAP7_75t_L g554 ( .A1(n_520), .A2(n_486), .B1(n_495), .B2(n_463), .Y(n_554) );
INVx2_ASAP7_75t_SL g555 ( .A(n_510), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_525), .B(n_457), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_516), .B(n_476), .Y(n_557) );
INVx2_ASAP7_75t_SL g558 ( .A(n_508), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_503), .B(n_472), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_503), .B(n_476), .Y(n_560) );
AO22x1_ASAP7_75t_L g561 ( .A1(n_548), .A2(n_506), .B1(n_528), .B2(n_511), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_545), .B(n_512), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_554), .A2(n_501), .B1(n_533), .B2(n_535), .Y(n_563) );
NAND3xp33_ASAP7_75t_L g564 ( .A(n_536), .B(n_526), .C(n_519), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_558), .B(n_523), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_551), .B(n_521), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_538), .B(n_507), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_536), .A2(n_498), .B1(n_504), .B2(n_511), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_542), .Y(n_569) );
AOI32xp33_ASAP7_75t_L g570 ( .A1(n_541), .A2(n_550), .A3(n_538), .B1(n_552), .B2(n_549), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_544), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_539), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_543), .B(n_540), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_537), .B(n_498), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_547), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_557), .A2(n_519), .B1(n_532), .B2(n_507), .Y(n_576) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_570), .B(n_555), .Y(n_577) );
INVxp67_ASAP7_75t_L g578 ( .A(n_565), .Y(n_578) );
INVx2_ASAP7_75t_SL g579 ( .A(n_572), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_564), .A2(n_556), .B1(n_553), .B2(n_546), .Y(n_580) );
AOI221xp5_ASAP7_75t_L g581 ( .A1(n_568), .A2(n_417), .B1(n_532), .B2(n_422), .C(n_493), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_567), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_569), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_571), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_573), .B(n_560), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_561), .B(n_514), .Y(n_586) );
OAI321xp33_ASAP7_75t_L g587 ( .A1(n_577), .A2(n_563), .A3(n_576), .B1(n_574), .B2(n_566), .C(n_562), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_583), .Y(n_588) );
AOI21xp33_ASAP7_75t_L g589 ( .A1(n_579), .A2(n_575), .B(n_530), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_586), .A2(n_559), .B1(n_514), .B2(n_518), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_580), .A2(n_518), .B1(n_493), .B2(n_480), .Y(n_591) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_582), .Y(n_592) );
AOI21xp5_ASAP7_75t_L g593 ( .A1(n_587), .A2(n_578), .B(n_580), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g594 ( .A1(n_590), .A2(n_584), .B1(n_585), .B2(n_581), .C(n_496), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_592), .Y(n_595) );
AOI221xp5_ASAP7_75t_L g596 ( .A1(n_589), .A2(n_496), .B1(n_409), .B2(n_489), .C(n_515), .Y(n_596) );
NAND4xp75_ASAP7_75t_L g597 ( .A(n_593), .B(n_591), .C(n_588), .D(n_402), .Y(n_597) );
NOR3x1_ASAP7_75t_L g598 ( .A(n_594), .B(n_462), .C(n_491), .Y(n_598) );
AND2x4_ASAP7_75t_L g599 ( .A(n_595), .B(n_464), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_599), .Y(n_600) );
AND5x1_ASAP7_75t_L g601 ( .A(n_597), .B(n_596), .C(n_491), .D(n_130), .E(n_131), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_600), .Y(n_602) );
NAND2x1p5_ASAP7_75t_L g603 ( .A(n_601), .B(n_598), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_602), .Y(n_604) );
AOI21xp5_ASAP7_75t_L g605 ( .A1(n_603), .A2(n_477), .B(n_464), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_604), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_605), .A2(n_402), .B1(n_477), .B2(n_390), .Y(n_607) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_606), .A2(n_402), .B(n_390), .Y(n_608) );
INVxp67_ASAP7_75t_L g609 ( .A(n_607), .Y(n_609) );
INVxp67_ASAP7_75t_L g610 ( .A(n_609), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_610), .A2(n_608), .B1(n_127), .B2(n_132), .Y(n_611) );
endmodule