module real_aes_4487_n_391 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_1302, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_388, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_1303, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_1301, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_1300, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_1299, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_391);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_1302;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_388;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_1303;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_1301;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_1300;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_1299;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_391;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_830;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_592;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_417;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_527;
wire n_552;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_859;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_954;
wire n_702;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1161;
wire n_686;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_837;
wire n_829;
wire n_1030;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1269;
wire n_677;
wire n_591;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_510;
wire n_550;
wire n_966;
wire n_994;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_807;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1194;
wire n_701;
wire n_809;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1120;
wire n_689;
wire n_946;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_739;
wire n_1162;
wire n_762;
wire n_442;
wire n_740;
wire n_639;
wire n_1186;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_414;
wire n_776;
wire n_1138;
wire n_890;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1055;
wire n_611;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_943;
wire n_977;
wire n_905;
wire n_878;
wire n_577;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1289;
wire n_937;
wire n_773;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_816;
wire n_625;
wire n_953;
wire n_716;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_443;
wire n_1029;
wire n_1207;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_1167;
wire n_609;
wire n_1006;
wire n_1259;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1054;
wire n_1050;
wire n_426;
wire n_1134;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1060;
wire n_1154;
wire n_632;
wire n_714;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1033;
wire n_1028;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_1139;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1127;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_1096;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1240;
wire n_987;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_555;
wire n_1295;
wire n_974;
wire n_857;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_666;
wire n_660;
wire n_886;
wire n_767;
wire n_889;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1198;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_449;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1273;
wire n_959;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_1183;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_698;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_855;
wire n_429;
AOI22xp5_ASAP7_75t_L g836 ( .A1(n_0), .A2(n_243), .B1(n_556), .B2(n_692), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_1), .A2(n_340), .B1(n_531), .B2(n_532), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_2), .A2(n_315), .B1(n_668), .B2(n_669), .Y(n_667) );
INVx1_ASAP7_75t_L g904 ( .A(n_3), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_4), .A2(n_268), .B1(n_525), .B2(n_531), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_5), .A2(n_320), .B1(n_860), .B2(n_861), .Y(n_859) );
INVx1_ASAP7_75t_L g1032 ( .A(n_6), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_7), .A2(n_201), .B1(n_495), .B2(n_661), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_8), .A2(n_317), .B1(n_558), .B2(n_630), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_9), .A2(n_233), .B1(n_416), .B2(n_640), .Y(n_671) );
INVx1_ASAP7_75t_L g486 ( .A(n_10), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_11), .A2(n_130), .B1(n_459), .B2(n_466), .Y(n_458) );
AOI22xp33_ASAP7_75t_SL g805 ( .A1(n_12), .A2(n_306), .B1(n_636), .B2(n_806), .Y(n_805) );
INVx1_ASAP7_75t_SL g950 ( .A(n_13), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_14), .A2(n_151), .B1(n_619), .B2(n_730), .Y(n_913) );
AOI221xp5_ASAP7_75t_L g900 ( .A1(n_15), .A2(n_296), .B1(n_596), .B2(n_901), .C(n_903), .Y(n_900) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_16), .A2(n_74), .B1(n_582), .B2(n_583), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_17), .A2(n_247), .B1(n_519), .B2(n_528), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_18), .A2(n_308), .B1(n_554), .B2(n_582), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_19), .A2(n_21), .B1(n_554), .B2(n_556), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g934 ( .A1(n_20), .A2(n_71), .B1(n_634), .B2(n_635), .Y(n_934) );
NAND2xp5_ASAP7_75t_SL g431 ( .A(n_22), .B(n_421), .Y(n_431) );
AOI21xp33_ASAP7_75t_L g567 ( .A1(n_23), .A2(n_495), .B(n_568), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g838 ( .A1(n_24), .A2(n_252), .B1(n_551), .B2(n_839), .Y(n_838) );
AOI22xp5_ASAP7_75t_L g1080 ( .A1(n_25), .A2(n_359), .B1(n_1075), .B2(n_1081), .Y(n_1080) );
INVx1_ASAP7_75t_L g845 ( .A(n_26), .Y(n_845) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_27), .A2(n_165), .B1(n_416), .B2(n_439), .Y(n_415) );
AOI221x1_ASAP7_75t_L g800 ( .A1(n_28), .A2(n_96), .B1(n_660), .B2(n_801), .C(n_802), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_29), .A2(n_372), .B1(n_454), .B2(n_632), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g1280 ( .A1(n_30), .A2(n_300), .B1(n_466), .B2(n_634), .Y(n_1280) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_31), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_32), .A2(n_37), .B1(n_556), .B2(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g948 ( .A(n_33), .Y(n_948) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_34), .A2(n_223), .B1(n_621), .B2(n_623), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_35), .A2(n_388), .B1(n_510), .B2(n_782), .Y(n_846) );
AOI22xp5_ASAP7_75t_L g875 ( .A1(n_36), .A2(n_182), .B1(n_876), .B2(n_877), .Y(n_875) );
INVx1_ASAP7_75t_L g884 ( .A(n_38), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_39), .A2(n_209), .B1(n_663), .B2(n_664), .Y(n_662) );
INVx1_ASAP7_75t_L g541 ( .A(n_40), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_41), .A2(n_157), .B1(n_734), .B2(n_841), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_42), .A2(n_80), .B1(n_454), .B2(n_632), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_43), .A2(n_259), .B1(n_501), .B2(n_566), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_44), .A2(n_120), .B1(n_521), .B2(n_522), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_45), .A2(n_339), .B1(n_466), .B2(n_634), .Y(n_955) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_46), .B(n_682), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_47), .A2(n_319), .B1(n_471), .B2(n_558), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_48), .A2(n_234), .B1(n_454), .B2(n_551), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_49), .A2(n_309), .B1(n_679), .B2(n_680), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_50), .A2(n_140), .B1(n_521), .B2(n_522), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_51), .A2(n_257), .B1(n_471), .B2(n_558), .Y(n_557) );
AOI22xp5_ASAP7_75t_L g1010 ( .A1(n_52), .A2(n_239), .B1(n_554), .B2(n_1011), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_53), .A2(n_390), .B1(n_617), .B2(n_619), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_54), .A2(n_358), .B1(n_537), .B2(n_709), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_55), .A2(n_115), .B1(n_454), .B2(n_632), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_56), .B(n_728), .Y(n_946) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_57), .A2(n_386), .B1(n_459), .B2(n_549), .Y(n_586) );
OA22x2_ASAP7_75t_L g426 ( .A1(n_58), .A2(n_168), .B1(n_421), .B2(n_425), .Y(n_426) );
INVx1_ASAP7_75t_L g446 ( .A(n_58), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_59), .A2(n_202), .B1(n_561), .B2(n_591), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_60), .A2(n_212), .B1(n_1065), .B2(n_1067), .Y(n_1064) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_61), .A2(n_336), .B1(n_527), .B2(n_528), .Y(n_526) );
CKINVDCx5p33_ASAP7_75t_R g813 ( .A(n_62), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_63), .A2(n_200), .B1(n_1055), .B2(n_1062), .Y(n_1110) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_64), .A2(n_274), .B1(n_497), .B2(n_857), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_65), .A2(n_262), .B1(n_454), .B2(n_551), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_66), .A2(n_156), .B1(n_510), .B2(n_726), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_67), .A2(n_379), .B1(n_518), .B2(n_551), .Y(n_798) );
INVx1_ASAP7_75t_L g853 ( .A(n_68), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_69), .B(n_591), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_70), .A2(n_326), .B1(n_549), .B2(n_634), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_72), .A2(n_328), .B1(n_558), .B2(n_786), .Y(n_785) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_73), .B(n_192), .Y(n_401) );
INVx1_ASAP7_75t_L g424 ( .A(n_73), .Y(n_424) );
OAI21xp33_ASAP7_75t_L g447 ( .A1(n_73), .A2(n_168), .B(n_448), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g790 ( .A1(n_75), .A2(n_354), .B1(n_459), .B2(n_549), .Y(n_790) );
AO221x2_ASAP7_75t_L g1084 ( .A1(n_76), .A2(n_360), .B1(n_1055), .B2(n_1073), .C(n_1085), .Y(n_1084) );
AOI21xp5_ASAP7_75t_L g862 ( .A1(n_77), .A2(n_863), .B(n_866), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_78), .A2(n_345), .B1(n_872), .B2(n_874), .Y(n_871) );
AOI22xp5_ASAP7_75t_L g1008 ( .A1(n_79), .A2(n_269), .B1(n_582), .B2(n_786), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_81), .A2(n_277), .B1(n_459), .B2(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g754 ( .A(n_82), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_83), .A2(n_224), .B1(n_459), .B2(n_734), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_84), .A2(n_193), .B1(n_596), .B2(n_940), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_85), .A2(n_249), .B1(n_680), .B2(n_728), .Y(n_992) );
AOI22xp5_ASAP7_75t_L g1087 ( .A1(n_86), .A2(n_348), .B1(n_1062), .B2(n_1088), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_87), .A2(n_368), .B1(n_473), .B2(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g1035 ( .A(n_88), .Y(n_1035) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_89), .A2(n_365), .B1(n_1067), .B2(n_1075), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_90), .A2(n_230), .B1(n_473), .B2(n_668), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_91), .A2(n_112), .B1(n_634), .B2(n_635), .Y(n_633) );
AOI21xp33_ASAP7_75t_L g595 ( .A1(n_92), .A2(n_596), .B(n_597), .Y(n_595) );
XOR2x2_ASAP7_75t_L g1021 ( .A(n_93), .B(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_L g1059 ( .A(n_94), .Y(n_1059) );
AND2x4_ASAP7_75t_L g1066 ( .A(n_94), .B(n_287), .Y(n_1066) );
HB1xp67_ASAP7_75t_L g1296 ( .A(n_94), .Y(n_1296) );
INVx1_ASAP7_75t_L g867 ( .A(n_95), .Y(n_867) );
AO22x1_ASAP7_75t_L g1085 ( .A1(n_97), .A2(n_199), .B1(n_1065), .B2(n_1081), .Y(n_1085) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_98), .A2(n_303), .B1(n_459), .B2(n_549), .Y(n_693) );
INVx1_ASAP7_75t_L g982 ( .A(n_99), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_100), .A2(n_161), .B1(n_510), .B2(n_680), .Y(n_1014) );
INVx1_ASAP7_75t_L g1038 ( .A(n_101), .Y(n_1038) );
AOI22xp33_ASAP7_75t_SL g638 ( .A1(n_102), .A2(n_176), .B1(n_639), .B2(n_640), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_103), .A2(n_375), .B1(n_549), .B2(n_634), .Y(n_995) );
AO22x1_ASAP7_75t_L g581 ( .A1(n_104), .A2(n_333), .B1(n_582), .B2(n_583), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g1090 ( .A1(n_105), .A2(n_138), .B1(n_1076), .B2(n_1091), .Y(n_1090) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_106), .A2(n_191), .B1(n_609), .B2(n_728), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_107), .A2(n_153), .B1(n_510), .B2(n_593), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g1288 ( .A1(n_108), .A2(n_1289), .B1(n_1290), .B2(n_1291), .Y(n_1288) );
INVx1_ASAP7_75t_L g1289 ( .A(n_108), .Y(n_1289) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_109), .A2(n_227), .B1(n_510), .B2(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_110), .B(n_563), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_111), .A2(n_124), .B1(n_663), .B2(n_679), .Y(n_912) );
INVx1_ASAP7_75t_L g1004 ( .A(n_113), .Y(n_1004) );
AOI22xp33_ASAP7_75t_SL g631 ( .A1(n_114), .A2(n_119), .B1(n_454), .B2(n_632), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_116), .A2(n_196), .B1(n_439), .B2(n_639), .Y(n_956) );
AOI22xp5_ASAP7_75t_L g1012 ( .A1(n_117), .A2(n_134), .B1(n_471), .B2(n_669), .Y(n_1012) );
INVx1_ASAP7_75t_L g1057 ( .A(n_118), .Y(n_1057) );
AND2x4_ASAP7_75t_L g1063 ( .A(n_118), .B(n_397), .Y(n_1063) );
INVx1_ASAP7_75t_SL g1089 ( .A(n_118), .Y(n_1089) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_121), .A2(n_370), .B1(n_669), .B2(n_908), .Y(n_907) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_122), .B(n_563), .Y(n_599) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_123), .A2(n_608), .B(n_611), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_125), .A2(n_264), .B1(n_668), .B2(n_669), .Y(n_763) );
AOI22xp33_ASAP7_75t_SL g998 ( .A1(n_126), .A2(n_128), .B1(n_473), .B2(n_668), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_127), .B(n_534), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g777 ( .A1(n_129), .A2(n_481), .B(n_778), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g1109 ( .A1(n_131), .A2(n_160), .B1(n_1075), .B2(n_1081), .Y(n_1109) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_132), .A2(n_256), .B1(n_495), .B2(n_497), .Y(n_494) );
AOI33xp33_ASAP7_75t_R g737 ( .A1(n_133), .A2(n_266), .A3(n_418), .B1(n_442), .B2(n_738), .B3(n_1299), .Y(n_737) );
INVx1_ASAP7_75t_L g545 ( .A(n_135), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_136), .A2(n_343), .B1(n_525), .B2(n_528), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_137), .A2(n_280), .B1(n_524), .B2(n_525), .Y(n_523) );
AO22x1_ASAP7_75t_L g909 ( .A1(n_139), .A2(n_335), .B1(n_632), .B2(n_639), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_141), .A2(n_347), .B1(n_596), .B2(n_657), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g1274 ( .A1(n_142), .A2(n_273), .B1(n_660), .B2(n_661), .Y(n_1274) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_143), .A2(n_241), .B1(n_841), .B2(n_879), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_144), .A2(n_172), .B1(n_630), .B2(n_736), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_145), .A2(n_276), .B1(n_519), .B2(n_524), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_146), .A2(n_206), .B1(n_661), .B2(n_682), .Y(n_947) );
AOI22xp5_ASAP7_75t_L g1272 ( .A1(n_147), .A2(n_246), .B1(n_1037), .B2(n_1273), .Y(n_1272) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_148), .A2(n_283), .B1(n_450), .B2(n_454), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_149), .B(n_759), .Y(n_758) );
AOI221xp5_ASAP7_75t_L g843 ( .A1(n_150), .A2(n_312), .B1(n_536), .B2(n_539), .C(n_844), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_152), .A2(n_301), .B1(n_684), .B2(n_724), .Y(n_723) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_154), .A2(n_605), .B1(n_641), .B2(n_642), .Y(n_604) );
INVx1_ASAP7_75t_L g641 ( .A(n_154), .Y(n_641) );
AOI22x1_ASAP7_75t_L g643 ( .A1(n_154), .A2(n_605), .B1(n_641), .B2(n_642), .Y(n_643) );
INVx1_ASAP7_75t_L g612 ( .A(n_155), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_158), .B(n_563), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_159), .A2(n_238), .B1(n_660), .B2(n_661), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_162), .A2(n_183), .B1(n_454), .B2(n_582), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_163), .A2(n_374), .B1(n_668), .B2(n_669), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_164), .A2(n_353), .B1(n_686), .B2(n_687), .Y(n_685) );
CKINVDCx6p67_ASAP7_75t_R g978 ( .A(n_166), .Y(n_978) );
INVx1_ASAP7_75t_L g438 ( .A(n_167), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_167), .B(n_444), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_167), .B(n_221), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_168), .B(n_295), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_169), .A2(n_237), .B1(n_1053), .B2(n_1060), .Y(n_1052) );
XNOR2x1_ASAP7_75t_L g514 ( .A(n_170), .B(n_515), .Y(n_514) );
XNOR2x2_ASAP7_75t_SL g542 ( .A(n_170), .B(n_515), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g1278 ( .A1(n_171), .A2(n_181), .B1(n_632), .B2(n_908), .Y(n_1278) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_173), .A2(n_355), .B1(n_454), .B2(n_632), .Y(n_666) );
INVx1_ASAP7_75t_L g959 ( .A(n_174), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_175), .A2(n_189), .B1(n_630), .B2(n_736), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_177), .B(n_536), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_178), .A2(n_198), .B1(n_518), .B2(n_527), .Y(n_894) );
INVx1_ASAP7_75t_L g960 ( .A(n_179), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_180), .A2(n_272), .B1(n_632), .B2(n_639), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_184), .A2(n_291), .B1(n_554), .B2(n_556), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_185), .B(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g748 ( .A(n_186), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_187), .A2(n_235), .B1(n_416), .B2(n_439), .Y(n_764) );
INVx1_ASAP7_75t_L g1030 ( .A(n_188), .Y(n_1030) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_190), .A2(n_204), .B1(n_663), .B2(n_711), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_192), .B(n_430), .Y(n_429) );
AOI22x1_ASAP7_75t_L g500 ( .A1(n_194), .A2(n_385), .B1(n_501), .B2(n_510), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_195), .A2(n_211), .B1(n_454), .B2(n_473), .Y(n_1045) );
AOI22xp5_ASAP7_75t_L g937 ( .A1(n_197), .A2(n_361), .B1(n_639), .B2(n_640), .Y(n_937) );
XNOR2x1_ASAP7_75t_L g1268 ( .A(n_200), .B(n_1269), .Y(n_1268) );
AOI22xp33_ASAP7_75t_L g1287 ( .A1(n_200), .A2(n_1288), .B1(n_1292), .B2(n_1294), .Y(n_1287) );
AOI22xp5_ASAP7_75t_L g996 ( .A1(n_203), .A2(n_316), .B1(n_639), .B2(n_640), .Y(n_996) );
CKINVDCx5p33_ASAP7_75t_R g818 ( .A(n_205), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_207), .A2(n_245), .B1(n_459), .B2(n_549), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_208), .A2(n_378), .B1(n_518), .B2(n_519), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_210), .A2(n_381), .B1(n_536), .B2(n_711), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_213), .A2(n_377), .B1(n_471), .B2(n_473), .Y(n_470) );
INVx1_ASAP7_75t_L g752 ( .A(n_214), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_215), .A2(n_334), .B1(n_439), .B2(n_668), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_216), .A2(n_292), .B1(n_524), .B2(n_527), .Y(n_810) );
XOR2x2_ASAP7_75t_L g720 ( .A(n_217), .B(n_721), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g1072 ( .A1(n_217), .A2(n_253), .B1(n_1055), .B2(n_1073), .Y(n_1072) );
AOI22xp5_ASAP7_75t_L g1043 ( .A1(n_218), .A2(n_307), .B1(n_466), .B2(n_1044), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_219), .A2(n_290), .B1(n_518), .B2(n_539), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_220), .A2(n_373), .B1(n_521), .B2(n_522), .Y(n_895) );
INVx1_ASAP7_75t_L g422 ( .A(n_221), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g781 ( .A1(n_222), .A2(n_351), .B1(n_510), .B2(n_782), .Y(n_781) );
CKINVDCx5p33_ASAP7_75t_R g820 ( .A(n_225), .Y(n_820) );
INVx1_ASAP7_75t_L g898 ( .A(n_226), .Y(n_898) );
OAI222xp33_ASAP7_75t_L g910 ( .A1(n_226), .A2(n_911), .B1(n_914), .B2(n_915), .C1(n_1302), .C2(n_1303), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_226), .B(n_915), .Y(n_919) );
INVx1_ASAP7_75t_L g833 ( .A(n_228), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g1102 ( .A1(n_228), .A2(n_330), .B1(n_1055), .B2(n_1062), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_229), .A2(n_371), .B1(n_524), .B2(n_525), .Y(n_893) );
INVx1_ASAP7_75t_L g964 ( .A(n_231), .Y(n_964) );
INVx1_ASAP7_75t_L g757 ( .A(n_232), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g1281 ( .A1(n_236), .A2(n_263), .B1(n_639), .B2(n_1282), .Y(n_1281) );
AOI22x1_ASAP7_75t_L g741 ( .A1(n_237), .A2(n_742), .B1(n_743), .B2(n_765), .Y(n_741) );
INVx1_ASAP7_75t_L g765 ( .A(n_237), .Y(n_765) );
AOI22xp5_ASAP7_75t_L g1082 ( .A1(n_240), .A2(n_279), .B1(n_1055), .B2(n_1062), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_242), .A2(n_278), .B1(n_466), .B2(n_634), .Y(n_670) );
INVx1_ASAP7_75t_L g945 ( .A(n_244), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g1271 ( .A(n_248), .B(n_654), .Y(n_1271) );
AOI22xp33_ASAP7_75t_SL g787 ( .A1(n_250), .A2(n_302), .B1(n_471), .B2(n_788), .Y(n_787) );
AOI221xp5_ASAP7_75t_L g1016 ( .A1(n_251), .A2(n_270), .B1(n_596), .B2(n_801), .C(n_1017), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g1096 ( .A1(n_254), .A2(n_322), .B1(n_1055), .B2(n_1060), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g1101 ( .A1(n_255), .A2(n_313), .B1(n_1065), .B2(n_1081), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_258), .A2(n_376), .B1(n_536), .B2(n_537), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g1074 ( .A1(n_260), .A2(n_356), .B1(n_1075), .B2(n_1076), .Y(n_1074) );
OAI21x1_ASAP7_75t_L g576 ( .A1(n_261), .A2(n_577), .B(n_600), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_261), .B(n_580), .Y(n_603) );
INVx1_ASAP7_75t_L g968 ( .A(n_265), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_267), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g988 ( .A(n_271), .Y(n_988) );
INVx1_ASAP7_75t_L g569 ( .A(n_275), .Y(n_569) );
INVx1_ASAP7_75t_L g1025 ( .A(n_281), .Y(n_1025) );
INVx1_ASAP7_75t_L g1018 ( .A(n_282), .Y(n_1018) );
INVx1_ASAP7_75t_L g773 ( .A(n_284), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_284), .B(n_789), .Y(n_793) );
AOI21xp5_ASAP7_75t_L g941 ( .A1(n_285), .A2(n_942), .B(n_944), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g1279 ( .A1(n_286), .A2(n_327), .B1(n_668), .B2(n_669), .Y(n_1279) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_287), .Y(n_402) );
AND2x4_ASAP7_75t_L g1058 ( .A(n_287), .B(n_1059), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_288), .A2(n_294), .B1(n_527), .B2(n_528), .Y(n_716) );
CKINVDCx5p33_ASAP7_75t_R g815 ( .A(n_289), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_293), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g436 ( .A(n_295), .Y(n_436) );
INVxp67_ASAP7_75t_L g509 ( .A(n_295), .Y(n_509) );
INVx1_ASAP7_75t_L g598 ( .A(n_297), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_298), .B(n_682), .Y(n_750) );
INVx1_ASAP7_75t_L g983 ( .A(n_299), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_304), .A2(n_349), .B1(n_466), .B2(n_634), .Y(n_914) );
INVx2_ASAP7_75t_L g397 ( .A(n_305), .Y(n_397) );
INVx1_ASAP7_75t_SL g799 ( .A(n_310), .Y(n_799) );
NOR3xp33_ASAP7_75t_L g826 ( .A(n_310), .B(n_827), .C(n_828), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_311), .A2(n_363), .B1(n_495), .B2(n_497), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_314), .A2(n_380), .B1(n_711), .B2(n_782), .Y(n_969) );
AOI21xp5_ASAP7_75t_SL g480 ( .A1(n_318), .A2(n_481), .B(n_485), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_321), .A2(n_324), .B1(n_531), .B2(n_537), .Y(n_888) );
XNOR2x2_ASAP7_75t_L g650 ( .A(n_322), .B(n_651), .Y(n_650) );
XOR2xp5_ASAP7_75t_L g695 ( .A(n_322), .B(n_651), .Y(n_695) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_323), .Y(n_512) );
AOI21xp33_ASAP7_75t_L g538 ( .A1(n_325), .A2(n_539), .B(n_540), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_329), .A2(n_342), .B1(n_556), .B2(n_639), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_331), .A2(n_350), .B1(n_561), .B2(n_684), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_332), .A2(n_346), .B1(n_539), .B2(n_709), .Y(n_887) );
INVx1_ASAP7_75t_L g779 ( .A(n_337), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_338), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g985 ( .A(n_341), .Y(n_985) );
AOI21xp5_ASAP7_75t_L g746 ( .A1(n_344), .A2(n_477), .B(n_747), .Y(n_746) );
XOR2xp5_ASAP7_75t_L g703 ( .A(n_348), .B(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_352), .B(n_664), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_357), .A2(n_362), .B1(n_561), .B2(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g694 ( .A(n_360), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_364), .A2(n_387), .B1(n_534), .B2(n_728), .Y(n_889) );
AND2x2_ASAP7_75t_L g802 ( .A(n_366), .B(n_614), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_367), .A2(n_383), .B1(n_629), .B2(n_640), .Y(n_1041) );
INVx1_ASAP7_75t_L g966 ( .A(n_369), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g1275 ( .A1(n_382), .A2(n_389), .B1(n_501), .B2(n_1276), .Y(n_1275) );
INVx1_ASAP7_75t_L g990 ( .A(n_384), .Y(n_990) );
AOI21xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_403), .B(n_1048), .Y(n_391) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
BUFx4_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
NAND3xp33_ASAP7_75t_L g394 ( .A(n_395), .B(n_398), .C(n_402), .Y(n_394) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_395), .B(n_1285), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_395), .B(n_1286), .Y(n_1293) );
AOI21xp5_ASAP7_75t_L g1297 ( .A1(n_395), .A2(n_402), .B(n_1089), .Y(n_1297) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AO21x1_ASAP7_75t_L g1295 ( .A1(n_396), .A2(n_1296), .B(n_1297), .Y(n_1295) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_397), .B(n_1057), .Y(n_1056) );
AND3x4_ASAP7_75t_L g1088 ( .A(n_397), .B(n_1058), .C(n_1089), .Y(n_1088) );
NOR2xp33_ASAP7_75t_L g1285 ( .A(n_398), .B(n_1286), .Y(n_1285) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AO21x2_ASAP7_75t_L g489 ( .A1(n_399), .A2(n_490), .B(n_492), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
INVx1_ASAP7_75t_L g1286 ( .A(n_402), .Y(n_1286) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B1(n_767), .B2(n_1047), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AOI22x1_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_408), .B1(n_646), .B2(n_647), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AO22x2_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_572), .B1(n_573), .B2(n_645), .Y(n_408) );
INVx2_ASAP7_75t_L g645 ( .A(n_409), .Y(n_645) );
XOR2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_543), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_412), .B1(n_513), .B2(n_542), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
XNOR2xp5_ASAP7_75t_L g412 ( .A(n_413), .B(n_512), .Y(n_412) );
NOR3xp33_ASAP7_75t_SL g413 ( .A(n_414), .B(n_457), .C(n_475), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_415), .B(n_449), .Y(n_414) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx8_ASAP7_75t_L g639 ( .A(n_417), .Y(n_639) );
AND2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_427), .Y(n_417) );
AND2x4_ASAP7_75t_L g451 ( .A(n_418), .B(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g479 ( .A(n_418), .B(n_468), .Y(n_479) );
AND2x2_ASAP7_75t_L g511 ( .A(n_418), .B(n_464), .Y(n_511) );
AND2x4_ASAP7_75t_L g518 ( .A(n_418), .B(n_427), .Y(n_518) );
AND2x4_ASAP7_75t_L g519 ( .A(n_418), .B(n_456), .Y(n_519) );
AND2x4_ASAP7_75t_L g531 ( .A(n_418), .B(n_464), .Y(n_531) );
AND2x2_ASAP7_75t_L g536 ( .A(n_418), .B(n_468), .Y(n_536) );
AND2x2_ASAP7_75t_L g555 ( .A(n_418), .B(n_427), .Y(n_555) );
AND2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_426), .Y(n_418) );
INVx1_ASAP7_75t_L g462 ( .A(n_419), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_423), .Y(n_419) );
NAND2xp33_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
INVx2_ASAP7_75t_L g425 ( .A(n_421), .Y(n_425) );
INVx3_ASAP7_75t_L g430 ( .A(n_421), .Y(n_430) );
NAND2xp33_ASAP7_75t_L g437 ( .A(n_421), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g448 ( .A(n_421), .Y(n_448) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_421), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_422), .B(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_424), .A2(n_448), .B(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g463 ( .A(n_426), .Y(n_463) );
AND2x2_ASAP7_75t_L g484 ( .A(n_426), .B(n_462), .Y(n_484) );
AND2x2_ASAP7_75t_L g507 ( .A(n_426), .B(n_508), .Y(n_507) );
AND2x4_ASAP7_75t_L g441 ( .A(n_427), .B(n_442), .Y(n_441) );
AND2x4_ASAP7_75t_L g472 ( .A(n_427), .B(n_461), .Y(n_472) );
AND2x4_ASAP7_75t_L g524 ( .A(n_427), .B(n_461), .Y(n_524) );
AND2x4_ASAP7_75t_L g527 ( .A(n_427), .B(n_442), .Y(n_527) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_427), .Y(n_738) );
AND2x4_ASAP7_75t_L g427 ( .A(n_428), .B(n_432), .Y(n_427) );
OR2x2_ASAP7_75t_L g453 ( .A(n_428), .B(n_433), .Y(n_453) );
AND2x4_ASAP7_75t_L g464 ( .A(n_428), .B(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g469 ( .A(n_428), .Y(n_469) );
AND2x2_ASAP7_75t_L g504 ( .A(n_428), .B(n_505), .Y(n_504) );
AND2x4_ASAP7_75t_L g428 ( .A(n_429), .B(n_431), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_430), .B(n_436), .Y(n_435) );
INVxp67_ASAP7_75t_L g444 ( .A(n_430), .Y(n_444) );
NAND3xp33_ASAP7_75t_L g492 ( .A(n_431), .B(n_443), .C(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g465 ( .A(n_434), .Y(n_465) );
AND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_437), .Y(n_434) );
INVx4_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx4_ASAP7_75t_L g556 ( .A(n_440), .Y(n_556) );
INVx4_ASAP7_75t_L g640 ( .A(n_440), .Y(n_640) );
INVx1_ASAP7_75t_L g788 ( .A(n_440), .Y(n_788) );
INVx2_ASAP7_75t_SL g1011 ( .A(n_440), .Y(n_1011) );
INVx1_ASAP7_75t_L g1282 ( .A(n_440), .Y(n_1282) );
INVx8_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AND2x4_ASAP7_75t_L g455 ( .A(n_442), .B(n_456), .Y(n_455) );
AND2x4_ASAP7_75t_L g499 ( .A(n_442), .B(n_468), .Y(n_499) );
AND2x4_ASAP7_75t_L g528 ( .A(n_442), .B(n_456), .Y(n_528) );
AND2x4_ASAP7_75t_L g537 ( .A(n_442), .B(n_468), .Y(n_537) );
AND2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_447), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
BUFx12f_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_451), .Y(n_551) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_451), .Y(n_582) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_451), .Y(n_632) );
BUFx3_ASAP7_75t_L g876 ( .A(n_451), .Y(n_876) );
AND2x4_ASAP7_75t_L g525 ( .A(n_452), .B(n_461), .Y(n_525) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g456 ( .A(n_453), .Y(n_456) );
BUFx12f_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx6_ASAP7_75t_L g584 ( .A(n_455), .Y(n_584) );
AND2x4_ASAP7_75t_L g474 ( .A(n_456), .B(n_461), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_470), .Y(n_457) );
BUFx12f_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_460), .Y(n_634) );
INVx3_ASAP7_75t_L g807 ( .A(n_460), .Y(n_807) );
AND2x4_ASAP7_75t_L g460 ( .A(n_461), .B(n_464), .Y(n_460) );
AND2x2_ASAP7_75t_L g467 ( .A(n_461), .B(n_468), .Y(n_467) );
AND2x4_ASAP7_75t_L g521 ( .A(n_461), .B(n_464), .Y(n_521) );
AND2x4_ASAP7_75t_L g522 ( .A(n_461), .B(n_468), .Y(n_522) );
AND2x4_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
AND2x4_ASAP7_75t_L g483 ( .A(n_464), .B(n_484), .Y(n_483) );
AND2x4_ASAP7_75t_L g539 ( .A(n_464), .B(n_484), .Y(n_539) );
AND2x4_ASAP7_75t_L g468 ( .A(n_465), .B(n_469), .Y(n_468) );
BUFx5_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_467), .Y(n_549) );
INVx1_ASAP7_75t_L g637 ( .A(n_467), .Y(n_637) );
BUFx3_ASAP7_75t_L g734 ( .A(n_467), .Y(n_734) );
AND2x4_ASAP7_75t_L g496 ( .A(n_468), .B(n_484), .Y(n_496) );
AND2x2_ASAP7_75t_L g534 ( .A(n_468), .B(n_484), .Y(n_534) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx12f_ASAP7_75t_L g630 ( .A(n_472), .Y(n_630) );
BUFx6f_ASAP7_75t_L g668 ( .A(n_472), .Y(n_668) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_474), .Y(n_558) );
BUFx6f_ASAP7_75t_L g669 ( .A(n_474), .Y(n_669) );
BUFx6f_ASAP7_75t_L g736 ( .A(n_474), .Y(n_736) );
NAND4xp25_ASAP7_75t_L g475 ( .A(n_476), .B(n_480), .C(n_494), .D(n_500), .Y(n_475) );
INVx3_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g563 ( .A(n_478), .Y(n_563) );
INVx2_ASAP7_75t_L g801 ( .A(n_478), .Y(n_801) );
INVx2_ASAP7_75t_L g865 ( .A(n_478), .Y(n_865) );
INVx3_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g610 ( .A(n_479), .Y(n_610) );
BUFx3_ASAP7_75t_L g686 ( .A(n_479), .Y(n_686) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g1037 ( .A(n_482), .Y(n_1037) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx3_ASAP7_75t_L g566 ( .A(n_483), .Y(n_566) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_483), .Y(n_596) );
BUFx3_ASAP7_75t_L g684 ( .A(n_483), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_487), .B(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g687 ( .A(n_487), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g778 ( .A(n_487), .B(n_779), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g844 ( .A(n_487), .B(n_845), .Y(n_844) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_488), .B(n_541), .Y(n_540) );
INVx2_ASAP7_75t_SL g711 ( .A(n_488), .Y(n_711) );
INVx2_ASAP7_75t_L g728 ( .A(n_488), .Y(n_728) );
BUFx6f_ASAP7_75t_L g1019 ( .A(n_488), .Y(n_1019) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx3_ASAP7_75t_L g571 ( .A(n_489), .Y(n_571) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_491), .B(n_506), .Y(n_505) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_496), .Y(n_591) );
INVx2_ASAP7_75t_L g618 ( .A(n_496), .Y(n_618) );
BUFx8_ASAP7_75t_SL g660 ( .A(n_496), .Y(n_660) );
BUFx3_ASAP7_75t_L g730 ( .A(n_496), .Y(n_730) );
INVx2_ASAP7_75t_L g965 ( .A(n_496), .Y(n_965) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx3_ASAP7_75t_L g661 ( .A(n_498), .Y(n_661) );
INVx2_ASAP7_75t_L g724 ( .A(n_498), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_498), .A2(n_985), .B1(n_986), .B2(n_988), .Y(n_984) );
INVx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_499), .Y(n_561) );
BUFx6f_ASAP7_75t_L g619 ( .A(n_499), .Y(n_619) );
INVx4_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
OAI21xp33_ASAP7_75t_L g611 ( .A1(n_502), .A2(n_612), .B(n_613), .Y(n_611) );
INVx2_ASAP7_75t_L g663 ( .A(n_502), .Y(n_663) );
INVx3_ASAP7_75t_L g759 ( .A(n_502), .Y(n_759) );
INVx2_ASAP7_75t_L g782 ( .A(n_502), .Y(n_782) );
OAI21xp5_ASAP7_75t_L g944 ( .A1(n_502), .A2(n_945), .B(n_946), .Y(n_944) );
INVx5_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx4f_ASAP7_75t_L g593 ( .A(n_503), .Y(n_593) );
BUFx2_ASAP7_75t_L g680 ( .A(n_503), .Y(n_680) );
BUFx2_ASAP7_75t_L g726 ( .A(n_503), .Y(n_726) );
AND2x4_ASAP7_75t_L g503 ( .A(n_504), .B(n_507), .Y(n_503) );
AND2x4_ASAP7_75t_L g532 ( .A(n_504), .B(n_507), .Y(n_532) );
AND2x2_ASAP7_75t_L g709 ( .A(n_504), .B(n_507), .Y(n_709) );
BUFx3_ASAP7_75t_L g861 ( .A(n_510), .Y(n_861) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g626 ( .A(n_511), .Y(n_626) );
BUFx3_ASAP7_75t_L g679 ( .A(n_511), .Y(n_679) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
OR2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_529), .Y(n_515) );
NAND4xp25_ASAP7_75t_L g516 ( .A(n_517), .B(n_520), .C(n_523), .D(n_526), .Y(n_516) );
NAND4xp25_ASAP7_75t_L g529 ( .A(n_530), .B(n_533), .C(n_535), .D(n_538), .Y(n_529) );
INVx2_ASAP7_75t_L g821 ( .A(n_531), .Y(n_821) );
INVx4_ASAP7_75t_L g814 ( .A(n_532), .Y(n_814) );
INVx2_ASAP7_75t_L g816 ( .A(n_537), .Y(n_816) );
INVx2_ASAP7_75t_L g819 ( .A(n_539), .Y(n_819) );
BUFx3_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
XNOR2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
NOR4xp75_ASAP7_75t_L g546 ( .A(n_547), .B(n_552), .C(n_559), .D(n_564), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_557), .Y(n_552) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
BUFx4f_ASAP7_75t_L g692 ( .A(n_555), .Y(n_692) );
BUFx3_ASAP7_75t_L g874 ( .A(n_558), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_562), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_565), .B(n_567), .Y(n_564) );
INVx2_ASAP7_75t_L g622 ( .A(n_566), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
INVx1_ASAP7_75t_L g664 ( .A(n_570), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g903 ( .A(n_570), .B(n_904), .Y(n_903) );
INVx4_ASAP7_75t_L g1276 ( .A(n_570), .Y(n_1276) );
INVx4_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx3_ASAP7_75t_L g615 ( .A(n_571), .Y(n_615) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_604), .B1(n_643), .B2(n_644), .Y(n_573) );
INVx1_ASAP7_75t_L g644 ( .A(n_574), .Y(n_644) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_588), .Y(n_577) );
NOR3xp33_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .C(n_585), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NOR3xp33_ASAP7_75t_L g602 ( .A(n_581), .B(n_594), .C(n_603), .Y(n_602) );
INVx5_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g786 ( .A(n_584), .Y(n_786) );
INVx3_ASAP7_75t_L g839 ( .A(n_584), .Y(n_839) );
INVx1_ASAP7_75t_L g908 ( .A(n_584), .Y(n_908) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_585), .B(n_589), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_589), .B(n_594), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_592), .Y(n_589) );
INVx2_ASAP7_75t_L g858 ( .A(n_591), .Y(n_858) );
INVx2_ASAP7_75t_SL g868 ( .A(n_593), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_599), .Y(n_594) );
INVx4_ASAP7_75t_L g753 ( .A(n_596), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx2_ASAP7_75t_L g642 ( .A(n_605), .Y(n_642) );
OR2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_627), .Y(n_605) );
NAND3xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_616), .C(n_620), .Y(n_606) );
BUFx3_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
BUFx6f_ASAP7_75t_L g655 ( .A(n_610), .Y(n_655) );
INVx4_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx3_ASAP7_75t_L g682 ( .A(n_618), .Y(n_682) );
INVx4_ASAP7_75t_L g1033 ( .A(n_619), .Y(n_1033) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
BUFx6f_ASAP7_75t_L g658 ( .A(n_626), .Y(n_658) );
INVx1_ASAP7_75t_L g962 ( .A(n_626), .Y(n_962) );
NAND4xp25_ASAP7_75t_SL g627 ( .A(n_628), .B(n_631), .C(n_633), .D(n_638), .Y(n_627) );
BUFx12f_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g873 ( .A(n_630), .Y(n_873) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
XNOR2x1_ASAP7_75t_L g647 ( .A(n_648), .B(n_698), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_672), .B1(n_695), .B2(n_696), .Y(n_649) );
OR2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_665), .Y(n_651) );
NAND4xp25_ASAP7_75t_L g652 ( .A(n_653), .B(n_656), .C(n_659), .D(n_662), .Y(n_652) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_L g1027 ( .A(n_655), .Y(n_1027) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
OAI21xp33_ASAP7_75t_L g756 ( .A1(n_658), .A2(n_757), .B(n_758), .Y(n_756) );
INVx2_ASAP7_75t_L g940 ( .A(n_658), .Y(n_940) );
INVx2_ASAP7_75t_L g1273 ( .A(n_658), .Y(n_1273) );
INVx1_ASAP7_75t_L g755 ( .A(n_661), .Y(n_755) );
NAND4xp25_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .C(n_670), .D(n_671), .Y(n_665) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g697 ( .A(n_673), .Y(n_697) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
XOR2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_694), .Y(n_675) );
NOR2x1_ASAP7_75t_L g676 ( .A(n_677), .B(n_688), .Y(n_676) );
NAND4xp25_ASAP7_75t_L g677 ( .A(n_678), .B(n_681), .C(n_683), .D(n_685), .Y(n_677) );
INVx2_ASAP7_75t_L g1039 ( .A(n_679), .Y(n_1039) );
BUFx2_ASAP7_75t_L g860 ( .A(n_684), .Y(n_860) );
INVx2_ASAP7_75t_L g902 ( .A(n_686), .Y(n_902) );
NAND4xp25_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .C(n_691), .D(n_693), .Y(n_688) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
XNOR2x1_ASAP7_75t_L g698 ( .A(n_699), .B(n_717), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
XNOR2x1_ASAP7_75t_L g831 ( .A(n_702), .B(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
OR2x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_712), .Y(n_704) );
NAND4xp25_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .C(n_708), .D(n_710), .Y(n_705) );
NAND4xp25_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .C(n_715), .D(n_716), .Y(n_712) );
OAI21x1_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_739), .B(n_766), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_720), .B(n_741), .Y(n_766) );
NOR2x1_ASAP7_75t_L g721 ( .A(n_722), .B(n_731), .Y(n_721) );
NAND4xp25_ASAP7_75t_L g722 ( .A(n_723), .B(n_725), .C(n_727), .D(n_729), .Y(n_722) );
INVx3_ASAP7_75t_L g749 ( .A(n_728), .Y(n_749) );
INVx2_ASAP7_75t_L g1031 ( .A(n_730), .Y(n_1031) );
NAND4xp25_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .C(n_735), .D(n_737), .Y(n_731) );
BUFx2_ASAP7_75t_L g879 ( .A(n_734), .Y(n_879) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
AND2x2_ASAP7_75t_L g743 ( .A(n_744), .B(n_760), .Y(n_743) );
NOR3xp33_ASAP7_75t_L g744 ( .A(n_745), .B(n_751), .C(n_756), .Y(n_744) );
NAND2xp5_ASAP7_75t_SL g745 ( .A(n_746), .B(n_750), .Y(n_745) );
NOR2xp33_ASAP7_75t_SL g747 ( .A(n_748), .B(n_749), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_753), .B1(n_754), .B2(n_755), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g958 ( .A1(n_753), .A2(n_959), .B1(n_960), .B2(n_961), .Y(n_958) );
OAI22xp5_ASAP7_75t_L g981 ( .A1(n_753), .A2(n_961), .B1(n_982), .B2(n_983), .Y(n_981) );
OAI22xp5_ASAP7_75t_L g963 ( .A1(n_755), .A2(n_964), .B1(n_965), .B2(n_966), .Y(n_963) );
AND4x1_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .C(n_763), .D(n_764), .Y(n_760) );
INVx1_ASAP7_75t_L g1047 ( .A(n_767), .Y(n_1047) );
XNOR2xp5_ASAP7_75t_L g767 ( .A(n_768), .B(n_926), .Y(n_767) );
AOI22xp5_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_850), .B1(n_924), .B2(n_925), .Y(n_768) );
INVx1_ASAP7_75t_L g924 ( .A(n_769), .Y(n_924) );
AOI22xp5_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_829), .B1(n_848), .B2(n_849), .Y(n_769) );
INVx2_ASAP7_75t_SL g849 ( .A(n_770), .Y(n_849) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
XNOR2xp5_ASAP7_75t_L g771 ( .A(n_772), .B(n_795), .Y(n_771) );
OAI21x1_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_774), .B(n_792), .Y(n_772) );
AND2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_783), .Y(n_774) );
NAND3xp33_ASAP7_75t_L g792 ( .A(n_775), .B(n_793), .C(n_794), .Y(n_792) );
AND4x1_ASAP7_75t_L g775 ( .A(n_776), .B(n_777), .C(n_780), .D(n_781), .Y(n_775) );
NOR2xp33_ASAP7_75t_L g783 ( .A(n_784), .B(n_789), .Y(n_783) );
INVxp67_ASAP7_75t_SL g794 ( .A(n_784), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_785), .B(n_787), .Y(n_784) );
BUFx2_ASAP7_75t_L g877 ( .A(n_786), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
INVx1_ASAP7_75t_L g972 ( .A(n_795), .Y(n_972) );
NAND2x1_ASAP7_75t_L g795 ( .A(n_796), .B(n_822), .Y(n_795) );
NOR3xp33_ASAP7_75t_L g796 ( .A(n_797), .B(n_803), .C(n_809), .Y(n_796) );
OAI22xp33_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_799), .B1(n_800), .B2(n_1300), .Y(n_797) );
INVx1_ASAP7_75t_L g827 ( .A(n_798), .Y(n_827) );
NOR2xp67_ASAP7_75t_L g803 ( .A(n_799), .B(n_804), .Y(n_803) );
OAI22xp5_ASAP7_75t_L g809 ( .A1(n_799), .A2(n_810), .B1(n_811), .B2(n_1301), .Y(n_809) );
INVx1_ASAP7_75t_L g824 ( .A(n_800), .Y(n_824) );
INVx1_ASAP7_75t_L g943 ( .A(n_801), .Y(n_943) );
INVx1_ASAP7_75t_L g991 ( .A(n_801), .Y(n_991) );
NAND3xp33_ASAP7_75t_L g822 ( .A(n_804), .B(n_823), .C(n_826), .Y(n_822) );
AND2x2_ASAP7_75t_L g804 ( .A(n_805), .B(n_808), .Y(n_804) );
BUFx4f_ASAP7_75t_L g1044 ( .A(n_806), .Y(n_1044) );
INVx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g841 ( .A(n_807), .Y(n_841) );
INVx1_ASAP7_75t_L g828 ( .A(n_810), .Y(n_828) );
INVx1_ASAP7_75t_L g825 ( .A(n_811), .Y(n_825) );
NOR2x1_ASAP7_75t_L g811 ( .A(n_812), .B(n_817), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_813), .A2(n_814), .B1(n_815), .B2(n_816), .Y(n_812) );
OAI22xp5_ASAP7_75t_L g817 ( .A1(n_818), .A2(n_819), .B1(n_820), .B2(n_821), .Y(n_817) );
NOR2xp33_ASAP7_75t_L g823 ( .A(n_824), .B(n_825), .Y(n_823) );
HB1xp67_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g848 ( .A(n_830), .Y(n_848) );
HB1xp67_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
XNOR2x1_ASAP7_75t_L g832 ( .A(n_833), .B(n_834), .Y(n_832) );
NOR2x1_ASAP7_75t_L g834 ( .A(n_835), .B(n_842), .Y(n_834) );
NAND4xp25_ASAP7_75t_SL g835 ( .A(n_836), .B(n_837), .C(n_838), .D(n_840), .Y(n_835) );
NAND3xp33_ASAP7_75t_L g842 ( .A(n_843), .B(n_846), .C(n_847), .Y(n_842) );
INVx2_ASAP7_75t_SL g925 ( .A(n_850), .Y(n_925) );
AO22x2_ASAP7_75t_L g850 ( .A1(n_851), .A2(n_852), .B1(n_881), .B2(n_923), .Y(n_850) );
INVx2_ASAP7_75t_SL g851 ( .A(n_852), .Y(n_851) );
XNOR2x1_ASAP7_75t_L g852 ( .A(n_853), .B(n_854), .Y(n_852) );
OR2x2_ASAP7_75t_L g854 ( .A(n_855), .B(n_870), .Y(n_854) );
NAND3xp33_ASAP7_75t_SL g855 ( .A(n_856), .B(n_859), .C(n_862), .Y(n_855) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
OAI21xp33_ASAP7_75t_L g967 ( .A1(n_864), .A2(n_968), .B(n_969), .Y(n_967) );
INVx2_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
OAI21xp33_ASAP7_75t_L g866 ( .A1(n_867), .A2(n_868), .B(n_869), .Y(n_866) );
NAND4xp25_ASAP7_75t_L g870 ( .A(n_871), .B(n_875), .C(n_878), .D(n_880), .Y(n_870) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g923 ( .A(n_881), .Y(n_923) );
XNOR2xp5_ASAP7_75t_L g881 ( .A(n_882), .B(n_896), .Y(n_881) );
INVx3_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
XNOR2x1_ASAP7_75t_L g883 ( .A(n_884), .B(n_885), .Y(n_883) );
OR2x2_ASAP7_75t_L g885 ( .A(n_886), .B(n_891), .Y(n_885) );
NAND4xp25_ASAP7_75t_L g886 ( .A(n_887), .B(n_888), .C(n_889), .D(n_890), .Y(n_886) );
NAND4xp25_ASAP7_75t_L g891 ( .A(n_892), .B(n_893), .C(n_894), .D(n_895), .Y(n_891) );
NAND2xp5_ASAP7_75t_SL g896 ( .A(n_897), .B(n_916), .Y(n_896) );
AOI21x1_ASAP7_75t_L g897 ( .A1(n_898), .A2(n_899), .B(n_910), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_900), .B(n_905), .Y(n_899) );
BUFx2_ASAP7_75t_L g917 ( .A(n_900), .Y(n_917) );
INVx2_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
NOR2xp33_ASAP7_75t_L g905 ( .A(n_906), .B(n_909), .Y(n_905) );
INVxp67_ASAP7_75t_SL g906 ( .A(n_907), .Y(n_906) );
AND2x2_ASAP7_75t_L g921 ( .A(n_907), .B(n_914), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_909), .Y(n_922) );
INVx1_ASAP7_75t_L g920 ( .A(n_911), .Y(n_920) );
AND2x2_ASAP7_75t_L g911 ( .A(n_912), .B(n_913), .Y(n_911) );
NAND4xp75_ASAP7_75t_L g916 ( .A(n_917), .B(n_918), .C(n_921), .D(n_922), .Y(n_916) );
NOR2x1_ASAP7_75t_L g918 ( .A(n_919), .B(n_920), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g926 ( .A1(n_927), .A2(n_928), .B1(n_973), .B2(n_974), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
AOI22x1_ASAP7_75t_L g928 ( .A1(n_929), .A2(n_930), .B1(n_970), .B2(n_971), .Y(n_928) );
INVx2_ASAP7_75t_SL g929 ( .A(n_930), .Y(n_929) );
XOR2x2_ASAP7_75t_L g930 ( .A(n_931), .B(n_949), .Y(n_930) );
XOR2x2_ASAP7_75t_L g931 ( .A(n_932), .B(n_948), .Y(n_931) );
NOR2x1_ASAP7_75t_L g932 ( .A(n_933), .B(n_938), .Y(n_932) );
NAND4xp25_ASAP7_75t_L g933 ( .A(n_934), .B(n_935), .C(n_936), .D(n_937), .Y(n_933) );
NAND3xp33_ASAP7_75t_L g938 ( .A(n_939), .B(n_941), .C(n_947), .Y(n_938) );
INVx1_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
XNOR2x1_ASAP7_75t_L g949 ( .A(n_950), .B(n_951), .Y(n_949) );
AND2x2_ASAP7_75t_L g951 ( .A(n_952), .B(n_957), .Y(n_951) );
AND4x1_ASAP7_75t_L g952 ( .A(n_953), .B(n_954), .C(n_955), .D(n_956), .Y(n_952) );
NOR3xp33_ASAP7_75t_L g957 ( .A(n_958), .B(n_963), .C(n_967), .Y(n_957) );
INVx2_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
INVx2_ASAP7_75t_SL g987 ( .A(n_965), .Y(n_987) );
INVx2_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
BUFx3_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
INVx1_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
XNOR2xp5_ASAP7_75t_L g974 ( .A(n_975), .B(n_1000), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_976), .Y(n_975) );
HB1xp67_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
XNOR2x1_ASAP7_75t_L g977 ( .A(n_978), .B(n_979), .Y(n_977) );
NAND2x1_ASAP7_75t_L g979 ( .A(n_980), .B(n_993), .Y(n_979) );
NOR3xp33_ASAP7_75t_SL g980 ( .A(n_981), .B(n_984), .C(n_989), .Y(n_980) );
INVx2_ASAP7_75t_L g986 ( .A(n_987), .Y(n_986) );
OAI21xp5_ASAP7_75t_L g989 ( .A1(n_990), .A2(n_991), .B(n_992), .Y(n_989) );
NOR2x1_ASAP7_75t_L g993 ( .A(n_994), .B(n_997), .Y(n_993) );
NAND2xp5_ASAP7_75t_L g994 ( .A(n_995), .B(n_996), .Y(n_994) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_998), .B(n_999), .Y(n_997) );
OAI22xp33_ASAP7_75t_SL g1000 ( .A1(n_1001), .A2(n_1020), .B1(n_1021), .B2(n_1046), .Y(n_1000) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1001), .Y(n_1046) );
INVx1_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
INVx1_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
XNOR2x1_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1005), .Y(n_1003) );
NAND4xp75_ASAP7_75t_L g1005 ( .A(n_1006), .B(n_1009), .C(n_1013), .D(n_1016), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_1007), .B(n_1008), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1012), .Y(n_1009) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1015), .Y(n_1013) );
NOR2xp33_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1019), .Y(n_1017) );
INVx1_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
NAND2x1_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1040), .Y(n_1022) );
NOR3xp33_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1029), .C(n_1034), .Y(n_1023) );
OAI21xp5_ASAP7_75t_L g1024 ( .A1(n_1025), .A2(n_1026), .B(n_1028), .Y(n_1024) );
INVx2_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
OAI22xp5_ASAP7_75t_L g1029 ( .A1(n_1030), .A2(n_1031), .B1(n_1032), .B2(n_1033), .Y(n_1029) );
OAI22xp33_ASAP7_75t_L g1034 ( .A1(n_1035), .A2(n_1036), .B1(n_1038), .B2(n_1039), .Y(n_1034) );
INVx2_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
AND4x1_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1042), .C(n_1043), .D(n_1045), .Y(n_1040) );
OAI221xp5_ASAP7_75t_L g1048 ( .A1(n_1049), .A2(n_1264), .B1(n_1266), .B2(n_1283), .C(n_1287), .Y(n_1048) );
AND5x1_ASAP7_75t_L g1049 ( .A(n_1050), .B(n_1200), .C(n_1229), .D(n_1244), .E(n_1251), .Y(n_1049) );
AOI211xp5_ASAP7_75t_L g1050 ( .A1(n_1051), .A2(n_1068), .B(n_1159), .C(n_1176), .Y(n_1050) );
NOR2xp33_ASAP7_75t_L g1162 ( .A(n_1051), .B(n_1095), .Y(n_1162) );
CKINVDCx5p33_ASAP7_75t_R g1195 ( .A(n_1051), .Y(n_1195) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_1052), .B(n_1064), .Y(n_1051) );
HB1xp67_ASAP7_75t_L g1265 ( .A(n_1053), .Y(n_1265) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
INVx3_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
AND2x4_ASAP7_75t_L g1055 ( .A(n_1056), .B(n_1058), .Y(n_1055) );
AND2x4_ASAP7_75t_L g1065 ( .A(n_1056), .B(n_1066), .Y(n_1065) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1056), .B(n_1066), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_1056), .B(n_1066), .Y(n_1091) );
AND2x4_ASAP7_75t_L g1062 ( .A(n_1058), .B(n_1063), .Y(n_1062) );
AND2x4_ASAP7_75t_L g1073 ( .A(n_1058), .B(n_1063), .Y(n_1073) );
INVx2_ASAP7_75t_L g1060 ( .A(n_1061), .Y(n_1060) );
INVx2_ASAP7_75t_SL g1061 ( .A(n_1062), .Y(n_1061) );
AND2x4_ASAP7_75t_L g1067 ( .A(n_1063), .B(n_1066), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1063), .B(n_1066), .Y(n_1076) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_1063), .B(n_1066), .Y(n_1081) );
NAND5xp2_ASAP7_75t_L g1068 ( .A(n_1069), .B(n_1126), .C(n_1137), .D(n_1141), .E(n_1154), .Y(n_1068) );
AOI21xp5_ASAP7_75t_L g1069 ( .A1(n_1070), .A2(n_1092), .B(n_1103), .Y(n_1069) );
OAI21xp5_ASAP7_75t_L g1174 ( .A1(n_1070), .A2(n_1140), .B(n_1175), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1077), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_1071), .B(n_1113), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_1071), .B(n_1120), .Y(n_1119) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_1071), .B(n_1086), .Y(n_1125) );
CKINVDCx6p67_ASAP7_75t_R g1129 ( .A(n_1071), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1071), .B(n_1118), .Y(n_1136) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_1071), .B(n_1146), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1071), .B(n_1145), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1071), .B(n_1083), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1071), .B(n_1155), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_1072), .B(n_1074), .Y(n_1071) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1077), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1083), .Y(n_1077) );
INVx3_ASAP7_75t_L g1120 ( .A(n_1078), .Y(n_1120) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_1078), .B(n_1157), .Y(n_1156) );
INVx3_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
NAND2xp5_ASAP7_75t_L g1111 ( .A(n_1079), .B(n_1112), .Y(n_1111) );
INVx2_ASAP7_75t_L g1124 ( .A(n_1079), .Y(n_1124) );
INVx2_ASAP7_75t_L g1135 ( .A(n_1079), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1079), .B(n_1129), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1181 ( .A(n_1079), .B(n_1158), .Y(n_1181) );
NOR2xp33_ASAP7_75t_L g1216 ( .A(n_1079), .B(n_1108), .Y(n_1216) );
NAND2xp5_ASAP7_75t_L g1238 ( .A(n_1079), .B(n_1115), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1082), .Y(n_1079) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1083), .Y(n_1148) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1083), .B(n_1129), .Y(n_1197) );
NAND2xp5_ASAP7_75t_L g1220 ( .A(n_1083), .B(n_1169), .Y(n_1220) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_1084), .B(n_1086), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_1084), .B(n_1113), .Y(n_1118) );
OR2x2_ASAP7_75t_L g1131 ( .A(n_1084), .B(n_1086), .Y(n_1131) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1084), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1084), .B(n_1129), .Y(n_1185) );
INVx1_ASAP7_75t_L g1113 ( .A(n_1086), .Y(n_1113) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1086), .B(n_1146), .Y(n_1145) );
AOI31xp33_ASAP7_75t_L g1236 ( .A1(n_1086), .A2(n_1186), .A3(n_1237), .B(n_1239), .Y(n_1236) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_1087), .B(n_1090), .Y(n_1086) );
NAND2xp5_ASAP7_75t_L g1242 ( .A(n_1092), .B(n_1223), .Y(n_1242) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
NOR3xp33_ASAP7_75t_L g1259 ( .A(n_1093), .B(n_1117), .C(n_1166), .Y(n_1259) );
OR2x2_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1098), .Y(n_1093) );
NOR2xp33_ASAP7_75t_L g1142 ( .A(n_1094), .B(n_1133), .Y(n_1142) );
INVx2_ASAP7_75t_L g1186 ( .A(n_1094), .Y(n_1186) );
NOR2xp33_ASAP7_75t_L g1194 ( .A(n_1094), .B(n_1195), .Y(n_1194) );
AND2x2_ASAP7_75t_L g1230 ( .A(n_1094), .B(n_1099), .Y(n_1230) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_1094), .B(n_1172), .Y(n_1256) );
INVx4_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_1095), .B(n_1106), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_1095), .B(n_1139), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_1095), .B(n_1100), .Y(n_1153) );
NAND3xp33_ASAP7_75t_L g1243 ( .A(n_1095), .B(n_1145), .C(n_1216), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1097), .Y(n_1095) );
INVxp67_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_1099), .B(n_1108), .Y(n_1115) );
OR2x2_ASAP7_75t_L g1140 ( .A(n_1099), .B(n_1107), .Y(n_1140) );
OR2x2_ASAP7_75t_L g1158 ( .A(n_1099), .B(n_1108), .Y(n_1158) );
INVx2_ASAP7_75t_L g1172 ( .A(n_1099), .Y(n_1172) );
INVx2_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
OR2x2_ASAP7_75t_L g1133 ( .A(n_1100), .B(n_1108), .Y(n_1133) );
NAND2xp5_ASAP7_75t_L g1100 ( .A(n_1101), .B(n_1102), .Y(n_1100) );
OAI211xp5_ASAP7_75t_SL g1103 ( .A1(n_1104), .A2(n_1111), .B(n_1114), .C(n_1121), .Y(n_1103) );
A2O1A1O1Ixp25_ASAP7_75t_L g1231 ( .A1(n_1104), .A2(n_1211), .B(n_1232), .C(n_1233), .D(n_1236), .Y(n_1231) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1105), .Y(n_1104) );
AOI211xp5_ASAP7_75t_L g1222 ( .A1(n_1106), .A2(n_1170), .B(n_1211), .C(n_1223), .Y(n_1222) );
INVx2_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1107), .Y(n_1152) );
INVx4_ASAP7_75t_L g1107 ( .A(n_1108), .Y(n_1107) );
NAND2xp5_ASAP7_75t_L g1123 ( .A(n_1108), .B(n_1124), .Y(n_1123) );
NOR2xp33_ASAP7_75t_L g1263 ( .A(n_1108), .B(n_1124), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1109), .B(n_1110), .Y(n_1108) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1113), .B(n_1129), .Y(n_1199) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_1115), .B(n_1116), .Y(n_1114) );
AOI22xp5_ASAP7_75t_L g1126 ( .A1(n_1115), .A2(n_1127), .B1(n_1132), .B2(n_1134), .Y(n_1126) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1115), .Y(n_1175) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
NAND2xp5_ASAP7_75t_L g1117 ( .A(n_1118), .B(n_1119), .Y(n_1117) );
NAND2xp5_ASAP7_75t_L g1137 ( .A(n_1118), .B(n_1138), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1118), .B(n_1169), .Y(n_1168) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1118), .Y(n_1180) );
AOI322xp5_ASAP7_75t_L g1177 ( .A1(n_1119), .A2(n_1132), .A3(n_1136), .B1(n_1156), .B2(n_1178), .C1(n_1181), .C2(n_1182), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_1119), .B(n_1155), .Y(n_1254) );
NOR2x1_ASAP7_75t_L g1130 ( .A(n_1120), .B(n_1131), .Y(n_1130) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_1120), .B(n_1145), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1120), .B(n_1226), .Y(n_1225) );
NOR2x1_ASAP7_75t_L g1247 ( .A(n_1120), .B(n_1227), .Y(n_1247) );
NAND2xp5_ASAP7_75t_L g1121 ( .A(n_1122), .B(n_1125), .Y(n_1121) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1124), .B(n_1185), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1124), .B(n_1235), .Y(n_1234) );
NAND2xp5_ASAP7_75t_L g1241 ( .A(n_1125), .B(n_1135), .Y(n_1241) );
NAND2xp5_ASAP7_75t_L g1249 ( .A(n_1127), .B(n_1250), .Y(n_1249) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
NOR2xp33_ASAP7_75t_L g1201 ( .A(n_1128), .B(n_1202), .Y(n_1201) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_1129), .B(n_1130), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1129), .B(n_1155), .Y(n_1192) );
NAND2xp5_ASAP7_75t_L g1227 ( .A(n_1129), .B(n_1145), .Y(n_1227) );
NAND2xp5_ASAP7_75t_L g1262 ( .A(n_1129), .B(n_1146), .Y(n_1262) );
OAI21xp5_ASAP7_75t_L g1228 ( .A1(n_1130), .A2(n_1132), .B(n_1226), .Y(n_1228) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1131), .Y(n_1155) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1133), .Y(n_1132) );
AND2x2_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1136), .Y(n_1134) );
NOR2xp33_ASAP7_75t_L g1147 ( .A(n_1135), .B(n_1148), .Y(n_1147) );
NOR2xp33_ASAP7_75t_L g1198 ( .A(n_1135), .B(n_1199), .Y(n_1198) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1136), .Y(n_1160) );
OAI21xp5_ASAP7_75t_L g1196 ( .A1(n_1138), .A2(n_1197), .B(n_1198), .Y(n_1196) );
NAND2xp5_ASAP7_75t_L g1207 ( .A(n_1139), .B(n_1208), .Y(n_1207) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g1141 ( .A1(n_1142), .A2(n_1143), .B1(n_1147), .B2(n_1149), .Y(n_1141) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
OAI21xp33_ASAP7_75t_L g1252 ( .A1(n_1144), .A2(n_1211), .B(n_1253), .Y(n_1252) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1145), .Y(n_1179) );
OAI211xp5_ASAP7_75t_L g1260 ( .A1(n_1145), .A2(n_1162), .B(n_1261), .C(n_1263), .Y(n_1260) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1147), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1150), .B(n_1153), .Y(n_1149) );
HB1xp67_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1151), .Y(n_1167) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1152), .Y(n_1190) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1153), .Y(n_1240) );
AOI221xp5_ASAP7_75t_L g1251 ( .A1(n_1153), .A2(n_1247), .B1(n_1252), .B2(n_1255), .C(n_1257), .Y(n_1251) );
NAND2xp5_ASAP7_75t_L g1154 ( .A(n_1155), .B(n_1156), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1155), .B(n_1169), .Y(n_1173) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
OAI22xp5_ASAP7_75t_L g1163 ( .A1(n_1158), .A2(n_1164), .B1(n_1170), .B2(n_1173), .Y(n_1163) );
O2A1O1Ixp33_ASAP7_75t_SL g1159 ( .A1(n_1160), .A2(n_1161), .B(n_1163), .C(n_1174), .Y(n_1159) );
NOR2xp33_ASAP7_75t_L g1214 ( .A(n_1160), .B(n_1215), .Y(n_1214) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
OAI211xp5_ASAP7_75t_L g1209 ( .A1(n_1165), .A2(n_1171), .B(n_1210), .C(n_1211), .Y(n_1209) );
NAND2xp5_ASAP7_75t_L g1165 ( .A(n_1166), .B(n_1168), .Y(n_1165) );
HB1xp67_ASAP7_75t_L g1202 ( .A(n_1166), .Y(n_1202) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1167), .Y(n_1166) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1167), .Y(n_1219) );
O2A1O1Ixp33_ASAP7_75t_L g1229 ( .A1(n_1168), .A2(n_1201), .B(n_1230), .C(n_1231), .Y(n_1229) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
INVx3_ASAP7_75t_SL g1171 ( .A(n_1172), .Y(n_1171) );
OAI221xp5_ASAP7_75t_L g1203 ( .A1(n_1172), .A2(n_1175), .B1(n_1204), .B2(n_1206), .C(n_1207), .Y(n_1203) );
NAND2xp5_ASAP7_75t_L g1221 ( .A(n_1172), .B(n_1195), .Y(n_1221) );
NOR4xp25_ASAP7_75t_L g1213 ( .A(n_1173), .B(n_1214), .C(n_1217), .D(n_1221), .Y(n_1213) );
OAI221xp5_ASAP7_75t_L g1176 ( .A1(n_1177), .A2(n_1186), .B1(n_1187), .B2(n_1193), .C(n_1196), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1180), .Y(n_1178) );
NAND2xp5_ASAP7_75t_L g1182 ( .A(n_1183), .B(n_1184), .Y(n_1182) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1185), .Y(n_1184) );
A2O1A1Ixp33_ASAP7_75t_SL g1244 ( .A1(n_1186), .A2(n_1245), .B(n_1247), .C(n_1248), .Y(n_1244) );
INVxp67_ASAP7_75t_SL g1187 ( .A(n_1188), .Y(n_1187) );
NOR2xp33_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1191), .Y(n_1188) );
OAI221xp5_ASAP7_75t_L g1212 ( .A1(n_1189), .A2(n_1213), .B1(n_1222), .B2(n_1224), .C(n_1228), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g1253 ( .A(n_1189), .B(n_1254), .Y(n_1253) );
INVx2_ASAP7_75t_L g1189 ( .A(n_1190), .Y(n_1189) );
HB1xp67_ASAP7_75t_L g1246 ( .A(n_1190), .Y(n_1246) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
NOR2xp33_ASAP7_75t_L g1204 ( .A(n_1192), .B(n_1205), .Y(n_1204) );
OAI311xp33_ASAP7_75t_L g1200 ( .A1(n_1193), .A2(n_1201), .A3(n_1203), .B1(n_1209), .C1(n_1212), .Y(n_1200) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
INVx2_ASAP7_75t_L g1211 ( .A(n_1195), .Y(n_1211) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1197), .Y(n_1206) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1216), .Y(n_1215) );
NOR2xp33_ASAP7_75t_L g1217 ( .A(n_1218), .B(n_1220), .Y(n_1217) );
HB1xp67_ASAP7_75t_L g1250 ( .A(n_1218), .Y(n_1250) );
HB1xp67_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1227), .Y(n_1226) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
OAI211xp5_ASAP7_75t_L g1239 ( .A1(n_1240), .A2(n_1241), .B(n_1242), .C(n_1243), .Y(n_1239) );
CKINVDCx16_ASAP7_75t_R g1245 ( .A(n_1246), .Y(n_1245) );
INVxp67_ASAP7_75t_L g1248 ( .A(n_1249), .Y(n_1248) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
NAND2xp5_ASAP7_75t_L g1257 ( .A(n_1258), .B(n_1260), .Y(n_1257) );
INVxp67_ASAP7_75t_L g1258 ( .A(n_1259), .Y(n_1258) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1262), .Y(n_1261) );
CKINVDCx20_ASAP7_75t_R g1264 ( .A(n_1265), .Y(n_1264) );
INVxp33_ASAP7_75t_SL g1266 ( .A(n_1267), .Y(n_1266) );
INVx2_ASAP7_75t_L g1267 ( .A(n_1268), .Y(n_1267) );
HB1xp67_ASAP7_75t_L g1290 ( .A(n_1269), .Y(n_1290) );
OR2x2_ASAP7_75t_L g1269 ( .A(n_1270), .B(n_1277), .Y(n_1269) );
NAND4xp25_ASAP7_75t_L g1270 ( .A(n_1271), .B(n_1272), .C(n_1274), .D(n_1275), .Y(n_1270) );
NAND4xp25_ASAP7_75t_L g1277 ( .A(n_1278), .B(n_1279), .C(n_1280), .D(n_1281), .Y(n_1277) );
CKINVDCx16_ASAP7_75t_R g1283 ( .A(n_1284), .Y(n_1283) );
INVxp67_ASAP7_75t_SL g1291 ( .A(n_1290), .Y(n_1291) );
BUFx2_ASAP7_75t_SL g1292 ( .A(n_1293), .Y(n_1292) );
BUFx2_ASAP7_75t_L g1294 ( .A(n_1295), .Y(n_1294) );
endmodule