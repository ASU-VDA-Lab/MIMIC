module real_jpeg_31176_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_0),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_0),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g201 ( 
.A(n_0),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_L g178 ( 
.A1(n_1),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_1),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_3),
.Y(n_74)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_4),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_4),
.Y(n_127)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_4),
.Y(n_131)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_4),
.Y(n_140)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

AO22x1_ASAP7_75t_SL g61 ( 
.A1(n_5),
.A2(n_56),
.B1(n_62),
.B2(n_64),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_5),
.A2(n_56),
.B1(n_136),
.B2(n_138),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_5),
.A2(n_56),
.B1(n_155),
.B2(n_158),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_5),
.B(n_239),
.Y(n_238)
);

OAI32xp33_ASAP7_75t_L g259 ( 
.A1(n_5),
.A2(n_260),
.A3(n_262),
.B1(n_265),
.B2(n_271),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_5),
.B(n_66),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_5),
.B(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_5),
.B(n_145),
.Y(n_325)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_6),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_6),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_6),
.Y(n_276)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_8),
.Y(n_149)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_8),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_9),
.A2(n_189),
.B1(n_190),
.B2(n_193),
.Y(n_188)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_9),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_9),
.A2(n_193),
.B1(n_365),
.B2(n_367),
.Y(n_364)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_10),
.Y(n_104)
);

AOI22x1_ASAP7_75t_L g44 ( 
.A1(n_11),
.A2(n_45),
.B1(n_47),
.B2(n_50),
.Y(n_44)
);

INVx2_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_11),
.A2(n_50),
.B1(n_125),
.B2(n_128),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_11),
.A2(n_50),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_348),
.Y(n_12)
);

INVxp67_ASAP7_75t_SL g13 ( 
.A(n_14),
.Y(n_13)
);

AOI21x1_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_247),
.B(n_344),
.Y(n_14)
);

INVxp33_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_226),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_17),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_213),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_18),
.B(n_213),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_141),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_19),
.B(n_375),
.C(n_376),
.Y(n_374)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

MAJx2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_59),
.C(n_98),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp33_ASAP7_75t_L g215 ( 
.A1(n_22),
.A2(n_23),
.B1(n_59),
.B2(n_216),
.Y(n_215)
);

AOI22x1_ASAP7_75t_L g373 ( 
.A1(n_22),
.A2(n_23),
.B1(n_219),
.B2(n_230),
.Y(n_373)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OA22x2_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_44),
.B1(n_51),
.B2(n_52),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_25),
.B(n_53),
.Y(n_208)
);

NOR2x1_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_34),
.Y(n_25)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_26),
.Y(n_239)
);

AO22x1_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_31),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

AOI22x1_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_38),
.B1(n_41),
.B2(n_42),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_40),
.Y(n_112)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_43),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_44),
.A2(n_51),
.B(n_208),
.Y(n_207)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_50),
.A2(n_84),
.B(n_87),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_88),
.Y(n_87)
);

INVxp33_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21x1_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_56),
.B(n_57),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_56),
.B(n_272),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_56),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_56),
.B(n_311),
.Y(n_310)
);

OAI32xp33_ASAP7_75t_L g99 ( 
.A1(n_57),
.A2(n_100),
.A3(n_105),
.B1(n_108),
.B2(n_110),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_59),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_59),
.A2(n_216),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

OA21x2_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_65),
.B(n_82),
.Y(n_59)
);

AOI21x1_ASAP7_75t_L g210 ( 
.A1(n_60),
.A2(n_65),
.B(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_61),
.B(n_90),
.Y(n_221)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_66),
.B(n_83),
.Y(n_220)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_91),
.Y(n_90)
);

AOI22x1_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_72),
.B1(n_75),
.B2(n_79),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_70),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_71),
.Y(n_160)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_81),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_81),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g369 ( 
.A(n_81),
.Y(n_369)
);

NAND2xp33_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_90),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_90),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_94),
.B1(n_95),
.B2(n_97),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_96),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_98),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_115),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_99),
.A2(n_115),
.B1(n_116),
.B2(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_99),
.Y(n_235)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_104),
.Y(n_261)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_113),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_114),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_115),
.B(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_116),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_116),
.B(n_325),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_116),
.B(n_325),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_124),
.B1(n_132),
.B2(n_135),
.Y(n_116)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_117),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_117),
.B(n_135),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_120),
.Y(n_281)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_123),
.Y(n_317)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_124),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_127),
.Y(n_185)
);

INVx6_ASAP7_75t_L g301 ( 
.A(n_127),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx4f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_131),
.Y(n_180)
);

INVx3_ASAP7_75t_SL g132 ( 
.A(n_133),
.Y(n_132)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_135),
.B(n_278),
.Y(n_277)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_196),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_142),
.Y(n_375)
);

OAI22x1_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_175),
.B1(n_176),
.B2(n_195),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_143),
.A2(n_195),
.B1(n_258),
.B2(n_338),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_144),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_144),
.B(n_291),
.Y(n_330)
);

NAND2x1_ASAP7_75t_L g372 ( 
.A(n_144),
.B(n_176),
.Y(n_372)
);

AO22x2_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_153),
.B1(n_161),
.B2(n_167),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_145),
.B(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2x1p5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_146),
.B(n_162),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_146),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_146),
.B(n_169),
.Y(n_225)
);

OA22x2_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_150),
.B2(n_151),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_152),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_153),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2x1_ASAP7_75t_L g204 ( 
.A(n_154),
.B(n_168),
.Y(n_204)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_156),
.A2(n_170),
.B1(n_172),
.B2(n_174),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_157),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_157),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_157),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_157),
.Y(n_366)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVxp33_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVxp67_ASAP7_75t_SL g167 ( 
.A(n_168),
.Y(n_167)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22x1_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_186),
.B1(n_188),
.B2(n_194),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_178),
.B(n_278),
.Y(n_358)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_185),
.Y(n_189)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_187),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_188),
.A2(n_199),
.B(n_202),
.Y(n_198)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_194),
.B(n_279),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_195),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_195),
.B(n_290),
.C(n_291),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_196),
.Y(n_376)
);

XNOR2x1_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_206),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_197),
.Y(n_355)
);

AND2x4_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_203),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_203),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx4_ASAP7_75t_SL g323 ( 
.A(n_201),
.Y(n_323)
);

OA21x2_ASAP7_75t_L g241 ( 
.A1(n_202),
.A2(n_242),
.B(n_244),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_203),
.A2(n_219),
.B1(n_230),
.B2(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_203),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_203),
.B(n_296),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_204),
.Y(n_362)
);

OA22x2_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_209),
.B1(n_210),
.B2(n_212),
.Y(n_206)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_207),
.Y(n_212)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_210),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_217),
.C(n_218),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_246),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_237),
.C(n_240),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_218),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_222),
.C(n_223),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_219),
.A2(n_223),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_219),
.Y(n_230)
);

AND2x4_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_222),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_223),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_245),
.Y(n_226)
);

NOR2x1_ASAP7_75t_L g346 ( 
.A(n_227),
.B(n_245),
.Y(n_346)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_234),
.C(n_236),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_251),
.Y(n_250)
);

XNOR2x1_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_232),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_230),
.B(n_332),
.C(n_341),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_232),
.B(n_354),
.C(n_355),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_236),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_237),
.A2(n_238),
.B1(n_240),
.B2(n_241),
.Y(n_256)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_240),
.B(n_295),
.Y(n_294)
);

NAND2xp33_ASAP7_75t_SL g327 ( 
.A(n_240),
.B(n_295),
.Y(n_327)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_241),
.B(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_282),
.B(n_343),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_250),
.B(n_252),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_257),
.C(n_258),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_253),
.A2(n_254),
.B1(n_337),
.B2(n_339),
.Y(n_336)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_258),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_277),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_259),
.B(n_277),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_261),
.Y(n_260)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

BUFx4f_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx3_ASAP7_75t_SL g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

AOI21x1_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_335),
.B(n_342),
.Y(n_282)
);

OAI21x1_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_292),
.B(n_334),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_289),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_285),
.B(n_289),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_286),
.Y(n_341)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_288),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_328),
.B(n_333),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_318),
.B(n_327),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_296),
.B(n_332),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_297),
.A2(n_302),
.B1(n_310),
.B2(n_315),
.Y(n_296)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_306),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g311 ( 
.A(n_312),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_315),
.B(n_321),
.Y(n_320)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_324),
.B(n_326),
.Y(n_318)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_331),
.Y(n_328)
);

NOR2xp67_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_331),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_340),
.Y(n_335)
);

NOR2xp67_ASAP7_75t_L g342 ( 
.A(n_336),
.B(n_340),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_337),
.Y(n_339)
);

NAND2xp33_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_347),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_377),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_374),
.Y(n_351)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_352),
.B(n_374),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_356),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_371),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_359),
.B1(n_360),
.B2(n_370),
.Y(n_357)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_358),
.Y(n_370)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_361),
.B(n_363),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);


endmodule