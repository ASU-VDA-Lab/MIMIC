module real_aes_7316_n_367 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_367);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_367;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_1066;
wire n_684;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_1106;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_1067;
wire n_518;
wire n_673;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_1114;
wire n_580;
wire n_577;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_1113;
wire n_766;
wire n_852;
wire n_974;
wire n_919;
wire n_857;
wire n_1089;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_1034;
wire n_549;
wire n_376;
wire n_571;
wire n_491;
wire n_923;
wire n_894;
wire n_694;
wire n_1123;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_551;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_955;
wire n_889;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_932;
wire n_948;
wire n_399;
wire n_700;
wire n_1046;
wire n_677;
wire n_958;
wire n_1021;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_1040;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1099;
wire n_709;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_966;
wire n_1108;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_892;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_578;
wire n_370;
wire n_994;
wire n_384;
wire n_744;
wire n_938;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_1053;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_369;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_755;
wire n_1025;
wire n_532;
wire n_656;
wire n_746;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_523;
wire n_860;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_1049;
wire n_796;
wire n_874;
wire n_801;
wire n_1126;
wire n_383;
wire n_529;
wire n_1115;
wire n_725;
wire n_455;
wire n_504;
wire n_973;
wire n_1081;
wire n_671;
wire n_960;
wire n_1084;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_1121;
wire n_885;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_1017;
wire n_737;
wire n_1013;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_1063;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_867;
wire n_745;
wire n_398;
wire n_1100;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_947;
wire n_561;
wire n_970;
wire n_876;
wire n_1112;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_733;
wire n_617;
wire n_658;
wire n_676;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1103;
wire n_1037;
wire n_1031;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_1041;
wire n_501;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_713;
wire n_598;
wire n_404;
wire n_728;
wire n_735;
wire n_756;
wire n_997;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1028;
wire n_1000;
wire n_1003;
wire n_727;
wire n_1014;
wire n_397;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_637;
wire n_526;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_1071;
wire n_787;
wire n_1052;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_1090;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_1045;
wire n_837;
wire n_967;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_1088;
wire n_988;
wire n_1055;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1097;
wire n_500;
wire n_601;
wire n_1101;
wire n_1076;
wire n_463;
wire n_661;
wire n_396;
wire n_804;
wire n_1102;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_1039;
wire n_802;
wire n_868;
wire n_877;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1024;
wire n_1104;
wire n_842;
wire n_1061;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_SL g954 ( .A1(n_0), .A2(n_55), .B1(n_563), .B2(n_955), .Y(n_954) );
AOI22xp33_ASAP7_75t_SL g1004 ( .A1(n_1), .A2(n_275), .B1(n_579), .B2(n_580), .Y(n_1004) );
CKINVDCx20_ASAP7_75t_R g635 ( .A(n_2), .Y(n_635) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_3), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_4), .Y(n_808) );
CKINVDCx20_ASAP7_75t_R g992 ( .A(n_5), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_6), .A2(n_131), .B1(n_489), .B2(n_871), .Y(n_870) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_7), .Y(n_507) );
AO22x2_ASAP7_75t_L g389 ( .A1(n_8), .A2(n_214), .B1(n_390), .B2(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g1089 ( .A(n_8), .Y(n_1089) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_9), .A2(n_152), .B1(n_582), .B2(n_618), .Y(n_617) );
CKINVDCx20_ASAP7_75t_R g1026 ( .A(n_10), .Y(n_1026) );
CKINVDCx20_ASAP7_75t_R g1060 ( .A(n_11), .Y(n_1060) );
CKINVDCx20_ASAP7_75t_R g639 ( .A(n_12), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_13), .A2(n_279), .B1(n_736), .B2(n_748), .Y(n_1005) );
CKINVDCx20_ASAP7_75t_R g1044 ( .A(n_14), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_15), .A2(n_101), .B1(n_618), .B2(n_1012), .Y(n_1011) );
CKINVDCx20_ASAP7_75t_R g933 ( .A(n_16), .Y(n_933) );
AOI222xp33_ASAP7_75t_L g956 ( .A1(n_17), .A2(n_49), .B1(n_141), .B2(n_387), .C1(n_469), .C2(n_957), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_18), .A2(n_51), .B1(n_597), .B2(n_598), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_19), .A2(n_239), .B1(n_495), .B2(n_496), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_20), .A2(n_149), .B1(n_425), .B2(n_429), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_21), .B(n_637), .Y(n_864) );
CKINVDCx20_ASAP7_75t_R g998 ( .A(n_22), .Y(n_998) );
CKINVDCx20_ASAP7_75t_R g918 ( .A(n_23), .Y(n_918) );
CKINVDCx20_ASAP7_75t_R g898 ( .A(n_24), .Y(n_898) );
AOI222xp33_ASAP7_75t_L g760 ( .A1(n_25), .A2(n_54), .B1(n_327), .B2(n_563), .C1(n_630), .C2(n_761), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g928 ( .A(n_26), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_27), .A2(n_118), .B1(n_538), .B2(n_540), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_28), .A2(n_52), .B1(n_458), .B2(n_843), .Y(n_842) );
CKINVDCx20_ASAP7_75t_R g974 ( .A(n_29), .Y(n_974) );
AO22x2_ASAP7_75t_L g393 ( .A1(n_30), .A2(n_107), .B1(n_390), .B2(n_394), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_31), .A2(n_357), .B1(n_546), .B2(n_548), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_32), .A2(n_240), .B1(n_540), .B2(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g778 ( .A(n_33), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_34), .A2(n_110), .B1(n_490), .B2(n_576), .Y(n_575) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_35), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g885 ( .A1(n_36), .A2(n_264), .B1(n_542), .B2(n_871), .Y(n_885) );
CKINVDCx20_ASAP7_75t_R g863 ( .A(n_37), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_38), .B(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_39), .B(n_509), .Y(n_835) );
CKINVDCx20_ASAP7_75t_R g838 ( .A(n_40), .Y(n_838) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_41), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_42), .A2(n_282), .B1(n_402), .B2(n_407), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_43), .A2(n_320), .B1(n_695), .B2(n_786), .Y(n_785) );
AOI22xp5_ASAP7_75t_L g899 ( .A1(n_44), .A2(n_205), .B1(n_402), .B2(n_530), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_45), .B(n_413), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g632 ( .A(n_46), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g1051 ( .A(n_47), .Y(n_1051) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_48), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_50), .A2(n_119), .B1(n_1017), .B2(n_1020), .Y(n_1016) );
AOI22xp33_ASAP7_75t_SL g482 ( .A1(n_53), .A2(n_363), .B1(n_483), .B2(n_485), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_56), .A2(n_137), .B1(n_591), .B2(n_623), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_57), .A2(n_236), .B1(n_495), .B2(n_496), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_58), .A2(n_274), .B1(n_788), .B2(n_876), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_59), .B(n_637), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_60), .A2(n_103), .B1(n_447), .B2(n_675), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g854 ( .A1(n_61), .A2(n_855), .B1(n_878), .B2(n_879), .Y(n_854) );
INVx1_ASAP7_75t_L g878 ( .A(n_61), .Y(n_878) );
CKINVDCx20_ASAP7_75t_R g811 ( .A(n_62), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_63), .A2(n_329), .B1(n_495), .B2(n_496), .Y(n_845) );
CKINVDCx20_ASAP7_75t_R g1067 ( .A(n_64), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_65), .A2(n_288), .B1(n_788), .B2(n_791), .Y(n_787) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_66), .Y(n_771) );
AOI22xp33_ASAP7_75t_SL g488 ( .A1(n_67), .A2(n_179), .B1(n_489), .B2(n_491), .Y(n_488) );
INVx1_ASAP7_75t_L g1100 ( .A(n_68), .Y(n_1100) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_69), .A2(n_342), .B1(n_590), .B2(n_591), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_70), .A2(n_99), .B1(n_506), .B2(n_540), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g1108 ( .A1(n_71), .A2(n_326), .B1(n_485), .B2(n_591), .Y(n_1108) );
INVx1_ASAP7_75t_L g952 ( .A(n_72), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_73), .A2(n_94), .B1(n_980), .B2(n_982), .Y(n_979) );
AOI211xp5_ASAP7_75t_L g367 ( .A1(n_74), .A2(n_368), .B(n_377), .C(n_1091), .Y(n_367) );
AOI222xp33_ASAP7_75t_L g1068 ( .A1(n_75), .A2(n_268), .B1(n_325), .B2(n_630), .C1(n_637), .C2(n_1069), .Y(n_1068) );
NAND2xp5_ASAP7_75t_L g1030 ( .A(n_76), .B(n_957), .Y(n_1030) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_77), .A2(n_246), .B1(n_402), .B2(n_407), .Y(n_401) );
AOI22xp33_ASAP7_75t_SL g468 ( .A1(n_78), .A2(n_300), .B1(n_469), .B2(n_470), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_79), .A2(n_280), .B1(n_444), .B2(n_481), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g1032 ( .A(n_80), .Y(n_1032) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_81), .A2(n_202), .B1(n_470), .B2(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g882 ( .A(n_82), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_83), .A2(n_200), .B1(n_489), .B2(n_602), .Y(n_691) );
AO22x2_ASAP7_75t_L g399 ( .A1(n_84), .A2(n_241), .B1(n_390), .B2(n_391), .Y(n_399) );
INVx1_ASAP7_75t_L g1086 ( .A(n_84), .Y(n_1086) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_85), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_86), .A2(n_87), .B1(n_481), .B2(n_736), .Y(n_820) );
CKINVDCx20_ASAP7_75t_R g926 ( .A(n_88), .Y(n_926) );
AOI22xp5_ASAP7_75t_L g888 ( .A1(n_89), .A2(n_104), .B1(n_439), .B2(n_817), .Y(n_888) );
AOI22xp5_ASAP7_75t_L g995 ( .A1(n_90), .A2(n_219), .B1(n_403), .B2(n_407), .Y(n_995) );
OA22x2_ASAP7_75t_L g906 ( .A1(n_91), .A2(n_907), .B1(n_908), .B2(n_909), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_91), .Y(n_907) );
AOI22x1_ASAP7_75t_L g822 ( .A1(n_92), .A2(n_823), .B1(n_847), .B2(n_848), .Y(n_822) );
INVx1_ASAP7_75t_L g847 ( .A(n_92), .Y(n_847) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_93), .Y(n_522) );
INVx1_ASAP7_75t_L g641 ( .A(n_95), .Y(n_641) );
AOI221xp5_ASAP7_75t_L g1064 ( .A1(n_96), .A2(n_315), .B1(n_725), .B2(n_727), .C(n_1065), .Y(n_1064) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_97), .Y(n_812) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_98), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_100), .A2(n_175), .B1(n_429), .B2(n_755), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_102), .A2(n_348), .B1(n_543), .B2(n_604), .Y(n_603) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_105), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_106), .A2(n_142), .B1(n_458), .B2(n_459), .Y(n_457) );
INVx1_ASAP7_75t_L g1090 ( .A(n_107), .Y(n_1090) );
CKINVDCx20_ASAP7_75t_R g893 ( .A(n_108), .Y(n_893) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_109), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_111), .A2(n_208), .B1(n_459), .B2(n_548), .Y(n_680) );
CKINVDCx20_ASAP7_75t_R g1046 ( .A(n_112), .Y(n_1046) );
CKINVDCx20_ASAP7_75t_R g994 ( .A(n_113), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_114), .A2(n_278), .B1(n_444), .B2(n_447), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_115), .B(n_637), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_116), .A2(n_283), .B1(n_538), .B2(n_618), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_117), .A2(n_129), .B1(n_602), .B2(n_677), .Y(n_676) );
AOI22xp33_ASAP7_75t_SL g474 ( .A1(n_120), .A2(n_228), .B1(n_413), .B2(n_475), .Y(n_474) );
AOI22xp5_ASAP7_75t_L g1001 ( .A1(n_121), .A2(n_295), .B1(n_438), .B2(n_540), .Y(n_1001) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_122), .Y(n_510) );
AOI22xp33_ASAP7_75t_SL g729 ( .A1(n_123), .A2(n_168), .B1(n_425), .B2(n_730), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_124), .A2(n_201), .B1(n_484), .B2(n_485), .Y(n_1022) );
AOI22xp33_ASAP7_75t_SL g735 ( .A1(n_125), .A2(n_290), .B1(n_552), .B2(n_736), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_126), .A2(n_163), .B1(n_947), .B2(n_948), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_127), .A2(n_319), .B1(n_403), .B2(n_730), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g867 ( .A(n_128), .Y(n_867) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_130), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_132), .A2(n_316), .B1(n_590), .B2(n_733), .Y(n_746) );
AOI222xp33_ASAP7_75t_L g605 ( .A1(n_133), .A2(n_215), .B1(n_301), .B2(n_387), .C1(n_514), .C2(n_606), .Y(n_605) );
AOI22xp33_ASAP7_75t_SL g494 ( .A1(n_134), .A2(n_298), .B1(n_495), .B2(n_496), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_135), .A2(n_194), .B1(n_582), .B2(n_584), .Y(n_581) );
CKINVDCx20_ASAP7_75t_R g892 ( .A(n_136), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_138), .A2(n_191), .B1(n_542), .B2(n_543), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_139), .A2(n_232), .B1(n_576), .B2(n_944), .Y(n_943) );
AND2x6_ASAP7_75t_L g372 ( .A(n_140), .B(n_373), .Y(n_372) );
HB1xp67_ASAP7_75t_L g1083 ( .A(n_140), .Y(n_1083) );
AOI22xp33_ASAP7_75t_SL g478 ( .A1(n_143), .A2(n_160), .B1(n_479), .B2(n_481), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_144), .A2(n_229), .B1(n_489), .B2(n_675), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_145), .A2(n_166), .B1(n_444), .B2(n_549), .Y(n_819) );
INVx1_ASAP7_75t_L g670 ( .A(n_146), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_147), .A2(n_250), .B1(n_634), .B2(n_817), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_148), .A2(n_266), .B1(n_548), .B2(n_623), .Y(n_846) );
CKINVDCx20_ASAP7_75t_R g965 ( .A(n_150), .Y(n_965) );
AOI22xp5_ASAP7_75t_L g922 ( .A1(n_151), .A2(n_247), .B1(n_453), .B2(n_923), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_153), .A2(n_177), .B1(n_573), .B2(n_574), .Y(n_572) );
INVx1_ASAP7_75t_L g1121 ( .A(n_154), .Y(n_1121) );
AOI22xp5_ASAP7_75t_SL g1123 ( .A1(n_154), .A2(n_1093), .B1(n_1113), .B2(n_1121), .Y(n_1123) );
AOI22xp5_ASAP7_75t_L g886 ( .A1(n_155), .A2(n_294), .B1(n_549), .B2(n_584), .Y(n_886) );
NAND2xp5_ASAP7_75t_SL g726 ( .A(n_156), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g1096 ( .A(n_157), .Y(n_1096) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_158), .Y(n_709) );
AO22x2_ASAP7_75t_L g397 ( .A1(n_159), .A2(n_234), .B1(n_390), .B2(n_394), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g1087 ( .A(n_159), .B(n_1088), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_161), .A2(n_172), .B1(n_623), .B2(n_733), .Y(n_783) );
AOI22xp33_ASAP7_75t_SL g739 ( .A1(n_162), .A2(n_245), .B1(n_740), .B2(n_741), .Y(n_739) );
XNOR2x2_ASAP7_75t_L g586 ( .A(n_164), .B(n_587), .Y(n_586) );
CKINVDCx20_ASAP7_75t_R g1055 ( .A(n_165), .Y(n_1055) );
AOI22xp33_ASAP7_75t_SL g722 ( .A1(n_167), .A2(n_256), .B1(n_407), .B2(n_470), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g832 ( .A(n_169), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_170), .A2(n_178), .B1(n_786), .B2(n_942), .Y(n_941) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_171), .Y(n_400) );
CKINVDCx20_ASAP7_75t_R g966 ( .A(n_173), .Y(n_966) );
CKINVDCx20_ASAP7_75t_R g968 ( .A(n_174), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_176), .A2(n_309), .B1(n_459), .B2(n_582), .Y(n_592) );
CKINVDCx20_ASAP7_75t_R g991 ( .A(n_180), .Y(n_991) );
AOI22xp33_ASAP7_75t_SL g435 ( .A1(n_181), .A2(n_218), .B1(n_436), .B2(n_439), .Y(n_435) );
AOI22xp33_ASAP7_75t_SL g738 ( .A1(n_182), .A2(n_190), .B1(n_439), .B2(n_602), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g889 ( .A1(n_183), .A2(n_222), .B1(n_736), .B2(n_890), .Y(n_889) );
AOI22xp5_ASAP7_75t_L g765 ( .A1(n_184), .A2(n_766), .B1(n_792), .B2(n_793), .Y(n_765) );
INVx1_ASAP7_75t_L g792 ( .A(n_184), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_185), .A2(n_305), .B1(n_548), .B2(n_623), .Y(n_622) );
CKINVDCx20_ASAP7_75t_R g859 ( .A(n_186), .Y(n_859) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_187), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_188), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_189), .A2(n_351), .B1(n_736), .B2(n_748), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_192), .A2(n_281), .B1(n_493), .B2(n_748), .Y(n_924) );
AOI22xp33_ASAP7_75t_SL g452 ( .A1(n_193), .A2(n_289), .B1(n_453), .B2(n_454), .Y(n_452) );
AOI22xp33_ASAP7_75t_SL g732 ( .A1(n_195), .A2(n_340), .B1(n_546), .B2(n_733), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_196), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_197), .B(n_637), .Y(n_636) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_198), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g627 ( .A(n_199), .Y(n_627) );
CKINVDCx20_ASAP7_75t_R g660 ( .A(n_203), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_204), .A2(n_213), .B1(n_470), .B2(n_971), .Y(n_970) );
CKINVDCx20_ASAP7_75t_R g1057 ( .A(n_206), .Y(n_1057) );
XNOR2x2_ASAP7_75t_L g938 ( .A(n_207), .B(n_939), .Y(n_938) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_209), .A2(n_244), .B1(n_481), .B2(n_602), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_210), .A2(n_216), .B1(n_579), .B2(n_695), .Y(n_694) );
CKINVDCx20_ASAP7_75t_R g1066 ( .A(n_211), .Y(n_1066) );
CKINVDCx20_ASAP7_75t_R g861 ( .A(n_212), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_217), .A2(n_333), .B1(n_493), .B2(n_942), .Y(n_1110) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_220), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g1111 ( .A1(n_221), .A2(n_260), .B1(n_1017), .B2(n_1020), .Y(n_1111) );
OA22x2_ASAP7_75t_L g800 ( .A1(n_223), .A2(n_801), .B1(n_802), .B2(n_821), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_223), .Y(n_801) );
CKINVDCx20_ASAP7_75t_R g1028 ( .A(n_224), .Y(n_1028) );
CKINVDCx20_ASAP7_75t_R g828 ( .A(n_225), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_226), .A2(n_356), .B1(n_484), .B2(n_950), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_227), .B(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g376 ( .A(n_230), .Y(n_376) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_231), .A2(n_614), .B1(n_647), .B2(n_648), .Y(n_613) );
INVx1_ASAP7_75t_L g647 ( .A(n_231), .Y(n_647) );
CKINVDCx20_ASAP7_75t_R g1033 ( .A(n_233), .Y(n_1033) );
AOI22xp5_ASAP7_75t_L g984 ( .A1(n_235), .A2(n_243), .B1(n_538), .B2(n_788), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_237), .B(n_421), .Y(n_420) );
AOI22xp33_ASAP7_75t_SL g472 ( .A1(n_238), .A2(n_261), .B1(n_408), .B2(n_473), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_242), .A2(n_334), .B1(n_430), .B2(n_469), .Y(n_569) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_248), .A2(n_688), .B1(n_713), .B2(n_714), .Y(n_687) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_248), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g667 ( .A(n_249), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_251), .A2(n_292), .B1(n_453), .B2(n_496), .Y(n_679) );
CKINVDCx20_ASAP7_75t_R g913 ( .A(n_252), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_253), .A2(n_349), .B1(n_485), .B2(n_733), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_254), .B(n_566), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_255), .A2(n_355), .B1(n_543), .B2(n_740), .Y(n_978) );
AOI22xp5_ASAP7_75t_L g1040 ( .A1(n_257), .A2(n_1041), .B1(n_1071), .B2(n_1072), .Y(n_1040) );
CKINVDCx20_ASAP7_75t_R g1071 ( .A(n_257), .Y(n_1071) );
CKINVDCx20_ASAP7_75t_R g932 ( .A(n_258), .Y(n_932) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_259), .Y(n_805) );
OA22x2_ASAP7_75t_L g462 ( .A1(n_262), .A2(n_463), .B1(n_464), .B2(n_497), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_262), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g953 ( .A(n_263), .B(n_728), .Y(n_953) );
INVx1_ASAP7_75t_L g1099 ( .A(n_265), .Y(n_1099) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_267), .A2(n_291), .B1(n_551), .B2(n_552), .Y(n_550) );
INVx1_ASAP7_75t_L g1103 ( .A(n_269), .Y(n_1103) );
INVx1_ASAP7_75t_L g390 ( .A(n_270), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_270), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_271), .A2(n_353), .B1(n_540), .B2(n_817), .Y(n_985) );
CKINVDCx20_ASAP7_75t_R g919 ( .A(n_272), .Y(n_919) );
CKINVDCx20_ASAP7_75t_R g1029 ( .A(n_273), .Y(n_1029) );
AOI22xp5_ASAP7_75t_L g1092 ( .A1(n_276), .A2(n_1093), .B1(n_1112), .B2(n_1113), .Y(n_1092) );
INVx1_ASAP7_75t_L g1112 ( .A(n_276), .Y(n_1112) );
CKINVDCx20_ASAP7_75t_R g997 ( .A(n_277), .Y(n_997) );
CKINVDCx20_ASAP7_75t_R g657 ( .A(n_284), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g1063 ( .A(n_285), .Y(n_1063) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_286), .Y(n_553) );
INVx1_ASAP7_75t_L g626 ( .A(n_287), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_293), .B(n_566), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g912 ( .A(n_296), .Y(n_912) );
AOI22xp33_ASAP7_75t_SL g578 ( .A1(n_297), .A2(n_346), .B1(n_579), .B2(n_580), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_299), .A2(n_314), .B1(n_438), .B2(n_618), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_302), .A2(n_339), .B1(n_444), .B2(n_890), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_303), .A2(n_324), .B1(n_430), .B2(n_514), .Y(n_894) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_304), .Y(n_775) );
INVx1_ASAP7_75t_L g375 ( .A(n_306), .Y(n_375) );
INVx1_ASAP7_75t_L g779 ( .A(n_307), .Y(n_779) );
CKINVDCx20_ASAP7_75t_R g662 ( .A(n_308), .Y(n_662) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_310), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_311), .Y(n_742) );
INVx1_ASAP7_75t_L g373 ( .A(n_312), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_313), .A2(n_344), .B1(n_481), .B2(n_489), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_317), .A2(n_321), .B1(n_421), .B2(n_595), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_318), .A2(n_328), .B1(n_574), .B2(n_602), .Y(n_601) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_322), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g1101 ( .A(n_323), .B(n_957), .Y(n_1101) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_330), .Y(n_561) );
CKINVDCx20_ASAP7_75t_R g664 ( .A(n_331), .Y(n_664) );
INVx1_ASAP7_75t_L g986 ( .A(n_332), .Y(n_986) );
CKINVDCx20_ASAP7_75t_R g858 ( .A(n_335), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_336), .B(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g1097 ( .A(n_337), .Y(n_1097) );
CKINVDCx20_ASAP7_75t_R g973 ( .A(n_338), .Y(n_973) );
CKINVDCx20_ASAP7_75t_R g915 ( .A(n_341), .Y(n_915) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_343), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g1048 ( .A(n_345), .Y(n_1048) );
INVx1_ASAP7_75t_L g1006 ( .A(n_347), .Y(n_1006) );
CKINVDCx20_ASAP7_75t_R g585 ( .A(n_350), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_352), .B(n_470), .Y(n_776) );
CKINVDCx20_ASAP7_75t_R g1025 ( .A(n_354), .Y(n_1025) );
OA22x2_ASAP7_75t_SL g652 ( .A1(n_358), .A2(n_653), .B1(n_654), .B2(n_681), .Y(n_652) );
INVx1_ASAP7_75t_L g681 ( .A(n_358), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g1007 ( .A1(n_359), .A2(n_1008), .B1(n_1034), .B2(n_1035), .Y(n_1007) );
INVx1_ASAP7_75t_L g1034 ( .A(n_359), .Y(n_1034) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_360), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g866 ( .A(n_361), .Y(n_866) );
INVx1_ASAP7_75t_L g1104 ( .A(n_362), .Y(n_1104) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_364), .A2(n_366), .B1(n_582), .B2(n_843), .Y(n_1014) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_365), .Y(n_773) );
CKINVDCx20_ASAP7_75t_R g368 ( .A(n_369), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_370), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x4_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
HB1xp67_ASAP7_75t_L g1082 ( .A(n_373), .Y(n_1082) );
OAI21xp5_ASAP7_75t_L g1119 ( .A1(n_374), .A2(n_1081), .B(n_1120), .Y(n_1119) );
AND2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
AOI221xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_795), .B1(n_1076), .B2(n_1077), .C(n_1078), .Y(n_377) );
INVx1_ASAP7_75t_L g1076 ( .A(n_378), .Y(n_1076) );
XNOR2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_609), .Y(n_378) );
XNOR2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_499), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_382), .B1(n_462), .B2(n_498), .Y(n_380) );
INVx3_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
XOR2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_461), .Y(n_382) );
NAND2x1_ASAP7_75t_SL g383 ( .A(n_384), .B(n_433), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_385), .B(n_411), .Y(n_384) );
OAI21xp5_ASAP7_75t_SL g385 ( .A1(n_386), .A2(n_400), .B(n_401), .Y(n_385) );
OAI21xp5_ASAP7_75t_SL g466 ( .A1(n_386), .A2(n_467), .B(n_468), .Y(n_466) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_387), .Y(n_506) );
INVx4_ASAP7_75t_L g631 ( .A(n_387), .Y(n_631) );
INVx2_ASAP7_75t_L g704 ( .A(n_387), .Y(n_704) );
BUFx3_ASAP7_75t_L g897 ( .A(n_387), .Y(n_897) );
AND2x6_ASAP7_75t_L g387 ( .A(n_388), .B(n_395), .Y(n_387) );
AND2x4_ASAP7_75t_L g408 ( .A(n_388), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g645 ( .A(n_388), .Y(n_645) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_393), .Y(n_388) );
AND2x2_ASAP7_75t_L g406 ( .A(n_389), .B(n_397), .Y(n_406) );
INVx2_ASAP7_75t_L g419 ( .A(n_389), .Y(n_419) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g394 ( .A(n_392), .Y(n_394) );
OR2x2_ASAP7_75t_L g418 ( .A(n_393), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g423 ( .A(n_393), .B(n_419), .Y(n_423) );
INVx2_ASAP7_75t_L g428 ( .A(n_393), .Y(n_428) );
INVx1_ASAP7_75t_L g432 ( .A(n_393), .Y(n_432) );
AND2x6_ASAP7_75t_L g438 ( .A(n_395), .B(n_417), .Y(n_438) );
AND2x2_ASAP7_75t_L g446 ( .A(n_395), .B(n_442), .Y(n_446) );
AND2x4_ASAP7_75t_L g453 ( .A(n_395), .B(n_423), .Y(n_453) );
AND2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_398), .Y(n_395) );
AND2x2_ASAP7_75t_L g416 ( .A(n_396), .B(n_399), .Y(n_416) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g441 ( .A(n_397), .B(n_410), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_397), .B(n_399), .Y(n_450) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g405 ( .A(n_399), .Y(n_405) );
INVx1_ASAP7_75t_L g410 ( .A(n_399), .Y(n_410) );
BUFx4f_ASAP7_75t_SL g761 ( .A(n_402), .Y(n_761) );
BUFx12f_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_403), .Y(n_470) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_403), .Y(n_509) );
AND2x4_ASAP7_75t_L g403 ( .A(n_404), .B(n_406), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g427 ( .A(n_405), .B(n_428), .Y(n_427) );
AND2x4_ASAP7_75t_L g426 ( .A(n_406), .B(n_427), .Y(n_426) );
AND2x4_ASAP7_75t_L g430 ( .A(n_406), .B(n_431), .Y(n_430) );
NAND2x1p5_ASAP7_75t_L g533 ( .A(n_406), .B(n_534), .Y(n_533) );
BUFx2_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_408), .Y(n_514) );
BUFx2_ASAP7_75t_SL g563 ( .A(n_408), .Y(n_563) );
INVx1_ASAP7_75t_L g646 ( .A(n_409), .Y(n_646) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NAND3xp33_ASAP7_75t_L g411 ( .A(n_412), .B(n_420), .C(n_424), .Y(n_411) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g566 ( .A(n_414), .Y(n_566) );
INVx2_ASAP7_75t_L g595 ( .A(n_414), .Y(n_595) );
INVx5_ASAP7_75t_L g728 ( .A(n_414), .Y(n_728) );
INVx4_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
AND2x6_ASAP7_75t_L g422 ( .A(n_416), .B(n_423), .Y(n_422) );
AND2x4_ASAP7_75t_L g458 ( .A(n_416), .B(n_442), .Y(n_458) );
INVx1_ASAP7_75t_L g521 ( .A(n_416), .Y(n_521) );
NAND2x1p5_ASAP7_75t_L g526 ( .A(n_416), .B(n_423), .Y(n_526) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g520 ( .A(n_418), .B(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g442 ( .A(n_419), .B(n_428), .Y(n_442) );
BUFx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_SL g476 ( .A(n_422), .Y(n_476) );
BUFx4f_ASAP7_75t_L g568 ( .A(n_422), .Y(n_568) );
BUFx2_ASAP7_75t_L g725 ( .A(n_422), .Y(n_725) );
AND2x2_ASAP7_75t_L g456 ( .A(n_423), .B(n_441), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g1050 ( .A(n_423), .B(n_441), .Y(n_1050) );
INVx2_ASAP7_75t_L g663 ( .A(n_425), .Y(n_663) );
BUFx2_ASAP7_75t_L g971 ( .A(n_425), .Y(n_971) );
INVx4_ASAP7_75t_L g1070 ( .A(n_425), .Y(n_1070) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx4f_ASAP7_75t_SL g469 ( .A(n_426), .Y(n_469) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_426), .Y(n_530) );
BUFx2_ASAP7_75t_L g634 ( .A(n_426), .Y(n_634) );
BUFx6f_ASAP7_75t_L g755 ( .A(n_426), .Y(n_755) );
INVx1_ASAP7_75t_L g534 ( .A(n_428), .Y(n_534) );
BUFx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx2_ASAP7_75t_L g473 ( .A(n_430), .Y(n_473) );
INVx1_ASAP7_75t_L g599 ( .A(n_430), .Y(n_599) );
BUFx2_ASAP7_75t_L g730 ( .A(n_430), .Y(n_730) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OR2x6_ASAP7_75t_L g460 ( .A(n_432), .B(n_450), .Y(n_460) );
NOR2x1_ASAP7_75t_L g433 ( .A(n_434), .B(n_451), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_443), .Y(n_434) );
INVx1_ASAP7_75t_L g1013 ( .A(n_436), .Y(n_1013) );
HB1xp67_ASAP7_75t_L g1062 ( .A(n_436), .Y(n_1062) );
INVx5_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_437), .Y(n_480) );
INVx4_ASAP7_75t_L g573 ( .A(n_437), .Y(n_573) );
INVx1_ASAP7_75t_L g758 ( .A(n_437), .Y(n_758) );
INVx2_ASAP7_75t_L g942 ( .A(n_437), .Y(n_942) );
INVx11_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx11_ASAP7_75t_L g539 ( .A(n_438), .Y(n_539) );
BUFx3_ASAP7_75t_L g496 ( .A(n_439), .Y(n_496) );
BUFx3_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx3_ASAP7_75t_L g540 ( .A(n_440), .Y(n_540) );
BUFx3_ASAP7_75t_L g574 ( .A(n_440), .Y(n_574) );
BUFx3_ASAP7_75t_L g948 ( .A(n_440), .Y(n_948) );
AND2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_441), .B(n_442), .Y(n_936) );
AND2x4_ASAP7_75t_L g448 ( .A(n_442), .B(n_449), .Y(n_448) );
INVx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx3_ASAP7_75t_L g542 ( .A(n_445), .Y(n_542) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_446), .Y(n_490) );
BUFx2_ASAP7_75t_SL g604 ( .A(n_446), .Y(n_604) );
BUFx2_ASAP7_75t_SL g740 ( .A(n_446), .Y(n_740) );
BUFx2_ASAP7_75t_L g843 ( .A(n_447), .Y(n_843) );
BUFx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx3_ASAP7_75t_L g481 ( .A(n_448), .Y(n_481) );
BUFx2_ASAP7_75t_SL g543 ( .A(n_448), .Y(n_543) );
BUFx3_ASAP7_75t_L g576 ( .A(n_448), .Y(n_576) );
BUFx3_ASAP7_75t_L g677 ( .A(n_448), .Y(n_677) );
BUFx2_ASAP7_75t_SL g741 ( .A(n_448), .Y(n_741) );
BUFx2_ASAP7_75t_L g890 ( .A(n_448), .Y(n_890) );
AND2x2_ASAP7_75t_L g584 ( .A(n_449), .B(n_534), .Y(n_584) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_457), .Y(n_451) );
BUFx3_ASAP7_75t_L g495 ( .A(n_453), .Y(n_495) );
INVx6_ASAP7_75t_L g547 ( .A(n_453), .Y(n_547) );
BUFx3_ASAP7_75t_L g817 ( .A(n_453), .Y(n_817) );
BUFx3_ASAP7_75t_L g1019 ( .A(n_453), .Y(n_1019) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_454), .Y(n_591) );
INVx2_ASAP7_75t_L g981 ( .A(n_454), .Y(n_981) );
INVx4_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g484 ( .A(n_455), .Y(n_484) );
INVx5_ASAP7_75t_L g549 ( .A(n_455), .Y(n_549) );
INVx3_ASAP7_75t_L g580 ( .A(n_455), .Y(n_580) );
BUFx3_ASAP7_75t_L g734 ( .A(n_455), .Y(n_734) );
INVx1_ASAP7_75t_L g923 ( .A(n_455), .Y(n_923) );
INVx8_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx3_ASAP7_75t_L g493 ( .A(n_458), .Y(n_493) );
BUFx3_ASAP7_75t_L g551 ( .A(n_458), .Y(n_551) );
INVx2_ASAP7_75t_L g583 ( .A(n_458), .Y(n_583) );
BUFx3_ASAP7_75t_L g736 ( .A(n_458), .Y(n_736) );
BUFx6f_ASAP7_75t_L g790 ( .A(n_458), .Y(n_790) );
INVx1_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
INVx6_ASAP7_75t_SL g486 ( .A(n_460), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g810 ( .A1(n_460), .A2(n_644), .B1(n_811), .B2(n_812), .Y(n_810) );
INVx1_ASAP7_75t_L g982 ( .A(n_460), .Y(n_982) );
INVx1_ASAP7_75t_L g498 ( .A(n_462), .Y(n_498) );
INVx1_ASAP7_75t_SL g497 ( .A(n_464), .Y(n_497) );
NAND3x1_ASAP7_75t_L g464 ( .A(n_465), .B(n_477), .C(n_487), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_471), .Y(n_465) );
INVx1_ASAP7_75t_L g833 ( .A(n_469), .Y(n_833) );
INVx2_ASAP7_75t_L g607 ( .A(n_470), .Y(n_607) );
BUFx3_ASAP7_75t_L g637 ( .A(n_470), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_474), .Y(n_471) );
INVx1_ASAP7_75t_SL g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_482), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVxp67_ASAP7_75t_L g1052 ( .A(n_485), .Y(n_1052) );
BUFx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx2_ASAP7_75t_L g552 ( .A(n_486), .Y(n_552) );
BUFx4f_ASAP7_75t_SL g623 ( .A(n_486), .Y(n_623) );
BUFx2_ASAP7_75t_L g748 ( .A(n_486), .Y(n_748) );
BUFx2_ASAP7_75t_L g950 ( .A(n_486), .Y(n_950) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_494), .Y(n_487) );
BUFx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx3_ASAP7_75t_L g618 ( .A(n_490), .Y(n_618) );
BUFx6f_ASAP7_75t_L g947 ( .A(n_490), .Y(n_947) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g1059 ( .A1(n_492), .A2(n_1060), .B1(n_1061), .B2(n_1063), .Y(n_1059) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
BUFx2_ASAP7_75t_L g675 ( .A(n_493), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_501), .B1(n_554), .B2(n_555), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
XOR2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_553), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_535), .Y(n_502) );
NOR3xp33_ASAP7_75t_L g503 ( .A(n_504), .B(n_515), .C(n_527), .Y(n_503) );
OAI221xp5_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_507), .B1(n_508), .B2(n_510), .C(n_511), .Y(n_504) );
OAI21xp5_ASAP7_75t_L g560 ( .A1(n_505), .A2(n_561), .B(n_562), .Y(n_560) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_SL g831 ( .A(n_506), .Y(n_831) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx4f_ASAP7_75t_L g957 ( .A(n_509), .Y(n_957) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_517), .B1(n_522), .B2(n_523), .Y(n_515) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_519), .A2(n_525), .B1(n_626), .B2(n_627), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g1024 ( .A1(n_519), .A2(n_751), .B1(n_1025), .B2(n_1026), .Y(n_1024) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g659 ( .A(n_520), .Y(n_659) );
BUFx3_ASAP7_75t_L g770 ( .A(n_520), .Y(n_770) );
OAI221xp5_ASAP7_75t_L g891 ( .A1(n_520), .A2(n_525), .B1(n_892), .B2(n_893), .C(n_894), .Y(n_891) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_523), .A2(n_657), .B1(n_658), .B2(n_660), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_523), .A2(n_769), .B1(n_770), .B2(n_771), .Y(n_768) );
OAI22xp5_ASAP7_75t_L g857 ( .A1(n_523), .A2(n_827), .B1(n_858), .B2(n_859), .Y(n_857) );
OAI22xp5_ASAP7_75t_SL g911 ( .A1(n_523), .A2(n_827), .B1(n_912), .B2(n_913), .Y(n_911) );
OAI22xp5_ASAP7_75t_L g964 ( .A1(n_523), .A2(n_710), .B1(n_965), .B2(n_966), .Y(n_964) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
BUFx3_ASAP7_75t_L g712 ( .A(n_525), .Y(n_712) );
BUFx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g752 ( .A(n_526), .Y(n_752) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_529), .B1(n_531), .B2(n_532), .Y(n_527) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_530), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g836 ( .A1(n_532), .A2(n_671), .B1(n_837), .B2(n_838), .Y(n_836) );
OAI22xp33_ASAP7_75t_L g917 ( .A1(n_532), .A2(n_862), .B1(n_918), .B2(n_919), .Y(n_917) );
OAI22xp5_ASAP7_75t_L g1031 ( .A1(n_532), .A2(n_671), .B1(n_1032), .B2(n_1033), .Y(n_1031) );
BUFx3_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_533), .Y(n_640) );
INVx4_ASAP7_75t_L g669 ( .A(n_533), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g996 ( .A1(n_533), .A2(n_774), .B1(n_997), .B2(n_998), .Y(n_996) );
OAI22xp5_ASAP7_75t_L g1065 ( .A1(n_533), .A2(n_644), .B1(n_1066), .B2(n_1067), .Y(n_1065) );
OAI22xp5_ASAP7_75t_L g1102 ( .A1(n_533), .A2(n_975), .B1(n_1103), .B2(n_1104), .Y(n_1102) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_536), .B(n_544), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_541), .Y(n_536) );
INVx2_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
INVx4_ASAP7_75t_L g602 ( .A(n_539), .Y(n_602) );
OAI21xp33_ASAP7_75t_SL g807 ( .A1(n_539), .A2(n_808), .B(n_809), .Y(n_807) );
INVx4_ASAP7_75t_L g871 ( .A(n_539), .Y(n_871) );
INVx1_ASAP7_75t_L g696 ( .A(n_540), .Y(n_696) );
INVxp67_ASAP7_75t_L g1045 ( .A(n_542), .Y(n_1045) );
INVx1_ASAP7_75t_SL g929 ( .A(n_543), .Y(n_929) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_550), .Y(n_544) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g579 ( .A(n_547), .Y(n_579) );
INVx2_ASAP7_75t_L g590 ( .A(n_547), .Y(n_590) );
INVx3_ASAP7_75t_L g786 ( .A(n_547), .Y(n_786) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .B1(n_586), .B2(n_608), .Y(n_555) );
OAI22xp5_ASAP7_75t_SL g650 ( .A1(n_556), .A2(n_651), .B1(n_652), .B2(n_682), .Y(n_650) );
INVx2_ASAP7_75t_SL g682 ( .A(n_556), .Y(n_682) );
INVx3_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
XOR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_585), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_559), .B(n_570), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_560), .B(n_564), .Y(n_559) );
NAND3xp33_ASAP7_75t_L g564 ( .A(n_565), .B(n_567), .C(n_569), .Y(n_564) );
NOR2x1_ASAP7_75t_L g570 ( .A(n_571), .B(n_577), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_575), .Y(n_571) );
INVx1_ASAP7_75t_L g1021 ( .A(n_574), .Y(n_1021) );
HB1xp67_ASAP7_75t_L g791 ( .A(n_576), .Y(n_791) );
INVx2_ASAP7_75t_L g877 ( .A(n_576), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_581), .Y(n_577) );
INVxp67_ASAP7_75t_L g1056 ( .A(n_579), .Y(n_1056) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g608 ( .A(n_586), .Y(n_608) );
NAND4xp75_ASAP7_75t_L g587 ( .A(n_588), .B(n_593), .C(n_600), .D(n_605), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_592), .Y(n_588) );
AND2x2_ASAP7_75t_SL g593 ( .A(n_594), .B(n_596), .Y(n_593) );
INVx2_ASAP7_75t_SL g774 ( .A(n_597), .Y(n_774) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g955 ( .A(n_599), .Y(n_955) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_611), .B1(n_683), .B2(n_684), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_613), .B1(n_649), .B2(n_650), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g648 ( .A(n_614), .Y(n_648) );
AND2x2_ASAP7_75t_SL g614 ( .A(n_615), .B(n_624), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_616), .B(n_620), .Y(n_615) );
NAND2xp33_ASAP7_75t_SL g616 ( .A(n_617), .B(n_619), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
NOR3xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_628), .C(n_638), .Y(n_624) );
OAI221xp5_ASAP7_75t_SL g628 ( .A1(n_629), .A2(n_632), .B1(n_633), .B2(n_635), .C(n_636), .Y(n_628) );
OAI221xp5_ASAP7_75t_L g661 ( .A1(n_629), .A2(n_662), .B1(n_663), .B2(n_664), .C(n_665), .Y(n_661) );
OAI221xp5_ASAP7_75t_SL g860 ( .A1(n_629), .A2(n_861), .B1(n_862), .B2(n_863), .C(n_864), .Y(n_860) );
OAI221xp5_ASAP7_75t_L g1027 ( .A1(n_629), .A2(n_663), .B1(n_1028), .B2(n_1029), .C(n_1030), .Y(n_1027) );
OAI221xp5_ASAP7_75t_SL g1098 ( .A1(n_629), .A2(n_633), .B1(n_1099), .B2(n_1100), .C(n_1101), .Y(n_1098) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx4_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
BUFx2_ASAP7_75t_L g969 ( .A(n_631), .Y(n_969) );
OAI21xp5_ASAP7_75t_SL g993 ( .A1(n_631), .A2(n_994), .B(n_995), .Y(n_993) );
OAI221xp5_ASAP7_75t_SL g703 ( .A1(n_633), .A2(n_704), .B1(n_705), .B2(n_706), .C(n_707), .Y(n_703) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_640), .B1(n_641), .B2(n_642), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_642), .A2(n_700), .B1(n_701), .B2(n_702), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g865 ( .A1(n_642), .A2(n_701), .B1(n_866), .B2(n_867), .Y(n_865) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g975 ( .A(n_643), .Y(n_975) );
CKINVDCx16_ASAP7_75t_R g643 ( .A(n_644), .Y(n_643) );
BUFx2_ASAP7_75t_L g671 ( .A(n_644), .Y(n_671) );
OR2x6_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_SL g654 ( .A(n_655), .B(n_672), .Y(n_654) );
NOR3xp33_ASAP7_75t_L g655 ( .A(n_656), .B(n_661), .C(n_666), .Y(n_655) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_SL g710 ( .A(n_659), .Y(n_710) );
INVx2_ASAP7_75t_L g827 ( .A(n_659), .Y(n_827) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .B1(n_670), .B2(n_671), .Y(n_666) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx3_ASAP7_75t_SL g701 ( .A(n_669), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_671), .A2(n_701), .B1(n_778), .B2(n_779), .Y(n_777) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_678), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g673 ( .A(n_674), .B(n_676), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
OAI22xp5_ASAP7_75t_SL g684 ( .A1(n_685), .A2(n_764), .B1(n_765), .B2(n_794), .Y(n_684) );
INVx1_ASAP7_75t_L g794 ( .A(n_685), .Y(n_794) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_715), .B1(n_716), .B2(n_763), .Y(n_686) );
INVx1_ASAP7_75t_L g763 ( .A(n_687), .Y(n_763) );
INVx1_ASAP7_75t_SL g714 ( .A(n_688), .Y(n_714) );
AND2x2_ASAP7_75t_SL g688 ( .A(n_689), .B(n_698), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_693), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_697), .Y(n_693) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NOR3xp33_ASAP7_75t_SL g698 ( .A(n_699), .B(n_703), .C(n_708), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g972 ( .A1(n_701), .A2(n_973), .B1(n_974), .B2(n_975), .Y(n_972) );
OAI21xp5_ASAP7_75t_SL g720 ( .A1(n_704), .A2(n_721), .B(n_722), .Y(n_720) );
OAI221xp5_ASAP7_75t_L g772 ( .A1(n_704), .A2(n_773), .B1(n_774), .B2(n_775), .C(n_776), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_710), .B1(n_711), .B2(n_712), .Y(n_708) );
INVx2_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
XNOR2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_743), .Y(n_716) );
XOR2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_742), .Y(n_717) );
NAND3x1_ASAP7_75t_L g718 ( .A(n_719), .B(n_731), .C(n_737), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_723), .Y(n_719) );
NAND3xp33_ASAP7_75t_L g723 ( .A(n_724), .B(n_726), .C(n_729), .Y(n_723) );
BUFx6f_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_735), .Y(n_731) );
INVx3_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
INVx1_ASAP7_75t_L g927 ( .A(n_740), .Y(n_927) );
XOR2x2_ASAP7_75t_L g743 ( .A(n_744), .B(n_762), .Y(n_743) );
NAND4xp75_ASAP7_75t_L g744 ( .A(n_745), .B(n_749), .C(n_756), .D(n_760), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
OA211x2_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_751), .B(n_753), .C(n_754), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g804 ( .A1(n_751), .A2(n_770), .B1(n_805), .B2(n_806), .Y(n_804) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g829 ( .A(n_752), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g862 ( .A(n_755), .Y(n_862) );
AND2x2_ASAP7_75t_L g756 ( .A(n_757), .B(n_759), .Y(n_756) );
INVx2_ASAP7_75t_L g931 ( .A(n_758), .Y(n_931) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx2_ASAP7_75t_L g793 ( .A(n_766), .Y(n_793) );
AND2x2_ASAP7_75t_SL g766 ( .A(n_767), .B(n_780), .Y(n_766) );
NOR3xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_772), .C(n_777), .Y(n_767) );
OAI22xp5_ASAP7_75t_L g990 ( .A1(n_770), .A2(n_829), .B1(n_991), .B2(n_992), .Y(n_990) );
NOR2xp33_ASAP7_75t_L g780 ( .A(n_781), .B(n_784), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_782), .B(n_783), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_785), .B(n_787), .Y(n_784) );
INVx4_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx3_ASAP7_75t_L g944 ( .A(n_789), .Y(n_944) );
INVx4_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g1077 ( .A(n_795), .Y(n_1077) );
AOI22xp5_ASAP7_75t_SL g795 ( .A1(n_796), .A2(n_1039), .B1(n_1074), .B2(n_1075), .Y(n_795) );
INVx1_ASAP7_75t_L g1074 ( .A(n_796), .Y(n_1074) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_901), .B1(n_1037), .B2(n_1038), .Y(n_796) );
INVx1_ASAP7_75t_L g1037 ( .A(n_797), .Y(n_1037) );
AOI22xp5_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_851), .B1(n_852), .B2(n_900), .Y(n_797) );
INVx1_ASAP7_75t_L g900 ( .A(n_798), .Y(n_900) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_822), .B1(n_849), .B2(n_850), .Y(n_798) );
INVx1_ASAP7_75t_L g849 ( .A(n_799), .Y(n_849) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx2_ASAP7_75t_L g821 ( .A(n_802), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_803), .B(n_813), .Y(n_802) );
NOR3xp33_ASAP7_75t_L g803 ( .A(n_804), .B(n_807), .C(n_810), .Y(n_803) );
NOR2xp33_ASAP7_75t_L g813 ( .A(n_814), .B(n_818), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .Y(n_818) );
INVx2_ASAP7_75t_L g850 ( .A(n_822), .Y(n_850) );
INVx2_ASAP7_75t_SL g848 ( .A(n_823), .Y(n_848) );
AND2x2_ASAP7_75t_L g823 ( .A(n_824), .B(n_839), .Y(n_823) );
NOR3xp33_ASAP7_75t_L g824 ( .A(n_825), .B(n_830), .C(n_836), .Y(n_824) );
OAI22xp5_ASAP7_75t_L g825 ( .A1(n_826), .A2(n_827), .B1(n_828), .B2(n_829), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g1095 ( .A1(n_827), .A2(n_829), .B1(n_1096), .B2(n_1097), .Y(n_1095) );
OA211x2_ASAP7_75t_L g951 ( .A1(n_829), .A2(n_952), .B(n_953), .C(n_954), .Y(n_951) );
OAI221xp5_ASAP7_75t_SL g830 ( .A1(n_831), .A2(n_832), .B1(n_833), .B2(n_834), .C(n_835), .Y(n_830) );
NOR2xp33_ASAP7_75t_L g839 ( .A(n_840), .B(n_844), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_841), .B(n_842), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_845), .B(n_846), .Y(n_844) );
INVx2_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
OAI22xp5_ASAP7_75t_SL g852 ( .A1(n_853), .A2(n_854), .B1(n_880), .B2(n_881), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx2_ASAP7_75t_L g879 ( .A(n_855), .Y(n_879) );
AND2x2_ASAP7_75t_L g855 ( .A(n_856), .B(n_868), .Y(n_855) );
NOR3xp33_ASAP7_75t_L g856 ( .A(n_857), .B(n_860), .C(n_865), .Y(n_856) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_869), .B(n_873), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_870), .B(n_872), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_874), .B(n_875), .Y(n_873) );
INVx2_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g1043 ( .A1(n_877), .A2(n_1044), .B1(n_1045), .B2(n_1046), .Y(n_1043) );
AOI22xp5_ASAP7_75t_L g1039 ( .A1(n_880), .A2(n_881), .B1(n_1040), .B2(n_1073), .Y(n_1039) );
INVx2_ASAP7_75t_SL g880 ( .A(n_881), .Y(n_880) );
XNOR2x2_ASAP7_75t_L g881 ( .A(n_882), .B(n_883), .Y(n_881) );
NOR4xp75_ASAP7_75t_L g883 ( .A(n_884), .B(n_887), .C(n_891), .D(n_895), .Y(n_883) );
NAND2xp5_ASAP7_75t_SL g884 ( .A(n_885), .B(n_886), .Y(n_884) );
NAND2xp5_ASAP7_75t_SL g887 ( .A(n_888), .B(n_889), .Y(n_887) );
OAI21xp5_ASAP7_75t_SL g895 ( .A1(n_896), .A2(n_898), .B(n_899), .Y(n_895) );
OAI21xp33_ASAP7_75t_L g914 ( .A1(n_896), .A2(n_915), .B(n_916), .Y(n_914) );
INVx3_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
INVx1_ASAP7_75t_L g1038 ( .A(n_901), .Y(n_1038) );
XOR2xp5_ASAP7_75t_L g901 ( .A(n_902), .B(n_958), .Y(n_901) );
HB1xp67_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
OAI22xp5_ASAP7_75t_L g904 ( .A1(n_905), .A2(n_906), .B1(n_937), .B2(n_938), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx2_ASAP7_75t_SL g908 ( .A(n_909), .Y(n_908) );
AND2x2_ASAP7_75t_L g909 ( .A(n_910), .B(n_920), .Y(n_909) );
NOR3xp33_ASAP7_75t_L g910 ( .A(n_911), .B(n_914), .C(n_917), .Y(n_910) );
NOR3xp33_ASAP7_75t_L g920 ( .A(n_921), .B(n_925), .C(n_930), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_922), .B(n_924), .Y(n_921) );
OAI22xp5_ASAP7_75t_L g925 ( .A1(n_926), .A2(n_927), .B1(n_928), .B2(n_929), .Y(n_925) );
OAI22xp5_ASAP7_75t_L g930 ( .A1(n_931), .A2(n_932), .B1(n_933), .B2(n_934), .Y(n_930) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g1058 ( .A(n_935), .Y(n_1058) );
INVx1_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
NAND4xp75_ASAP7_75t_L g939 ( .A(n_940), .B(n_945), .C(n_951), .D(n_956), .Y(n_939) );
AND2x2_ASAP7_75t_L g940 ( .A(n_941), .B(n_943), .Y(n_940) );
AND2x2_ASAP7_75t_L g945 ( .A(n_946), .B(n_949), .Y(n_945) );
AOI22xp5_ASAP7_75t_L g958 ( .A1(n_959), .A2(n_960), .B1(n_1007), .B2(n_1036), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
XNOR2xp5_ASAP7_75t_L g960 ( .A(n_961), .B(n_987), .Y(n_960) );
XOR2x2_ASAP7_75t_L g961 ( .A(n_962), .B(n_986), .Y(n_961) );
NAND2xp5_ASAP7_75t_L g962 ( .A(n_963), .B(n_976), .Y(n_962) );
NOR3xp33_ASAP7_75t_L g963 ( .A(n_964), .B(n_967), .C(n_972), .Y(n_963) );
OAI21xp33_ASAP7_75t_L g967 ( .A1(n_968), .A2(n_969), .B(n_970), .Y(n_967) );
NOR2xp33_ASAP7_75t_L g976 ( .A(n_977), .B(n_983), .Y(n_976) );
NAND2xp5_ASAP7_75t_L g977 ( .A(n_978), .B(n_979), .Y(n_977) );
INVx3_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g983 ( .A(n_984), .B(n_985), .Y(n_983) );
XOR2x2_ASAP7_75t_L g987 ( .A(n_988), .B(n_1006), .Y(n_987) );
NAND2xp5_ASAP7_75t_L g988 ( .A(n_989), .B(n_999), .Y(n_988) );
NOR3xp33_ASAP7_75t_L g989 ( .A(n_990), .B(n_993), .C(n_996), .Y(n_989) );
NOR2xp33_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1003), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1002), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1005), .Y(n_1003) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1007), .Y(n_1036) );
INVx2_ASAP7_75t_L g1035 ( .A(n_1008), .Y(n_1035) );
AND2x2_ASAP7_75t_SL g1008 ( .A(n_1009), .B(n_1023), .Y(n_1008) );
NOR2xp33_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1015), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1014), .Y(n_1010) );
INVx2_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_1016), .B(n_1022), .Y(n_1015) );
INVx2_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
INVx3_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
INVx1_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
NOR3xp33_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1027), .C(n_1031), .Y(n_1023) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1039), .Y(n_1075) );
INVx1_ASAP7_75t_L g1073 ( .A(n_1040), .Y(n_1073) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1041), .Y(n_1072) );
AND4x1_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1053), .C(n_1064), .D(n_1068), .Y(n_1041) );
NOR2xp33_ASAP7_75t_SL g1042 ( .A(n_1043), .B(n_1047), .Y(n_1042) );
OAI22xp5_ASAP7_75t_L g1047 ( .A1(n_1048), .A2(n_1049), .B1(n_1051), .B2(n_1052), .Y(n_1047) );
BUFx2_ASAP7_75t_R g1049 ( .A(n_1050), .Y(n_1049) );
NOR2xp33_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1059), .Y(n_1053) );
OAI22xp5_ASAP7_75t_L g1054 ( .A1(n_1055), .A2(n_1056), .B1(n_1057), .B2(n_1058), .Y(n_1054) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
INVx3_ASAP7_75t_L g1069 ( .A(n_1070), .Y(n_1069) );
INVx2_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
NOR2x1_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1084), .Y(n_1079) );
OR2x2_ASAP7_75t_SL g1126 ( .A(n_1080), .B(n_1085), .Y(n_1126) );
NAND2xp5_ASAP7_75t_L g1080 ( .A(n_1081), .B(n_1083), .Y(n_1080) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
HB1xp67_ASAP7_75t_L g1114 ( .A(n_1082), .Y(n_1114) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_1082), .B(n_1117), .Y(n_1120) );
CKINVDCx16_ASAP7_75t_R g1117 ( .A(n_1083), .Y(n_1117) );
CKINVDCx20_ASAP7_75t_R g1084 ( .A(n_1085), .Y(n_1084) );
NAND2xp5_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1087), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1088 ( .A(n_1089), .B(n_1090), .Y(n_1088) );
OAI322xp33_ASAP7_75t_L g1091 ( .A1(n_1092), .A2(n_1114), .A3(n_1115), .B1(n_1118), .B2(n_1121), .C1(n_1122), .C2(n_1124), .Y(n_1091) );
INVx1_ASAP7_75t_SL g1113 ( .A(n_1093), .Y(n_1113) );
AND2x2_ASAP7_75t_SL g1093 ( .A(n_1094), .B(n_1105), .Y(n_1093) );
NOR3xp33_ASAP7_75t_L g1094 ( .A(n_1095), .B(n_1098), .C(n_1102), .Y(n_1094) );
NOR2xp33_ASAP7_75t_L g1105 ( .A(n_1106), .B(n_1109), .Y(n_1105) );
NAND2xp5_ASAP7_75t_L g1106 ( .A(n_1107), .B(n_1108), .Y(n_1106) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1111), .Y(n_1109) );
HB1xp67_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
CKINVDCx16_ASAP7_75t_R g1118 ( .A(n_1119), .Y(n_1118) );
HB1xp67_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
CKINVDCx20_ASAP7_75t_R g1124 ( .A(n_1125), .Y(n_1124) );
CKINVDCx20_ASAP7_75t_R g1125 ( .A(n_1126), .Y(n_1125) );
endmodule