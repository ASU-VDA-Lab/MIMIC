module real_aes_9237_n_234 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_234);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_234;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_239;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1346;
wire n_552;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_238;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_246;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_337;
wire n_247;
wire n_264;
wire n_237;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_245;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_248;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_1404;
wire n_402;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1145;
wire n_645;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_265;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1403;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_249;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_1175;
wire n_778;
wire n_1170;
wire n_522;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_243;
wire n_692;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_1343;
wire n_719;
wire n_465;
wire n_1156;
wire n_988;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_241;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_892;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_236;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_244;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_314;
wire n_283;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_240;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVx1_ASAP7_75t_L g1146 ( .A(n_0), .Y(n_1146) );
CKINVDCx5p33_ASAP7_75t_R g870 ( .A(n_1), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_2), .A2(n_226), .B1(n_779), .B2(n_780), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_2), .A2(n_226), .B1(n_791), .B2(n_792), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_3), .A2(n_207), .B1(n_689), .B2(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g709 ( .A(n_3), .Y(n_709) );
AO22x2_ASAP7_75t_L g928 ( .A1(n_4), .A2(n_929), .B1(n_971), .B2(n_972), .Y(n_928) );
INVxp67_ASAP7_75t_L g971 ( .A(n_4), .Y(n_971) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_5), .Y(n_247) );
AND2x2_ASAP7_75t_L g275 ( .A(n_5), .B(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_5), .B(n_179), .Y(n_304) );
INVx1_ASAP7_75t_L g357 ( .A(n_5), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g740 ( .A(n_6), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g1365 ( .A1(n_7), .A2(n_143), .B1(n_791), .B2(n_994), .Y(n_1365) );
INVx1_ASAP7_75t_L g1397 ( .A(n_7), .Y(n_1397) );
INVxp67_ASAP7_75t_SL g472 ( .A(n_8), .Y(n_472) );
AOI221xp5_ASAP7_75t_L g510 ( .A1(n_8), .A2(n_223), .B1(n_511), .B2(n_513), .C(n_515), .Y(n_510) );
INVx1_ASAP7_75t_L g817 ( .A(n_9), .Y(n_817) );
OAI22xp33_ASAP7_75t_L g845 ( .A1(n_9), .A2(n_129), .B1(n_731), .B2(n_737), .Y(n_845) );
INVx1_ASAP7_75t_L g644 ( .A(n_10), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_10), .A2(n_62), .B1(n_702), .B2(n_704), .Y(n_701) );
INVx1_ASAP7_75t_L g1258 ( .A(n_11), .Y(n_1258) );
INVxp33_ASAP7_75t_SL g456 ( .A(n_12), .Y(n_456) );
AOI221xp5_ASAP7_75t_L g495 ( .A1(n_12), .A2(n_66), .B1(n_421), .B2(n_496), .C(n_498), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_13), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g441 ( .A(n_14), .Y(n_441) );
INVxp67_ASAP7_75t_SL g809 ( .A(n_15), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_15), .A2(n_215), .B1(n_423), .B2(n_798), .Y(n_840) );
OAI221xp5_ASAP7_75t_L g295 ( .A1(n_16), .A2(n_84), .B1(n_296), .B2(n_305), .C(n_309), .Y(n_295) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_16), .A2(n_84), .B1(n_399), .B2(n_406), .Y(n_398) );
XNOR2xp5_ASAP7_75t_L g975 ( .A(n_17), .B(n_976), .Y(n_975) );
AO221x2_ASAP7_75t_L g1167 ( .A1(n_17), .A2(n_49), .B1(n_1144), .B2(n_1166), .C(n_1168), .Y(n_1167) );
INVx1_ASAP7_75t_L g1043 ( .A(n_18), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_18), .A2(n_177), .B1(n_519), .B2(n_692), .Y(n_1063) );
OR2x2_ASAP7_75t_L g371 ( .A(n_19), .B(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g389 ( .A(n_19), .Y(n_389) );
INVx1_ASAP7_75t_L g1169 ( .A(n_20), .Y(n_1169) );
AOI22xp33_ASAP7_75t_SL g826 ( .A1(n_21), .A2(n_68), .B1(n_773), .B2(n_827), .Y(n_826) );
INVxp33_ASAP7_75t_L g850 ( .A(n_21), .Y(n_850) );
INVx1_ASAP7_75t_L g1185 ( .A(n_22), .Y(n_1185) );
INVx1_ASAP7_75t_L g880 ( .A(n_23), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_23), .A2(n_157), .B1(n_913), .B2(n_916), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_24), .A2(n_87), .B1(n_666), .B2(n_668), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_24), .A2(n_87), .B1(n_685), .B2(n_686), .Y(n_684) );
INVx1_ASAP7_75t_L g522 ( .A(n_25), .Y(n_522) );
INVx1_ASAP7_75t_L g274 ( .A(n_26), .Y(n_274) );
OR2x2_ASAP7_75t_L g303 ( .A(n_26), .B(n_304), .Y(n_303) );
BUFx2_ASAP7_75t_L g315 ( .A(n_26), .Y(n_315) );
BUFx2_ASAP7_75t_L g447 ( .A(n_26), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g1360 ( .A(n_27), .Y(n_1360) );
INVx1_ASAP7_75t_L g988 ( .A(n_28), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g996 ( .A1(n_28), .A2(n_176), .B1(n_773), .B2(n_997), .Y(n_996) );
INVx1_ASAP7_75t_L g872 ( .A(n_29), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_29), .A2(n_133), .B1(n_693), .B2(n_922), .Y(n_921) );
INVx1_ASAP7_75t_L g1256 ( .A(n_30), .Y(n_1256) );
INVx1_ASAP7_75t_L g815 ( .A(n_31), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_31), .A2(n_54), .B1(n_583), .B2(n_838), .Y(n_837) );
OAI221xp5_ASAP7_75t_L g937 ( .A1(n_32), .A2(n_203), .B1(n_737), .B2(n_938), .C(n_939), .Y(n_937) );
INVx1_ASAP7_75t_L g946 ( .A(n_32), .Y(n_946) );
OAI221xp5_ASAP7_75t_L g460 ( .A1(n_33), .A2(n_48), .B1(n_296), .B2(n_309), .C(n_461), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_33), .A2(n_48), .B1(n_399), .B2(n_507), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g1106 ( .A(n_34), .Y(n_1106) );
CKINVDCx16_ASAP7_75t_R g1182 ( .A(n_35), .Y(n_1182) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_36), .A2(n_197), .B1(n_787), .B2(n_789), .Y(n_991) );
AOI22xp33_ASAP7_75t_SL g1003 ( .A1(n_36), .A2(n_197), .B1(n_770), .B2(n_821), .Y(n_1003) );
INVx1_ASAP7_75t_L g1252 ( .A(n_37), .Y(n_1252) );
CKINVDCx5p33_ASAP7_75t_R g1073 ( .A(n_38), .Y(n_1073) );
AOI22xp33_ASAP7_75t_L g1050 ( .A1(n_39), .A2(n_232), .B1(n_671), .B2(n_672), .Y(n_1050) );
AOI22xp33_ASAP7_75t_SL g1056 ( .A1(n_39), .A2(n_232), .B1(n_412), .B2(n_1057), .Y(n_1056) );
INVx1_ASAP7_75t_L g655 ( .A(n_40), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_40), .A2(n_214), .B1(n_675), .B2(n_677), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_41), .A2(n_69), .B1(n_773), .B2(n_824), .Y(n_823) );
AOI22xp33_ASAP7_75t_SL g834 ( .A1(n_41), .A2(n_69), .B1(n_798), .B2(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g1028 ( .A(n_42), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_42), .A2(n_137), .B1(n_675), .B2(n_677), .Y(n_1051) );
OAI22xp5_ASAP7_75t_L g981 ( .A1(n_43), .A2(n_200), .B1(n_737), .B2(n_982), .Y(n_981) );
OAI22xp33_ASAP7_75t_L g1012 ( .A1(n_43), .A2(n_200), .B1(n_755), .B2(n_1013), .Y(n_1012) );
AOI221xp5_ASAP7_75t_L g569 ( .A1(n_44), .A2(n_61), .B1(n_313), .B2(n_570), .C(n_571), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_44), .A2(n_61), .B1(n_583), .B2(n_584), .Y(n_582) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_45), .Y(n_347) );
INVx1_ASAP7_75t_L g482 ( .A(n_46), .Y(n_482) );
INVx1_ASAP7_75t_L g1356 ( .A(n_47), .Y(n_1356) );
AOI221xp5_ASAP7_75t_L g1385 ( .A1(n_47), .A2(n_50), .B1(n_549), .B2(n_768), .C(n_783), .Y(n_1385) );
INVx1_ASAP7_75t_L g1354 ( .A(n_50), .Y(n_1354) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_51), .A2(n_80), .B1(n_821), .B2(n_830), .Y(n_829) );
INVxp67_ASAP7_75t_SL g843 ( .A(n_51), .Y(n_843) );
INVx1_ASAP7_75t_L g1033 ( .A(n_52), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_52), .A2(n_105), .B1(n_752), .B2(n_1053), .Y(n_1052) );
AO22x2_ASAP7_75t_L g624 ( .A1(n_53), .A2(n_625), .B1(n_719), .B2(n_720), .Y(n_624) );
INVxp67_ASAP7_75t_SL g719 ( .A(n_53), .Y(n_719) );
INVxp33_ASAP7_75t_L g811 ( .A(n_54), .Y(n_811) );
INVx1_ASAP7_75t_L g1194 ( .A(n_55), .Y(n_1194) );
CKINVDCx16_ASAP7_75t_R g1199 ( .A(n_56), .Y(n_1199) );
AOI21xp5_ASAP7_75t_L g893 ( .A1(n_57), .A2(n_667), .B(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g897 ( .A(n_57), .Y(n_897) );
INVx1_ASAP7_75t_L g748 ( .A(n_58), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_58), .A2(n_123), .B1(n_792), .B2(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g1066 ( .A(n_59), .Y(n_1066) );
INVx1_ASAP7_75t_L g944 ( .A(n_60), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_60), .A2(n_185), .B1(n_607), .B2(n_689), .Y(n_970) );
INVx1_ASAP7_75t_L g649 ( .A(n_62), .Y(n_649) );
INVx1_ASAP7_75t_L g751 ( .A(n_63), .Y(n_751) );
AOI22xp33_ASAP7_75t_SL g795 ( .A1(n_63), .A2(n_181), .B1(n_789), .B2(n_796), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_64), .A2(n_194), .B1(n_773), .B2(n_957), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_64), .A2(n_194), .B1(n_689), .B2(n_798), .Y(n_966) );
INVx1_ASAP7_75t_L g1086 ( .A(n_65), .Y(n_1086) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_65), .A2(n_85), .B1(n_421), .B2(n_689), .Y(n_1125) );
INVxp33_ASAP7_75t_L g458 ( .A(n_66), .Y(n_458) );
INVx1_ASAP7_75t_L g1152 ( .A(n_67), .Y(n_1152) );
INVxp67_ASAP7_75t_SL g851 ( .A(n_68), .Y(n_851) );
INVx1_ASAP7_75t_L g743 ( .A(n_70), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_70), .A2(n_113), .B1(n_773), .B2(n_775), .Y(n_772) );
XNOR2x2_ASAP7_75t_L g1023 ( .A(n_71), .B(n_1024), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g1370 ( .A1(n_72), .A2(n_150), .B1(n_792), .B2(n_993), .Y(n_1370) );
OAI22xp5_ASAP7_75t_L g1401 ( .A1(n_72), .A2(n_150), .B1(n_1402), .B2(n_1403), .Y(n_1401) );
INVxp33_ASAP7_75t_L g464 ( .A(n_73), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_73), .A2(n_114), .B1(n_517), .B2(n_519), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g1159 ( .A1(n_74), .A2(n_134), .B1(n_1160), .B2(n_1163), .Y(n_1159) );
AOI221xp5_ASAP7_75t_L g543 ( .A1(n_75), .A2(n_89), .B1(n_544), .B2(n_546), .C(n_549), .Y(n_543) );
INVx1_ASAP7_75t_L g596 ( .A(n_75), .Y(n_596) );
OAI222xp33_ASAP7_75t_L g730 ( .A1(n_76), .A2(n_162), .B1(n_192), .B2(n_731), .C1(n_734), .C2(n_737), .Y(n_730) );
INVx1_ASAP7_75t_L g753 ( .A(n_76), .Y(n_753) );
AO22x2_ASAP7_75t_L g725 ( .A1(n_77), .A2(n_726), .B1(n_727), .B2(n_801), .Y(n_725) );
INVxp67_ASAP7_75t_SL g726 ( .A(n_77), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_78), .A2(n_95), .B1(n_768), .B2(n_783), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_78), .A2(n_95), .B1(n_787), .B2(n_789), .Y(n_786) );
INVx1_ASAP7_75t_L g372 ( .A(n_79), .Y(n_372) );
INVx1_ASAP7_75t_L g390 ( .A(n_79), .Y(n_390) );
INVxp33_ASAP7_75t_L g847 ( .A(n_80), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_81), .A2(n_147), .B1(n_789), .B2(n_1006), .Y(n_1005) );
INVx1_ASAP7_75t_L g1018 ( .A(n_81), .Y(n_1018) );
CKINVDCx16_ASAP7_75t_R g1201 ( .A(n_82), .Y(n_1201) );
AOI22xp33_ASAP7_75t_SL g992 ( .A1(n_83), .A2(n_124), .B1(n_993), .B2(n_994), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_83), .A2(n_124), .B1(n_779), .B2(n_1001), .Y(n_1000) );
INVx1_ASAP7_75t_L g1095 ( .A(n_85), .Y(n_1095) );
AOI221xp5_ASAP7_75t_L g889 ( .A1(n_86), .A2(n_211), .B1(n_779), .B2(n_890), .C(n_891), .Y(n_889) );
INVx1_ASAP7_75t_L g898 ( .A(n_86), .Y(n_898) );
INVx1_ASAP7_75t_L g739 ( .A(n_88), .Y(n_739) );
AOI22xp33_ASAP7_75t_SL g767 ( .A1(n_88), .A2(n_192), .B1(n_768), .B2(n_770), .Y(n_767) );
INVx1_ASAP7_75t_L g602 ( .A(n_89), .Y(n_602) );
XNOR2xp5_ASAP7_75t_L g1409 ( .A(n_90), .B(n_1410), .Y(n_1409) );
INVx1_ASAP7_75t_L g1184 ( .A(n_91), .Y(n_1184) );
INVx1_ASAP7_75t_L g1091 ( .A(n_92), .Y(n_1091) );
AOI221xp5_ASAP7_75t_L g1122 ( .A1(n_92), .A2(n_201), .B1(n_366), .B2(n_496), .C(n_1123), .Y(n_1122) );
CKINVDCx5p33_ASAP7_75t_R g341 ( .A(n_93), .Y(n_341) );
INVx1_ASAP7_75t_L g561 ( .A(n_94), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_94), .A2(n_209), .B1(n_366), .B2(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g277 ( .A(n_96), .Y(n_277) );
AOI221xp5_ASAP7_75t_L g373 ( .A1(n_96), .A2(n_196), .B1(n_374), .B2(n_381), .C(n_385), .Y(n_373) );
INVx1_ASAP7_75t_L g488 ( .A(n_97), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_98), .A2(n_193), .B1(n_541), .B2(n_573), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_98), .A2(n_193), .B1(n_366), .B2(n_394), .Y(n_581) );
INVx1_ASAP7_75t_L g979 ( .A(n_99), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_99), .A2(n_172), .B1(n_571), .B2(n_821), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_100), .A2(n_228), .B1(n_821), .B2(n_822), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_100), .A2(n_228), .B1(n_382), .B2(n_787), .Y(n_836) );
AO221x2_ASAP7_75t_L g1137 ( .A1(n_101), .A2(n_166), .B1(n_1138), .B2(n_1144), .C(n_1145), .Y(n_1137) );
CKINVDCx5p33_ASAP7_75t_R g1362 ( .A(n_102), .Y(n_1362) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_103), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_104), .A2(n_213), .B1(n_671), .B2(n_672), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_104), .A2(n_213), .B1(n_392), .B2(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g1027 ( .A(n_105), .Y(n_1027) );
INVx1_ASAP7_75t_L g239 ( .A(n_106), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g887 ( .A(n_107), .Y(n_887) );
CKINVDCx5p33_ASAP7_75t_R g985 ( .A(n_108), .Y(n_985) );
CKINVDCx5p33_ASAP7_75t_R g633 ( .A(n_109), .Y(n_633) );
AOI21xp33_ASAP7_75t_L g878 ( .A1(n_110), .A2(n_313), .B(n_570), .Y(n_878) );
INVx1_ASAP7_75t_L g910 ( .A(n_110), .Y(n_910) );
XOR2xp5_ASAP7_75t_L g261 ( .A(n_111), .B(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g940 ( .A(n_112), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_112), .A2(n_132), .B1(n_821), .B2(n_959), .Y(n_964) );
INVx1_ASAP7_75t_L g742 ( .A(n_113), .Y(n_742) );
INVxp67_ASAP7_75t_SL g474 ( .A(n_114), .Y(n_474) );
CKINVDCx5p33_ASAP7_75t_R g1105 ( .A(n_115), .Y(n_1105) );
AOI22xp5_ASAP7_75t_L g1165 ( .A1(n_116), .A2(n_161), .B1(n_1144), .B2(n_1166), .Y(n_1165) );
AOI222xp33_ASAP7_75t_L g1345 ( .A1(n_116), .A2(n_1346), .B1(n_1404), .B2(n_1408), .C1(n_1411), .C2(n_1415), .Y(n_1345) );
XNOR2xp5_ASAP7_75t_L g1347 ( .A(n_116), .B(n_1348), .Y(n_1347) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_117), .A2(n_195), .B1(n_541), .B2(n_542), .Y(n_540) );
INVx1_ASAP7_75t_L g605 ( .A(n_117), .Y(n_605) );
INVx1_ASAP7_75t_L g320 ( .A(n_118), .Y(n_320) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_118), .A2(n_156), .B1(n_412), .B2(n_414), .C(n_416), .Y(n_411) );
INVx1_ASAP7_75t_L g335 ( .A(n_119), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_119), .A2(n_148), .B1(n_421), .B2(n_423), .Y(n_420) );
INVx1_ASAP7_75t_L g1040 ( .A(n_120), .Y(n_1040) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_120), .A2(n_180), .B1(n_421), .B2(n_1060), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_121), .A2(n_216), .B1(n_421), .B2(n_686), .Y(n_690) );
INVx1_ASAP7_75t_L g715 ( .A(n_121), .Y(n_715) );
CKINVDCx5p33_ASAP7_75t_R g869 ( .A(n_122), .Y(n_869) );
INVx1_ASAP7_75t_L g747 ( .A(n_123), .Y(n_747) );
CKINVDCx5p33_ASAP7_75t_R g1099 ( .A(n_125), .Y(n_1099) );
INVx1_ASAP7_75t_L g288 ( .A(n_126), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_126), .A2(n_229), .B1(n_392), .B2(n_393), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g867 ( .A(n_127), .Y(n_867) );
INVx1_ASAP7_75t_L g1170 ( .A(n_128), .Y(n_1170) );
INVxp67_ASAP7_75t_SL g816 ( .A(n_129), .Y(n_816) );
INVx1_ASAP7_75t_L g953 ( .A(n_130), .Y(n_953) );
AOI22xp33_ASAP7_75t_SL g969 ( .A1(n_130), .A2(n_135), .B1(n_789), .B2(n_796), .Y(n_969) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_131), .A2(n_190), .B1(n_556), .B2(n_558), .Y(n_555) );
INVx1_ASAP7_75t_L g618 ( .A(n_131), .Y(n_618) );
INVx1_ASAP7_75t_L g932 ( .A(n_132), .Y(n_932) );
INVx1_ASAP7_75t_L g873 ( .A(n_133), .Y(n_873) );
INVx1_ASAP7_75t_L g948 ( .A(n_135), .Y(n_948) );
INVx1_ASAP7_75t_L g1071 ( .A(n_136), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1117 ( .A1(n_136), .A2(n_219), .B1(n_413), .B2(n_589), .Y(n_1117) );
INVx1_ASAP7_75t_L g1031 ( .A(n_137), .Y(n_1031) );
INVx1_ASAP7_75t_L g622 ( .A(n_138), .Y(n_622) );
CKINVDCx5p33_ASAP7_75t_R g1030 ( .A(n_139), .Y(n_1030) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_140), .A2(n_205), .B1(n_792), .B2(n_1008), .Y(n_1007) );
INVx1_ASAP7_75t_L g1015 ( .A(n_140), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_141), .A2(n_168), .B1(n_768), .B2(n_959), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_141), .A2(n_168), .B1(n_787), .B2(n_789), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g1049 ( .A1(n_142), .A2(n_165), .B1(n_666), .B2(n_668), .Y(n_1049) );
AOI22xp33_ASAP7_75t_SL g1059 ( .A1(n_142), .A2(n_165), .B1(n_685), .B2(n_1060), .Y(n_1059) );
INVx1_ASAP7_75t_L g1399 ( .A(n_143), .Y(n_1399) );
AOI22xp5_ASAP7_75t_L g1173 ( .A1(n_144), .A2(n_153), .B1(n_1160), .B2(n_1163), .Y(n_1173) );
CKINVDCx5p33_ASAP7_75t_R g884 ( .A(n_145), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g1366 ( .A1(n_146), .A2(n_187), .B1(n_583), .B2(n_1367), .Y(n_1366) );
INVx1_ASAP7_75t_L g1390 ( .A(n_146), .Y(n_1390) );
INVx1_ASAP7_75t_L g1011 ( .A(n_147), .Y(n_1011) );
INVx1_ASAP7_75t_L g317 ( .A(n_148), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g1101 ( .A(n_149), .Y(n_1101) );
INVx1_ASAP7_75t_L g486 ( .A(n_151), .Y(n_486) );
CKINVDCx5p33_ASAP7_75t_R g1357 ( .A(n_152), .Y(n_1357) );
AOI22xp5_ASAP7_75t_L g1174 ( .A1(n_154), .A2(n_184), .B1(n_1138), .B2(n_1175), .Y(n_1174) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_155), .Y(n_241) );
AND3x2_ASAP7_75t_L g1142 ( .A(n_155), .B(n_239), .C(n_1143), .Y(n_1142) );
NAND2xp5_ASAP7_75t_L g1149 ( .A(n_155), .B(n_239), .Y(n_1149) );
INVx1_ASAP7_75t_L g328 ( .A(n_156), .Y(n_328) );
INVx1_ASAP7_75t_L g877 ( .A(n_157), .Y(n_877) );
CKINVDCx5p33_ASAP7_75t_R g892 ( .A(n_158), .Y(n_892) );
INVx2_ASAP7_75t_L g252 ( .A(n_159), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g935 ( .A(n_160), .Y(n_935) );
INVx1_ASAP7_75t_L g756 ( .A(n_162), .Y(n_756) );
CKINVDCx5p33_ASAP7_75t_R g882 ( .A(n_163), .Y(n_882) );
XOR2xp5_ASAP7_75t_L g449 ( .A(n_164), .B(n_450), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g1211 ( .A1(n_167), .A2(n_171), .B1(n_1144), .B2(n_1166), .Y(n_1211) );
INVx1_ASAP7_75t_L g1143 ( .A(n_169), .Y(n_1143) );
INVx1_ASAP7_75t_L g1035 ( .A(n_170), .Y(n_1035) );
OAI22xp5_ASAP7_75t_L g1041 ( .A1(n_170), .A2(n_189), .B1(n_702), .B2(n_1013), .Y(n_1041) );
INVx1_ASAP7_75t_L g984 ( .A(n_172), .Y(n_984) );
CKINVDCx16_ASAP7_75t_R g804 ( .A(n_173), .Y(n_804) );
INVx1_ASAP7_75t_L g1254 ( .A(n_174), .Y(n_1254) );
INVx1_ASAP7_75t_L g1375 ( .A(n_175), .Y(n_1375) );
INVx1_ASAP7_75t_L g987 ( .A(n_176), .Y(n_987) );
INVx1_ASAP7_75t_L g1044 ( .A(n_177), .Y(n_1044) );
OAI221xp5_ASAP7_75t_L g1078 ( .A1(n_178), .A2(n_182), .B1(n_296), .B2(n_305), .C(n_1079), .Y(n_1078) );
OAI221xp5_ASAP7_75t_L g1111 ( .A1(n_178), .A2(n_182), .B1(n_406), .B2(n_1112), .C(n_1114), .Y(n_1111) );
INVx1_ASAP7_75t_L g254 ( .A(n_179), .Y(n_254) );
INVx2_ASAP7_75t_L g276 ( .A(n_179), .Y(n_276) );
INVx1_ASAP7_75t_L g1046 ( .A(n_180), .Y(n_1046) );
INVx1_ASAP7_75t_L g761 ( .A(n_181), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g1210 ( .A1(n_183), .A2(n_208), .B1(n_1160), .B2(n_1163), .Y(n_1210) );
AO22x2_ASAP7_75t_L g862 ( .A1(n_184), .A2(n_863), .B1(n_925), .B2(n_926), .Y(n_862) );
INVxp67_ASAP7_75t_SL g925 ( .A(n_184), .Y(n_925) );
INVx1_ASAP7_75t_L g943 ( .A(n_185), .Y(n_943) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_186), .B(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g1393 ( .A(n_187), .Y(n_1393) );
INVx1_ASAP7_75t_L g491 ( .A(n_188), .Y(n_491) );
INVx1_ASAP7_75t_L g1037 ( .A(n_189), .Y(n_1037) );
INVx1_ASAP7_75t_L g613 ( .A(n_190), .Y(n_613) );
INVx1_ASAP7_75t_L g652 ( .A(n_191), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_191), .A2(n_198), .B1(n_666), .B2(n_668), .Y(n_678) );
INVx1_ASAP7_75t_L g592 ( .A(n_195), .Y(n_592) );
INVx1_ASAP7_75t_L g283 ( .A(n_196), .Y(n_283) );
INVx1_ASAP7_75t_L g642 ( .A(n_198), .Y(n_642) );
INVx1_ASAP7_75t_L g812 ( .A(n_199), .Y(n_812) );
INVx1_ASAP7_75t_L g1089 ( .A(n_201), .Y(n_1089) );
INVx1_ASAP7_75t_L g1195 ( .A(n_202), .Y(n_1195) );
INVx1_ASAP7_75t_L g947 ( .A(n_203), .Y(n_947) );
INVxp33_ASAP7_75t_SL g459 ( .A(n_204), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_204), .A2(n_210), .B1(n_502), .B2(n_504), .Y(n_501) );
INVx1_ASAP7_75t_L g1016 ( .A(n_205), .Y(n_1016) );
INVx1_ASAP7_75t_L g1141 ( .A(n_206), .Y(n_1141) );
NAND2xp5_ASAP7_75t_L g1154 ( .A(n_206), .B(n_1151), .Y(n_1154) );
INVx1_ASAP7_75t_L g712 ( .A(n_207), .Y(n_712) );
INVx1_ASAP7_75t_L g565 ( .A(n_209), .Y(n_565) );
INVxp33_ASAP7_75t_SL g454 ( .A(n_210), .Y(n_454) );
INVx1_ASAP7_75t_L g900 ( .A(n_211), .Y(n_900) );
CKINVDCx5p33_ASAP7_75t_R g1353 ( .A(n_212), .Y(n_1353) );
INVx1_ASAP7_75t_L g637 ( .A(n_214), .Y(n_637) );
INVx1_ASAP7_75t_L g808 ( .A(n_215), .Y(n_808) );
INVx1_ASAP7_75t_L g697 ( .A(n_216), .Y(n_697) );
INVx1_ASAP7_75t_L g1075 ( .A(n_217), .Y(n_1075) );
AOI21xp33_ASAP7_75t_L g1118 ( .A1(n_217), .A2(n_1119), .B(n_1120), .Y(n_1118) );
INVx2_ASAP7_75t_L g251 ( .A(n_218), .Y(n_251) );
INVx1_ASAP7_75t_L g1076 ( .A(n_219), .Y(n_1076) );
AOI22xp33_ASAP7_75t_L g1368 ( .A1(n_220), .A2(n_221), .B1(n_1367), .B2(n_1369), .Y(n_1368) );
OAI211xp5_ASAP7_75t_SL g1377 ( .A1(n_220), .A2(n_1378), .B(n_1379), .C(n_1386), .Y(n_1377) );
OAI221xp5_ASAP7_75t_L g1387 ( .A1(n_221), .A2(n_1388), .B1(n_1389), .B2(n_1396), .C(n_1400), .Y(n_1387) );
INVx1_ASAP7_75t_L g554 ( .A(n_222), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_222), .A2(n_233), .B1(n_514), .B2(n_587), .Y(n_586) );
INVxp33_ASAP7_75t_SL g468 ( .A(n_223), .Y(n_468) );
INVx1_ASAP7_75t_L g936 ( .A(n_224), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_224), .A2(n_227), .B1(n_773), .B2(n_963), .Y(n_962) );
CKINVDCx5p33_ASAP7_75t_R g1108 ( .A(n_225), .Y(n_1108) );
INVx1_ASAP7_75t_L g933 ( .A(n_227), .Y(n_933) );
INVx1_ASAP7_75t_L g266 ( .A(n_229), .Y(n_266) );
INVx1_ASAP7_75t_L g368 ( .A(n_230), .Y(n_368) );
BUFx3_ASAP7_75t_L g380 ( .A(n_230), .Y(n_380) );
BUFx3_ASAP7_75t_L g369 ( .A(n_231), .Y(n_369) );
INVx1_ASAP7_75t_L g397 ( .A(n_231), .Y(n_397) );
INVx1_ASAP7_75t_L g568 ( .A(n_233), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_255), .B(n_1129), .Y(n_234) );
BUFx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x4_ASAP7_75t_L g236 ( .A(n_237), .B(n_242), .Y(n_236) );
AND2x4_ASAP7_75t_L g1407 ( .A(n_237), .B(n_243), .Y(n_1407) );
NOR2xp33_ASAP7_75t_SL g237 ( .A(n_238), .B(n_240), .Y(n_237) );
INVx1_ASAP7_75t_SL g1414 ( .A(n_238), .Y(n_1414) );
NAND2xp5_ASAP7_75t_L g1419 ( .A(n_238), .B(n_240), .Y(n_1419) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g1413 ( .A(n_240), .B(n_1414), .Y(n_1413) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_244), .B(n_248), .Y(n_243) );
INVxp67_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
OR2x2_ASAP7_75t_L g718 ( .A(n_245), .B(n_447), .Y(n_718) );
OR2x6_ASAP7_75t_L g764 ( .A(n_245), .B(n_447), .Y(n_764) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g664 ( .A(n_246), .B(n_254), .Y(n_664) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g313 ( .A(n_247), .B(n_314), .Y(n_313) );
INVx8_ASAP7_75t_L g714 ( .A(n_248), .Y(n_714) );
OR2x6_ASAP7_75t_L g248 ( .A(n_249), .B(n_253), .Y(n_248) );
INVx1_ASAP7_75t_L g319 ( .A(n_249), .Y(n_319) );
OR2x2_ASAP7_75t_L g444 ( .A(n_249), .B(n_303), .Y(n_444) );
INVx2_ASAP7_75t_SL g467 ( .A(n_249), .Y(n_467) );
OR2x6_ASAP7_75t_L g717 ( .A(n_249), .B(n_708), .Y(n_717) );
INVx2_ASAP7_75t_SL g1085 ( .A(n_249), .Y(n_1085) );
BUFx6f_ASAP7_75t_L g1104 ( .A(n_249), .Y(n_1104) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
AND2x4_ASAP7_75t_L g271 ( .A(n_251), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g281 ( .A(n_251), .Y(n_281) );
AND2x2_ASAP7_75t_L g287 ( .A(n_251), .B(n_252), .Y(n_287) );
INVx2_ASAP7_75t_L g292 ( .A(n_251), .Y(n_292) );
INVx1_ASAP7_75t_L g326 ( .A(n_251), .Y(n_326) );
INVx2_ASAP7_75t_L g272 ( .A(n_252), .Y(n_272) );
INVx1_ASAP7_75t_L g294 ( .A(n_252), .Y(n_294) );
INVx1_ASAP7_75t_L g301 ( .A(n_252), .Y(n_301) );
INVx1_ASAP7_75t_L g325 ( .A(n_252), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_252), .B(n_292), .Y(n_334) );
AND2x4_ASAP7_75t_L g703 ( .A(n_253), .B(n_301), .Y(n_703) );
INVx2_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g704 ( .A(n_254), .B(n_705), .Y(n_704) );
OR2x2_ASAP7_75t_L g1013 ( .A(n_254), .B(n_705), .Y(n_1013) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_257), .B1(n_857), .B2(n_858), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
XNOR2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_524), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AO22x2_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_261), .B1(n_449), .B2(n_523), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_358), .Y(n_262) );
NOR3xp33_ASAP7_75t_L g263 ( .A(n_264), .B(n_295), .C(n_311), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_282), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_267), .B1(n_277), .B2(n_278), .Y(n_265) );
BUFx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
BUFx2_ASAP7_75t_L g455 ( .A(n_268), .Y(n_455) );
BUFx2_ASAP7_75t_L g1072 ( .A(n_268), .Y(n_1072) );
AND2x4_ASAP7_75t_L g268 ( .A(n_269), .B(n_273), .Y(n_268) );
INVx2_ASAP7_75t_L g781 ( .A(n_269), .Y(n_781) );
INVx1_ASAP7_75t_L g881 ( .A(n_269), .Y(n_881) );
INVx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx3_ASAP7_75t_L g478 ( .A(n_270), .Y(n_478) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_270), .Y(n_485) );
INVx3_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g339 ( .A(n_271), .Y(n_339) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_271), .Y(n_343) );
INVx1_ASAP7_75t_L g564 ( .A(n_271), .Y(n_564) );
AND2x4_ASAP7_75t_L g280 ( .A(n_272), .B(n_281), .Y(n_280) );
AND2x6_ASAP7_75t_L g278 ( .A(n_273), .B(n_279), .Y(n_278) );
AND2x4_ASAP7_75t_L g284 ( .A(n_273), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g289 ( .A(n_273), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_273), .B(n_290), .Y(n_1077) );
AND2x4_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx1_ASAP7_75t_L g354 ( .A(n_274), .Y(n_354) );
OR2x2_ASAP7_75t_L g595 ( .A(n_274), .B(n_371), .Y(n_595) );
INVx2_ASAP7_75t_L g553 ( .A(n_275), .Y(n_553) );
AND2x2_ASAP7_75t_L g560 ( .A(n_275), .B(n_291), .Y(n_560) );
AND2x4_ASAP7_75t_L g567 ( .A(n_275), .B(n_545), .Y(n_567) );
INVx1_ASAP7_75t_L g314 ( .A(n_276), .Y(n_314) );
INVx1_ASAP7_75t_L g356 ( .A(n_276), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_278), .A2(n_454), .B1(n_455), .B2(n_456), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_278), .A2(n_1071), .B1(n_1072), .B2(n_1073), .Y(n_1070) );
NAND2x1p5_ASAP7_75t_L g310 ( .A(n_279), .B(n_302), .Y(n_310) );
BUFx3_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
BUFx3_ASAP7_75t_L g548 ( .A(n_280), .Y(n_548) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_280), .Y(n_571) );
AND2x4_ASAP7_75t_L g698 ( .A(n_280), .B(n_699), .Y(n_698) );
BUFx6f_ASAP7_75t_L g771 ( .A(n_280), .Y(n_771) );
BUFx2_ASAP7_75t_L g951 ( .A(n_280), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_284), .B1(n_288), .B2(n_289), .Y(n_282) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_284), .A2(n_289), .B1(n_458), .B2(n_459), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_284), .A2(n_1075), .B1(n_1076), .B2(n_1077), .Y(n_1074) );
INVx2_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
INVx2_ASAP7_75t_SL g537 ( .A(n_286), .Y(n_537) );
INVx2_ASAP7_75t_L g667 ( .A(n_286), .Y(n_667) );
INVx3_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_287), .Y(n_545) );
INVx2_ASAP7_75t_SL g676 ( .A(n_290), .Y(n_676) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_291), .Y(n_541) );
BUFx2_ASAP7_75t_L g671 ( .A(n_291), .Y(n_671) );
AND2x4_ASAP7_75t_L g707 ( .A(n_291), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g774 ( .A(n_291), .Y(n_774) );
BUFx2_ASAP7_75t_L g779 ( .A(n_291), .Y(n_779) );
AND2x4_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
INVx1_ASAP7_75t_L g308 ( .A(n_292), .Y(n_308) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2x1_ASAP7_75t_SL g298 ( .A(n_299), .B(n_302), .Y(n_298) );
NAND2x1p5_ASAP7_75t_L g556 ( .A(n_299), .B(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
HB1xp67_ASAP7_75t_L g886 ( .A(n_301), .Y(n_886) );
NAND2x1p5_ASAP7_75t_L g306 ( .A(n_302), .B(n_307), .Y(n_306) );
INVx3_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g536 ( .A(n_304), .Y(n_536) );
BUFx4f_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx4f_ASAP7_75t_L g461 ( .A(n_306), .Y(n_461) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x6_ASAP7_75t_L g558 ( .A(n_308), .B(n_535), .Y(n_558) );
BUFx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx2_ASAP7_75t_L g1079 ( .A(n_310), .Y(n_1079) );
OAI33xp33_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_316), .A3(n_327), .B1(n_340), .B2(n_345), .B3(n_351), .Y(n_311) );
OAI33xp33_ASAP7_75t_L g462 ( .A1(n_312), .A2(n_351), .A3(n_463), .B1(n_471), .B2(n_479), .B3(n_487), .Y(n_462) );
INVx1_ASAP7_75t_L g1082 ( .A(n_312), .Y(n_1082) );
OR2x6_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
INVx1_ASAP7_75t_L g708 ( .A(n_314), .Y(n_708) );
INVx2_ASAP7_75t_L g362 ( .A(n_315), .Y(n_362) );
BUFx2_ASAP7_75t_L g659 ( .A(n_315), .Y(n_659) );
OAI22xp33_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_318), .B1(n_320), .B2(n_321), .Y(n_316) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g346 ( .A(n_319), .Y(n_346) );
BUFx3_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OAI21xp5_ASAP7_75t_L g876 ( .A1(n_322), .A2(n_877), .B(n_878), .Y(n_876) );
BUFx3_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g490 ( .A(n_323), .Y(n_490) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
AND2x2_ASAP7_75t_L g349 ( .A(n_325), .B(n_326), .Y(n_349) );
INVx1_ASAP7_75t_L g705 ( .A(n_326), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_329), .B1(n_335), .B2(n_336), .Y(n_327) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_329), .A2(n_341), .B1(n_342), .B2(n_344), .Y(n_340) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g473 ( .A(n_332), .Y(n_473) );
BUFx3_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g1094 ( .A(n_333), .Y(n_1094) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx2_ASAP7_75t_L g481 ( .A(n_334), .Y(n_481) );
INVx1_ASAP7_75t_L g1382 ( .A(n_334), .Y(n_1382) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OAI22xp5_ASAP7_75t_L g1396 ( .A1(n_338), .A2(n_1397), .B1(n_1398), .B2(n_1399), .Y(n_1396) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g711 ( .A(n_339), .Y(n_711) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_341), .A2(n_365), .B1(n_373), .B2(n_391), .C(n_398), .Y(n_364) );
INVx2_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
INVx4_ASAP7_75t_L g673 ( .A(n_343), .Y(n_673) );
BUFx3_ASAP7_75t_L g677 ( .A(n_343), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_344), .A2(n_347), .B1(n_433), .B2(n_438), .Y(n_432) );
OAI22xp33_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_347), .B1(n_348), .B2(n_350), .Y(n_345) );
OAI21xp5_ASAP7_75t_SL g891 ( .A1(n_348), .A2(n_892), .B(n_893), .Y(n_891) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g470 ( .A(n_349), .Y(n_470) );
BUFx2_ASAP7_75t_L g1088 ( .A(n_349), .Y(n_1088) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_350), .A2(n_411), .B1(n_420), .B2(n_425), .C(n_428), .Y(n_410) );
OAI33xp33_ASAP7_75t_L g1080 ( .A1(n_351), .A2(n_1081), .A3(n_1083), .B1(n_1090), .B2(n_1098), .B3(n_1102), .Y(n_1080) );
CKINVDCx8_ASAP7_75t_R g351 ( .A(n_352), .Y(n_351) );
NAND3xp33_ASAP7_75t_L g766 ( .A(n_352), .B(n_767), .C(n_772), .Y(n_766) );
NAND3xp33_ASAP7_75t_L g961 ( .A(n_352), .B(n_962), .C(n_964), .Y(n_961) );
NAND3xp33_ASAP7_75t_L g995 ( .A(n_352), .B(n_996), .C(n_998), .Y(n_995) );
INVx5_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx6_ASAP7_75t_L g679 ( .A(n_353), .Y(n_679) );
OR2x6_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
NAND2x1p5_ASAP7_75t_L g612 ( .A(n_354), .B(n_401), .Y(n_612) );
INVx2_ASAP7_75t_L g550 ( .A(n_355), .Y(n_550) );
BUFx2_ASAP7_75t_L g894 ( .A(n_355), .Y(n_894) );
NAND2x1p5_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_L g700 ( .A(n_356), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_363), .B1(n_441), .B2(n_442), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_359), .A2(n_442), .B1(n_493), .B2(n_522), .Y(n_492) );
AOI31xp33_ASAP7_75t_L g538 ( .A1(n_359), .A2(n_539), .A3(n_559), .B(n_566), .Y(n_538) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NOR2xp67_ASAP7_75t_L g532 ( .A(n_361), .B(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g579 ( .A(n_362), .B(n_580), .Y(n_579) );
AND2x4_ASAP7_75t_L g663 ( .A(n_362), .B(n_664), .Y(n_663) );
OR2x6_ASAP7_75t_L g682 ( .A(n_362), .B(n_683), .Y(n_682) );
AND2x4_ASAP7_75t_L g784 ( .A(n_362), .B(n_664), .Y(n_784) );
OR2x2_ASAP7_75t_L g833 ( .A(n_362), .B(n_683), .Y(n_833) );
BUFx2_ASAP7_75t_L g864 ( .A(n_362), .Y(n_864) );
NAND3xp33_ASAP7_75t_L g363 ( .A(n_364), .B(n_410), .C(n_432), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g494 ( .A1(n_365), .A2(n_482), .B1(n_495), .B2(n_501), .C(n_506), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g1110 ( .A1(n_365), .A2(n_1099), .B(n_1111), .Y(n_1110) );
AND2x4_ASAP7_75t_L g365 ( .A(n_366), .B(n_370), .Y(n_365) );
BUFx3_ASAP7_75t_L g392 ( .A(n_366), .Y(n_392) );
INVx1_ASAP7_75t_L g503 ( .A(n_366), .Y(n_503) );
INVx2_ASAP7_75t_SL g512 ( .A(n_366), .Y(n_512) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_367), .Y(n_413) );
INVx2_ASAP7_75t_SL g608 ( .A(n_367), .Y(n_608) );
AND2x6_ASAP7_75t_L g656 ( .A(n_367), .B(n_630), .Y(n_656) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_367), .Y(n_693) );
BUFx2_ASAP7_75t_L g791 ( .A(n_367), .Y(n_791) );
BUFx2_ASAP7_75t_L g798 ( .A(n_367), .Y(n_798) );
BUFx6f_ASAP7_75t_L g915 ( .A(n_367), .Y(n_915) );
AND2x4_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx1_ASAP7_75t_L g437 ( .A(n_368), .Y(n_437) );
INVx2_ASAP7_75t_L g378 ( .A(n_369), .Y(n_378) );
AND2x2_ASAP7_75t_L g384 ( .A(n_369), .B(n_380), .Y(n_384) );
AND2x4_ASAP7_75t_L g426 ( .A(n_370), .B(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
OR2x2_ASAP7_75t_L g434 ( .A(n_371), .B(n_435), .Y(n_434) );
OR2x2_ASAP7_75t_L g439 ( .A(n_371), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g402 ( .A(n_372), .Y(n_402) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g1006 ( .A(n_375), .Y(n_1006) );
INVx4_ASAP7_75t_L g1369 ( .A(n_375), .Y(n_1369) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g518 ( .A(n_376), .Y(n_518) );
INVx2_ASAP7_75t_L g654 ( .A(n_376), .Y(n_654) );
INVx2_ASAP7_75t_L g788 ( .A(n_376), .Y(n_788) );
INVx1_ASAP7_75t_L g796 ( .A(n_376), .Y(n_796) );
INVx2_ASAP7_75t_SL g1119 ( .A(n_376), .Y(n_1119) );
INVx6_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g422 ( .A(n_377), .Y(n_422) );
AND2x2_ASAP7_75t_L g448 ( .A(n_377), .B(n_401), .Y(n_448) );
BUFx2_ASAP7_75t_L g583 ( .A(n_377), .Y(n_583) );
AND2x4_ASAP7_75t_L g634 ( .A(n_377), .B(n_635), .Y(n_634) );
AND2x4_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx1_ASAP7_75t_L g409 ( .A(n_378), .Y(n_409) );
INVx1_ASAP7_75t_L g405 ( .A(n_379), .Y(n_405) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x4_ASAP7_75t_L g396 ( .A(n_380), .B(n_397), .Y(n_396) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_382), .Y(n_643) );
AND2x2_ASAP7_75t_L g844 ( .A(n_382), .B(n_630), .Y(n_844) );
HB1xp67_ASAP7_75t_L g980 ( .A(n_382), .Y(n_980) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g415 ( .A(n_383), .Y(n_415) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_383), .Y(n_431) );
INVx2_ASAP7_75t_L g585 ( .A(n_383), .Y(n_585) );
AND2x4_ASAP7_75t_L g628 ( .A(n_383), .B(n_629), .Y(n_628) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_384), .Y(n_427) );
BUFx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx2_ASAP7_75t_SL g500 ( .A(n_387), .Y(n_500) );
AND2x4_ASAP7_75t_L g590 ( .A(n_387), .B(n_447), .Y(n_590) );
AND2x4_ASAP7_75t_L g694 ( .A(n_387), .B(n_447), .Y(n_694) );
CKINVDCx5p33_ASAP7_75t_R g1120 ( .A(n_387), .Y(n_1120) );
AND2x4_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
AND2x4_ASAP7_75t_L g401 ( .A(n_388), .B(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g419 ( .A(n_389), .B(n_390), .Y(n_419) );
INVx1_ASAP7_75t_L g631 ( .A(n_389), .Y(n_631) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_389), .Y(n_636) );
INVx1_ASAP7_75t_L g640 ( .A(n_389), .Y(n_640) );
INVx1_ASAP7_75t_L g658 ( .A(n_390), .Y(n_658) );
BUFx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
OR2x6_ASAP7_75t_L g594 ( .A(n_395), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_396), .Y(n_424) );
INVx2_ASAP7_75t_L g440 ( .A(n_396), .Y(n_440) );
INVx1_ASAP7_75t_L g520 ( .A(n_396), .Y(n_520) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_396), .Y(n_589) );
INVx1_ASAP7_75t_L g436 ( .A(n_397), .Y(n_436) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x4_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
AND2x2_ASAP7_75t_L g407 ( .A(n_401), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g430 ( .A(n_401), .Y(n_430) );
AND2x4_ASAP7_75t_L g1113 ( .A(n_401), .B(n_403), .Y(n_1113) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g616 ( .A(n_404), .Y(n_616) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g648 ( .A(n_405), .Y(n_648) );
INVx2_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g508 ( .A(n_408), .Y(n_508) );
BUFx3_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AND2x6_ASAP7_75t_L g650 ( .A(n_409), .B(n_631), .Y(n_650) );
BUFx3_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g620 ( .A(n_415), .Y(n_620) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g515 ( .A(n_419), .Y(n_515) );
INVx1_ASAP7_75t_L g580 ( .A(n_419), .Y(n_580) );
INVx2_ASAP7_75t_L g683 ( .A(n_419), .Y(n_683) );
BUFx3_ASAP7_75t_L g1124 ( .A(n_419), .Y(n_1124) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_SL g587 ( .A(n_422), .Y(n_587) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AND2x6_ASAP7_75t_L g638 ( .A(n_424), .B(n_639), .Y(n_638) );
HB1xp67_ASAP7_75t_L g835 ( .A(n_424), .Y(n_835) );
INVx2_ASAP7_75t_L g1058 ( .A(n_424), .Y(n_1058) );
AOI221xp5_ASAP7_75t_L g509 ( .A1(n_425), .A2(n_428), .B1(n_491), .B2(n_510), .C(n_516), .Y(n_509) );
AOI221xp5_ASAP7_75t_L g1121 ( .A1(n_425), .A2(n_428), .B1(n_1106), .B2(n_1122), .C(n_1125), .Y(n_1121) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_427), .Y(n_514) );
INVx1_ASAP7_75t_L g839 ( .A(n_427), .Y(n_839) );
INVx1_ASAP7_75t_L g903 ( .A(n_427), .Y(n_903) );
BUFx4f_ASAP7_75t_L g1034 ( .A(n_427), .Y(n_1034) );
INVx2_ASAP7_75t_SL g1061 ( .A(n_427), .Y(n_1061) );
AND2x4_ASAP7_75t_L g428 ( .A(n_429), .B(n_431), .Y(n_428) );
INVx1_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g507 ( .A(n_430), .B(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g497 ( .A(n_431), .Y(n_497) );
INVx1_ASAP7_75t_L g687 ( .A(n_431), .Y(n_687) );
OAI21xp33_ASAP7_75t_L g939 ( .A1(n_431), .A2(n_629), .B(n_940), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_433), .A2(n_438), .B1(n_486), .B2(n_488), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_433), .A2(n_438), .B1(n_1101), .B2(n_1105), .Y(n_1126) );
INVx6_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g909 ( .A(n_435), .Y(n_909) );
OR2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
AND2x2_ASAP7_75t_L g600 ( .A(n_436), .B(n_437), .Y(n_600) );
INVx4_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g505 ( .A(n_440), .Y(n_505) );
AOI21xp33_ASAP7_75t_L g1107 ( .A1(n_442), .A2(n_1108), .B(n_1109), .Y(n_1107) );
INVx5_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AND2x4_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OR2x6_ASAP7_75t_L g531 ( .A(n_446), .B(n_532), .Y(n_531) );
AND2x4_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
INVx1_ASAP7_75t_L g523 ( .A(n_449), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_492), .Y(n_450) );
NOR3xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_460), .C(n_462), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_457), .Y(n_452) );
OAI22xp33_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B1(n_468), .B2(n_469), .Y(n_463) );
OAI22xp33_ASAP7_75t_L g487 ( .A1(n_465), .A2(n_488), .B1(n_489), .B2(n_491), .Y(n_487) );
BUFx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
OR2x6_ASAP7_75t_L g575 ( .A(n_470), .B(n_535), .Y(n_575) );
OR2x2_ASAP7_75t_L g1400 ( .A(n_470), .B(n_535), .Y(n_1400) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B1(n_474), .B2(n_475), .Y(n_471) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_478), .Y(n_542) );
INVx2_ASAP7_75t_L g776 ( .A(n_478), .Y(n_776) );
INVx2_ASAP7_75t_L g825 ( .A(n_478), .Y(n_825) );
INVx2_ASAP7_75t_L g828 ( .A(n_478), .Y(n_828) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_482), .B1(n_483), .B2(n_486), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g879 ( .A1(n_480), .A2(n_880), .B1(n_881), .B2(n_882), .Y(n_879) );
BUFx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g963 ( .A(n_485), .Y(n_963) );
INVx2_ASAP7_75t_SL g1097 ( .A(n_485), .Y(n_1097) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NAND3xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_509), .C(n_521), .Y(n_493) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g793 ( .A(n_505), .Y(n_793) );
OR2x6_ASAP7_75t_L g611 ( .A(n_508), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
BUFx2_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
HB1xp67_ASAP7_75t_L g916 ( .A(n_514), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g1373 ( .A(n_514), .B(n_621), .Y(n_1373) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
BUFx3_ASAP7_75t_L g685 ( .A(n_518), .Y(n_685) );
INVx1_ASAP7_75t_L g911 ( .A(n_519), .Y(n_911) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g922 ( .A(n_520), .Y(n_922) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_722), .B1(n_855), .B2(n_856), .Y(n_524) );
INVx2_ASAP7_75t_L g856 ( .A(n_525), .Y(n_856) );
AOI21x1_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_623), .B(n_721), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g721 ( .A(n_527), .B(n_624), .Y(n_721) );
XOR2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_622), .Y(n_527) );
NOR3xp33_ASAP7_75t_L g528 ( .A(n_529), .B(n_538), .C(n_576), .Y(n_528) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g1374 ( .A(n_531), .B(n_1375), .Y(n_1374) );
INVx1_ASAP7_75t_L g868 ( .A(n_533), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_537), .Y(n_533) );
AND2x2_ASAP7_75t_L g885 ( .A(n_534), .B(n_886), .Y(n_885) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g557 ( .A(n_535), .Y(n_557) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx2_ASAP7_75t_L g821 ( .A(n_537), .Y(n_821) );
AOI221xp5_ASAP7_75t_SL g539 ( .A1(n_540), .A2(n_543), .B1(n_551), .B2(n_554), .C(n_555), .Y(n_539) );
BUFx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_545), .Y(n_570) );
INVx3_ASAP7_75t_L g769 ( .A(n_545), .Y(n_769) );
AOI211xp5_ASAP7_75t_L g696 ( .A1(n_546), .A2(n_697), .B(n_698), .C(n_701), .Y(n_696) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g783 ( .A(n_547), .Y(n_783) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x4_ASAP7_75t_L g551 ( .A(n_548), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
AOI222xp33_ASAP7_75t_L g866 ( .A1(n_551), .A2(n_567), .B1(n_867), .B2(n_868), .C1(n_869), .C2(n_870), .Y(n_866) );
INVx8_ASAP7_75t_L g1378 ( .A(n_551), .Y(n_1378) );
AND2x4_ASAP7_75t_L g562 ( .A(n_552), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
CKINVDCx11_ASAP7_75t_R g888 ( .A(n_558), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_561), .B1(n_562), .B2(n_565), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_560), .A2(n_562), .B1(n_872), .B2(n_873), .Y(n_871) );
INVx3_ASAP7_75t_L g1402 ( .A(n_560), .Y(n_1402) );
INVx3_ASAP7_75t_L g1403 ( .A(n_562), .Y(n_1403) );
INVx1_ASAP7_75t_L g1002 ( .A(n_563), .Y(n_1002) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g573 ( .A(n_564), .Y(n_573) );
AOI221xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_568), .B1(n_569), .B2(n_572), .C(n_574), .Y(n_566) );
CKINVDCx6p67_ASAP7_75t_R g1388 ( .A(n_567), .Y(n_1388) );
INVx1_ASAP7_75t_L g1054 ( .A(n_570), .Y(n_1054) );
INVx2_ASAP7_75t_SL g669 ( .A(n_571), .Y(n_669) );
BUFx6f_ASAP7_75t_L g822 ( .A(n_571), .Y(n_822) );
NOR3xp33_ASAP7_75t_L g874 ( .A(n_574), .B(n_875), .C(n_889), .Y(n_874) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND4xp25_ASAP7_75t_L g576 ( .A(n_577), .B(n_591), .C(n_601), .D(n_609), .Y(n_576) );
AOI33xp33_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_581), .A3(n_582), .B1(n_586), .B2(n_588), .B3(n_590), .Y(n_577) );
NAND3xp33_ASAP7_75t_L g785 ( .A(n_578), .B(n_786), .C(n_790), .Y(n_785) );
NAND3xp33_ASAP7_75t_L g965 ( .A(n_578), .B(n_966), .C(n_967), .Y(n_965) );
NAND3xp33_ASAP7_75t_L g990 ( .A(n_578), .B(n_991), .C(n_992), .Y(n_990) );
INVx3_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx3_ASAP7_75t_L g789 ( .A(n_585), .Y(n_789) );
AND2x2_ASAP7_75t_L g603 ( .A(n_587), .B(n_604), .Y(n_603) );
BUFx6f_ASAP7_75t_L g689 ( .A(n_589), .Y(n_689) );
INVx1_ASAP7_75t_L g800 ( .A(n_590), .Y(n_800) );
AOI33xp33_ASAP7_75t_L g831 ( .A1(n_590), .A2(n_832), .A3(n_834), .B1(n_836), .B2(n_837), .B3(n_840), .Y(n_831) );
NAND3xp33_ASAP7_75t_L g968 ( .A(n_590), .B(n_969), .C(n_970), .Y(n_968) );
NAND3xp33_ASAP7_75t_L g1004 ( .A(n_590), .B(n_1005), .C(n_1007), .Y(n_1004) );
AOI33xp33_ASAP7_75t_L g1363 ( .A1(n_590), .A2(n_1364), .A3(n_1365), .B1(n_1366), .B2(n_1368), .B3(n_1370), .Y(n_1363) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_593), .B1(n_596), .B2(n_597), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g1352 ( .A1(n_593), .A2(n_597), .B1(n_1353), .B2(n_1354), .Y(n_1352) );
CKINVDCx6p67_ASAP7_75t_R g593 ( .A(n_594), .Y(n_593) );
OR2x6_ASAP7_75t_L g598 ( .A(n_595), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g604 ( .A(n_595), .Y(n_604) );
CKINVDCx6p67_ASAP7_75t_R g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g736 ( .A(n_600), .Y(n_736) );
INVx1_ASAP7_75t_L g920 ( .A(n_600), .Y(n_920) );
BUFx4f_ASAP7_75t_L g1116 ( .A(n_600), .Y(n_1116) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_603), .B1(n_605), .B2(n_606), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g1355 ( .A1(n_603), .A2(n_606), .B1(n_1356), .B2(n_1357), .Y(n_1355) );
AND2x2_ASAP7_75t_L g606 ( .A(n_604), .B(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g1008 ( .A(n_608), .Y(n_1008) );
AOI221xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_613), .B1(n_614), .B2(n_618), .C(n_619), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g1359 ( .A1(n_610), .A2(n_1360), .B1(n_1361), .B2(n_1362), .Y(n_1359) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx2_ASAP7_75t_SL g617 ( .A(n_612), .Y(n_617) );
INVx1_ASAP7_75t_L g621 ( .A(n_612), .Y(n_621) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g1361 ( .A(n_615), .Y(n_1361) );
NAND2x1p5_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g720 ( .A(n_625), .Y(n_720) );
AOI211x1_ASAP7_75t_SL g625 ( .A1(n_626), .A2(n_657), .B(n_660), .C(n_695), .Y(n_625) );
NAND4xp25_ASAP7_75t_L g626 ( .A(n_627), .B(n_632), .C(n_641), .D(n_651), .Y(n_626) );
BUFx2_ASAP7_75t_L g904 ( .A(n_627), .Y(n_904) );
NAND4xp25_ASAP7_75t_SL g1025 ( .A(n_627), .B(n_1026), .C(n_1029), .D(n_1032), .Y(n_1025) );
INVx5_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_628), .B(n_730), .Y(n_729) );
AOI211xp5_ASAP7_75t_L g842 ( .A1(n_628), .A2(n_843), .B(n_844), .C(n_845), .Y(n_842) );
AOI211xp5_ASAP7_75t_L g978 ( .A1(n_628), .A2(n_979), .B(n_980), .C(n_981), .Y(n_978) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B1(n_637), .B2(n_638), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_633), .A2(n_714), .B1(n_715), .B2(n_716), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_634), .A2(n_653), .B1(n_739), .B2(n_740), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_634), .A2(n_812), .B1(n_847), .B2(n_848), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_634), .A2(n_638), .B1(n_867), .B2(n_900), .Y(n_899) );
AOI221xp5_ASAP7_75t_L g934 ( .A1(n_634), .A2(n_656), .B1(n_935), .B2(n_936), .C(n_937), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_634), .A2(n_653), .B1(n_984), .B2(n_985), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_634), .A2(n_638), .B1(n_1030), .B2(n_1031), .Y(n_1029) );
AND2x4_ASAP7_75t_L g646 ( .A(n_635), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_638), .A2(n_656), .B1(n_742), .B2(n_743), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_638), .A2(n_656), .B1(n_850), .B2(n_851), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_638), .A2(n_653), .B1(n_932), .B2(n_933), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g986 ( .A1(n_638), .A2(n_656), .B1(n_987), .B2(n_988), .Y(n_986) );
AND2x4_ASAP7_75t_L g653 ( .A(n_639), .B(n_654), .Y(n_653) );
AND2x4_ASAP7_75t_L g848 ( .A(n_639), .B(n_654), .Y(n_848) );
INVx1_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g732 ( .A(n_640), .B(n_733), .Y(n_732) );
AOI222xp33_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_643), .B1(n_644), .B2(n_645), .C1(n_649), .C2(n_650), .Y(n_641) );
AOI222xp33_ASAP7_75t_L g901 ( .A1(n_645), .A2(n_650), .B1(n_884), .B2(n_887), .C1(n_892), .C2(n_902), .Y(n_901) );
BUFx4f_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g982 ( .A(n_646), .Y(n_982) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g733 ( .A(n_648), .Y(n_733) );
INVx3_ASAP7_75t_L g737 ( .A(n_650), .Y(n_737) );
AOI222xp33_ASAP7_75t_L g1032 ( .A1(n_650), .A2(n_1033), .B1(n_1034), .B2(n_1035), .C1(n_1036), .C2(n_1037), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B1(n_655), .B2(n_656), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g896 ( .A1(n_653), .A2(n_656), .B1(n_897), .B2(n_898), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_653), .A2(n_656), .B1(n_1027), .B2(n_1028), .Y(n_1026) );
BUFx6f_ASAP7_75t_L g744 ( .A(n_657), .Y(n_744) );
AO211x2_ASAP7_75t_L g976 ( .A1(n_657), .A2(n_977), .B(n_989), .C(n_1009), .Y(n_976) );
AND2x4_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
AND2x4_ASAP7_75t_L g853 ( .A(n_658), .B(n_659), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_680), .Y(n_660) );
AOI33xp33_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_665), .A3(n_670), .B1(n_674), .B2(n_678), .B3(n_679), .Y(n_661) );
AOI33xp33_ASAP7_75t_L g1048 ( .A1(n_662), .A2(n_679), .A3(n_1049), .B1(n_1050), .B2(n_1051), .B3(n_1052), .Y(n_1048) );
BUFx3_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NAND3xp33_ASAP7_75t_L g999 ( .A(n_663), .B(n_1000), .C(n_1003), .Y(n_999) );
INVx1_ASAP7_75t_L g1395 ( .A(n_664), .Y(n_1395) );
BUFx3_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AOI211xp5_ASAP7_75t_L g1010 ( .A1(n_668), .A2(n_698), .B(n_1011), .C(n_1012), .Y(n_1010) );
INVx2_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g752 ( .A(n_669), .Y(n_752) );
INVx2_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g890 ( .A(n_673), .Y(n_890) );
INVx3_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g1100 ( .A(n_677), .Y(n_1100) );
AOI33xp33_ASAP7_75t_L g819 ( .A1(n_679), .A2(n_784), .A3(n_820), .B1(n_823), .B2(n_826), .B3(n_829), .Y(n_819) );
AOI33xp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_684), .A3(n_688), .B1(n_690), .B2(n_691), .B3(n_694), .Y(n_680) );
AOI33xp33_ASAP7_75t_L g1055 ( .A1(n_681), .A2(n_1056), .A3(n_1059), .B1(n_1062), .B2(n_1063), .B3(n_1064), .Y(n_1055) );
CKINVDCx5p33_ASAP7_75t_R g681 ( .A(n_682), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g905 ( .A1(n_682), .A2(n_906), .B1(n_917), .B2(n_923), .Y(n_905) );
INVx2_ASAP7_75t_L g1364 ( .A(n_682), .Y(n_1364) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
BUFx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
BUFx4f_ASAP7_75t_L g993 ( .A(n_693), .Y(n_993) );
BUFx4f_ASAP7_75t_L g924 ( .A(n_694), .Y(n_924) );
BUFx4f_ASAP7_75t_L g1064 ( .A(n_694), .Y(n_1064) );
AOI31xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_706), .A3(n_713), .B(n_718), .Y(n_695) );
CKINVDCx11_ASAP7_75t_R g762 ( .A(n_698), .Y(n_762) );
AOI211xp5_ASAP7_75t_L g1039 ( .A1(n_698), .A2(n_959), .B(n_1040), .C(n_1041), .Y(n_1039) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVxp67_ASAP7_75t_L g759 ( .A(n_700), .Y(n_759) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g755 ( .A(n_703), .Y(n_755) );
AOI222xp33_ASAP7_75t_L g945 ( .A1(n_703), .A2(n_757), .B1(n_946), .B2(n_947), .C1(n_948), .C2(n_949), .Y(n_945) );
INVx1_ASAP7_75t_L g758 ( .A(n_705), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_709), .B1(n_710), .B2(n_712), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_707), .A2(n_747), .B1(n_748), .B2(n_749), .Y(n_746) );
AOI22xp5_ASAP7_75t_L g807 ( .A1(n_707), .A2(n_749), .B1(n_808), .B2(n_809), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_707), .A2(n_749), .B1(n_943), .B2(n_944), .Y(n_942) );
AOI22xp33_ASAP7_75t_SL g1014 ( .A1(n_707), .A2(n_710), .B1(n_1015), .B2(n_1016), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_707), .A2(n_749), .B1(n_1043), .B2(n_1044), .Y(n_1042) );
AND2x4_ASAP7_75t_L g710 ( .A(n_708), .B(n_711), .Y(n_710) );
AND2x4_ASAP7_75t_L g749 ( .A(n_708), .B(n_711), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_714), .A2(n_716), .B1(n_740), .B2(n_761), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_714), .A2(n_811), .B1(n_812), .B2(n_813), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_714), .A2(n_813), .B1(n_935), .B2(n_953), .Y(n_952) );
AOI22xp33_ASAP7_75t_SL g1017 ( .A1(n_714), .A2(n_716), .B1(n_985), .B2(n_1018), .Y(n_1017) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_714), .A2(n_813), .B1(n_1030), .B2(n_1046), .Y(n_1045) );
INVx5_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx4_ASAP7_75t_L g813 ( .A(n_717), .Y(n_813) );
INVx1_ASAP7_75t_L g855 ( .A(n_722), .Y(n_855) );
AO22x1_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_724), .B1(n_802), .B2(n_854), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g801 ( .A(n_727), .Y(n_801) );
AOI221x1_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_744), .B1(n_745), .B2(n_763), .C(n_765), .Y(n_727) );
NAND3xp33_ASAP7_75t_L g728 ( .A(n_729), .B(n_738), .C(n_741), .Y(n_728) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g938 ( .A(n_732), .Y(n_938) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
AOI221x1_ASAP7_75t_SL g863 ( .A1(n_744), .A2(n_864), .B1(n_865), .B2(n_895), .C(n_905), .Y(n_863) );
AOI221x1_ASAP7_75t_L g929 ( .A1(n_744), .A2(n_763), .B1(n_930), .B2(n_941), .C(n_954), .Y(n_929) );
AOI211x1_ASAP7_75t_L g1024 ( .A1(n_744), .A2(n_1025), .B(n_1038), .C(n_1047), .Y(n_1024) );
NAND4xp25_ASAP7_75t_SL g745 ( .A(n_746), .B(n_750), .C(n_760), .D(n_762), .Y(n_745) );
AOI222xp33_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_752), .B1(n_753), .B2(n_754), .C1(n_756), .C2(n_757), .Y(n_750) );
AOI222xp33_ASAP7_75t_L g814 ( .A1(n_752), .A2(n_754), .B1(n_757), .B2(n_815), .C1(n_816), .C2(n_817), .Y(n_814) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
AND2x4_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
NAND4xp25_ASAP7_75t_SL g806 ( .A(n_762), .B(n_807), .C(n_810), .D(n_814), .Y(n_806) );
NAND4xp25_ASAP7_75t_SL g941 ( .A(n_762), .B(n_942), .C(n_945), .D(n_952), .Y(n_941) );
AOI211xp5_ASAP7_75t_L g805 ( .A1(n_763), .A2(n_806), .B(n_818), .C(n_841), .Y(n_805) );
CKINVDCx16_ASAP7_75t_R g763 ( .A(n_764), .Y(n_763) );
AOI31xp33_ASAP7_75t_L g1009 ( .A1(n_764), .A2(n_1010), .A3(n_1014), .B(n_1017), .Y(n_1009) );
AOI31xp33_ASAP7_75t_L g1038 ( .A1(n_764), .A2(n_1039), .A3(n_1042), .B(n_1045), .Y(n_1038) );
NAND4xp25_ASAP7_75t_L g765 ( .A(n_766), .B(n_777), .C(n_785), .D(n_794), .Y(n_765) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
HB1xp67_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
BUFx2_ASAP7_75t_L g830 ( .A(n_771), .Y(n_830) );
INVx2_ASAP7_75t_SL g960 ( .A(n_771), .Y(n_960) );
INVx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
NAND3xp33_ASAP7_75t_L g777 ( .A(n_778), .B(n_782), .C(n_784), .Y(n_777) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
NAND3xp33_ASAP7_75t_L g955 ( .A(n_784), .B(n_956), .C(n_958), .Y(n_955) );
BUFx6f_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g994 ( .A(n_793), .Y(n_994) );
NAND3xp33_ASAP7_75t_L g794 ( .A(n_795), .B(n_797), .C(n_799), .Y(n_794) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g854 ( .A(n_802), .Y(n_854) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
XNOR2xp5_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .Y(n_803) );
OAI22xp5_ASAP7_75t_L g1179 ( .A1(n_804), .A2(n_1180), .B1(n_1181), .B2(n_1182), .Y(n_1179) );
NAND2xp5_ASAP7_75t_SL g818 ( .A(n_819), .B(n_831), .Y(n_818) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx2_ASAP7_75t_L g997 ( .A(n_825), .Y(n_997) );
INVx2_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx2_ASAP7_75t_SL g957 ( .A(n_828), .Y(n_957) );
INVx1_ASAP7_75t_SL g832 ( .A(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
AOI31xp33_ASAP7_75t_SL g841 ( .A1(n_842), .A2(n_846), .A3(n_849), .B(n_852), .Y(n_841) );
INVx1_ASAP7_75t_SL g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
XNOR2xp5_ASAP7_75t_L g858 ( .A(n_859), .B(n_1021), .Y(n_858) );
AOI22xp5_ASAP7_75t_L g859 ( .A1(n_860), .A2(n_974), .B1(n_1019), .B2(n_1020), .Y(n_859) );
INVx1_ASAP7_75t_L g1019 ( .A(n_860), .Y(n_1019) );
AOI22xp5_ASAP7_75t_L g860 ( .A1(n_861), .A2(n_862), .B1(n_927), .B2(n_973), .Y(n_860) );
INVx2_ASAP7_75t_SL g861 ( .A(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g926 ( .A(n_863), .Y(n_926) );
CKINVDCx8_ASAP7_75t_R g1128 ( .A(n_864), .Y(n_1128) );
NAND3xp33_ASAP7_75t_L g865 ( .A(n_866), .B(n_871), .C(n_874), .Y(n_865) );
OAI221xp5_ASAP7_75t_L g917 ( .A1(n_869), .A2(n_870), .B1(n_908), .B2(n_918), .C(n_921), .Y(n_917) );
OAI21xp5_ASAP7_75t_SL g875 ( .A1(n_876), .A2(n_879), .B(n_883), .Y(n_875) );
OAI221xp5_ASAP7_75t_L g906 ( .A1(n_882), .A2(n_907), .B1(n_910), .B2(n_911), .C(n_912), .Y(n_906) );
AOI22xp5_ASAP7_75t_L g883 ( .A1(n_884), .A2(n_885), .B1(n_887), .B2(n_888), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g1386 ( .A1(n_885), .A2(n_888), .B1(n_1360), .B2(n_1362), .Y(n_1386) );
NAND4xp25_ASAP7_75t_SL g895 ( .A(n_896), .B(n_899), .C(n_901), .D(n_904), .Y(n_895) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
BUFx2_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
INVx2_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx2_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
INVx2_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
CKINVDCx5p33_ASAP7_75t_R g923 ( .A(n_924), .Y(n_923) );
HB1xp67_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
INVx1_ASAP7_75t_L g973 ( .A(n_928), .Y(n_973) );
INVx1_ASAP7_75t_L g972 ( .A(n_929), .Y(n_972) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_931), .B(n_934), .Y(n_930) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
NAND4xp25_ASAP7_75t_L g954 ( .A(n_955), .B(n_961), .C(n_965), .D(n_968), .Y(n_954) );
INVx2_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
INVx1_ASAP7_75t_L g1020 ( .A(n_974), .Y(n_1020) );
HB1xp67_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
NAND3xp33_ASAP7_75t_L g977 ( .A(n_978), .B(n_983), .C(n_986), .Y(n_977) );
INVx1_ASAP7_75t_L g1036 ( .A(n_982), .Y(n_1036) );
NAND4xp25_ASAP7_75t_L g989 ( .A(n_990), .B(n_995), .C(n_999), .D(n_1004), .Y(n_989) );
INVx1_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1002), .Y(n_1384) );
HB1xp67_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
XNOR2xp5_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1065), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_1048), .B(n_1055), .Y(n_1047) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
INVx2_ASAP7_75t_L g1060 ( .A(n_1061), .Y(n_1060) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1061), .Y(n_1367) );
XNOR2x1_ASAP7_75t_L g1065 ( .A(n_1066), .B(n_1067), .Y(n_1065) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1107), .Y(n_1067) );
NOR3xp33_ASAP7_75t_SL g1068 ( .A(n_1069), .B(n_1078), .C(n_1080), .Y(n_1068) );
NAND2xp5_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1074), .Y(n_1069) );
OAI211xp5_ASAP7_75t_L g1114 ( .A1(n_1073), .A2(n_1115), .B(n_1117), .C(n_1118), .Y(n_1114) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
OAI22xp33_ASAP7_75t_L g1083 ( .A1(n_1084), .A2(n_1086), .B1(n_1087), .B2(n_1089), .Y(n_1083) );
INVx3_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
OAI22xp33_ASAP7_75t_L g1102 ( .A1(n_1087), .A2(n_1103), .B1(n_1105), .B2(n_1106), .Y(n_1102) );
OAI221xp5_ASAP7_75t_L g1389 ( .A1(n_1087), .A2(n_1390), .B1(n_1391), .B2(n_1393), .C(n_1394), .Y(n_1389) );
INVx2_ASAP7_75t_L g1087 ( .A(n_1088), .Y(n_1087) );
OAI22xp5_ASAP7_75t_L g1090 ( .A1(n_1091), .A2(n_1092), .B1(n_1095), .B2(n_1096), .Y(n_1090) );
OAI22xp5_ASAP7_75t_L g1098 ( .A1(n_1092), .A2(n_1099), .B1(n_1100), .B2(n_1101), .Y(n_1098) );
INVx2_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
INVx2_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
BUFx2_ASAP7_75t_L g1103 ( .A(n_1104), .Y(n_1103) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1104), .Y(n_1392) );
AOI31xp33_ASAP7_75t_L g1109 ( .A1(n_1110), .A2(n_1121), .A3(n_1126), .B(n_1127), .Y(n_1109) );
INVx1_ASAP7_75t_SL g1112 ( .A(n_1113), .Y(n_1112) );
INVx2_ASAP7_75t_SL g1115 ( .A(n_1116), .Y(n_1115) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
OAI31xp33_ASAP7_75t_L g1376 ( .A1(n_1127), .A2(n_1377), .A3(n_1387), .B(n_1401), .Y(n_1376) );
INVx2_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
OAI21xp33_ASAP7_75t_SL g1129 ( .A1(n_1130), .A2(n_1343), .B(n_1345), .Y(n_1129) );
NOR2x1_ASAP7_75t_L g1130 ( .A(n_1131), .B(n_1309), .Y(n_1130) );
NAND2xp5_ASAP7_75t_L g1131 ( .A(n_1132), .B(n_1260), .Y(n_1131) );
NOR4xp25_ASAP7_75t_L g1132 ( .A(n_1133), .B(n_1202), .C(n_1222), .D(n_1238), .Y(n_1132) );
AOI21xp33_ASAP7_75t_L g1133 ( .A1(n_1134), .A2(n_1186), .B(n_1190), .Y(n_1133) );
OR2x2_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1155), .Y(n_1134) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_1135), .B(n_1187), .Y(n_1266) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1135), .Y(n_1304) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1136), .Y(n_1264) );
NAND2xp5_ASAP7_75t_L g1267 ( .A(n_1136), .B(n_1268), .Y(n_1267) );
NAND2xp5_ASAP7_75t_L g1323 ( .A(n_1136), .B(n_1324), .Y(n_1323) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1136), .Y(n_1334) );
HB1xp67_ASAP7_75t_L g1136 ( .A(n_1137), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1137), .B(n_1209), .Y(n_1208) );
INVx2_ASAP7_75t_SL g1221 ( .A(n_1137), .Y(n_1221) );
OR2x2_ASAP7_75t_L g1236 ( .A(n_1137), .B(n_1209), .Y(n_1236) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1138), .Y(n_1200) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1138), .Y(n_1253) );
BUFx3_ASAP7_75t_L g1344 ( .A(n_1138), .Y(n_1344) );
AND2x4_ASAP7_75t_L g1138 ( .A(n_1139), .B(n_1142), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1139), .B(n_1142), .Y(n_1166) );
HB1xp67_ASAP7_75t_L g1418 ( .A(n_1139), .Y(n_1418) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
AND2x4_ASAP7_75t_L g1144 ( .A(n_1140), .B(n_1142), .Y(n_1144) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1141), .Y(n_1140) );
NAND2xp5_ASAP7_75t_L g1150 ( .A(n_1141), .B(n_1151), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1143), .Y(n_1151) );
INVx2_ASAP7_75t_L g1176 ( .A(n_1144), .Y(n_1176) );
INVx1_ASAP7_75t_SL g1181 ( .A(n_1144), .Y(n_1181) );
OAI22xp33_ASAP7_75t_L g1145 ( .A1(n_1146), .A2(n_1147), .B1(n_1152), .B2(n_1153), .Y(n_1145) );
OAI22xp5_ASAP7_75t_L g1183 ( .A1(n_1147), .A2(n_1153), .B1(n_1184), .B2(n_1185), .Y(n_1183) );
OAI22xp33_ASAP7_75t_L g1193 ( .A1(n_1147), .A2(n_1194), .B1(n_1195), .B2(n_1196), .Y(n_1193) );
BUFx3_ASAP7_75t_L g1257 ( .A(n_1147), .Y(n_1257) );
BUFx6f_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
OAI22xp5_ASAP7_75t_L g1168 ( .A1(n_1148), .A2(n_1153), .B1(n_1169), .B2(n_1170), .Y(n_1168) );
OR2x2_ASAP7_75t_L g1148 ( .A(n_1149), .B(n_1150), .Y(n_1148) );
OR2x2_ASAP7_75t_L g1153 ( .A(n_1149), .B(n_1154), .Y(n_1153) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1149), .Y(n_1162) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1150), .Y(n_1161) );
HB1xp67_ASAP7_75t_L g1417 ( .A(n_1151), .Y(n_1417) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1153), .Y(n_1197) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1154), .Y(n_1164) );
A2O1A1Ixp33_ASAP7_75t_L g1202 ( .A1(n_1155), .A2(n_1203), .B(n_1207), .C(n_1212), .Y(n_1202) );
NAND2xp5_ASAP7_75t_L g1155 ( .A(n_1156), .B(n_1171), .Y(n_1155) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_1156), .B(n_1206), .Y(n_1205) );
OAI21xp5_ASAP7_75t_L g1231 ( .A1(n_1156), .A2(n_1232), .B(n_1233), .Y(n_1231) );
NAND3xp33_ASAP7_75t_L g1286 ( .A(n_1156), .B(n_1244), .C(n_1287), .Y(n_1286) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
OR2x2_ASAP7_75t_L g1293 ( .A(n_1157), .B(n_1172), .Y(n_1293) );
OR2x2_ASAP7_75t_L g1314 ( .A(n_1157), .B(n_1178), .Y(n_1314) );
OR2x2_ASAP7_75t_L g1157 ( .A(n_1158), .B(n_1167), .Y(n_1157) );
AND2x2_ASAP7_75t_L g1189 ( .A(n_1158), .B(n_1167), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1158), .B(n_1215), .Y(n_1214) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1158), .Y(n_1226) );
O2A1O1Ixp33_ASAP7_75t_SL g1238 ( .A1(n_1158), .A2(n_1239), .B(n_1242), .C(n_1249), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1158), .B(n_1178), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_1159), .B(n_1165), .Y(n_1158) );
AND2x4_ASAP7_75t_L g1160 ( .A(n_1161), .B(n_1162), .Y(n_1160) );
AND2x4_ASAP7_75t_L g1163 ( .A(n_1162), .B(n_1164), .Y(n_1163) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1166), .Y(n_1180) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1167), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1167), .B(n_1177), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1248 ( .A(n_1167), .B(n_1226), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1167), .B(n_1171), .Y(n_1265) );
AOI32xp33_ASAP7_75t_L g1296 ( .A1(n_1167), .A2(n_1228), .A3(n_1280), .B1(n_1297), .B2(n_1298), .Y(n_1296) );
A2O1A1Ixp33_ASAP7_75t_L g1300 ( .A1(n_1167), .A2(n_1172), .B(n_1235), .C(n_1270), .Y(n_1300) );
NAND2xp5_ASAP7_75t_L g1316 ( .A(n_1171), .B(n_1189), .Y(n_1316) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1172), .B(n_1177), .Y(n_1171) );
NAND2xp5_ASAP7_75t_L g1188 ( .A(n_1172), .B(n_1189), .Y(n_1188) );
NOR2xp33_ASAP7_75t_L g1206 ( .A(n_1172), .B(n_1177), .Y(n_1206) );
INVx2_ASAP7_75t_L g1217 ( .A(n_1172), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1172), .B(n_1192), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_1172), .B(n_1241), .Y(n_1240) );
INVx4_ASAP7_75t_L g1278 ( .A(n_1172), .Y(n_1278) );
OR2x2_ASAP7_75t_L g1281 ( .A(n_1172), .B(n_1282), .Y(n_1281) );
NAND2xp5_ASAP7_75t_L g1288 ( .A(n_1172), .B(n_1283), .Y(n_1288) );
OR2x2_ASAP7_75t_L g1337 ( .A(n_1172), .B(n_1314), .Y(n_1337) );
AND2x6_ASAP7_75t_L g1172 ( .A(n_1173), .B(n_1174), .Y(n_1172) );
INVx2_ASAP7_75t_L g1175 ( .A(n_1176), .Y(n_1175) );
OAI22xp5_ASAP7_75t_L g1251 ( .A1(n_1176), .A2(n_1252), .B1(n_1253), .B2(n_1254), .Y(n_1251) );
NOR2xp33_ASAP7_75t_L g1187 ( .A(n_1177), .B(n_1188), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1177), .B(n_1214), .Y(n_1213) );
OR2x2_ASAP7_75t_L g1272 ( .A(n_1177), .B(n_1215), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1177), .B(n_1248), .Y(n_1306) );
CKINVDCx6p67_ASAP7_75t_R g1177 ( .A(n_1178), .Y(n_1177) );
OR2x2_ASAP7_75t_L g1225 ( .A(n_1178), .B(n_1226), .Y(n_1225) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1178), .B(n_1226), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1263 ( .A(n_1178), .B(n_1214), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1178), .B(n_1248), .Y(n_1270) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1178), .B(n_1189), .Y(n_1291) );
OAI211xp5_ASAP7_75t_SL g1295 ( .A1(n_1178), .A2(n_1223), .B(n_1296), .C(n_1300), .Y(n_1295) );
NAND2xp5_ASAP7_75t_L g1302 ( .A(n_1178), .B(n_1303), .Y(n_1302) );
OR2x6_ASAP7_75t_SL g1178 ( .A(n_1179), .B(n_1183), .Y(n_1178) );
OAI22xp5_ASAP7_75t_L g1198 ( .A1(n_1181), .A2(n_1199), .B1(n_1200), .B2(n_1201), .Y(n_1198) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_1189), .B(n_1278), .Y(n_1303) );
INVx1_ASAP7_75t_SL g1280 ( .A(n_1190), .Y(n_1280) );
INVx3_ASAP7_75t_L g1190 ( .A(n_1191), .Y(n_1190) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1191), .Y(n_1224) );
OR2x2_ASAP7_75t_L g1230 ( .A(n_1191), .B(n_1209), .Y(n_1230) );
NAND2xp5_ASAP7_75t_L g1249 ( .A(n_1191), .B(n_1250), .Y(n_1249) );
OAI211xp5_ASAP7_75t_L g1261 ( .A1(n_1191), .A2(n_1262), .B(n_1266), .C(n_1267), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1274 ( .A(n_1191), .B(n_1208), .Y(n_1274) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1191), .B(n_1221), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1191), .B(n_1244), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_1191), .B(n_1283), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1338 ( .A(n_1191), .B(n_1209), .Y(n_1338) );
INVx3_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1192), .B(n_1209), .Y(n_1308) );
OR2x2_ASAP7_75t_L g1341 ( .A(n_1192), .B(n_1236), .Y(n_1341) );
OR2x2_ASAP7_75t_L g1192 ( .A(n_1193), .B(n_1198), .Y(n_1192) );
HB1xp67_ASAP7_75t_L g1259 ( .A(n_1196), .Y(n_1259) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1204), .Y(n_1203) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
NOR2xp33_ASAP7_75t_L g1333 ( .A(n_1205), .B(n_1334), .Y(n_1333) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1208), .Y(n_1207) );
AOI221xp5_ASAP7_75t_L g1275 ( .A1(n_1208), .A2(n_1276), .B1(n_1279), .B2(n_1284), .C(n_1285), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1208), .B(n_1277), .Y(n_1297) );
OAI22xp5_ASAP7_75t_L g1310 ( .A1(n_1208), .A2(n_1311), .B1(n_1317), .B2(n_1320), .Y(n_1310) );
OR2x2_ASAP7_75t_L g1220 ( .A(n_1209), .B(n_1221), .Y(n_1220) );
AND2x2_ASAP7_75t_L g1241 ( .A(n_1209), .B(n_1221), .Y(n_1241) );
INVx2_ASAP7_75t_L g1244 ( .A(n_1209), .Y(n_1244) );
AND2x4_ASAP7_75t_L g1209 ( .A(n_1210), .B(n_1211), .Y(n_1209) );
OAI21xp5_ASAP7_75t_L g1212 ( .A1(n_1213), .A2(n_1216), .B(n_1219), .Y(n_1212) );
OAI22xp5_ASAP7_75t_L g1305 ( .A1(n_1213), .A2(n_1269), .B1(n_1278), .B2(n_1306), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1331 ( .A(n_1213), .B(n_1278), .Y(n_1331) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1214), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1276 ( .A(n_1214), .B(n_1277), .Y(n_1276) );
O2A1O1Ixp33_ASAP7_75t_L g1332 ( .A1(n_1216), .A2(n_1263), .B(n_1324), .C(n_1333), .Y(n_1332) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1217), .B(n_1218), .Y(n_1216) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1217), .B(n_1229), .Y(n_1228) );
NOR2xp33_ASAP7_75t_L g1243 ( .A(n_1217), .B(n_1244), .Y(n_1243) );
INVx2_ASAP7_75t_L g1269 ( .A(n_1217), .Y(n_1269) );
NAND2xp5_ASAP7_75t_L g1223 ( .A(n_1219), .B(n_1224), .Y(n_1223) );
INVx2_ASAP7_75t_L g1219 ( .A(n_1220), .Y(n_1219) );
INVx2_ASAP7_75t_SL g1283 ( .A(n_1221), .Y(n_1283) );
OAI221xp5_ASAP7_75t_L g1222 ( .A1(n_1223), .A2(n_1225), .B1(n_1227), .B2(n_1230), .C(n_1231), .Y(n_1222) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1225), .Y(n_1229) );
OAI211xp5_ASAP7_75t_SL g1285 ( .A1(n_1225), .A2(n_1230), .B(n_1286), .C(n_1289), .Y(n_1285) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1228), .Y(n_1227) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
NAND2xp5_ASAP7_75t_L g1234 ( .A(n_1235), .B(n_1237), .Y(n_1234) );
AND2x2_ASAP7_75t_L g1320 ( .A(n_1235), .B(n_1278), .Y(n_1320) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1236), .Y(n_1235) );
AOI22xp33_ASAP7_75t_L g1262 ( .A1(n_1236), .A2(n_1263), .B1(n_1264), .B2(n_1265), .Y(n_1262) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1241), .Y(n_1327) );
NAND2xp5_ASAP7_75t_L g1242 ( .A(n_1243), .B(n_1245), .Y(n_1242) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1244), .Y(n_1299) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_1246), .B(n_1247), .Y(n_1245) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1248), .Y(n_1247) );
CKINVDCx5p33_ASAP7_75t_R g1289 ( .A(n_1250), .Y(n_1289) );
OR2x6_ASAP7_75t_SL g1250 ( .A(n_1251), .B(n_1255), .Y(n_1250) );
OAI22xp5_ASAP7_75t_L g1255 ( .A1(n_1256), .A2(n_1257), .B1(n_1258), .B2(n_1259), .Y(n_1255) );
OAI32xp33_ASAP7_75t_L g1260 ( .A1(n_1261), .A2(n_1271), .A3(n_1289), .B1(n_1295), .B2(n_1301), .Y(n_1260) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1263), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1269), .B(n_1270), .Y(n_1268) );
OAI211xp5_ASAP7_75t_SL g1271 ( .A1(n_1272), .A2(n_1273), .B(n_1275), .C(n_1290), .Y(n_1271) );
OAI21xp33_ASAP7_75t_L g1336 ( .A1(n_1272), .A2(n_1278), .B(n_1337), .Y(n_1336) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1274), .Y(n_1273) );
NAND2xp5_ASAP7_75t_L g1342 ( .A(n_1274), .B(n_1291), .Y(n_1342) );
NAND2xp5_ASAP7_75t_L g1340 ( .A(n_1277), .B(n_1284), .Y(n_1340) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
NOR2xp33_ASAP7_75t_L g1279 ( .A(n_1280), .B(n_1281), .Y(n_1279) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1281), .Y(n_1325) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1288), .Y(n_1287) );
A2O1A1Ixp33_ASAP7_75t_SL g1309 ( .A1(n_1289), .A2(n_1310), .B(n_1321), .C(n_1335), .Y(n_1309) );
OAI21xp5_ASAP7_75t_L g1290 ( .A1(n_1291), .A2(n_1292), .B(n_1294), .Y(n_1290) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1293), .Y(n_1292) );
A2O1A1Ixp33_ASAP7_75t_L g1339 ( .A1(n_1293), .A2(n_1340), .B(n_1341), .C(n_1342), .Y(n_1339) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1299), .Y(n_1298) );
O2A1O1Ixp33_ASAP7_75t_SL g1301 ( .A1(n_1302), .A2(n_1304), .B(n_1305), .C(n_1307), .Y(n_1301) );
O2A1O1Ixp33_ASAP7_75t_L g1321 ( .A1(n_1306), .A2(n_1322), .B(n_1325), .C(n_1326), .Y(n_1321) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1308), .Y(n_1307) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
NOR2xp33_ASAP7_75t_L g1312 ( .A(n_1313), .B(n_1315), .Y(n_1312) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1314), .Y(n_1313) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1316), .Y(n_1315) );
NOR2xp33_ASAP7_75t_L g1317 ( .A(n_1318), .B(n_1319), .Y(n_1317) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1320), .Y(n_1319) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
A2O1A1Ixp33_ASAP7_75t_L g1326 ( .A1(n_1327), .A2(n_1328), .B(n_1330), .C(n_1332), .Y(n_1326) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1331), .Y(n_1330) );
AOI21xp5_ASAP7_75t_L g1335 ( .A1(n_1336), .A2(n_1338), .B(n_1339), .Y(n_1335) );
CKINVDCx5p33_ASAP7_75t_R g1343 ( .A(n_1344), .Y(n_1343) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1347), .Y(n_1346) );
HB1xp67_ASAP7_75t_L g1410 ( .A(n_1348), .Y(n_1410) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1349), .Y(n_1348) );
NAND3xp33_ASAP7_75t_L g1349 ( .A(n_1350), .B(n_1374), .C(n_1376), .Y(n_1349) );
NOR2xp33_ASAP7_75t_L g1350 ( .A(n_1351), .B(n_1358), .Y(n_1350) );
NAND2xp5_ASAP7_75t_L g1351 ( .A(n_1352), .B(n_1355), .Y(n_1351) );
OAI221xp5_ASAP7_75t_L g1379 ( .A1(n_1353), .A2(n_1357), .B1(n_1380), .B2(n_1383), .C(n_1385), .Y(n_1379) );
NAND3xp33_ASAP7_75t_L g1358 ( .A(n_1359), .B(n_1363), .C(n_1371), .Y(n_1358) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1372), .Y(n_1371) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1373), .Y(n_1372) );
BUFx2_ASAP7_75t_L g1380 ( .A(n_1381), .Y(n_1380) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1382), .Y(n_1381) );
INVx2_ASAP7_75t_L g1398 ( .A(n_1382), .Y(n_1398) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1384), .Y(n_1383) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1392), .Y(n_1391) );
INVx2_ASAP7_75t_L g1394 ( .A(n_1395), .Y(n_1394) );
BUFx2_ASAP7_75t_L g1404 ( .A(n_1405), .Y(n_1404) );
INVx1_ASAP7_75t_L g1405 ( .A(n_1406), .Y(n_1405) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1407), .Y(n_1406) );
INVxp67_ASAP7_75t_L g1408 ( .A(n_1409), .Y(n_1408) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1412), .Y(n_1411) );
CKINVDCx5p33_ASAP7_75t_R g1412 ( .A(n_1413), .Y(n_1412) );
A2O1A1Ixp33_ASAP7_75t_L g1415 ( .A1(n_1414), .A2(n_1416), .B(n_1418), .C(n_1419), .Y(n_1415) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
endmodule