module fake_jpeg_5185_n_261 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_261);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_261;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx2_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx11_ASAP7_75t_SL g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_38),
.Y(n_45)
);

INVx2_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_32),
.B(n_18),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_40),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_37),
.B(n_18),
.Y(n_61)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_39),
.B(n_20),
.Y(n_87)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_17),
.Y(n_51)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_29),
.B1(n_28),
.B2(n_27),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_47),
.A2(n_70),
.B1(n_17),
.B2(n_20),
.Y(n_93)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_50),
.Y(n_92)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_32),
.A2(n_29),
.B1(n_13),
.B2(n_28),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_52),
.A2(n_63),
.B(n_69),
.Y(n_98)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_57),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

CKINVDCx9p33_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g103 ( 
.A(n_56),
.Y(n_103)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_59),
.B(n_62),
.Y(n_114)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_64),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_65),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_40),
.B(n_30),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_25),
.B(n_27),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_25),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_66),
.B(n_81),
.Y(n_116)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_74),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_39),
.A2(n_12),
.B1(n_16),
.B2(n_19),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_41),
.A2(n_12),
.B1(n_16),
.B2(n_22),
.Y(n_70)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_37),
.B(n_22),
.Y(n_76)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_82),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_37),
.B(n_21),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_78),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_32),
.A2(n_21),
.B1(n_19),
.B2(n_30),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_1),
.B(n_4),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_37),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_80),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_32),
.B(n_30),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_37),
.B(n_30),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_85),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_37),
.B(n_24),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_23),
.Y(n_101)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_93),
.A2(n_107),
.B1(n_110),
.B2(n_79),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_81),
.A2(n_30),
.B1(n_17),
.B2(n_24),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_54),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_62),
.A2(n_24),
.B1(n_23),
.B2(n_3),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_102),
.A2(n_52),
.B1(n_69),
.B2(n_49),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_62),
.A2(n_24),
.B1(n_2),
.B2(n_3),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_81),
.A2(n_23),
.B1(n_2),
.B2(n_4),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_58),
.Y(n_122)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_125),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_121),
.A2(n_124),
.B1(n_127),
.B2(n_131),
.Y(n_163)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_45),
.B(n_59),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_123),
.A2(n_132),
.B(n_117),
.Y(n_154)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_48),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_129),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_98),
.A2(n_68),
.B1(n_73),
.B2(n_71),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_84),
.Y(n_128)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_128),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_84),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_130),
.B(n_145),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_93),
.A2(n_73),
.B1(n_71),
.B2(n_65),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_66),
.B(n_23),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_116),
.A2(n_88),
.B1(n_57),
.B2(n_46),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_134),
.A2(n_142),
.B1(n_144),
.B2(n_96),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_90),
.B(n_1),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_135),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_23),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_139),
.Y(n_158)
);

MAJx2_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_72),
.C(n_89),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_105),
.C(n_111),
.Y(n_168)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_97),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_140),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_72),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_103),
.Y(n_140)
);

NOR3xp33_ASAP7_75t_SL g141 ( 
.A(n_109),
.B(n_72),
.C(n_89),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_143),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_116),
.A2(n_46),
.B1(n_55),
.B2(n_7),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_100),
.A2(n_11),
.B1(n_6),
.B2(n_7),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_95),
.B(n_5),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_95),
.B(n_5),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_148),
.Y(n_162)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_92),
.Y(n_147)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_96),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_151),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_117),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_157),
.C(n_164),
.Y(n_187)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_154),
.A2(n_158),
.B(n_171),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_102),
.Y(n_157)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_167),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_105),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_90),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_125),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_103),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_172),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_144),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_132),
.A2(n_118),
.B(n_113),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_171),
.A2(n_120),
.B(n_133),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_111),
.C(n_96),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_133),
.A2(n_113),
.B1(n_91),
.B2(n_112),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_173),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_124),
.A2(n_91),
.B1(n_94),
.B2(n_108),
.Y(n_174)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_165),
.B(n_142),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_179),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_152),
.B(n_129),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_153),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_193),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_181),
.A2(n_190),
.B1(n_191),
.B2(n_184),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_152),
.B(n_129),
.Y(n_183)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_184),
.A2(n_186),
.B(n_188),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_127),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_172),
.C(n_163),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_154),
.A2(n_120),
.B(n_141),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_138),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_189),
.B(n_195),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

INVx3_ASAP7_75t_SL g212 ( 
.A(n_191),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_147),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_194),
.A2(n_150),
.B(n_162),
.Y(n_210)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_160),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_192),
.A2(n_163),
.B1(n_169),
.B2(n_174),
.Y(n_196)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_196),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_210),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_192),
.A2(n_131),
.B1(n_167),
.B2(n_158),
.Y(n_199)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_190),
.A2(n_168),
.B1(n_175),
.B2(n_155),
.Y(n_201)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_202),
.B(n_205),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_178),
.A2(n_175),
.B1(n_156),
.B2(n_159),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_195),
.B(n_156),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_207),
.B(n_211),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g208 ( 
.A(n_176),
.Y(n_208)
);

INVx13_ASAP7_75t_L g217 ( 
.A(n_208),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_194),
.C(n_183),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_187),
.C(n_179),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_185),
.A2(n_162),
.B1(n_155),
.B2(n_151),
.Y(n_211)
);

NAND3xp33_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_170),
.C(n_103),
.Y(n_213)
);

AO21x1_ASAP7_75t_L g216 ( 
.A1(n_213),
.A2(n_186),
.B(n_180),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_224),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_219),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_182),
.C(n_193),
.Y(n_219)
);

XNOR2x1_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_198),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_197),
.Y(n_232)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_212),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_225),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_214),
.A2(n_196),
.B1(n_200),
.B2(n_177),
.Y(n_227)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_224),
.B(n_204),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_233),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_225),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_232),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_214),
.A2(n_201),
.B1(n_199),
.B2(n_212),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_182),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_218),
.C(n_220),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_222),
.A2(n_215),
.B(n_226),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_200),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_234),
.A2(n_222),
.B1(n_226),
.B2(n_221),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_237),
.B(n_170),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_240),
.A2(n_217),
.B(n_208),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_208),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_243),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_217),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_219),
.C(n_210),
.Y(n_243)
);

AOI21xp33_ASAP7_75t_L g245 ( 
.A1(n_239),
.A2(n_206),
.B(n_230),
.Y(n_245)
);

AOI21x1_ASAP7_75t_L g251 ( 
.A1(n_245),
.A2(n_243),
.B(n_237),
.Y(n_251)
);

AOI322xp5_ASAP7_75t_L g246 ( 
.A1(n_244),
.A2(n_223),
.A3(n_236),
.B1(n_216),
.B2(n_232),
.C1(n_235),
.C2(n_206),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_250),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_249),
.C(n_238),
.Y(n_252)
);

AOI21x1_ASAP7_75t_L g256 ( 
.A1(n_251),
.A2(n_249),
.B(n_208),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_252),
.A2(n_242),
.B1(n_253),
.B2(n_247),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_149),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_115),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_255),
.A2(n_256),
.B(n_252),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_257),
.B(n_115),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_258),
.B(n_259),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_104),
.Y(n_261)
);


endmodule