module fake_jpeg_4045_n_326 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_48),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_16),
.Y(n_41)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_42),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_8),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_43),
.B(n_55),
.Y(n_100)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_0),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_52),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_57),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_24),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_28),
.B(n_0),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_17),
.B(n_8),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_17),
.B(n_7),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_56),
.B(n_23),
.Y(n_104)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_46),
.A2(n_21),
.B1(n_31),
.B2(n_35),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_59),
.A2(n_64),
.B1(n_83),
.B2(n_33),
.Y(n_133)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx5_ASAP7_75t_SL g123 ( 
.A(n_60),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_24),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_61),
.B(n_68),
.Y(n_129)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_63),
.B(n_71),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_39),
.A2(n_27),
.B1(n_21),
.B2(n_31),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_57),
.A2(n_21),
.B1(n_31),
.B2(n_20),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_69),
.A2(n_81),
.B1(n_85),
.B2(n_105),
.Y(n_114)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

CKINVDCx12_ASAP7_75t_R g72 ( 
.A(n_45),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_38),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_91),
.Y(n_107)
);

CKINVDCx12_ASAP7_75t_R g77 ( 
.A(n_41),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_77),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_41),
.B(n_30),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_78),
.B(n_88),
.Y(n_115)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_80),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_37),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_57),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_39),
.A2(n_26),
.B1(n_34),
.B2(n_22),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_86),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_48),
.A2(n_23),
.B1(n_20),
.B2(n_22),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_89),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_55),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_37),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_95),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_18),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_47),
.B(n_34),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_94),
.Y(n_111)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_35),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_97),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_53),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_101),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_51),
.B(n_26),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_38),
.Y(n_116)
);

AO22x2_ASAP7_75t_L g105 ( 
.A1(n_54),
.A2(n_19),
.B1(n_33),
.B2(n_36),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_105),
.A2(n_25),
.B1(n_30),
.B2(n_28),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_106),
.A2(n_121),
.B(n_127),
.C(n_87),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_38),
.B(n_18),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_108),
.A2(n_75),
.B(n_68),
.Y(n_142)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_113),
.Y(n_153)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_116),
.B(n_90),
.Y(n_151)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_118),
.B(n_135),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_105),
.A2(n_25),
.B1(n_18),
.B2(n_36),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_65),
.B(n_0),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_125),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_65),
.B(n_0),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g126 ( 
.A(n_105),
.B(n_1),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_132),
.C(n_83),
.Y(n_146)
);

NAND2xp33_ASAP7_75t_L g127 ( 
.A(n_65),
.B(n_36),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g130 ( 
.A1(n_99),
.A2(n_36),
.B1(n_33),
.B2(n_19),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_130),
.A2(n_99),
.B1(n_74),
.B2(n_73),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_76),
.B(n_33),
.C(n_3),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_137),
.B1(n_96),
.B2(n_80),
.Y(n_154)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_62),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_136),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_73),
.A2(n_15),
.B1(n_9),
.B2(n_10),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_141),
.Y(n_177)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_142),
.A2(n_170),
.B(n_115),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_123),
.Y(n_143)
);

CKINVDCx10_ASAP7_75t_R g191 ( 
.A(n_143),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_129),
.B(n_100),
.Y(n_144)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_145),
.A2(n_154),
.B1(n_155),
.B2(n_163),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_146),
.B(n_152),
.Y(n_196)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_148),
.B(n_150),
.Y(n_192)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_149),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_112),
.Y(n_150)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

OAI21xp33_ASAP7_75t_SL g152 ( 
.A1(n_127),
.A2(n_126),
.B(n_122),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_133),
.A2(n_60),
.B1(n_74),
.B2(n_102),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_156),
.Y(n_189)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_112),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_158),
.Y(n_178)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_107),
.B(n_78),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_161),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_160),
.A2(n_174),
.B1(n_128),
.B2(n_119),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_107),
.B(n_78),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_120),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_168),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_114),
.A2(n_102),
.B1(n_82),
.B2(n_92),
.Y(n_163)
);

INVx3_ASAP7_75t_SL g164 ( 
.A(n_130),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_164),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_126),
.A2(n_90),
.B1(n_103),
.B2(n_95),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_134),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_106),
.A2(n_103),
.B1(n_93),
.B2(n_98),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_121),
.A2(n_93),
.B1(n_70),
.B2(n_97),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_173),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_128),
.A2(n_62),
.B(n_86),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_138),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_115),
.A2(n_84),
.B1(n_9),
.B2(n_12),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_129),
.B(n_15),
.Y(n_175)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_175),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_182),
.A2(n_200),
.B1(n_156),
.B2(n_147),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_186),
.B(n_201),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_148),
.A2(n_125),
.B(n_126),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_187),
.B(n_193),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_190),
.B1(n_194),
.B2(n_198),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_142),
.A2(n_134),
.B(n_119),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_160),
.A2(n_130),
.B1(n_132),
.B2(n_111),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_130),
.B(n_138),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_195),
.A2(n_139),
.B(n_173),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_131),
.C(n_117),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_168),
.C(n_139),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_171),
.A2(n_111),
.B1(n_117),
.B2(n_113),
.Y(n_198)
);

AND2x6_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_131),
.Y(n_199)
);

XNOR2x1_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_140),
.Y(n_229)
);

OAI21x1_ASAP7_75t_R g200 ( 
.A1(n_164),
.A2(n_113),
.B(n_135),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_153),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_204),
.Y(n_223)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

NOR2x1p5_ASAP7_75t_SL g205 ( 
.A(n_164),
.B(n_1),
.Y(n_205)
);

OAI32xp33_ASAP7_75t_L g230 ( 
.A1(n_205),
.A2(n_157),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_146),
.A2(n_110),
.B1(n_118),
.B2(n_109),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_208),
.A2(n_163),
.B1(n_166),
.B2(n_167),
.Y(n_218)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_151),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_210),
.Y(n_226)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_161),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_211),
.B(n_214),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_196),
.C(n_180),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_203),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_215),
.B(n_216),
.Y(n_251)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_178),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_189),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_217),
.B(n_220),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_218),
.A2(n_219),
.B1(n_236),
.B2(n_207),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_190),
.A2(n_194),
.B1(n_179),
.B2(n_182),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_178),
.Y(n_220)
);

AO21x1_ASAP7_75t_L g244 ( 
.A1(n_221),
.A2(n_230),
.B(n_237),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_181),
.B(n_150),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_193),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

A2O1A1O1Ixp25_ASAP7_75t_L g227 ( 
.A1(n_187),
.A2(n_145),
.B(n_162),
.C(n_158),
.D(n_141),
.Y(n_227)
);

A2O1A1O1Ixp25_ASAP7_75t_L g257 ( 
.A1(n_227),
.A2(n_221),
.B(n_195),
.C(n_223),
.D(n_226),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_177),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_228),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_229),
.A2(n_199),
.B(n_206),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_149),
.Y(n_231)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_231),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_191),
.Y(n_232)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_191),
.B(n_147),
.Y(n_233)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_233),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_200),
.Y(n_235)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_192),
.A2(n_143),
.B(n_4),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_205),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_238),
.A2(n_257),
.B(n_259),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_239),
.A2(n_247),
.B1(n_220),
.B2(n_216),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_250),
.C(n_258),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_230),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_219),
.A2(n_179),
.B1(n_207),
.B2(n_184),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_213),
.B(n_196),
.C(n_180),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_234),
.A2(n_229),
.B(n_212),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_252),
.A2(n_253),
.B(n_237),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_234),
.A2(n_212),
.B(n_206),
.Y(n_253)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_218),
.B(n_197),
.C(n_208),
.Y(n_258)
);

NOR2xp67_ASAP7_75t_SL g259 ( 
.A(n_211),
.B(n_200),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_215),
.Y(n_260)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_260),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_222),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_264),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_263),
.A2(n_270),
.B1(n_261),
.B2(n_276),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_267),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_232),
.Y(n_267)
);

INVx13_ASAP7_75t_L g268 ( 
.A(n_248),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_240),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_217),
.Y(n_269)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_259),
.A2(n_235),
.B(n_184),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_270),
.A2(n_272),
.B(n_256),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_242),
.B(n_224),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_273),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_256),
.A2(n_186),
.B(n_225),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_258),
.C(n_243),
.Y(n_273)
);

NOR2xp67_ASAP7_75t_SL g274 ( 
.A(n_257),
.B(n_228),
.Y(n_274)
);

NOR3xp33_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_238),
.C(n_244),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_239),
.B(n_176),
.C(n_183),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_247),
.Y(n_287)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_277),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_241),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_285),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_280),
.A2(n_246),
.B(n_244),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_287),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_249),
.Y(n_285)
);

MAJx2_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_238),
.C(n_244),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_286),
.A2(n_261),
.B(n_263),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_268),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_254),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_290),
.B(n_265),
.C(n_273),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_293),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_265),
.C(n_271),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_294),
.A2(n_298),
.B(n_300),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_287),
.A2(n_266),
.B1(n_245),
.B2(n_246),
.Y(n_295)
);

AOI322xp5_ASAP7_75t_L g305 ( 
.A1(n_295),
.A2(n_280),
.A3(n_290),
.B1(n_278),
.B2(n_283),
.C1(n_275),
.C2(n_136),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_288),
.B(n_245),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_301),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_278),
.C(n_267),
.Y(n_298)
);

NAND4xp25_ASAP7_75t_SL g302 ( 
.A(n_282),
.B(n_214),
.C(n_240),
.D(n_249),
.Y(n_302)
);

INVx6_ASAP7_75t_L g307 ( 
.A(n_302),
.Y(n_307)
);

NOR2x1_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_286),
.Y(n_303)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_303),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_305),
.A2(n_308),
.B(n_294),
.Y(n_315)
);

AOI21x1_ASAP7_75t_L g308 ( 
.A1(n_293),
.A2(n_283),
.B(n_136),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_3),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_310),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_299),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_296),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_312),
.A2(n_313),
.B(n_318),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_305),
.A2(n_291),
.B1(n_298),
.B2(n_292),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_314),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_316),
.C(n_317),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_307),
.A2(n_13),
.B1(n_14),
.B2(n_136),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_13),
.Y(n_317)
);

AOI322xp5_ASAP7_75t_L g324 ( 
.A1(n_320),
.A2(n_322),
.A3(n_3),
.B1(n_4),
.B2(n_6),
.C1(n_297),
.C2(n_303),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_313),
.A2(n_309),
.B1(n_306),
.B2(n_304),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_319),
.A2(n_321),
.B1(n_14),
.B2(n_5),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_323),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_324),
.Y(n_326)
);


endmodule