module fake_aes_3558_n_32 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_32);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_32;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NAND2xp5_ASAP7_75t_L g11 ( .A(n_5), .B(n_9), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_3), .Y(n_12) );
NOR2xp33_ASAP7_75t_R g13 ( .A(n_2), .B(n_6), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_4), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_8), .B(n_7), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_12), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_14), .B(n_0), .Y(n_17) );
NOR3xp33_ASAP7_75t_SL g18 ( .A(n_15), .B(n_0), .C(n_1), .Y(n_18) );
BUFx8_ASAP7_75t_L g19 ( .A(n_16), .Y(n_19) );
INVx6_ASAP7_75t_L g20 ( .A(n_17), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
NAND2xp5_ASAP7_75t_SL g22 ( .A(n_20), .B(n_18), .Y(n_22) );
INVx1_ASAP7_75t_SL g23 ( .A(n_21), .Y(n_23) );
OR2x2_ASAP7_75t_L g24 ( .A(n_22), .B(n_19), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
INVxp33_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
NAND2xp5_ASAP7_75t_L g27 ( .A(n_25), .B(n_1), .Y(n_27) );
OAI21xp5_ASAP7_75t_L g28 ( .A1(n_25), .A2(n_11), .B(n_13), .Y(n_28) );
INVx1_ASAP7_75t_SL g29 ( .A(n_27), .Y(n_29) );
AND2x4_ASAP7_75t_L g30 ( .A(n_28), .B(n_2), .Y(n_30) );
CKINVDCx20_ASAP7_75t_R g31 ( .A(n_29), .Y(n_31) );
AOI322xp5_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_3), .A3(n_10), .B1(n_13), .B2(n_26), .C1(n_30), .C2(n_29), .Y(n_32) );
endmodule