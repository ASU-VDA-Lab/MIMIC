module fake_aes_391_n_26 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_26);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_26;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
NAND2xp5_ASAP7_75t_L g13 ( .A(n_4), .B(n_7), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_12), .Y(n_14) );
CKINVDCx20_ASAP7_75t_R g15 ( .A(n_6), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_3), .Y(n_16) );
AO21x2_ASAP7_75t_L g17 ( .A1(n_1), .A2(n_2), .B(n_10), .Y(n_17) );
OR2x2_ASAP7_75t_L g18 ( .A(n_17), .B(n_0), .Y(n_18) );
NOR2xp33_ASAP7_75t_L g19 ( .A(n_14), .B(n_0), .Y(n_19) );
NOR2xp33_ASAP7_75t_R g20 ( .A(n_18), .B(n_15), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
NOR4xp25_ASAP7_75t_L g22 ( .A(n_21), .B(n_19), .C(n_13), .D(n_17), .Y(n_22) );
AOI221xp5_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_16), .B1(n_1), .B2(n_8), .C(n_9), .Y(n_23) );
BUFx12f_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
NOR2x1p5_ASAP7_75t_L g25 ( .A(n_24), .B(n_5), .Y(n_25) );
NAND3xp33_ASAP7_75t_L g26 ( .A(n_25), .B(n_24), .C(n_11), .Y(n_26) );
endmodule