module fake_netlist_6_1199_n_1144 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1144);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1144;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_462;
wire n_1033;
wire n_607;
wire n_671;
wire n_726;
wire n_1052;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_988;
wire n_969;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_1132;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_1138;
wire n_893;
wire n_925;
wire n_485;
wire n_1099;
wire n_1026;
wire n_443;
wire n_1101;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_1127;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_1139;
wire n_222;
wire n_248;
wire n_300;
wire n_517;
wire n_718;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_544;
wire n_468;
wire n_1078;
wire n_504;
wire n_923;
wire n_314;
wire n_1140;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_1015;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_360;
wire n_977;
wire n_945;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_1143;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_761;
wire n_428;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_842;
wire n_525;
wire n_1116;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_886;
wire n_448;
wire n_844;
wire n_1017;
wire n_1004;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_901;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_1084;
wire n_460;
wire n_929;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_1121;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_962;
wire n_824;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_1142;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_981;
wire n_476;
wire n_880;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_409;
wire n_345;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_1141;
wire n_249;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_1125;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_518;
wire n_299;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1131;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_928;
wire n_835;
wire n_690;
wire n_850;
wire n_1089;
wire n_1135;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_1124;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_869;
wire n_351;
wire n_437;
wire n_1082;
wire n_259;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_1001;
wire n_827;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_1134;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_1129;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g218 ( 
.A(n_32),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_197),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_170),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_177),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_216),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_212),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_96),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_110),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_39),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_81),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_121),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_135),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_156),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_217),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_26),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_211),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_2),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_123),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_12),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_127),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_206),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_19),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_43),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_209),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_114),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_47),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_30),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_132),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_179),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_58),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_61),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_124),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_128),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_42),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_28),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_76),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_147),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_65),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_164),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_103),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_166),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_149),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_105),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_98),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_194),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_118),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_40),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_154),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_60),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_21),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_138),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_141),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_1),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_125),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_168),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_213),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_109),
.Y(n_274)
);

BUFx5_ASAP7_75t_L g275 ( 
.A(n_104),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_69),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_195),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_63),
.Y(n_278)
);

BUFx10_ASAP7_75t_L g279 ( 
.A(n_178),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_205),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_68),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_4),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_173),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_54),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_15),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_78),
.Y(n_286)
);

BUFx5_ASAP7_75t_L g287 ( 
.A(n_167),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_234),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_267),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_267),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_220),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_222),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_236),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_283),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_283),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_218),
.Y(n_296)
);

INVxp33_ASAP7_75t_SL g297 ( 
.A(n_232),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_221),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_279),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_270),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_279),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_282),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_223),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_224),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_226),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_235),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_242),
.Y(n_307)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_248),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_243),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_285),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_245),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_246),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_228),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_239),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_230),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_219),
.Y(n_316)
);

BUFx5_ASAP7_75t_L g317 ( 
.A(n_255),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_225),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_275),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_256),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_244),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_257),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_262),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_269),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_274),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_247),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_280),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_278),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_284),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_275),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_231),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_252),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_252),
.Y(n_333)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_241),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_227),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_287),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_229),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_324),
.B(n_241),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_332),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_333),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_318),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_318),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_318),
.Y(n_343)
);

OA21x2_ASAP7_75t_L g344 ( 
.A1(n_319),
.A2(n_336),
.B(n_330),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_318),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_319),
.Y(n_346)
);

OAI21x1_ASAP7_75t_L g347 ( 
.A1(n_330),
.A2(n_287),
.B(n_275),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_296),
.B(n_253),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_321),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_336),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_298),
.B(n_233),
.Y(n_351)
);

OA21x2_ASAP7_75t_L g352 ( 
.A1(n_337),
.A2(n_238),
.B(n_237),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_288),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_317),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_304),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_290),
.A2(n_240),
.B1(n_249),
.B2(n_250),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_305),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_317),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_317),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_290),
.A2(n_251),
.B1(n_254),
.B2(n_258),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_317),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_317),
.Y(n_362)
);

INVx2_ASAP7_75t_SL g363 ( 
.A(n_299),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_306),
.Y(n_364)
);

INVx5_ASAP7_75t_L g365 ( 
.A(n_317),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_307),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_317),
.Y(n_367)
);

INVxp33_ASAP7_75t_SL g368 ( 
.A(n_291),
.Y(n_368)
);

OA21x2_ASAP7_75t_L g369 ( 
.A1(n_309),
.A2(n_260),
.B(n_259),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_293),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_294),
.B(n_261),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_311),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_295),
.B(n_263),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_312),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_320),
.B(n_264),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_322),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_302),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_323),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_325),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_327),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_300),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_299),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_329),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_335),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_308),
.B(n_265),
.Y(n_385)
);

OA21x2_ASAP7_75t_L g386 ( 
.A1(n_289),
.A2(n_268),
.B(n_266),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_314),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_334),
.B(n_271),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_292),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_302),
.A2(n_276),
.B1(n_286),
.B2(n_281),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_310),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_301),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_349),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_344),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_344),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_390),
.B(n_303),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_344),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_338),
.B(n_334),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_373),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_344),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_346),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_341),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_377),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_338),
.B(n_313),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_346),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_350),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_341),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_390),
.B(n_315),
.Y(n_408)
);

CKINVDCx6p67_ASAP7_75t_R g409 ( 
.A(n_377),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_363),
.B(n_331),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_346),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_350),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_350),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_350),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_374),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_363),
.B(n_297),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_374),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_389),
.Y(n_418)
);

OR2x6_ASAP7_75t_L g419 ( 
.A(n_385),
.B(n_301),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_379),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_379),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_379),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_341),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_379),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_374),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_376),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_376),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_341),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_385),
.B(n_310),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_376),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_378),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_392),
.B(n_272),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_368),
.B(n_273),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_392),
.B(n_375),
.Y(n_434)
);

INVx2_ASAP7_75t_SL g435 ( 
.A(n_371),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_341),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_356),
.B(n_326),
.Y(n_437)
);

AOI21x1_ASAP7_75t_L g438 ( 
.A1(n_347),
.A2(n_287),
.B(n_275),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_378),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_378),
.Y(n_440)
);

BUFx10_ASAP7_75t_L g441 ( 
.A(n_375),
.Y(n_441)
);

BUFx10_ASAP7_75t_L g442 ( 
.A(n_375),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_391),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_383),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_383),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_383),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_356),
.B(n_316),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_341),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_372),
.Y(n_449)
);

NAND2xp33_ASAP7_75t_SL g450 ( 
.A(n_360),
.B(n_381),
.Y(n_450)
);

BUFx10_ASAP7_75t_L g451 ( 
.A(n_375),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_342),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_392),
.B(n_277),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_373),
.B(n_275),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g455 ( 
.A(n_387),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_372),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_342),
.Y(n_457)
);

INVxp33_ASAP7_75t_L g458 ( 
.A(n_387),
.Y(n_458)
);

OAI22xp33_ASAP7_75t_L g459 ( 
.A1(n_387),
.A2(n_328),
.B1(n_316),
.B2(n_2),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_380),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_380),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_342),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_355),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_392),
.B(n_275),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_342),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_342),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_355),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_342),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_458),
.B(n_386),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_455),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_455),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_435),
.B(n_360),
.Y(n_472)
);

AND2x6_ASAP7_75t_L g473 ( 
.A(n_394),
.B(n_359),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_418),
.B(n_328),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_449),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_449),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_399),
.B(n_384),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_394),
.A2(n_347),
.B(n_369),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_456),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_399),
.Y(n_480)
);

NOR2xp67_ASAP7_75t_L g481 ( 
.A(n_393),
.B(n_382),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_456),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_460),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_460),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_461),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_461),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_404),
.B(n_386),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_402),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_418),
.B(n_391),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_420),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_429),
.B(n_386),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_412),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_412),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_413),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_398),
.B(n_386),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_435),
.B(n_384),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_420),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_421),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_409),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_421),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_403),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_422),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_422),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_424),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_413),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_424),
.Y(n_506)
);

XNOR2x2_ASAP7_75t_L g507 ( 
.A(n_447),
.B(n_384),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_454),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_395),
.B(n_359),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_415),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_454),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_415),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_395),
.B(n_359),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_409),
.Y(n_514)
);

NAND2x1p5_ASAP7_75t_L g515 ( 
.A(n_397),
.B(n_347),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_417),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_443),
.Y(n_517)
);

INVxp33_ASAP7_75t_L g518 ( 
.A(n_437),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_414),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_397),
.B(n_359),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_414),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_417),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_419),
.B(n_416),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_400),
.B(n_369),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_425),
.Y(n_525)
);

NOR2xp67_ASAP7_75t_L g526 ( 
.A(n_433),
.B(n_388),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_406),
.Y(n_527)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_419),
.B(n_351),
.Y(n_528)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_450),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_396),
.B(n_351),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_408),
.B(n_388),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_SL g532 ( 
.A(n_459),
.B(n_287),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_419),
.B(n_364),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_425),
.Y(n_534)
);

XOR2x2_ASAP7_75t_L g535 ( 
.A(n_410),
.B(n_0),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_426),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_426),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_427),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_419),
.B(n_364),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_434),
.B(n_364),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_427),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_431),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_430),
.Y(n_543)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_419),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_453),
.B(n_369),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_430),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_440),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_440),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_441),
.B(n_353),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_432),
.B(n_369),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_444),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_444),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_400),
.B(n_431),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_445),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_508),
.B(n_441),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_517),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_490),
.Y(n_557)
);

INVx1_ASAP7_75t_SL g558 ( 
.A(n_501),
.Y(n_558)
);

AND2x2_ASAP7_75t_SL g559 ( 
.A(n_532),
.B(n_352),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_501),
.Y(n_560)
);

BUFx8_ASAP7_75t_L g561 ( 
.A(n_523),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_511),
.B(n_441),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_477),
.B(n_441),
.Y(n_563)
);

AND2x6_ASAP7_75t_SL g564 ( 
.A(n_530),
.B(n_353),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_497),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_530),
.B(n_442),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_480),
.B(n_442),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_496),
.B(n_442),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_480),
.B(n_442),
.Y(n_569)
);

A2O1A1Ixp33_ASAP7_75t_SL g570 ( 
.A1(n_491),
.A2(n_423),
.B(n_436),
.C(n_428),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_542),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_487),
.A2(n_451),
.B1(n_352),
.B2(n_439),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_495),
.A2(n_352),
.B1(n_439),
.B2(n_445),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_487),
.A2(n_451),
.B1(n_352),
.B2(n_464),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_481),
.B(n_451),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_507),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_470),
.B(n_370),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_SL g578 ( 
.A(n_532),
.B(n_451),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_475),
.B(n_406),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_469),
.A2(n_467),
.B1(n_463),
.B2(n_446),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_476),
.B(n_479),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_518),
.B(n_348),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_529),
.B(n_446),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_SL g584 ( 
.A1(n_529),
.A2(n_287),
.B1(n_348),
.B2(n_370),
.Y(n_584)
);

NAND3xp33_ASAP7_75t_L g585 ( 
.A(n_472),
.B(n_340),
.C(n_339),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_549),
.B(n_406),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_482),
.B(n_463),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_SL g588 ( 
.A(n_544),
.B(n_287),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_483),
.B(n_467),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_471),
.B(n_402),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_469),
.A2(n_457),
.B1(n_466),
.B2(n_465),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_498),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_528),
.B(n_402),
.Y(n_593)
);

NAND3xp33_ASAP7_75t_SL g594 ( 
.A(n_514),
.B(n_340),
.C(n_339),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_484),
.B(n_485),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_526),
.B(n_402),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_533),
.B(n_355),
.Y(n_597)
);

INVx1_ASAP7_75t_SL g598 ( 
.A(n_489),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_486),
.B(n_448),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_540),
.B(n_405),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_540),
.A2(n_405),
.B1(n_411),
.B2(n_401),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_500),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_539),
.B(n_402),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_SL g604 ( 
.A1(n_474),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_502),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_531),
.B(n_345),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_553),
.B(n_411),
.Y(n_607)
);

NAND2x1_ASAP7_75t_L g608 ( 
.A(n_473),
.B(n_423),
.Y(n_608)
);

INVx8_ASAP7_75t_L g609 ( 
.A(n_473),
.Y(n_609)
);

INVx5_ASAP7_75t_L g610 ( 
.A(n_473),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_544),
.B(n_423),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_550),
.A2(n_366),
.B1(n_357),
.B2(n_355),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_545),
.A2(n_401),
.B1(n_366),
.B2(n_357),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g614 ( 
.A(n_535),
.B(n_345),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_527),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_524),
.A2(n_452),
.B1(n_466),
.B2(n_465),
.Y(n_616)
);

AND2x6_ASAP7_75t_SL g617 ( 
.A(n_499),
.B(n_3),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_503),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_504),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_506),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_524),
.A2(n_448),
.B1(n_462),
.B2(n_457),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_553),
.B(n_428),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_509),
.B(n_428),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_510),
.A2(n_357),
.B1(n_355),
.B2(n_366),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_557),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_605),
.Y(n_626)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_560),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g628 ( 
.A(n_558),
.Y(n_628)
);

INVx5_ASAP7_75t_L g629 ( 
.A(n_609),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_609),
.Y(n_630)
);

OR2x2_ASAP7_75t_L g631 ( 
.A(n_558),
.B(n_492),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_571),
.B(n_493),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_L g633 ( 
.A1(n_559),
.A2(n_478),
.B(n_509),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_556),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_576),
.A2(n_516),
.B1(n_522),
.B2(n_512),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_578),
.A2(n_520),
.B(n_513),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_599),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_577),
.B(n_494),
.Y(n_638)
);

NAND2xp33_ASAP7_75t_SL g639 ( 
.A(n_575),
.B(n_488),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_599),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_577),
.B(n_505),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_578),
.A2(n_534),
.B1(n_536),
.B2(n_525),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_565),
.Y(n_643)
);

NAND2x2_ASAP7_75t_L g644 ( 
.A(n_614),
.B(n_438),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_582),
.B(n_513),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_592),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_561),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_566),
.B(n_520),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_602),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_606),
.B(n_478),
.Y(n_650)
);

NOR2x1_ASAP7_75t_L g651 ( 
.A(n_568),
.B(n_537),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_619),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_609),
.Y(n_653)
);

AND2x6_ASAP7_75t_L g654 ( 
.A(n_563),
.B(n_488),
.Y(n_654)
);

AND3x2_ASAP7_75t_SL g655 ( 
.A(n_604),
.B(n_521),
.C(n_519),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_581),
.A2(n_554),
.B1(n_552),
.B2(n_551),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_618),
.B(n_597),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_584),
.A2(n_548),
.B1(n_547),
.B2(n_546),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_608),
.Y(n_659)
);

INVxp67_ASAP7_75t_SL g660 ( 
.A(n_600),
.Y(n_660)
);

AND2x4_ASAP7_75t_L g661 ( 
.A(n_620),
.B(n_538),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_595),
.Y(n_662)
);

BUFx2_ASAP7_75t_L g663 ( 
.A(n_561),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_587),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_610),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_615),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_607),
.B(n_473),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_585),
.B(n_541),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_567),
.B(n_543),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_589),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_615),
.Y(n_671)
);

INVx3_ASAP7_75t_SL g672 ( 
.A(n_598),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_622),
.B(n_515),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_610),
.Y(n_674)
);

NOR3xp33_ASAP7_75t_SL g675 ( 
.A(n_594),
.B(n_4),
.C(n_5),
.Y(n_675)
);

NAND2xp33_ASAP7_75t_SL g676 ( 
.A(n_569),
.B(n_488),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_583),
.B(n_515),
.Y(n_677)
);

BUFx8_ASAP7_75t_L g678 ( 
.A(n_617),
.Y(n_678)
);

BUFx2_ASAP7_75t_L g679 ( 
.A(n_564),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_598),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_579),
.Y(n_681)
);

INVx4_ASAP7_75t_L g682 ( 
.A(n_610),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_610),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_623),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_586),
.B(n_452),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_580),
.B(n_462),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_588),
.A2(n_355),
.B1(n_357),
.B2(n_366),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_593),
.Y(n_688)
);

HB1xp67_ASAP7_75t_L g689 ( 
.A(n_628),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_645),
.B(n_662),
.Y(n_690)
);

OAI21x1_ASAP7_75t_L g691 ( 
.A1(n_636),
.A2(n_621),
.B(n_616),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_643),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_664),
.B(n_670),
.Y(n_693)
);

AOI21xp33_ASAP7_75t_L g694 ( 
.A1(n_650),
.A2(n_588),
.B(n_572),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_625),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_657),
.B(n_611),
.Y(n_696)
);

AO21x1_ASAP7_75t_L g697 ( 
.A1(n_676),
.A2(n_603),
.B(n_574),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_646),
.Y(n_698)
);

OAI21x1_ASAP7_75t_L g699 ( 
.A1(n_673),
.A2(n_591),
.B(n_573),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_648),
.A2(n_562),
.B(n_555),
.Y(n_700)
);

OAI21x1_ASAP7_75t_L g701 ( 
.A1(n_673),
.A2(n_438),
.B(n_596),
.Y(n_701)
);

OAI21xp5_ASAP7_75t_L g702 ( 
.A1(n_648),
.A2(n_612),
.B(n_613),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_657),
.B(n_660),
.Y(n_703)
);

NAND2xp33_ASAP7_75t_L g704 ( 
.A(n_630),
.B(n_601),
.Y(n_704)
);

OAI21x1_ASAP7_75t_L g705 ( 
.A1(n_685),
.A2(n_590),
.B(n_624),
.Y(n_705)
);

AO21x2_ASAP7_75t_L g706 ( 
.A1(n_633),
.A2(n_570),
.B(n_358),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_684),
.B(n_436),
.Y(n_707)
);

OAI21xp5_ASAP7_75t_L g708 ( 
.A1(n_633),
.A2(n_468),
.B(n_436),
.Y(n_708)
);

AOI21xp33_ASAP7_75t_L g709 ( 
.A1(n_651),
.A2(n_681),
.B(n_635),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_638),
.B(n_468),
.Y(n_710)
);

OAI21x1_ASAP7_75t_L g711 ( 
.A1(n_685),
.A2(n_468),
.B(n_358),
.Y(n_711)
);

AOI21xp33_ASAP7_75t_L g712 ( 
.A1(n_627),
.A2(n_366),
.B(n_357),
.Y(n_712)
);

OAI21x1_ASAP7_75t_L g713 ( 
.A1(n_686),
.A2(n_358),
.B(n_354),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_638),
.B(n_357),
.Y(n_714)
);

AO31x2_ASAP7_75t_L g715 ( 
.A1(n_686),
.A2(n_367),
.A3(n_362),
.B(n_361),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_680),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_641),
.B(n_366),
.Y(n_717)
);

AND3x4_ASAP7_75t_L g718 ( 
.A(n_647),
.B(n_5),
.C(n_6),
.Y(n_718)
);

INVx4_ASAP7_75t_L g719 ( 
.A(n_629),
.Y(n_719)
);

OAI21xp5_ASAP7_75t_L g720 ( 
.A1(n_667),
.A2(n_677),
.B(n_642),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_631),
.B(n_6),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_641),
.B(n_407),
.Y(n_722)
);

INVx4_ASAP7_75t_L g723 ( 
.A(n_629),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_665),
.Y(n_724)
);

AOI21x1_ASAP7_75t_SL g725 ( 
.A1(n_667),
.A2(n_7),
.B(n_8),
.Y(n_725)
);

AO31x2_ASAP7_75t_L g726 ( 
.A1(n_677),
.A2(n_367),
.A3(n_362),
.B(n_361),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_649),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_652),
.Y(n_728)
);

OAI21x1_ASAP7_75t_L g729 ( 
.A1(n_651),
.A2(n_361),
.B(n_354),
.Y(n_729)
);

AO31x2_ASAP7_75t_L g730 ( 
.A1(n_688),
.A2(n_367),
.A3(n_362),
.B(n_354),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_630),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_626),
.B(n_407),
.Y(n_732)
);

OAI21xp5_ASAP7_75t_L g733 ( 
.A1(n_642),
.A2(n_365),
.B(n_407),
.Y(n_733)
);

OAI21x1_ASAP7_75t_L g734 ( 
.A1(n_659),
.A2(n_407),
.B(n_343),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_639),
.A2(n_407),
.B(n_343),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_661),
.B(n_7),
.Y(n_736)
);

AND2x4_ASAP7_75t_L g737 ( 
.A(n_629),
.B(n_31),
.Y(n_737)
);

OAI21x1_ASAP7_75t_L g738 ( 
.A1(n_659),
.A2(n_343),
.B(n_34),
.Y(n_738)
);

A2O1A1Ixp33_ASAP7_75t_L g739 ( 
.A1(n_635),
.A2(n_343),
.B(n_9),
.C(n_10),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_682),
.A2(n_343),
.B(n_365),
.Y(n_740)
);

OAI21x1_ASAP7_75t_L g741 ( 
.A1(n_674),
.A2(n_343),
.B(n_35),
.Y(n_741)
);

INVx4_ASAP7_75t_L g742 ( 
.A(n_630),
.Y(n_742)
);

INVx1_ASAP7_75t_SL g743 ( 
.A(n_672),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_679),
.B(n_8),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_682),
.A2(n_365),
.B(n_36),
.Y(n_745)
);

AOI21xp33_ASAP7_75t_L g746 ( 
.A1(n_637),
.A2(n_9),
.B(n_10),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_634),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_658),
.A2(n_365),
.B(n_37),
.Y(n_748)
);

OAI21x1_ASAP7_75t_L g749 ( 
.A1(n_674),
.A2(n_38),
.B(n_33),
.Y(n_749)
);

OAI21x1_ASAP7_75t_L g750 ( 
.A1(n_711),
.A2(n_656),
.B(n_687),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_731),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_692),
.Y(n_752)
);

A2O1A1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_748),
.A2(n_675),
.B(n_669),
.C(n_661),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_716),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_695),
.Y(n_755)
);

A2O1A1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_702),
.A2(n_669),
.B(n_668),
.C(n_640),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_727),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_747),
.Y(n_758)
);

OAI21xp5_ASAP7_75t_L g759 ( 
.A1(n_700),
.A2(n_656),
.B(n_668),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_690),
.B(n_632),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_728),
.Y(n_761)
);

CKINVDCx20_ASAP7_75t_R g762 ( 
.A(n_743),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_SL g763 ( 
.A1(n_702),
.A2(n_683),
.B(n_665),
.Y(n_763)
);

AO31x2_ASAP7_75t_L g764 ( 
.A1(n_697),
.A2(n_671),
.A3(n_666),
.B(n_644),
.Y(n_764)
);

O2A1O1Ixp33_ASAP7_75t_L g765 ( 
.A1(n_739),
.A2(n_663),
.B(n_655),
.C(n_632),
.Y(n_765)
);

AO21x2_ASAP7_75t_L g766 ( 
.A1(n_694),
.A2(n_654),
.B(n_665),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_743),
.A2(n_654),
.B1(n_678),
.B2(n_653),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_694),
.A2(n_733),
.B(n_704),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_733),
.A2(n_683),
.B(n_654),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_696),
.B(n_653),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_731),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_703),
.A2(n_654),
.B1(n_678),
.B2(n_653),
.Y(n_772)
);

OR2x6_ASAP7_75t_L g773 ( 
.A(n_737),
.B(n_683),
.Y(n_773)
);

BUFx12f_ASAP7_75t_L g774 ( 
.A(n_731),
.Y(n_774)
);

OAI21xp33_ASAP7_75t_L g775 ( 
.A1(n_693),
.A2(n_11),
.B(n_12),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_721),
.B(n_11),
.Y(n_776)
);

AND2x4_ASAP7_75t_L g777 ( 
.A(n_742),
.B(n_41),
.Y(n_777)
);

OAI21xp5_ASAP7_75t_L g778 ( 
.A1(n_709),
.A2(n_365),
.B(n_13),
.Y(n_778)
);

NOR4xp25_ASAP7_75t_L g779 ( 
.A(n_746),
.B(n_13),
.C(n_14),
.D(n_15),
.Y(n_779)
);

INVx5_ASAP7_75t_L g780 ( 
.A(n_719),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_720),
.A2(n_365),
.B(n_45),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_689),
.B(n_14),
.Y(n_782)
);

OAI21x1_ASAP7_75t_L g783 ( 
.A1(n_713),
.A2(n_46),
.B(n_44),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_698),
.B(n_16),
.Y(n_784)
);

AO31x2_ASAP7_75t_L g785 ( 
.A1(n_735),
.A2(n_120),
.A3(n_215),
.B(n_214),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_736),
.B(n_16),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_724),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_L g788 ( 
.A1(n_718),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_788)
);

OA21x2_ASAP7_75t_L g789 ( 
.A1(n_691),
.A2(n_49),
.B(n_48),
.Y(n_789)
);

INVxp67_ASAP7_75t_SL g790 ( 
.A(n_722),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_720),
.A2(n_365),
.B(n_51),
.Y(n_791)
);

AOI21x1_ASAP7_75t_L g792 ( 
.A1(n_699),
.A2(n_126),
.B(n_210),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_709),
.A2(n_122),
.B(n_208),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_714),
.B(n_17),
.Y(n_794)
);

BUFx8_ASAP7_75t_L g795 ( 
.A(n_737),
.Y(n_795)
);

NAND3xp33_ASAP7_75t_SL g796 ( 
.A(n_744),
.B(n_18),
.C(n_20),
.Y(n_796)
);

BUFx2_ASAP7_75t_L g797 ( 
.A(n_724),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_707),
.Y(n_798)
);

AOI221xp5_ASAP7_75t_L g799 ( 
.A1(n_712),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.C(n_23),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_SL g800 ( 
.A1(n_719),
.A2(n_130),
.B(n_207),
.Y(n_800)
);

OAI21x1_ASAP7_75t_L g801 ( 
.A1(n_729),
.A2(n_129),
.B(n_204),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_742),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_732),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_717),
.B(n_22),
.Y(n_804)
);

AO31x2_ASAP7_75t_L g805 ( 
.A1(n_745),
.A2(n_119),
.A3(n_203),
.B(n_202),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_710),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_806)
);

OAI21xp33_ASAP7_75t_L g807 ( 
.A1(n_708),
.A2(n_24),
.B(n_25),
.Y(n_807)
);

OAI21xp5_ASAP7_75t_L g808 ( 
.A1(n_705),
.A2(n_26),
.B(n_27),
.Y(n_808)
);

OAI21x1_ASAP7_75t_L g809 ( 
.A1(n_734),
.A2(n_133),
.B(n_201),
.Y(n_809)
);

A2O1A1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_738),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_810)
);

OAI21xp5_ASAP7_75t_L g811 ( 
.A1(n_701),
.A2(n_29),
.B(n_30),
.Y(n_811)
);

INVx3_ASAP7_75t_L g812 ( 
.A(n_723),
.Y(n_812)
);

AO31x2_ASAP7_75t_L g813 ( 
.A1(n_706),
.A2(n_50),
.A3(n_52),
.B(n_53),
.Y(n_813)
);

A2O1A1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_749),
.A2(n_55),
.B(n_56),
.C(n_57),
.Y(n_814)
);

AO31x2_ASAP7_75t_L g815 ( 
.A1(n_706),
.A2(n_59),
.A3(n_62),
.B(n_64),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_772),
.A2(n_723),
.B1(n_708),
.B2(n_740),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_754),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_796),
.A2(n_741),
.B1(n_725),
.B2(n_726),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_775),
.A2(n_807),
.B1(n_799),
.B2(n_788),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_751),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_755),
.Y(n_821)
);

INVx4_ASAP7_75t_SL g822 ( 
.A(n_774),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_762),
.A2(n_66),
.B1(n_67),
.B2(n_70),
.Y(n_823)
);

INVx4_ASAP7_75t_SL g824 ( 
.A(n_802),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_752),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_SL g826 ( 
.A1(n_778),
.A2(n_715),
.B1(n_726),
.B2(n_730),
.Y(n_826)
);

BUFx4f_ASAP7_75t_SL g827 ( 
.A(n_795),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_757),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_761),
.Y(n_829)
);

INVx5_ASAP7_75t_L g830 ( 
.A(n_780),
.Y(n_830)
);

BUFx2_ASAP7_75t_L g831 ( 
.A(n_797),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_790),
.Y(n_832)
);

INVx2_ASAP7_75t_SL g833 ( 
.A(n_751),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_758),
.Y(n_834)
);

INVx6_ASAP7_75t_L g835 ( 
.A(n_771),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_771),
.Y(n_836)
);

CKINVDCx11_ASAP7_75t_R g837 ( 
.A(n_773),
.Y(n_837)
);

OAI22xp5_ASAP7_75t_L g838 ( 
.A1(n_767),
.A2(n_715),
.B1(n_726),
.B2(n_730),
.Y(n_838)
);

OAI22xp33_ASAP7_75t_L g839 ( 
.A1(n_760),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_753),
.A2(n_715),
.B1(n_730),
.B2(n_77),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_765),
.A2(n_74),
.B1(n_75),
.B2(n_79),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_SL g842 ( 
.A1(n_779),
.A2(n_80),
.B1(n_82),
.B2(n_83),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_803),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_794),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_813),
.Y(n_845)
);

BUFx8_ASAP7_75t_SL g846 ( 
.A(n_770),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_787),
.Y(n_847)
);

OAI22xp33_ASAP7_75t_L g848 ( 
.A1(n_786),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_798),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_764),
.Y(n_850)
);

BUFx5_ASAP7_75t_L g851 ( 
.A(n_792),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_804),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_806),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_764),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_811),
.A2(n_97),
.B1(n_99),
.B2(n_100),
.Y(n_855)
);

OAI22xp33_ASAP7_75t_L g856 ( 
.A1(n_776),
.A2(n_101),
.B1(n_102),
.B2(n_106),
.Y(n_856)
);

INVx1_ASAP7_75t_SL g857 ( 
.A(n_782),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_773),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_780),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_764),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_781),
.A2(n_107),
.B1(n_108),
.B2(n_111),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_756),
.B(n_112),
.Y(n_862)
);

BUFx2_ASAP7_75t_L g863 ( 
.A(n_812),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_780),
.Y(n_864)
);

CKINVDCx6p67_ASAP7_75t_R g865 ( 
.A(n_777),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_784),
.Y(n_866)
);

BUFx3_ASAP7_75t_L g867 ( 
.A(n_777),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_SL g868 ( 
.A1(n_768),
.A2(n_113),
.B1(n_115),
.B2(n_116),
.Y(n_868)
);

OAI22xp33_ASAP7_75t_L g869 ( 
.A1(n_791),
.A2(n_117),
.B1(n_131),
.B2(n_134),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_759),
.A2(n_136),
.B1(n_137),
.B2(n_139),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_766),
.Y(n_871)
);

AOI22xp5_ASAP7_75t_L g872 ( 
.A1(n_793),
.A2(n_140),
.B1(n_142),
.B2(n_143),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_821),
.Y(n_873)
);

CKINVDCx20_ASAP7_75t_R g874 ( 
.A(n_846),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_828),
.Y(n_875)
);

CKINVDCx6p67_ASAP7_75t_R g876 ( 
.A(n_834),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_850),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_829),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_845),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_854),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_845),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_860),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_843),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_832),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_871),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_849),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_830),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_825),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_866),
.B(n_808),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_830),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_831),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_851),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_859),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_851),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_851),
.Y(n_895)
);

INVx1_ASAP7_75t_SL g896 ( 
.A(n_817),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_857),
.B(n_763),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_851),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_838),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_851),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_847),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_859),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_826),
.Y(n_903)
);

AO21x2_ASAP7_75t_L g904 ( 
.A1(n_840),
.A2(n_769),
.B(n_810),
.Y(n_904)
);

AOI21x1_ASAP7_75t_L g905 ( 
.A1(n_862),
.A2(n_789),
.B(n_783),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_818),
.B(n_815),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_830),
.Y(n_907)
);

HB1xp67_ASAP7_75t_L g908 ( 
.A(n_863),
.Y(n_908)
);

OR2x6_ASAP7_75t_L g909 ( 
.A(n_816),
.B(n_800),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_859),
.Y(n_910)
);

OAI21x1_ASAP7_75t_L g911 ( 
.A1(n_861),
.A2(n_750),
.B(n_801),
.Y(n_911)
);

OAI21x1_ASAP7_75t_L g912 ( 
.A1(n_841),
.A2(n_809),
.B(n_789),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_868),
.B(n_815),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_864),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_864),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_864),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_858),
.Y(n_917)
);

BUFx2_ASAP7_75t_L g918 ( 
.A(n_858),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_858),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_885),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_877),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_879),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_907),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_877),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_877),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_892),
.B(n_813),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_899),
.B(n_813),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_899),
.B(n_785),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_882),
.Y(n_929)
);

BUFx2_ASAP7_75t_L g930 ( 
.A(n_907),
.Y(n_930)
);

AO21x2_ASAP7_75t_L g931 ( 
.A1(n_892),
.A2(n_869),
.B(n_814),
.Y(n_931)
);

OA21x2_ASAP7_75t_L g932 ( 
.A1(n_912),
.A2(n_819),
.B(n_855),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_896),
.B(n_837),
.Y(n_933)
);

AO21x2_ASAP7_75t_L g934 ( 
.A1(n_892),
.A2(n_872),
.B(n_848),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_879),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_882),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_881),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_881),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_873),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_884),
.B(n_842),
.Y(n_940)
);

AO21x2_ASAP7_75t_L g941 ( 
.A1(n_894),
.A2(n_856),
.B(n_839),
.Y(n_941)
);

INVxp67_ASAP7_75t_L g942 ( 
.A(n_891),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_873),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_875),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_882),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_875),
.Y(n_946)
);

AO21x2_ASAP7_75t_L g947 ( 
.A1(n_894),
.A2(n_823),
.B(n_785),
.Y(n_947)
);

AO21x2_ASAP7_75t_L g948 ( 
.A1(n_894),
.A2(n_898),
.B(n_900),
.Y(n_948)
);

OR2x2_ASAP7_75t_L g949 ( 
.A(n_886),
.B(n_833),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_923),
.B(n_895),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_939),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_923),
.B(n_895),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_930),
.B(n_895),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_930),
.B(n_917),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_942),
.B(n_898),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_939),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_920),
.B(n_908),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_921),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_949),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_921),
.B(n_898),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_949),
.B(n_878),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_922),
.B(n_917),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_926),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_943),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_921),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_943),
.B(n_878),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_944),
.Y(n_967)
);

OR2x2_ASAP7_75t_L g968 ( 
.A(n_924),
.B(n_903),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_924),
.B(n_900),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_944),
.B(n_903),
.Y(n_970)
);

AOI221xp5_ASAP7_75t_L g971 ( 
.A1(n_940),
.A2(n_897),
.B1(n_889),
.B2(n_906),
.C(n_913),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_922),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_971),
.A2(n_909),
.B1(n_913),
.B2(n_932),
.Y(n_973)
);

OR2x2_ASAP7_75t_L g974 ( 
.A(n_968),
.B(n_946),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_963),
.B(n_948),
.Y(n_975)
);

NAND3xp33_ASAP7_75t_L g976 ( 
.A(n_970),
.B(n_932),
.C(n_928),
.Y(n_976)
);

INVx1_ASAP7_75t_SL g977 ( 
.A(n_957),
.Y(n_977)
);

BUFx2_ASAP7_75t_L g978 ( 
.A(n_954),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_972),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_958),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_951),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_956),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_964),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_967),
.Y(n_984)
);

BUFx2_ASAP7_75t_L g985 ( 
.A(n_954),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_963),
.B(n_948),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_966),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_981),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_978),
.B(n_963),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_985),
.B(n_963),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_977),
.B(n_963),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_987),
.B(n_933),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_982),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_979),
.B(n_983),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_984),
.B(n_959),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_974),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_974),
.B(n_955),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_980),
.Y(n_998)
);

OR2x2_ASAP7_75t_L g999 ( 
.A(n_973),
.B(n_968),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_991),
.B(n_955),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_989),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_988),
.B(n_980),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_992),
.B(n_876),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_991),
.B(n_954),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_989),
.B(n_950),
.Y(n_1005)
);

OR2x2_ASAP7_75t_L g1006 ( 
.A(n_999),
.B(n_976),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_993),
.Y(n_1007)
);

AO221x2_ASAP7_75t_L g1008 ( 
.A1(n_1001),
.A2(n_996),
.B1(n_998),
.B2(n_992),
.C(n_876),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_1004),
.Y(n_1009)
);

OR2x2_ASAP7_75t_L g1010 ( 
.A(n_1006),
.B(n_994),
.Y(n_1010)
);

OAI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_1003),
.A2(n_909),
.B1(n_990),
.B2(n_932),
.Y(n_1011)
);

AO221x2_ASAP7_75t_L g1012 ( 
.A1(n_1007),
.A2(n_1002),
.B1(n_1003),
.B2(n_998),
.C(n_874),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_1005),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_1000),
.Y(n_1014)
);

NOR2x1_ASAP7_75t_L g1015 ( 
.A(n_1002),
.B(n_994),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_1015),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1010),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_1014),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_1009),
.B(n_990),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_1013),
.B(n_994),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_1012),
.B(n_1008),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_1011),
.A2(n_995),
.B1(n_909),
.B2(n_932),
.Y(n_1022)
);

OAI21x1_ASAP7_75t_L g1023 ( 
.A1(n_1015),
.A2(n_997),
.B(n_986),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_1015),
.Y(n_1024)
);

INVx1_ASAP7_75t_SL g1025 ( 
.A(n_1010),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1015),
.Y(n_1026)
);

OAI211xp5_ASAP7_75t_L g1027 ( 
.A1(n_1024),
.A2(n_870),
.B(n_918),
.C(n_852),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_SL g1028 ( 
.A(n_1025),
.B(n_827),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1025),
.Y(n_1029)
);

AOI221xp5_ASAP7_75t_L g1030 ( 
.A1(n_1016),
.A2(n_986),
.B1(n_975),
.B2(n_906),
.C(n_961),
.Y(n_1030)
);

INVxp67_ASAP7_75t_L g1031 ( 
.A(n_1018),
.Y(n_1031)
);

OAI322xp33_ASAP7_75t_L g1032 ( 
.A1(n_1021),
.A2(n_975),
.A3(n_917),
.B1(n_919),
.B2(n_946),
.C1(n_937),
.C2(n_935),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_1026),
.A2(n_909),
.B1(n_918),
.B2(n_865),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1017),
.B(n_962),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1020),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1020),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_1029),
.B(n_1019),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1031),
.B(n_1023),
.Y(n_1038)
);

OAI31xp33_ASAP7_75t_L g1039 ( 
.A1(n_1028),
.A2(n_1027),
.A3(n_1033),
.B(n_1035),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_1036),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_1034),
.A2(n_1022),
.B1(n_909),
.B2(n_919),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_1030),
.B(n_822),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_1032),
.B(n_962),
.Y(n_1043)
);

OAI221xp5_ASAP7_75t_L g1044 ( 
.A1(n_1028),
.A2(n_844),
.B1(n_853),
.B2(n_867),
.C(n_919),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_1029),
.B(n_822),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1029),
.Y(n_1046)
);

AOI221xp5_ASAP7_75t_SL g1047 ( 
.A1(n_1038),
.A2(n_915),
.B1(n_910),
.B2(n_916),
.C(n_893),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1046),
.B(n_1045),
.Y(n_1048)
);

O2A1O1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_1039),
.A2(n_941),
.B(n_904),
.C(n_887),
.Y(n_1049)
);

NAND3xp33_ASAP7_75t_SL g1050 ( 
.A(n_1037),
.B(n_824),
.C(n_907),
.Y(n_1050)
);

A2O1A1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_1045),
.A2(n_902),
.B(n_890),
.C(n_887),
.Y(n_1051)
);

AOI221xp5_ASAP7_75t_L g1052 ( 
.A1(n_1040),
.A2(n_941),
.B1(n_916),
.B2(n_915),
.C(n_910),
.Y(n_1052)
);

NOR2x1_ASAP7_75t_L g1053 ( 
.A(n_1042),
.B(n_1043),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_1041),
.A2(n_941),
.B(n_934),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_1044),
.B(n_962),
.Y(n_1055)
);

INVx2_ASAP7_75t_SL g1056 ( 
.A(n_1048),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_1053),
.B(n_836),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_1055),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_1050),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1049),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1047),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_1051),
.B(n_950),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1054),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_1052),
.Y(n_1064)
);

INVx1_ASAP7_75t_SL g1065 ( 
.A(n_1048),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_1064),
.A2(n_890),
.B(n_902),
.C(n_914),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1056),
.Y(n_1067)
);

AOI211x1_ASAP7_75t_L g1068 ( 
.A1(n_1060),
.A2(n_953),
.B(n_952),
.C(n_969),
.Y(n_1068)
);

AND2x2_ASAP7_75t_SL g1069 ( 
.A(n_1057),
.B(n_1059),
.Y(n_1069)
);

NOR3xp33_ASAP7_75t_L g1070 ( 
.A(n_1065),
.B(n_1058),
.C(n_1059),
.Y(n_1070)
);

NOR3x1_ASAP7_75t_L g1071 ( 
.A(n_1063),
.B(n_824),
.C(n_937),
.Y(n_1071)
);

NOR2xp67_ASAP7_75t_L g1072 ( 
.A(n_1061),
.B(n_144),
.Y(n_1072)
);

NAND4xp75_ASAP7_75t_L g1073 ( 
.A(n_1062),
.B(n_914),
.C(n_952),
.D(n_953),
.Y(n_1073)
);

NAND3x1_ASAP7_75t_L g1074 ( 
.A(n_1070),
.B(n_1065),
.C(n_969),
.Y(n_1074)
);

NAND4xp25_ASAP7_75t_L g1075 ( 
.A(n_1072),
.B(n_1071),
.C(n_1067),
.D(n_1066),
.Y(n_1075)
);

NAND3xp33_ASAP7_75t_SL g1076 ( 
.A(n_1069),
.B(n_914),
.C(n_928),
.Y(n_1076)
);

NAND4xp75_ASAP7_75t_L g1077 ( 
.A(n_1068),
.B(n_960),
.C(n_927),
.D(n_835),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_1073),
.A2(n_902),
.B(n_965),
.C(n_958),
.Y(n_1078)
);

AOI221xp5_ASAP7_75t_L g1079 ( 
.A1(n_1070),
.A2(n_820),
.B1(n_893),
.B2(n_934),
.C(n_960),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1067),
.Y(n_1080)
);

AOI21xp33_ASAP7_75t_SL g1081 ( 
.A1(n_1080),
.A2(n_145),
.B(n_146),
.Y(n_1081)
);

NAND4xp25_ASAP7_75t_L g1082 ( 
.A(n_1075),
.B(n_888),
.C(n_927),
.D(n_900),
.Y(n_1082)
);

AOI211xp5_ASAP7_75t_L g1083 ( 
.A1(n_1076),
.A2(n_820),
.B(n_893),
.C(n_888),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_1078),
.B(n_893),
.Y(n_1084)
);

AND3x4_ASAP7_75t_L g1085 ( 
.A(n_1074),
.B(n_1077),
.C(n_1079),
.Y(n_1085)
);

NAND4xp25_ASAP7_75t_L g1086 ( 
.A(n_1075),
.B(n_901),
.C(n_883),
.D(n_886),
.Y(n_1086)
);

OAI321xp33_ASAP7_75t_L g1087 ( 
.A1(n_1075),
.A2(n_820),
.A3(n_893),
.B1(n_905),
.B2(n_938),
.C(n_935),
.Y(n_1087)
);

NOR3xp33_ASAP7_75t_L g1088 ( 
.A(n_1075),
.B(n_905),
.C(n_911),
.Y(n_1088)
);

NAND4xp75_ASAP7_75t_L g1089 ( 
.A(n_1080),
.B(n_835),
.C(n_938),
.D(n_151),
.Y(n_1089)
);

O2A1O1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_1080),
.A2(n_904),
.B(n_934),
.C(n_931),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1085),
.Y(n_1091)
);

NOR2xp67_ASAP7_75t_SL g1092 ( 
.A(n_1089),
.B(n_893),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_R g1093 ( 
.A(n_1081),
.B(n_148),
.Y(n_1093)
);

NOR2x1_ASAP7_75t_L g1094 ( 
.A(n_1084),
.B(n_150),
.Y(n_1094)
);

NAND2x1p5_ASAP7_75t_L g1095 ( 
.A(n_1083),
.B(n_1087),
.Y(n_1095)
);

INVxp33_ASAP7_75t_L g1096 ( 
.A(n_1086),
.Y(n_1096)
);

AND4x2_ASAP7_75t_L g1097 ( 
.A(n_1082),
.B(n_805),
.C(n_153),
.D(n_155),
.Y(n_1097)
);

NOR3xp33_ASAP7_75t_L g1098 ( 
.A(n_1088),
.B(n_911),
.C(n_912),
.Y(n_1098)
);

AOI221xp5_ASAP7_75t_L g1099 ( 
.A1(n_1090),
.A2(n_965),
.B1(n_926),
.B2(n_934),
.C(n_904),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1091),
.B(n_883),
.Y(n_1100)
);

INVxp67_ASAP7_75t_SL g1101 ( 
.A(n_1094),
.Y(n_1101)
);

NAND3xp33_ASAP7_75t_SL g1102 ( 
.A(n_1093),
.B(n_152),
.C(n_157),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1095),
.Y(n_1103)
);

NOR3xp33_ASAP7_75t_L g1104 ( 
.A(n_1096),
.B(n_158),
.C(n_159),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_1099),
.Y(n_1105)
);

NOR3xp33_ASAP7_75t_L g1106 ( 
.A(n_1098),
.B(n_160),
.C(n_161),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1097),
.Y(n_1107)
);

INVx1_ASAP7_75t_SL g1108 ( 
.A(n_1092),
.Y(n_1108)
);

NAND3xp33_ASAP7_75t_L g1109 ( 
.A(n_1091),
.B(n_886),
.C(n_901),
.Y(n_1109)
);

NAND4xp25_ASAP7_75t_L g1110 ( 
.A(n_1091),
.B(n_901),
.C(n_163),
.D(n_165),
.Y(n_1110)
);

NOR2xp67_ASAP7_75t_L g1111 ( 
.A(n_1091),
.B(n_162),
.Y(n_1111)
);

NAND4xp75_ASAP7_75t_L g1112 ( 
.A(n_1091),
.B(n_169),
.C(n_171),
.D(n_172),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1103),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1101),
.Y(n_1114)
);

NAND4xp75_ASAP7_75t_L g1115 ( 
.A(n_1111),
.B(n_174),
.C(n_175),
.D(n_176),
.Y(n_1115)
);

INVxp67_ASAP7_75t_SL g1116 ( 
.A(n_1104),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1107),
.Y(n_1117)
);

NAND4xp25_ASAP7_75t_L g1118 ( 
.A(n_1108),
.B(n_180),
.C(n_181),
.D(n_182),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_1112),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1100),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1105),
.Y(n_1121)
);

AOI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1113),
.A2(n_1102),
.B1(n_1110),
.B2(n_1106),
.Y(n_1122)
);

AOI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_1121),
.A2(n_1109),
.B1(n_947),
.B2(n_931),
.Y(n_1123)
);

INVx4_ASAP7_75t_L g1124 ( 
.A(n_1114),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_1117),
.Y(n_1125)
);

AO22x2_ASAP7_75t_L g1126 ( 
.A1(n_1120),
.A2(n_924),
.B1(n_945),
.B2(n_936),
.Y(n_1126)
);

OAI22x1_ASAP7_75t_L g1127 ( 
.A1(n_1119),
.A2(n_926),
.B1(n_925),
.B2(n_945),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1116),
.A2(n_947),
.B1(n_931),
.B2(n_926),
.Y(n_1128)
);

OAI22x1_ASAP7_75t_SL g1129 ( 
.A1(n_1124),
.A2(n_1115),
.B1(n_1118),
.B2(n_185),
.Y(n_1129)
);

INVx1_ASAP7_75t_SL g1130 ( 
.A(n_1125),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1122),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1130),
.A2(n_1123),
.B1(n_1126),
.B2(n_1128),
.Y(n_1132)
);

CKINVDCx20_ASAP7_75t_R g1133 ( 
.A(n_1132),
.Y(n_1133)
);

AOI22xp33_ASAP7_75t_L g1134 ( 
.A1(n_1133),
.A2(n_1131),
.B1(n_1127),
.B2(n_1129),
.Y(n_1134)
);

OAI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_1134),
.A2(n_880),
.B1(n_929),
.B2(n_945),
.Y(n_1135)
);

NAND4xp25_ASAP7_75t_L g1136 ( 
.A(n_1134),
.B(n_183),
.C(n_184),
.D(n_186),
.Y(n_1136)
);

AOI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1134),
.A2(n_947),
.B1(n_931),
.B2(n_948),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1136),
.A2(n_187),
.B(n_188),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_1135),
.B(n_189),
.Y(n_1139)
);

OR2x2_ASAP7_75t_L g1140 ( 
.A(n_1137),
.B(n_190),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1138),
.A2(n_191),
.B(n_192),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1139),
.B(n_193),
.Y(n_1142)
);

AO22x1_ASAP7_75t_L g1143 ( 
.A1(n_1141),
.A2(n_1140),
.B1(n_196),
.B2(n_198),
.Y(n_1143)
);

AOI211xp5_ASAP7_75t_L g1144 ( 
.A1(n_1143),
.A2(n_1142),
.B(n_199),
.C(n_200),
.Y(n_1144)
);


endmodule