module fake_jpeg_18731_n_175 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_175);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_33),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_18),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_40),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_39),
.Y(n_46)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_38),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_43),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_44),
.B(n_28),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_25),
.B1(n_21),
.B2(n_24),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_47),
.A2(n_53),
.B1(n_19),
.B2(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_18),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_49),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_18),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_18),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_25),
.B1(n_21),
.B2(n_29),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_16),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_60),
.B(n_62),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_39),
.B1(n_21),
.B2(n_31),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_61),
.A2(n_67),
.B(n_43),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_56),
.A2(n_22),
.B(n_19),
.C(n_18),
.Y(n_63)
);

NOR2x1_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_26),
.Y(n_87)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_70),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_0),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_15),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_69),
.B(n_76),
.Y(n_97)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_41),
.A2(n_26),
.B1(n_20),
.B2(n_27),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_72),
.A2(n_75),
.B1(n_46),
.B2(n_54),
.Y(n_85)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_26),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_67),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_49),
.A2(n_41),
.B1(n_46),
.B2(n_42),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_15),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_46),
.A2(n_27),
.B1(n_15),
.B2(n_20),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_77),
.A2(n_52),
.B1(n_50),
.B2(n_27),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_80),
.A2(n_86),
.B(n_96),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_43),
.C(n_50),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_61),
.C(n_71),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g82 ( 
.A(n_60),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_82),
.B(n_95),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_88),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_85),
.A2(n_90),
.B1(n_91),
.B2(n_73),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_87),
.B(n_3),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_50),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_68),
.A2(n_52),
.B1(n_1),
.B2(n_2),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_65),
.A2(n_74),
.B1(n_64),
.B2(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_2),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_57),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_103),
.Y(n_127)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_101),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_81),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_84),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_89),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_57),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_113),
.Y(n_130)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_110),
.C(n_90),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_61),
.C(n_63),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_94),
.A2(n_70),
.B1(n_66),
.B2(n_4),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_112),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_91),
.B(n_2),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_14),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_114),
.B(n_82),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_108),
.A2(n_80),
.B(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_117),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_108),
.A2(n_96),
.B(n_87),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_86),
.B(n_95),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_116),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_109),
.A2(n_95),
.B(n_96),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_122),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_105),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_121),
.B(n_123),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_100),
.A2(n_85),
.B1(n_84),
.B2(n_79),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_124),
.A2(n_110),
.B1(n_106),
.B2(n_101),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_102),
.C(n_112),
.Y(n_133)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_128),
.B(n_3),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_131),
.A2(n_140),
.B1(n_136),
.B2(n_137),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_136),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_107),
.C(n_103),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_141),
.C(n_120),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_124),
.Y(n_143)
);

OA21x2_ASAP7_75t_SL g138 ( 
.A1(n_123),
.A2(n_114),
.B(n_109),
.Y(n_138)
);

OA21x2_ASAP7_75t_SL g150 ( 
.A1(n_138),
.A2(n_117),
.B(n_129),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_126),
.A2(n_118),
.B1(n_119),
.B2(n_127),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_107),
.C(n_14),
.Y(n_141)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_143),
.A2(n_151),
.B(n_134),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_145),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_131),
.A2(n_129),
.B1(n_121),
.B2(n_127),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_147),
.C(n_150),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_130),
.Y(n_148)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_148),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_115),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_145),
.A2(n_132),
.B(n_115),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_152),
.A2(n_156),
.B(n_3),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_157),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_151),
.A2(n_128),
.B(n_141),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_133),
.B1(n_13),
.B2(n_12),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_147),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_161),
.Y(n_165)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_153),
.A2(n_146),
.B1(n_13),
.B2(n_6),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_163),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_158),
.A2(n_5),
.B(n_7),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_SL g168 ( 
.A1(n_164),
.A2(n_5),
.B(n_8),
.C(n_9),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_160),
.A2(n_159),
.B1(n_7),
.B2(n_8),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_166),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_168),
.Y(n_171)
);

NAND3xp33_ASAP7_75t_SL g170 ( 
.A(n_165),
.B(n_9),
.C(n_10),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_170),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_169),
.A2(n_167),
.B(n_168),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_172),
.A2(n_171),
.B(n_9),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_173),
.Y(n_175)
);


endmodule