module fake_aes_12752_n_882 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_237, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_242, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_882, n_880);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_237;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_242;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_882;
output n_880;
wire n_663;
wire n_707;
wire n_791;
wire n_513;
wire n_361;
wire n_838;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_878;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_564;
wire n_353;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_316;
wire n_545;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_789;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_384;
wire n_476;
wire n_617;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_567;
wire n_809;
wire n_580;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_490;
wire n_393;
wire n_247;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_415;
wire n_482;
wire n_394;
wire n_703;
wire n_442;
wire n_331;
wire n_485;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_729;
wire n_519;
wire n_338;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_876;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_621;
wire n_423;
wire n_342;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_716;
wire n_653;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_522;
wire n_264;
wire n_573;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_409;
wire n_363;
wire n_315;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_639;
wire n_376;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_498;
wire n_597;
wire n_349;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_837;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_581;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_515;
wire n_253;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_606;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_781;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_SL g244 ( .A(n_14), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_78), .Y(n_245) );
INVxp67_ASAP7_75t_L g246 ( .A(n_161), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_143), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_200), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_132), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_19), .Y(n_250) );
INVx2_ASAP7_75t_SL g251 ( .A(n_73), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_167), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_52), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_153), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_133), .Y(n_255) );
INVx1_ASAP7_75t_SL g256 ( .A(n_18), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_51), .Y(n_257) );
INVx2_ASAP7_75t_SL g258 ( .A(n_112), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_36), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_61), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_194), .Y(n_261) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_197), .Y(n_262) );
INVx1_ASAP7_75t_SL g263 ( .A(n_135), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_80), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g265 ( .A(n_184), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_115), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_84), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_100), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_168), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_214), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_139), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_19), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_242), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_65), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_221), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_38), .Y(n_276) );
BUFx3_ASAP7_75t_L g277 ( .A(n_95), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_92), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_190), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_91), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_32), .Y(n_281) );
CKINVDCx16_ASAP7_75t_R g282 ( .A(n_9), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_37), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_146), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_31), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_142), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_136), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_130), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_72), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_224), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_229), .Y(n_291) );
BUFx6f_ASAP7_75t_L g292 ( .A(n_71), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_56), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_99), .Y(n_294) );
INVxp67_ASAP7_75t_SL g295 ( .A(n_82), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_113), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_131), .Y(n_297) );
BUFx10_ASAP7_75t_L g298 ( .A(n_77), .Y(n_298) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_109), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_171), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_147), .Y(n_301) );
CKINVDCx20_ASAP7_75t_R g302 ( .A(n_110), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_30), .Y(n_303) );
INVxp67_ASAP7_75t_L g304 ( .A(n_185), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_182), .Y(n_305) );
CKINVDCx16_ASAP7_75t_R g306 ( .A(n_191), .Y(n_306) );
CKINVDCx16_ASAP7_75t_R g307 ( .A(n_63), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_204), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_7), .Y(n_309) );
BUFx10_ASAP7_75t_L g310 ( .A(n_85), .Y(n_310) );
INVxp67_ASAP7_75t_SL g311 ( .A(n_187), .Y(n_311) );
CKINVDCx16_ASAP7_75t_R g312 ( .A(n_216), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_96), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_18), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_231), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_230), .Y(n_316) );
BUFx8_ASAP7_75t_SL g317 ( .A(n_241), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_186), .Y(n_318) );
CKINVDCx20_ASAP7_75t_R g319 ( .A(n_86), .Y(n_319) );
CKINVDCx20_ASAP7_75t_R g320 ( .A(n_105), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_13), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_23), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_54), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_43), .Y(n_324) );
CKINVDCx16_ASAP7_75t_R g325 ( .A(n_53), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_88), .Y(n_326) );
INVx1_ASAP7_75t_SL g327 ( .A(n_90), .Y(n_327) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_164), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_106), .Y(n_329) );
INVx2_ASAP7_75t_SL g330 ( .A(n_127), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_151), .Y(n_331) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_7), .Y(n_332) );
CKINVDCx20_ASAP7_75t_R g333 ( .A(n_10), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_215), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_119), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_87), .Y(n_336) );
INVx1_ASAP7_75t_SL g337 ( .A(n_202), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_128), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_30), .Y(n_339) );
BUFx5_ASAP7_75t_L g340 ( .A(n_20), .Y(n_340) );
CKINVDCx5p33_ASAP7_75t_R g341 ( .A(n_219), .Y(n_341) );
INVx1_ASAP7_75t_SL g342 ( .A(n_26), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_222), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_159), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_210), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_180), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_25), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_162), .Y(n_348) );
INVx1_ASAP7_75t_SL g349 ( .A(n_163), .Y(n_349) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_145), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_193), .Y(n_351) );
BUFx10_ASAP7_75t_L g352 ( .A(n_83), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_172), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_43), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_46), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_239), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_176), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_188), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_81), .Y(n_359) );
INVx1_ASAP7_75t_SL g360 ( .A(n_68), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_123), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_67), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_24), .Y(n_363) );
BUFx8_ASAP7_75t_SL g364 ( .A(n_89), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_5), .Y(n_365) );
CKINVDCx5p33_ASAP7_75t_R g366 ( .A(n_98), .Y(n_366) );
INVx3_ASAP7_75t_L g367 ( .A(n_137), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_64), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_57), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_120), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_235), .Y(n_371) );
CKINVDCx20_ASAP7_75t_R g372 ( .A(n_218), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_58), .Y(n_373) );
BUFx3_ASAP7_75t_L g374 ( .A(n_32), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_74), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_62), .Y(n_376) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_292), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_367), .B(n_0), .Y(n_378) );
INVx5_ASAP7_75t_L g379 ( .A(n_367), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_282), .B(n_0), .Y(n_380) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_292), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_340), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_321), .Y(n_383) );
INVx3_ASAP7_75t_L g384 ( .A(n_298), .Y(n_384) );
BUFx3_ASAP7_75t_L g385 ( .A(n_277), .Y(n_385) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_292), .Y(n_386) );
AND2x4_ASAP7_75t_L g387 ( .A(n_321), .B(n_1), .Y(n_387) );
AND2x4_ASAP7_75t_L g388 ( .A(n_374), .B(n_1), .Y(n_388) );
INVx5_ASAP7_75t_L g389 ( .A(n_292), .Y(n_389) );
INVx3_ASAP7_75t_L g390 ( .A(n_298), .Y(n_390) );
AND2x6_ASAP7_75t_L g391 ( .A(n_277), .B(n_55), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_306), .B(n_2), .Y(n_392) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_299), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_251), .B(n_2), .Y(n_394) );
INVx3_ASAP7_75t_L g395 ( .A(n_298), .Y(n_395) );
BUFx8_ASAP7_75t_SL g396 ( .A(n_332), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_299), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_340), .Y(n_398) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_299), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_299), .Y(n_400) );
BUFx8_ASAP7_75t_L g401 ( .A(n_340), .Y(n_401) );
INVx5_ASAP7_75t_L g402 ( .A(n_258), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_330), .B(n_3), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_328), .B(n_3), .Y(n_404) );
BUFx8_ASAP7_75t_SL g405 ( .A(n_333), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_383), .B(n_307), .Y(n_406) );
OA22x2_ASAP7_75t_L g407 ( .A1(n_383), .A2(n_285), .B1(n_355), .B2(n_259), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_384), .A2(n_302), .B1(n_372), .B2(n_305), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_387), .A2(n_325), .B1(n_312), .B2(n_305), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_387), .A2(n_372), .B1(n_302), .B2(n_250), .Y(n_410) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_401), .Y(n_411) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_387), .A2(n_272), .B1(n_276), .B2(n_257), .Y(n_412) );
AND2x4_ASAP7_75t_L g413 ( .A(n_384), .B(n_390), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_382), .Y(n_414) );
AO22x2_ASAP7_75t_L g415 ( .A1(n_387), .A2(n_374), .B1(n_256), .B2(n_342), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_384), .B(n_350), .Y(n_416) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_377), .Y(n_417) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_388), .A2(n_283), .B1(n_303), .B2(n_281), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_384), .B(n_310), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_382), .Y(n_420) );
OAI22xp33_ASAP7_75t_L g421 ( .A1(n_380), .A2(n_244), .B1(n_314), .B2(n_309), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_390), .B(n_310), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_390), .B(n_310), .Y(n_423) );
OAI22xp5_ASAP7_75t_SL g424 ( .A1(n_396), .A2(n_319), .B1(n_320), .B2(n_265), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_388), .Y(n_425) );
OAI22xp33_ASAP7_75t_R g426 ( .A1(n_405), .A2(n_247), .B1(n_248), .B2(n_245), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_390), .B(n_352), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_398), .Y(n_428) );
OAI22xp5_ASAP7_75t_SL g429 ( .A1(n_404), .A2(n_324), .B1(n_339), .B2(n_322), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_423), .B(n_395), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_414), .Y(n_431) );
AOI21x1_ASAP7_75t_L g432 ( .A1(n_414), .A2(n_398), .B(n_394), .Y(n_432) );
AND2x4_ASAP7_75t_L g433 ( .A(n_423), .B(n_419), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_413), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_416), .B(n_395), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_420), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_425), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_413), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_413), .Y(n_439) );
INVxp67_ASAP7_75t_L g440 ( .A(n_408), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_411), .B(n_395), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_422), .B(n_395), .Y(n_442) );
AND2x4_ASAP7_75t_L g443 ( .A(n_427), .B(n_388), .Y(n_443) );
XOR2x2_ASAP7_75t_L g444 ( .A(n_410), .B(n_380), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_407), .Y(n_445) );
CKINVDCx5p33_ASAP7_75t_R g446 ( .A(n_424), .Y(n_446) );
XOR2xp5_ASAP7_75t_L g447 ( .A(n_409), .B(n_392), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_406), .B(n_401), .Y(n_448) );
BUFx6f_ASAP7_75t_SL g449 ( .A(n_426), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_420), .Y(n_450) );
AND2x4_ASAP7_75t_L g451 ( .A(n_411), .B(n_388), .Y(n_451) );
XNOR2x2_ASAP7_75t_L g452 ( .A(n_415), .B(n_378), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_428), .Y(n_453) );
INVx3_ASAP7_75t_L g454 ( .A(n_428), .Y(n_454) );
XOR2xp5_ASAP7_75t_L g455 ( .A(n_415), .B(n_392), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_407), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_415), .Y(n_457) );
AND2x4_ASAP7_75t_L g458 ( .A(n_433), .B(n_406), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_457), .A2(n_401), .B1(n_429), .B2(n_418), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_431), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_433), .B(n_412), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_433), .B(n_421), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_453), .Y(n_463) );
BUFx3_ASAP7_75t_L g464 ( .A(n_453), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_456), .B(n_379), .Y(n_465) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_432), .Y(n_466) );
INVx4_ASAP7_75t_L g467 ( .A(n_451), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_431), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_451), .B(n_379), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_451), .B(n_379), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_445), .B(n_379), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_443), .B(n_379), .Y(n_472) );
INVx1_ASAP7_75t_SL g473 ( .A(n_436), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_443), .B(n_379), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_437), .B(n_421), .Y(n_475) );
INVx3_ASAP7_75t_L g476 ( .A(n_454), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_435), .B(n_379), .Y(n_477) );
INVxp33_ASAP7_75t_L g478 ( .A(n_455), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_443), .B(n_385), .Y(n_479) );
OAI21xp5_ASAP7_75t_L g480 ( .A1(n_432), .A2(n_403), .B(n_394), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_448), .B(n_403), .Y(n_481) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_454), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_440), .B(n_385), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_447), .B(n_347), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_436), .Y(n_485) );
INVx2_ASAP7_75t_SL g486 ( .A(n_454), .Y(n_486) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_450), .Y(n_487) );
AND2x4_ASAP7_75t_L g488 ( .A(n_434), .B(n_295), .Y(n_488) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_458), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_458), .B(n_455), .Y(n_490) );
OR2x6_ASAP7_75t_L g491 ( .A(n_467), .B(n_438), .Y(n_491) );
OR2x6_ASAP7_75t_L g492 ( .A(n_467), .B(n_439), .Y(n_492) );
NOR2x1_ASAP7_75t_L g493 ( .A(n_464), .B(n_437), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_462), .B(n_430), .Y(n_494) );
NOR2xp33_ASAP7_75t_SL g495 ( .A(n_467), .B(n_446), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_462), .B(n_442), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_458), .B(n_444), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_461), .B(n_447), .Y(n_498) );
INVxp67_ASAP7_75t_SL g499 ( .A(n_464), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_458), .B(n_444), .Y(n_500) );
INVx3_ASAP7_75t_L g501 ( .A(n_464), .Y(n_501) );
INVx8_ASAP7_75t_L g502 ( .A(n_479), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_463), .B(n_450), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_460), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_463), .Y(n_505) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_466), .Y(n_506) );
INVx5_ASAP7_75t_L g507 ( .A(n_467), .Y(n_507) );
OR2x6_ASAP7_75t_L g508 ( .A(n_461), .B(n_441), .Y(n_508) );
BUFx3_ASAP7_75t_L g509 ( .A(n_460), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_481), .B(n_401), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_478), .B(n_446), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_460), .Y(n_512) );
INVx3_ASAP7_75t_L g513 ( .A(n_482), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_468), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_480), .B(n_385), .Y(n_515) );
AND2x6_ASAP7_75t_L g516 ( .A(n_473), .B(n_452), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_484), .B(n_449), .Y(n_517) );
AND2x2_ASAP7_75t_SL g518 ( .A(n_466), .B(n_452), .Y(n_518) );
INVx2_ASAP7_75t_SL g519 ( .A(n_469), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_468), .Y(n_520) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_466), .Y(n_521) );
INVx6_ASAP7_75t_SL g522 ( .A(n_488), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_468), .Y(n_523) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_466), .Y(n_524) );
NAND2x1p5_ASAP7_75t_L g525 ( .A(n_507), .B(n_473), .Y(n_525) );
BUFx2_ASAP7_75t_SL g526 ( .A(n_507), .Y(n_526) );
BUFx4_ASAP7_75t_SL g527 ( .A(n_491), .Y(n_527) );
BUFx12f_ASAP7_75t_L g528 ( .A(n_507), .Y(n_528) );
INVx3_ASAP7_75t_L g529 ( .A(n_501), .Y(n_529) );
INVx3_ASAP7_75t_L g530 ( .A(n_501), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_505), .Y(n_531) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_506), .Y(n_532) );
INVx5_ASAP7_75t_L g533 ( .A(n_507), .Y(n_533) );
BUFx4_ASAP7_75t_SL g534 ( .A(n_491), .Y(n_534) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_506), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_505), .Y(n_536) );
BUFx24_ASAP7_75t_L g537 ( .A(n_522), .Y(n_537) );
INVx2_ASAP7_75t_SL g538 ( .A(n_507), .Y(n_538) );
INVx5_ASAP7_75t_L g539 ( .A(n_507), .Y(n_539) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_506), .Y(n_540) );
BUFx2_ASAP7_75t_L g541 ( .A(n_499), .Y(n_541) );
BUFx3_ASAP7_75t_L g542 ( .A(n_509), .Y(n_542) );
INVx3_ASAP7_75t_SL g543 ( .A(n_502), .Y(n_543) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_522), .Y(n_544) );
INVx4_ASAP7_75t_L g545 ( .A(n_501), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_504), .Y(n_546) );
BUFx12f_ASAP7_75t_L g547 ( .A(n_497), .Y(n_547) );
INVx3_ASAP7_75t_SL g548 ( .A(n_502), .Y(n_548) );
BUFx3_ASAP7_75t_L g549 ( .A(n_509), .Y(n_549) );
BUFx5_ASAP7_75t_L g550 ( .A(n_523), .Y(n_550) );
INVx3_ASAP7_75t_SL g551 ( .A(n_502), .Y(n_551) );
BUFx8_ASAP7_75t_SL g552 ( .A(n_491), .Y(n_552) );
BUFx2_ASAP7_75t_SL g553 ( .A(n_504), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_500), .A2(n_449), .B1(n_459), .B2(n_483), .Y(n_554) );
NAND2x1p5_ASAP7_75t_L g555 ( .A(n_493), .B(n_523), .Y(n_555) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_512), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_498), .B(n_459), .Y(n_557) );
BUFx3_ASAP7_75t_L g558 ( .A(n_512), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_514), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_500), .A2(n_449), .B1(n_483), .B2(n_475), .Y(n_560) );
INVxp67_ASAP7_75t_SL g561 ( .A(n_514), .Y(n_561) );
INVx1_ASAP7_75t_SL g562 ( .A(n_522), .Y(n_562) );
INVx3_ASAP7_75t_L g563 ( .A(n_491), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_497), .B(n_475), .Y(n_564) );
INVx2_ASAP7_75t_SL g565 ( .A(n_502), .Y(n_565) );
BUFx2_ASAP7_75t_SL g566 ( .A(n_520), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_503), .Y(n_567) );
BUFx3_ASAP7_75t_L g568 ( .A(n_492), .Y(n_568) );
INVx3_ASAP7_75t_L g569 ( .A(n_492), .Y(n_569) );
BUFx12f_ASAP7_75t_L g570 ( .A(n_492), .Y(n_570) );
INVx1_ASAP7_75t_SL g571 ( .A(n_492), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_490), .B(n_485), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_489), .Y(n_573) );
NAND2x1p5_ASAP7_75t_L g574 ( .A(n_493), .B(n_482), .Y(n_574) );
OAI22xp33_ASAP7_75t_L g575 ( .A1(n_543), .A2(n_495), .B1(n_508), .B2(n_510), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_546), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_531), .Y(n_577) );
BUFx12f_ASAP7_75t_L g578 ( .A(n_528), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_554), .A2(n_508), .B1(n_518), .B2(n_516), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_546), .Y(n_580) );
BUFx2_ASAP7_75t_L g581 ( .A(n_528), .Y(n_581) );
OAI22xp33_ASAP7_75t_L g582 ( .A1(n_543), .A2(n_508), .B1(n_496), .B2(n_494), .Y(n_582) );
AOI21xp33_ASAP7_75t_L g583 ( .A1(n_557), .A2(n_515), .B(n_541), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_559), .Y(n_584) );
BUFx5_ASAP7_75t_L g585 ( .A(n_558), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_536), .Y(n_586) );
CKINVDCx20_ASAP7_75t_R g587 ( .A(n_552), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_553), .A2(n_518), .B1(n_515), .B2(n_466), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_566), .A2(n_466), .B1(n_480), .B2(n_485), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_547), .A2(n_516), .B1(n_519), .B2(n_517), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_564), .A2(n_511), .B1(n_519), .B2(n_483), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_572), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_560), .A2(n_516), .B1(n_479), .B2(n_488), .Y(n_593) );
INVx6_ASAP7_75t_L g594 ( .A(n_533), .Y(n_594) );
OAI22xp33_ASAP7_75t_L g595 ( .A1(n_548), .A2(n_466), .B1(n_486), .B2(n_487), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_556), .Y(n_596) );
INVx4_ASAP7_75t_L g597 ( .A(n_533), .Y(n_597) );
CKINVDCx11_ASAP7_75t_R g598 ( .A(n_548), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_550), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_570), .A2(n_524), .B1(n_506), .B2(n_521), .Y(n_600) );
CKINVDCx20_ASAP7_75t_R g601 ( .A(n_551), .Y(n_601) );
BUFx6f_ASAP7_75t_L g602 ( .A(n_533), .Y(n_602) );
INVxp67_ASAP7_75t_L g603 ( .A(n_526), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_570), .A2(n_524), .B1(n_506), .B2(n_521), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_550), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_567), .Y(n_606) );
INVx3_ASAP7_75t_L g607 ( .A(n_533), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_563), .A2(n_471), .B1(n_477), .B2(n_474), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_550), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_563), .A2(n_472), .B1(n_474), .B2(n_476), .Y(n_610) );
BUFx2_ASAP7_75t_L g611 ( .A(n_539), .Y(n_611) );
CKINVDCx11_ASAP7_75t_R g612 ( .A(n_551), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_565), .B(n_354), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_573), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_550), .Y(n_615) );
AOI22xp33_ASAP7_75t_SL g616 ( .A1(n_568), .A2(n_524), .B1(n_521), .B2(n_513), .Y(n_616) );
AOI22xp33_ASAP7_75t_SL g617 ( .A1(n_568), .A2(n_524), .B1(n_521), .B2(n_513), .Y(n_617) );
INVx3_ASAP7_75t_L g618 ( .A(n_539), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_550), .B(n_513), .Y(n_619) );
INVx3_ASAP7_75t_L g620 ( .A(n_539), .Y(n_620) );
AOI22xp33_ASAP7_75t_SL g621 ( .A1(n_569), .A2(n_521), .B1(n_524), .B2(n_352), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_550), .Y(n_622) );
INVx1_ASAP7_75t_SL g623 ( .A(n_541), .Y(n_623) );
BUFx3_ASAP7_75t_L g624 ( .A(n_539), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_544), .Y(n_625) );
BUFx12f_ASAP7_75t_L g626 ( .A(n_544), .Y(n_626) );
CKINVDCx11_ASAP7_75t_R g627 ( .A(n_562), .Y(n_627) );
BUFx4_ASAP7_75t_SL g628 ( .A(n_542), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_550), .Y(n_629) );
CKINVDCx5p33_ASAP7_75t_R g630 ( .A(n_527), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_569), .A2(n_472), .B1(n_474), .B2(n_476), .Y(n_631) );
INVx2_ASAP7_75t_SL g632 ( .A(n_534), .Y(n_632) );
CKINVDCx6p67_ASAP7_75t_R g633 ( .A(n_537), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_525), .A2(n_487), .B1(n_486), .B2(n_476), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_558), .B(n_465), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_569), .A2(n_472), .B1(n_476), .B2(n_352), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_565), .B(n_363), .Y(n_637) );
AOI22xp33_ASAP7_75t_SL g638 ( .A1(n_538), .A2(n_487), .B1(n_365), .B2(n_470), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_571), .A2(n_486), .B1(n_469), .B2(n_470), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_525), .A2(n_487), .B1(n_482), .B2(n_311), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_525), .A2(n_487), .B1(n_482), .B2(n_246), .Y(n_641) );
CKINVDCx11_ASAP7_75t_R g642 ( .A(n_542), .Y(n_642) );
BUFx6f_ASAP7_75t_L g643 ( .A(n_549), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_561), .B(n_487), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_529), .B(n_487), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_555), .Y(n_646) );
BUFx6f_ASAP7_75t_L g647 ( .A(n_549), .Y(n_647) );
CKINVDCx20_ASAP7_75t_R g648 ( .A(n_545), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_545), .A2(n_482), .B1(n_340), .B2(n_391), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_555), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_574), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_576), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_648), .A2(n_545), .B1(n_574), .B2(n_530), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_593), .A2(n_530), .B1(n_529), .B2(n_340), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_591), .A2(n_530), .B1(n_529), .B2(n_340), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_583), .A2(n_340), .B1(n_364), .B2(n_317), .Y(n_656) );
OAI222xp33_ASAP7_75t_L g657 ( .A1(n_623), .A2(n_574), .B1(n_253), .B2(n_255), .C1(n_373), .C2(n_318), .Y(n_657) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_623), .Y(n_658) );
INVx1_ASAP7_75t_SL g659 ( .A(n_598), .Y(n_659) );
CKINVDCx11_ASAP7_75t_R g660 ( .A(n_612), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_580), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_583), .A2(n_266), .B1(n_268), .B2(n_260), .Y(n_662) );
AOI22xp33_ASAP7_75t_SL g663 ( .A1(n_581), .A2(n_535), .B1(n_540), .B2(n_532), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_582), .A2(n_592), .B1(n_632), .B2(n_575), .Y(n_664) );
INVx4_ASAP7_75t_L g665 ( .A(n_633), .Y(n_665) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_615), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_579), .A2(n_269), .B1(n_289), .B2(n_287), .Y(n_667) );
CKINVDCx6p67_ASAP7_75t_R g668 ( .A(n_578), .Y(n_668) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_622), .Y(n_669) );
AOI22xp33_ASAP7_75t_SL g670 ( .A1(n_611), .A2(n_535), .B1(n_540), .B2(n_532), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_601), .B(n_304), .Y(n_671) );
BUFx6f_ASAP7_75t_L g672 ( .A(n_602), .Y(n_672) );
BUFx8_ASAP7_75t_SL g673 ( .A(n_587), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_590), .A2(n_326), .B1(n_336), .B2(n_290), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_596), .B(n_4), .Y(n_675) );
INVxp67_ASAP7_75t_L g676 ( .A(n_613), .Y(n_676) );
AOI22xp33_ASAP7_75t_SL g677 ( .A1(n_594), .A2(n_348), .B1(n_356), .B2(n_344), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_639), .A2(n_362), .B1(n_369), .B2(n_361), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_642), .B(n_4), .Y(n_679) );
AOI222xp33_ASAP7_75t_L g680 ( .A1(n_614), .A2(n_370), .B1(n_371), .B2(n_270), .C1(n_279), .C2(n_286), .Y(n_680) );
INVx2_ASAP7_75t_L g681 ( .A(n_584), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_608), .A2(n_270), .B1(n_286), .B2(n_279), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_638), .A2(n_300), .B1(n_371), .B2(n_327), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_606), .A2(n_397), .B1(n_400), .B2(n_391), .Y(n_684) );
INVx3_ASAP7_75t_L g685 ( .A(n_597), .Y(n_685) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_629), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_627), .A2(n_391), .B1(n_337), .B2(n_349), .Y(n_687) );
OAI21xp33_ASAP7_75t_L g688 ( .A1(n_637), .A2(n_400), .B(n_397), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_610), .A2(n_391), .B1(n_360), .B2(n_263), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_577), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_586), .B(n_5), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_631), .A2(n_391), .B1(n_402), .B2(n_381), .Y(n_692) );
AND2x2_ASAP7_75t_L g693 ( .A(n_603), .B(n_6), .Y(n_693) );
OAI21xp5_ASAP7_75t_L g694 ( .A1(n_641), .A2(n_391), .B(n_402), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_588), .A2(n_391), .B1(n_402), .B2(n_381), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_588), .A2(n_391), .B1(n_381), .B2(n_386), .Y(n_696) );
BUFx3_ASAP7_75t_L g697 ( .A(n_630), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_641), .A2(n_252), .B1(n_254), .B2(n_249), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_644), .Y(n_699) );
INVx5_ASAP7_75t_SL g700 ( .A(n_602), .Y(n_700) );
INVx4_ASAP7_75t_L g701 ( .A(n_602), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_635), .A2(n_381), .B1(n_386), .B2(n_377), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_628), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_625), .B(n_8), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_635), .A2(n_381), .B1(n_386), .B2(n_377), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_636), .A2(n_262), .B1(n_264), .B2(n_261), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_607), .A2(n_271), .B1(n_273), .B2(n_267), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_644), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_607), .B(n_8), .Y(n_709) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_626), .Y(n_710) );
BUFx12f_ASAP7_75t_L g711 ( .A(n_643), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_618), .Y(n_712) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_589), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_624), .A2(n_386), .B1(n_393), .B2(n_377), .Y(n_714) );
AOI21xp33_ASAP7_75t_L g715 ( .A1(n_646), .A2(n_402), .B(n_386), .Y(n_715) );
AOI222xp33_ASAP7_75t_L g716 ( .A1(n_620), .A2(n_650), .B1(n_640), .B2(n_589), .C1(n_600), .C2(n_604), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_620), .B(n_10), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_651), .Y(n_718) );
AOI22xp33_ASAP7_75t_SL g719 ( .A1(n_600), .A2(n_275), .B1(n_278), .B2(n_274), .Y(n_719) );
CKINVDCx5p33_ASAP7_75t_R g720 ( .A(n_643), .Y(n_720) );
AOI22xp33_ASAP7_75t_SL g721 ( .A1(n_604), .A2(n_284), .B1(n_288), .B2(n_280), .Y(n_721) );
AOI22xp33_ASAP7_75t_SL g722 ( .A1(n_640), .A2(n_293), .B1(n_294), .B2(n_291), .Y(n_722) );
OAI22xp33_ASAP7_75t_SL g723 ( .A1(n_599), .A2(n_297), .B1(n_301), .B2(n_296), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_647), .B(n_11), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_647), .A2(n_402), .B1(n_393), .B2(n_399), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_647), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_605), .A2(n_402), .B1(n_393), .B2(n_399), .Y(n_727) );
INVx3_ASAP7_75t_L g728 ( .A(n_609), .Y(n_728) );
OAI21xp5_ASAP7_75t_SL g729 ( .A1(n_621), .A2(n_11), .B(n_12), .Y(n_729) );
AOI22xp33_ASAP7_75t_SL g730 ( .A1(n_634), .A2(n_313), .B1(n_315), .B2(n_308), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_619), .A2(n_316), .B1(n_323), .B2(n_329), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_645), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_690), .B(n_585), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_664), .A2(n_585), .B1(n_645), .B2(n_617), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_664), .A2(n_585), .B1(n_616), .B2(n_595), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_656), .A2(n_649), .B1(n_358), .B2(n_357), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_652), .Y(n_737) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_656), .A2(n_331), .B1(n_334), .B2(n_335), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_676), .A2(n_377), .B1(n_399), .B2(n_393), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_667), .A2(n_393), .B1(n_399), .B2(n_359), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_729), .A2(n_338), .B1(n_341), .B2(n_343), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_682), .A2(n_345), .B1(n_346), .B2(n_351), .Y(n_742) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_682), .A2(n_353), .B1(n_366), .B2(n_368), .Y(n_743) );
INVx2_ASAP7_75t_L g744 ( .A(n_661), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_716), .A2(n_399), .B1(n_376), .B2(n_375), .Y(n_745) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_665), .A2(n_389), .B1(n_13), .B2(n_14), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_654), .A2(n_389), .B1(n_417), .B2(n_16), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_665), .A2(n_389), .B1(n_15), .B2(n_16), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_654), .A2(n_389), .B1(n_417), .B2(n_17), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_655), .A2(n_389), .B1(n_417), .B2(n_17), .Y(n_750) );
AOI222xp33_ASAP7_75t_L g751 ( .A1(n_679), .A2(n_12), .B1(n_15), .B2(n_20), .C1(n_21), .C2(n_22), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_658), .Y(n_752) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_671), .B(n_21), .Y(n_753) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_662), .A2(n_389), .B1(n_26), .B2(n_27), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_662), .A2(n_25), .B1(n_27), .B2(n_28), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_724), .A2(n_28), .B1(n_29), .B2(n_31), .Y(n_756) );
AOI22xp33_ASAP7_75t_SL g757 ( .A1(n_685), .A2(n_29), .B1(n_33), .B2(n_34), .Y(n_757) );
OAI222xp33_ASAP7_75t_L g758 ( .A1(n_653), .A2(n_33), .B1(n_34), .B2(n_35), .C1(n_36), .C2(n_37), .Y(n_758) );
AOI222xp33_ASAP7_75t_L g759 ( .A1(n_704), .A2(n_35), .B1(n_38), .B2(n_39), .C1(n_40), .C2(n_41), .Y(n_759) );
OAI21xp5_ASAP7_75t_L g760 ( .A1(n_657), .A2(n_39), .B(n_40), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_674), .A2(n_42), .B1(n_44), .B2(n_45), .Y(n_761) );
AOI22xp33_ASAP7_75t_SL g762 ( .A1(n_685), .A2(n_45), .B1(n_46), .B2(n_47), .Y(n_762) );
NAND3xp33_ASAP7_75t_L g763 ( .A(n_680), .B(n_677), .C(n_693), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_703), .A2(n_48), .B1(n_49), .B2(n_50), .Y(n_764) );
AOI22xp5_ASAP7_75t_L g765 ( .A1(n_683), .A2(n_59), .B1(n_60), .B2(n_66), .Y(n_765) );
AND2x2_ASAP7_75t_L g766 ( .A(n_658), .B(n_69), .Y(n_766) );
AND2x2_ASAP7_75t_L g767 ( .A(n_720), .B(n_70), .Y(n_767) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_719), .A2(n_75), .B1(n_76), .B2(n_79), .Y(n_768) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_721), .A2(n_93), .B1(n_94), .B2(n_97), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_678), .A2(n_732), .B1(n_675), .B2(n_688), .Y(n_770) );
AOI22xp33_ASAP7_75t_SL g771 ( .A1(n_726), .A2(n_101), .B1(n_102), .B2(n_103), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_691), .B(n_699), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_708), .A2(n_709), .B1(n_717), .B2(n_660), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_713), .A2(n_104), .B1(n_107), .B2(n_108), .Y(n_774) );
OAI222xp33_ASAP7_75t_L g775 ( .A1(n_659), .A2(n_111), .B1(n_114), .B2(n_116), .C1(n_117), .C2(n_118), .Y(n_775) );
AOI22xp33_ASAP7_75t_SL g776 ( .A1(n_701), .A2(n_121), .B1(n_122), .B2(n_124), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_712), .A2(n_125), .B1(n_126), .B2(n_129), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_713), .A2(n_134), .B1(n_138), .B2(n_140), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_666), .A2(n_141), .B1(n_144), .B2(n_148), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_666), .A2(n_149), .B1(n_150), .B2(n_152), .Y(n_780) );
AOI22xp5_ASAP7_75t_L g781 ( .A1(n_698), .A2(n_154), .B1(n_155), .B2(n_156), .Y(n_781) );
OAI21xp5_ASAP7_75t_SL g782 ( .A1(n_663), .A2(n_722), .B(n_730), .Y(n_782) );
OAI222xp33_ASAP7_75t_L g783 ( .A1(n_701), .A2(n_157), .B1(n_158), .B2(n_160), .C1(n_165), .C2(n_166), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_669), .A2(n_169), .B1(n_170), .B2(n_173), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_669), .A2(n_174), .B1(n_175), .B2(n_177), .Y(n_785) );
AO22x1_ASAP7_75t_L g786 ( .A1(n_697), .A2(n_178), .B1(n_179), .B2(n_181), .Y(n_786) );
NOR2xp67_ASAP7_75t_L g787 ( .A(n_711), .B(n_183), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g788 ( .A1(n_731), .A2(n_189), .B1(n_192), .B2(n_195), .Y(n_788) );
OA21x2_ASAP7_75t_L g789 ( .A1(n_696), .A2(n_196), .B(n_198), .Y(n_789) );
NOR3xp33_ASAP7_75t_SL g790 ( .A(n_782), .B(n_668), .C(n_673), .Y(n_790) );
NAND2xp5_ASAP7_75t_SL g791 ( .A(n_734), .B(n_670), .Y(n_791) );
OAI21xp33_ASAP7_75t_L g792 ( .A1(n_745), .A2(n_705), .B(n_702), .Y(n_792) );
AOI221xp5_ASAP7_75t_L g793 ( .A1(n_753), .A2(n_723), .B1(n_686), .B2(n_718), .C(n_702), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_772), .B(n_686), .Y(n_794) );
AND2x2_ASAP7_75t_L g795 ( .A(n_752), .B(n_737), .Y(n_795) );
OAI221xp5_ASAP7_75t_SL g796 ( .A1(n_773), .A2(n_705), .B1(n_696), .B2(n_687), .C(n_714), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_744), .B(n_681), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_733), .B(n_728), .Y(n_798) );
NAND3xp33_ASAP7_75t_L g799 ( .A(n_764), .B(n_695), .C(n_715), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_770), .B(n_672), .Y(n_800) );
NAND2xp5_ASAP7_75t_SL g801 ( .A(n_735), .B(n_672), .Y(n_801) );
NOR3xp33_ASAP7_75t_L g802 ( .A(n_758), .B(n_707), .C(n_706), .Y(n_802) );
OAI21xp5_ASAP7_75t_SL g803 ( .A1(n_775), .A2(n_694), .B(n_689), .Y(n_803) );
OAI21xp5_ASAP7_75t_L g804 ( .A1(n_760), .A2(n_710), .B(n_692), .Y(n_804) );
OAI22xp5_ASAP7_75t_L g805 ( .A1(n_763), .A2(n_700), .B1(n_672), .B2(n_727), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_766), .B(n_672), .Y(n_806) );
OAI221xp5_ASAP7_75t_SL g807 ( .A1(n_764), .A2(n_725), .B1(n_684), .B2(n_203), .C(n_205), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_735), .B(n_199), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_767), .B(n_201), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_751), .B(n_206), .Y(n_810) );
NAND3xp33_ASAP7_75t_L g811 ( .A(n_759), .B(n_207), .C(n_208), .Y(n_811) );
AND2x2_ASAP7_75t_L g812 ( .A(n_789), .B(n_209), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_754), .A2(n_746), .B1(n_748), .B2(n_756), .Y(n_813) );
NOR3xp33_ASAP7_75t_SL g814 ( .A(n_783), .B(n_243), .C(n_212), .Y(n_814) );
AND2x2_ASAP7_75t_L g815 ( .A(n_789), .B(n_211), .Y(n_815) );
AND2x2_ASAP7_75t_L g816 ( .A(n_757), .B(n_213), .Y(n_816) );
OAI22xp5_ASAP7_75t_L g817 ( .A1(n_762), .A2(n_217), .B1(n_220), .B2(n_223), .Y(n_817) );
OAI221xp5_ASAP7_75t_SL g818 ( .A1(n_755), .A2(n_225), .B1(n_226), .B2(n_227), .C(n_228), .Y(n_818) );
OAI21xp33_ASAP7_75t_SL g819 ( .A1(n_787), .A2(n_232), .B(n_233), .Y(n_819) );
OAI21xp5_ASAP7_75t_SL g820 ( .A1(n_771), .A2(n_234), .B(n_236), .Y(n_820) );
AND2x2_ASAP7_75t_L g821 ( .A(n_774), .B(n_240), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_761), .B(n_237), .Y(n_822) );
AOI21xp33_ASAP7_75t_SL g823 ( .A1(n_786), .A2(n_238), .B(n_769), .Y(n_823) );
OAI221xp5_ASAP7_75t_SL g824 ( .A1(n_750), .A2(n_749), .B1(n_747), .B2(n_774), .C(n_778), .Y(n_824) );
NAND3xp33_ASAP7_75t_L g825 ( .A(n_739), .B(n_778), .C(n_779), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_779), .B(n_780), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_795), .B(n_780), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_794), .B(n_765), .Y(n_828) );
XNOR2xp5_ASAP7_75t_L g829 ( .A(n_790), .B(n_768), .Y(n_829) );
AO21x2_ASAP7_75t_L g830 ( .A1(n_801), .A2(n_781), .B(n_788), .Y(n_830) );
OR2x2_ASAP7_75t_L g831 ( .A(n_795), .B(n_784), .Y(n_831) );
NOR2x1_ASAP7_75t_R g832 ( .A(n_791), .B(n_776), .Y(n_832) );
OR2x2_ASAP7_75t_L g833 ( .A(n_797), .B(n_785), .Y(n_833) );
HB1xp67_ASAP7_75t_L g834 ( .A(n_798), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_800), .B(n_740), .Y(n_835) );
AND2x2_ASAP7_75t_L g836 ( .A(n_806), .B(n_777), .Y(n_836) );
NAND2xp5_ASAP7_75t_SL g837 ( .A(n_823), .B(n_741), .Y(n_837) );
NOR2xp33_ASAP7_75t_L g838 ( .A(n_805), .B(n_736), .Y(n_838) );
AOI211x1_ASAP7_75t_L g839 ( .A1(n_804), .A2(n_738), .B(n_742), .C(n_743), .Y(n_839) );
BUFx3_ASAP7_75t_L g840 ( .A(n_812), .Y(n_840) );
INVx2_ASAP7_75t_SL g841 ( .A(n_815), .Y(n_841) );
INVx2_ASAP7_75t_L g842 ( .A(n_815), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_813), .A2(n_802), .B1(n_811), .B2(n_810), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g844 ( .A1(n_826), .A2(n_825), .B1(n_793), .B2(n_814), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_813), .B(n_792), .Y(n_845) );
XOR2xp5_ASAP7_75t_L g846 ( .A(n_829), .B(n_809), .Y(n_846) );
INVx2_ASAP7_75t_L g847 ( .A(n_834), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_834), .Y(n_848) );
INVx2_ASAP7_75t_SL g849 ( .A(n_840), .Y(n_849) );
NAND3xp33_ASAP7_75t_L g850 ( .A(n_839), .B(n_803), .C(n_796), .Y(n_850) );
INVx2_ASAP7_75t_L g851 ( .A(n_842), .Y(n_851) );
INVx3_ASAP7_75t_L g852 ( .A(n_840), .Y(n_852) );
NAND4xp75_ASAP7_75t_L g853 ( .A(n_845), .B(n_819), .C(n_821), .D(n_816), .Y(n_853) );
XNOR2xp5_ASAP7_75t_L g854 ( .A(n_843), .B(n_817), .Y(n_854) );
AND2x2_ASAP7_75t_L g855 ( .A(n_841), .B(n_821), .Y(n_855) );
NAND4xp75_ASAP7_75t_L g856 ( .A(n_837), .B(n_808), .C(n_822), .D(n_820), .Y(n_856) );
AND2x2_ASAP7_75t_L g857 ( .A(n_842), .B(n_799), .Y(n_857) );
NAND4xp75_ASAP7_75t_L g858 ( .A(n_838), .B(n_824), .C(n_807), .D(n_818), .Y(n_858) );
XNOR2xp5_ASAP7_75t_L g859 ( .A(n_846), .B(n_844), .Y(n_859) );
INVxp67_ASAP7_75t_L g860 ( .A(n_850), .Y(n_860) );
XOR2x2_ASAP7_75t_L g861 ( .A(n_854), .B(n_843), .Y(n_861) );
HB1xp67_ASAP7_75t_L g862 ( .A(n_847), .Y(n_862) );
INVx2_ASAP7_75t_L g863 ( .A(n_847), .Y(n_863) );
INVxp67_ASAP7_75t_L g864 ( .A(n_857), .Y(n_864) );
OA22x2_ASAP7_75t_L g865 ( .A1(n_860), .A2(n_849), .B1(n_852), .B2(n_857), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_862), .Y(n_866) );
INVx2_ASAP7_75t_L g867 ( .A(n_866), .Y(n_867) );
BUFx2_ASAP7_75t_L g868 ( .A(n_865), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_868), .A2(n_860), .B1(n_861), .B2(n_864), .Y(n_869) );
AOI22xp5_ASAP7_75t_L g870 ( .A1(n_869), .A2(n_859), .B1(n_864), .B2(n_858), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_870), .Y(n_871) );
NAND2xp5_ASAP7_75t_SL g872 ( .A(n_871), .B(n_867), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_872), .Y(n_873) );
INVx2_ASAP7_75t_L g874 ( .A(n_873), .Y(n_874) );
OAI22x1_ASAP7_75t_L g875 ( .A1(n_874), .A2(n_862), .B1(n_848), .B2(n_863), .Y(n_875) );
INVx2_ASAP7_75t_SL g876 ( .A(n_875), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_876), .A2(n_835), .B1(n_852), .B2(n_830), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_877), .Y(n_878) );
AOI22xp5_ASAP7_75t_L g879 ( .A1(n_878), .A2(n_853), .B1(n_856), .B2(n_828), .Y(n_879) );
UNKNOWN g880 ( );
AOI221xp5_ASAP7_75t_L g881 ( .A1(n_880), .A2(n_855), .B1(n_827), .B2(n_836), .C(n_851), .Y(n_881) );
AOI211xp5_ASAP7_75t_L g882 ( .A1(n_881), .A2(n_832), .B(n_833), .C(n_831), .Y(n_882) );
endmodule