module real_jpeg_6975_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_455;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_1),
.A2(n_109),
.B1(n_110),
.B2(n_113),
.Y(n_108)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_1),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_1),
.A2(n_77),
.B1(n_113),
.B2(n_171),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_L g229 ( 
.A1(n_1),
.A2(n_113),
.B1(n_230),
.B2(n_232),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g379 ( 
.A1(n_1),
.A2(n_71),
.B1(n_113),
.B2(n_380),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_2),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_2),
.Y(n_140)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_2),
.Y(n_143)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_2),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_2),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_2),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_2),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_3),
.A2(n_139),
.B1(n_141),
.B2(n_142),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_3),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_3),
.A2(n_122),
.B1(n_141),
.B2(n_278),
.Y(n_277)
);

OAI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_3),
.A2(n_141),
.B1(n_314),
.B2(n_319),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_3),
.A2(n_141),
.B1(n_218),
.B2(n_369),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_5),
.A2(n_140),
.B1(n_189),
.B2(n_191),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_5),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_5),
.A2(n_191),
.B1(n_330),
.B2(n_332),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_5),
.A2(n_191),
.B1(n_269),
.B2(n_314),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_5),
.A2(n_92),
.B1(n_191),
.B2(n_403),
.Y(n_402)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_6),
.A2(n_48),
.B1(n_52),
.B2(n_53),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_6),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_6),
.A2(n_52),
.B1(n_116),
.B2(n_121),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_6),
.A2(n_52),
.B1(n_269),
.B2(n_271),
.Y(n_268)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_7),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_8),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_8),
.Y(n_344)
);

OAI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_9),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_30)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_9),
.A2(n_34),
.B1(n_157),
.B2(n_161),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_10),
.A2(n_146),
.B1(n_147),
.B2(n_149),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_10),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_10),
.A2(n_136),
.B1(n_146),
.B2(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_10),
.A2(n_146),
.B1(n_297),
.B2(n_300),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g324 ( 
.A1(n_10),
.A2(n_31),
.B1(n_146),
.B2(n_325),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_11),
.A2(n_35),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_11),
.A2(n_43),
.B1(n_218),
.B2(n_220),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_12),
.A2(n_74),
.B1(n_75),
.B2(n_79),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_12),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_12),
.A2(n_74),
.B1(n_177),
.B2(n_181),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_12),
.A2(n_74),
.B1(n_209),
.B2(n_211),
.Y(n_208)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_13),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_14),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_14),
.Y(n_133)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_14),
.Y(n_256)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_14),
.Y(n_260)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_15),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_15),
.A2(n_220),
.B1(n_264),
.B2(n_293),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_15),
.B(n_307),
.C(n_310),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_15),
.B(n_101),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_15),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_15),
.B(n_82),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_15),
.B(n_375),
.Y(n_374)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_16),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_236),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_235),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_200),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_20),
.B(n_200),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_153),
.C(n_166),
.Y(n_20)
);

FAx1_ASAP7_75t_SL g282 ( 
.A(n_21),
.B(n_153),
.CI(n_166),
.CON(n_282),
.SN(n_282)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_83),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_22),
.B(n_84),
.C(n_124),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_46),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_23),
.B(n_46),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B1(n_37),
.B2(n_42),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_24),
.A2(n_39),
.B(n_42),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_24),
.A2(n_267),
.B1(n_272),
.B2(n_274),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_24),
.A2(n_313),
.B(n_321),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_24),
.A2(n_264),
.B(n_321),
.Y(n_345)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_25),
.A2(n_176),
.B1(n_183),
.B2(n_184),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_25),
.B(n_324),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_25),
.A2(n_350),
.B1(n_356),
.B2(n_357),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_25),
.A2(n_268),
.B1(n_379),
.B2(n_409),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_30),
.Y(n_183)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_32),
.Y(n_271)
);

INVx8_ASAP7_75t_L g320 ( 
.A(n_32),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_33),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_33),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g342 ( 
.A(n_35),
.Y(n_342)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_36),
.Y(n_182)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_41),
.Y(n_323)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_41),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g310 ( 
.A(n_45),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_57),
.B1(n_73),
.B2(n_82),
.Y(n_46)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_47),
.Y(n_174)
);

NAND2xp33_ASAP7_75t_SL g389 ( 
.A(n_48),
.B(n_390),
.Y(n_389)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_51),
.Y(n_334)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_55),
.Y(n_172)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_57),
.A2(n_73),
.B1(n_82),
.B2(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_57),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_57),
.A2(n_82),
.B1(n_156),
.B2(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_57),
.B(n_296),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_68),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_62),
.B1(n_64),
.B2(n_66),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_68),
.A2(n_329),
.B(n_335),
.Y(n_328)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_78),
.Y(n_160)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_78),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_78),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_78),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_78),
.Y(n_301)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_80),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_82),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_82),
.B(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_124),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_108),
.B1(n_114),
.B2(n_115),
.Y(n_84)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_85),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_85),
.A2(n_114),
.B1(n_277),
.B2(n_402),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_101),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_92),
.B1(n_96),
.B2(n_98),
.Y(n_86)
);

AOI32xp33_ASAP7_75t_L g385 ( 
.A1(n_87),
.A2(n_161),
.A3(n_374),
.B1(n_386),
.B2(n_389),
.Y(n_385)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_92),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_95),
.Y(n_198)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_95),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_97),
.Y(n_391)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_100),
.Y(n_213)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

AOI22x1_ASAP7_75t_L g193 ( 
.A1(n_101),
.A2(n_194),
.B1(n_195),
.B2(n_199),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_101),
.A2(n_194),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

AO22x2_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_104),
.B1(n_105),
.B2(n_107),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_108),
.Y(n_199)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_114),
.B(n_196),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_114),
.A2(n_402),
.B(n_405),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_115),
.Y(n_207)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_SL g372 ( 
.A1(n_117),
.A2(n_264),
.B(n_373),
.Y(n_372)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_120),
.Y(n_252)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_120),
.Y(n_262)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_120),
.Y(n_388)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_120),
.Y(n_404)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_123),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_138),
.B(n_144),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_125),
.A2(n_138),
.B1(n_188),
.B2(n_192),
.Y(n_187)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_126),
.B(n_145),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_126),
.A2(n_425),
.B(n_427),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_134),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_134)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_133),
.Y(n_137)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_142),
.Y(n_231)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_144),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_152),
.Y(n_144)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_150),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_150),
.B(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_152),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_152),
.B(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_164),
.B2(n_165),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_155),
.B(n_164),
.Y(n_224)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_160),
.Y(n_299)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_160),
.Y(n_305)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx5_ASAP7_75t_L g294 ( 
.A(n_163),
.Y(n_294)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_164),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_164),
.A2(n_165),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_186),
.C(n_193),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_167),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_175),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_168),
.B(n_175),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_173),
.B2(n_174),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_169),
.A2(n_292),
.B(n_295),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_169),
.A2(n_173),
.B1(n_329),
.B2(n_368),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_169),
.A2(n_295),
.B(n_368),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_170),
.A2(n_173),
.B(n_335),
.Y(n_430)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_171),
.Y(n_369)
);

INVx5_ASAP7_75t_SL g171 ( 
.A(n_172),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_176),
.Y(n_274)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_179),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_185),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_186),
.A2(n_187),
.B1(n_193),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_188),
.A2(n_192),
.B(n_234),
.Y(n_247)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_189),
.Y(n_426)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_192),
.B(n_264),
.Y(n_407)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_193),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_194),
.A2(n_276),
.B(n_281),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_194),
.A2(n_281),
.B(n_372),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_194),
.B(n_195),
.Y(n_405)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_222),
.B2(n_223),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_214),
.B(n_221),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_215),
.Y(n_221)
);

INVx4_ASAP7_75t_SL g209 ( 
.A(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_234),
.Y(n_227)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_283),
.B(n_455),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_282),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_239),
.B(n_282),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_244),
.C(n_245),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_240),
.A2(n_241),
.B1(n_244),
.B2(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_244),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_245),
.B(n_445),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_248),
.C(n_275),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_246),
.A2(n_247),
.B1(n_275),
.B2(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_248),
.B(n_439),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_265),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_249),
.A2(n_265),
.B1(n_266),
.B2(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_249),
.Y(n_418)
);

OAI32xp33_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_253),
.A3(n_255),
.B1(n_257),
.B2(n_263),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_261),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

OAI21xp33_ASAP7_75t_SL g425 ( 
.A1(n_263),
.A2(n_264),
.B(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_275),
.Y(n_440)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx24_ASAP7_75t_SL g457 ( 
.A(n_282),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_433),
.B(n_452),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

AOI21x1_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_413),
.B(n_432),
.Y(n_285)
);

AO21x1_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_393),
.B(n_412),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_362),
.B(n_392),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_338),
.B(n_361),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_311),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_290),
.B(n_311),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_302),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_291),
.A2(n_302),
.B1(n_303),
.B2(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_291),
.Y(n_359)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_294),
.Y(n_331)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_306),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_326),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_312),
.B(n_327),
.C(n_337),
.Y(n_363)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_313),
.Y(n_357)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_316),
.Y(n_325)
);

INVx6_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx5_ASAP7_75t_L g382 ( 
.A(n_318),
.Y(n_382)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_324),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_327),
.A2(n_328),
.B1(n_336),
.B2(n_337),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_354),
.B(n_360),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_346),
.B(n_353),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_345),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_344),
.Y(n_350)
);

INVx4_ASAP7_75t_L g384 ( 
.A(n_344),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_347),
.B(n_352),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_347),
.B(n_352),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_349),
.B(n_351),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_348),
.Y(n_356)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_351),
.A2(n_378),
.B(n_383),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_358),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_355),
.B(n_358),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_364),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_363),
.B(n_364),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_376),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_366),
.A2(n_367),
.B1(n_370),
.B2(n_371),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_367),
.B(n_370),
.C(n_376),
.Y(n_394)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVxp33_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_385),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_377),
.B(n_385),
.Y(n_399)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx3_ASAP7_75t_SL g383 ( 
.A(n_384),
.Y(n_383)
);

INVx5_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_395),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_394),
.B(n_395),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_397),
.B1(n_400),
.B2(n_411),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_398),
.B(n_399),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_398),
.B(n_399),
.C(n_411),
.Y(n_414)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_400),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_SL g400 ( 
.A(n_401),
.B(n_406),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_401),
.B(n_407),
.C(n_408),
.Y(n_419)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_408),
.Y(n_406)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_415),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_414),
.B(n_415),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_422),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_417),
.A2(n_419),
.B1(n_420),
.B2(n_421),
.Y(n_416)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_417),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_419),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_419),
.B(n_420),
.C(n_422),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_423),
.A2(n_424),
.B1(n_428),
.B2(n_431),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_423),
.B(n_429),
.C(n_430),
.Y(n_443)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_428),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g428 ( 
.A(n_429),
.B(n_430),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_435),
.B(n_447),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_436),
.A2(n_453),
.B(n_454),
.Y(n_452)
);

NOR2x1_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_444),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_437),
.B(n_444),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_441),
.C(n_443),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_438),
.B(n_450),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_441),
.A2(n_442),
.B1(n_443),
.B2(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_443),
.Y(n_451)
);

OR2x2_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_449),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_448),
.B(n_449),
.Y(n_453)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);


endmodule