module fake_jpeg_26669_n_291 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_291);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_291;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_11),
.B(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_38),
.Y(n_52)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_17),
.Y(n_39)
);

INVx5_ASAP7_75t_SL g45 ( 
.A(n_39),
.Y(n_45)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_50),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_22),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_43),
.B(n_48),
.Y(n_87)
);

OAI21xp33_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_17),
.B(n_30),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_44),
.A2(n_28),
.B(n_21),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_38),
.A2(n_30),
.B1(n_18),
.B2(n_29),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_41),
.B1(n_30),
.B2(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_26),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_26),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_39),
.B(n_27),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_53),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_28),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_55),
.Y(n_85)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_56),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_35),
.B(n_24),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_60),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_25),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_30),
.B1(n_21),
.B2(n_31),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_61),
.A2(n_47),
.B1(n_58),
.B2(n_28),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_64),
.A2(n_66),
.B1(n_45),
.B2(n_51),
.Y(n_97)
);

AOI32xp33_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_41),
.A3(n_37),
.B1(n_32),
.B2(n_27),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_79),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_18),
.B1(n_24),
.B2(n_31),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_22),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_73),
.B(n_61),
.Y(n_95)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_78),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_22),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_18),
.B1(n_32),
.B2(n_19),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_75),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_59),
.C(n_52),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_82),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_44),
.B(n_61),
.C(n_60),
.Y(n_93)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_45),
.A2(n_19),
.B1(n_25),
.B2(n_29),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_45),
.A2(n_31),
.B1(n_24),
.B2(n_21),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_86),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_22),
.Y(n_112)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_90),
.B(n_92),
.Y(n_125)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_SL g118 ( 
.A(n_93),
.B(n_66),
.C(n_81),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_99),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_70),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_96),
.B(n_70),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_97),
.A2(n_112),
.B1(n_89),
.B2(n_67),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_50),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_104),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_63),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_105),
.Y(n_134)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_63),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_62),
.Y(n_107)
);

FAx1_ASAP7_75t_SL g126 ( 
.A(n_107),
.B(n_113),
.CI(n_115),
.CON(n_126),
.SN(n_126)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_77),
.B(n_20),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_111),
.B(n_99),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_62),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_88),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_62),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_116),
.B(n_121),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_118),
.A2(n_124),
.B(n_135),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_108),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_119),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_SL g159 ( 
.A1(n_120),
.A2(n_142),
.B(n_115),
.Y(n_159)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

BUFx24_ASAP7_75t_SL g122 ( 
.A(n_99),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_122),
.B(n_123),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_76),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_112),
.A2(n_73),
.B1(n_67),
.B2(n_71),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_127),
.A2(n_110),
.B1(n_93),
.B2(n_112),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_114),
.A2(n_71),
.B1(n_67),
.B2(n_73),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_112),
.B1(n_97),
.B2(n_101),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_109),
.Y(n_129)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_100),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_94),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_138),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_69),
.Y(n_133)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

BUFx8_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

INVx3_ASAP7_75t_SL g156 ( 
.A(n_136),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_73),
.C(n_83),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_141),
.C(n_95),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_107),
.B(n_83),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_82),
.Y(n_139)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_33),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_95),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_80),
.C(n_55),
.Y(n_141)
);

NOR3xp33_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_42),
.C(n_46),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_151),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_127),
.C(n_126),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_94),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_147),
.A2(n_149),
.B(n_154),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_132),
.A2(n_110),
.B(n_93),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_157),
.Y(n_175)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_159),
.Y(n_181)
);

AND2x6_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_101),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_165),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_105),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_163),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_101),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_126),
.B1(n_130),
.B2(n_103),
.Y(n_183)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_132),
.A2(n_91),
.B(n_104),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_166),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_141),
.A2(n_119),
.B(n_137),
.C(n_124),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_167),
.A2(n_154),
.B1(n_163),
.B2(n_166),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_98),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_72),
.Y(n_188)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_125),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_57),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_128),
.A2(n_98),
.B1(n_103),
.B2(n_75),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_171),
.A2(n_75),
.B1(n_129),
.B2(n_109),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_173),
.B(n_177),
.C(n_185),
.Y(n_200)
);

INVxp33_ASAP7_75t_SL g174 ( 
.A(n_156),
.Y(n_174)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_155),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_178),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_126),
.C(n_121),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_147),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_161),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_186),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_183),
.A2(n_186),
.B1(n_191),
.B2(n_189),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_96),
.C(n_72),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_187),
.A2(n_196),
.B1(n_157),
.B2(n_153),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_188),
.B(n_189),
.Y(n_215)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_190),
.B(n_144),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_144),
.B(n_57),
.Y(n_191)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

A2O1A1O1Ixp25_ASAP7_75t_L g192 ( 
.A1(n_149),
.A2(n_136),
.B(n_33),
.C(n_20),
.D(n_4),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_192),
.B(n_164),
.Y(n_199)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_152),
.Y(n_207)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_178),
.B(n_150),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_198),
.Y(n_226)
);

NOR3xp33_ASAP7_75t_SL g237 ( 
.A(n_199),
.B(n_9),
.C(n_14),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_148),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_203),
.A2(n_213),
.B(n_8),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_167),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_218),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_205),
.A2(n_209),
.B1(n_183),
.B2(n_195),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_219),
.Y(n_228)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_175),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_217),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_196),
.A2(n_170),
.B1(n_160),
.B2(n_167),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_143),
.C(n_168),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_212),
.C(n_194),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_211),
.A2(n_172),
.B1(n_176),
.B2(n_187),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_170),
.C(n_151),
.Y(n_212)
);

AND2x6_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_158),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_145),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_214),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_20),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_136),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_216),
.A2(n_195),
.B(n_194),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_220),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_227),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_222),
.B(n_233),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_223),
.A2(n_224),
.B1(n_236),
.B2(n_213),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_205),
.A2(n_172),
.B1(n_182),
.B2(n_181),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_204),
.B(n_192),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_231),
.Y(n_239)
);

A2O1A1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_202),
.A2(n_193),
.B(n_156),
.C(n_10),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_20),
.C(n_9),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_210),
.C(n_201),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_212),
.B(n_8),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_209),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_7),
.Y(n_248)
);

FAx1_ASAP7_75t_SL g238 ( 
.A(n_225),
.B(n_200),
.CI(n_199),
.CON(n_238),
.SN(n_238)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_233),
.A2(n_216),
.B(n_203),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_222),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_246),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_218),
.C(n_215),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_230),
.C(n_224),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_206),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_248),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_244),
.A2(n_228),
.B1(n_10),
.B2(n_11),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_7),
.Y(n_246)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_234),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_249),
.A2(n_229),
.B1(n_237),
.B2(n_227),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_0),
.Y(n_250)
);

INVxp33_ASAP7_75t_L g258 ( 
.A(n_250),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_252),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_253),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_247),
.A2(n_226),
.B1(n_223),
.B2(n_220),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_254),
.A2(n_245),
.B1(n_239),
.B2(n_246),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_235),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_260),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_231),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_262),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_245),
.B(n_6),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_263),
.A2(n_250),
.B(n_239),
.Y(n_271)
);

NOR2xp67_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_240),
.Y(n_264)
);

A2O1A1O1Ixp25_ASAP7_75t_L g279 ( 
.A1(n_264),
.A2(n_266),
.B(n_269),
.C(n_268),
.D(n_267),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_241),
.C(n_242),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_270),
.Y(n_278)
);

OAI21xp33_ASAP7_75t_SL g269 ( 
.A1(n_255),
.A2(n_251),
.B(n_243),
.Y(n_269)
);

AOI322xp5_ASAP7_75t_L g277 ( 
.A1(n_269),
.A2(n_258),
.A3(n_5),
.B1(n_4),
.B2(n_12),
.C1(n_13),
.C2(n_15),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_257),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_249),
.C(n_11),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_256),
.C(n_260),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_276),
.C(n_1),
.Y(n_283)
);

OAI211xp5_ASAP7_75t_L g282 ( 
.A1(n_275),
.A2(n_277),
.B(n_279),
.C(n_0),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_258),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_265),
.B(n_15),
.Y(n_280)
);

INVxp33_ASAP7_75t_L g284 ( 
.A(n_280),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_278),
.A2(n_272),
.B(n_15),
.Y(n_281)
);

AOI21xp33_ASAP7_75t_L g287 ( 
.A1(n_281),
.A2(n_283),
.B(n_285),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_282),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_280),
.A2(n_1),
.B(n_2),
.Y(n_285)
);

BUFx24_ASAP7_75t_SL g288 ( 
.A(n_286),
.Y(n_288)
);

AOI322xp5_ASAP7_75t_L g289 ( 
.A1(n_288),
.A2(n_1),
.A3(n_2),
.B1(n_284),
.B2(n_287),
.C1(n_282),
.C2(n_213),
.Y(n_289)
);

BUFx24_ASAP7_75t_SL g290 ( 
.A(n_289),
.Y(n_290)
);

BUFx24_ASAP7_75t_SL g291 ( 
.A(n_290),
.Y(n_291)
);


endmodule