module fake_netlist_6_4393_n_200 (n_7, n_6, n_12, n_4, n_2, n_3, n_5, n_1, n_0, n_9, n_11, n_8, n_10, n_200);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_3;
input n_5;
input n_1;
input n_0;
input n_9;
input n_11;
input n_8;
input n_10;

output n_200;

wire n_52;
wire n_16;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_21;
wire n_18;
wire n_193;
wire n_147;
wire n_154;
wire n_191;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_199;
wire n_161;
wire n_22;
wire n_138;
wire n_68;
wire n_166;
wire n_28;
wire n_184;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_153;
wire n_168;
wire n_125;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_24;
wire n_131;
wire n_105;
wire n_54;
wire n_132;
wire n_188;
wire n_102;
wire n_186;
wire n_87;
wire n_195;
wire n_189;
wire n_32;
wire n_66;
wire n_85;
wire n_130;
wire n_78;
wire n_84;
wire n_99;
wire n_164;
wire n_100;
wire n_129;
wire n_13;
wire n_121;
wire n_197;
wire n_137;
wire n_23;
wire n_17;
wire n_142;
wire n_20;
wire n_143;
wire n_180;
wire n_19;
wire n_47;
wire n_62;
wire n_29;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_15;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_151;
wire n_110;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_181;
wire n_76;
wire n_36;
wire n_182;
wire n_26;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_108;
wire n_94;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_196;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_198;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_190;
wire n_14;
wire n_123;
wire n_136;
wire n_72;
wire n_187;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_35;
wire n_183;
wire n_115;
wire n_69;
wire n_128;
wire n_30;
wire n_79;
wire n_43;
wire n_194;
wire n_171;
wire n_31;
wire n_192;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVxp67_ASAP7_75t_SL g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_23),
.B(n_22),
.Y(n_27)
);

CKINVDCx5p33_ASAP7_75t_R g28 ( 
.A(n_23),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_20),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_25),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_33),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NAND2x1p5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_25),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_28),
.B(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_14),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_19),
.Y(n_44)
);

AND2x4_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_19),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_18),
.B1(n_17),
.B2(n_15),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_17),
.B(n_0),
.C(n_5),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_4),
.B(n_7),
.C(n_9),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_4),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_12),
.Y(n_51)
);

NOR2x1p5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_7),
.Y(n_52)
);

AOI22x1_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_38),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_37),
.Y(n_55)
);

NAND2x1p5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_35),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_35),
.Y(n_59)
);

OR2x6_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_44),
.Y(n_60)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

AOI21x1_ASAP7_75t_L g63 ( 
.A1(n_34),
.A2(n_35),
.B(n_37),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_39),
.B1(n_36),
.B2(n_40),
.Y(n_64)
);

OR2x6_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_42),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_34),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_43),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

AOI21x1_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_43),
.B(n_63),
.Y(n_70)
);

AOI21x1_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_51),
.B(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_55),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

AO21x1_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_56),
.B(n_64),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

AO21x2_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_48),
.B(n_61),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_SL g78 ( 
.A1(n_47),
.A2(n_48),
.B(n_57),
.C(n_53),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_52),
.Y(n_79)
);

OAI21x1_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_63),
.B(n_57),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

OAI21x1_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_63),
.B(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_54),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_50),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_59),
.Y(n_85)
);

AO21x2_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_51),
.B(n_49),
.Y(n_86)
);

AOI21x1_ASAP7_75t_L g87 ( 
.A1(n_50),
.A2(n_62),
.B(n_63),
.Y(n_87)
);

AND2x4_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_50),
.Y(n_88)
);

OAI21x1_ASAP7_75t_L g89 ( 
.A1(n_63),
.A2(n_57),
.B(n_56),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_72),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_85),
.Y(n_92)
);

OAI21x1_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_80),
.B(n_87),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_65),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_72),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_67),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_65),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_76),
.Y(n_102)
);

CKINVDCx12_ASAP7_75t_R g103 ( 
.A(n_65),
.Y(n_103)
);

AND2x4_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_81),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_76),
.A2(n_74),
.B1(n_88),
.B2(n_73),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_65),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_73),
.A2(n_79),
.B1(n_81),
.B2(n_84),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_73),
.A2(n_74),
.B1(n_76),
.B2(n_78),
.Y(n_111)
);

AND2x4_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_109),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

AO21x2_ASAP7_75t_L g114 ( 
.A1(n_111),
.A2(n_80),
.B(n_71),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

OA21x2_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_82),
.B(n_89),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_73),
.B1(n_111),
.B2(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

OAI21x1_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_82),
.B(n_71),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_97),
.A2(n_77),
.B1(n_68),
.B2(n_86),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_70),
.B(n_86),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_86),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_90),
.A2(n_70),
.B(n_77),
.C(n_95),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_90),
.A2(n_77),
.B1(n_95),
.B2(n_106),
.Y(n_127)
);

AO21x2_ASAP7_75t_L g128 ( 
.A1(n_93),
.A2(n_77),
.B(n_108),
.Y(n_128)
);

AND2x4_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_77),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

AND2x4_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_104),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_101),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_R g135 ( 
.A(n_124),
.B(n_92),
.Y(n_135)
);

AND2x4_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_104),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

AND2x4_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_104),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_94),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_112),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_109),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_96),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_107),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_133),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

AOI33xp33_ASAP7_75t_L g150 ( 
.A1(n_131),
.A2(n_127),
.A3(n_118),
.B1(n_121),
.B2(n_143),
.B3(n_141),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_94),
.Y(n_151)
);

AND2x4_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_129),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_151),
.A2(n_99),
.B1(n_106),
.B2(n_103),
.Y(n_153)
);

OAI31xp33_ASAP7_75t_L g154 ( 
.A1(n_145),
.A2(n_107),
.A3(n_118),
.B(n_108),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_134),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_152),
.A2(n_99),
.B1(n_103),
.B2(n_127),
.Y(n_159)
);

INVxp67_ASAP7_75t_SL g160 ( 
.A(n_149),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_161),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_157),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_150),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_157),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_128),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_155),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_153),
.Y(n_169)
);

AND4x1_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_154),
.C(n_159),
.D(n_126),
.Y(n_170)
);

AOI221xp5_ASAP7_75t_L g171 ( 
.A1(n_169),
.A2(n_160),
.B1(n_135),
.B2(n_158),
.C(n_147),
.Y(n_171)
);

OAI211xp5_ASAP7_75t_SL g172 ( 
.A1(n_168),
.A2(n_126),
.B(n_147),
.C(n_148),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_165),
.A2(n_152),
.B1(n_140),
.B2(n_138),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_167),
.Y(n_174)
);

AND2x4_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_152),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_166),
.B(n_138),
.Y(n_176)
);

OAI211xp5_ASAP7_75t_L g177 ( 
.A1(n_163),
.A2(n_121),
.B(n_105),
.C(n_142),
.Y(n_177)
);

OAI221xp5_ASAP7_75t_L g178 ( 
.A1(n_163),
.A2(n_142),
.B1(n_122),
.B2(n_137),
.C(n_119),
.Y(n_178)
);

NOR2x1p5_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_167),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_172),
.A2(n_128),
.B(n_122),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_171),
.A2(n_173),
.B1(n_176),
.B2(n_177),
.Y(n_181)
);

NAND3xp33_ASAP7_75t_SL g182 ( 
.A(n_170),
.B(n_166),
.C(n_137),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_128),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_128),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_181),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_138),
.Y(n_186)
);

CKINVDCx8_ASAP7_75t_R g187 ( 
.A(n_179),
.Y(n_187)
);

AND3x4_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_136),
.C(n_133),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_187),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_185),
.A2(n_180),
.B1(n_183),
.B2(n_128),
.Y(n_190)
);

OAI22x1_ASAP7_75t_L g191 ( 
.A1(n_188),
.A2(n_136),
.B1(n_116),
.B2(n_129),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_186),
.A2(n_120),
.B(n_136),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_187),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_114),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_193),
.A2(n_129),
.B1(n_119),
.B2(n_116),
.Y(n_195)
);

AO21x2_ASAP7_75t_L g196 ( 
.A1(n_189),
.A2(n_190),
.B(n_192),
.Y(n_196)
);

AOI221xp5_ASAP7_75t_SL g197 ( 
.A1(n_195),
.A2(n_191),
.B1(n_194),
.B2(n_190),
.C(n_115),
.Y(n_197)
);

NAND5xp2_ASAP7_75t_L g198 ( 
.A(n_196),
.B(n_110),
.C(n_104),
.D(n_114),
.E(n_112),
.Y(n_198)
);

XOR2x2_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_114),
.Y(n_199)
);

NOR4xp25_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_198),
.C(n_125),
.D(n_123),
.Y(n_200)
);


endmodule