module fake_netlist_1_9223_n_37 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_37);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_37;
wire n_20;
wire n_36;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_30;
wire n_26;
wire n_13;
wire n_16;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
INVx1_ASAP7_75t_L g11 ( .A(n_0), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_2), .Y(n_12) );
INVxp67_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_10), .B(n_6), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_10), .Y(n_15) );
NOR2x1p5_ASAP7_75t_L g16 ( .A(n_1), .B(n_2), .Y(n_16) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_9), .Y(n_17) );
INVx4_ASAP7_75t_L g18 ( .A(n_14), .Y(n_18) );
AOI21xp5_ASAP7_75t_L g19 ( .A1(n_12), .A2(n_0), .B(n_1), .Y(n_19) );
AOI21xp5_ASAP7_75t_L g20 ( .A1(n_12), .A2(n_3), .B(n_4), .Y(n_20) );
AOI22xp5_ASAP7_75t_L g21 ( .A1(n_14), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_21) );
NOR2xp33_ASAP7_75t_L g22 ( .A(n_13), .B(n_15), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_19), .Y(n_23) );
NAND2xp33_ASAP7_75t_R g24 ( .A(n_22), .B(n_14), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_18), .B(n_12), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_25), .B(n_13), .Y(n_26) );
NAND2xp5_ASAP7_75t_SL g27 ( .A(n_25), .B(n_20), .Y(n_27) );
AND2x4_ASAP7_75t_L g28 ( .A(n_25), .B(n_21), .Y(n_28) );
INVxp67_ASAP7_75t_L g29 ( .A(n_26), .Y(n_29) );
AND2x2_ASAP7_75t_L g30 ( .A(n_28), .B(n_23), .Y(n_30) );
O2A1O1Ixp33_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_27), .B(n_28), .C(n_23), .Y(n_31) );
AOI22xp5_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_24), .B1(n_17), .B2(n_16), .Y(n_32) );
INVxp67_ASAP7_75t_L g33 ( .A(n_32), .Y(n_33) );
NAND2xp5_ASAP7_75t_L g34 ( .A(n_31), .B(n_30), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_34), .Y(n_35) );
OAI22xp5_ASAP7_75t_SL g36 ( .A1(n_33), .A2(n_11), .B1(n_6), .B2(n_7), .Y(n_36) );
AOI22xp33_ASAP7_75t_L g37 ( .A1(n_35), .A2(n_5), .B1(n_9), .B2(n_36), .Y(n_37) );
endmodule