module fake_jpeg_22461_n_276 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_276);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_276;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_30),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_38),
.B(n_22),
.Y(n_59)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx2_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_28),
.B1(n_18),
.B2(n_22),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_23),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_43),
.Y(n_77)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_47),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_59),
.Y(n_69)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

INVxp67_ASAP7_75t_SL g87 ( 
.A(n_49),
.Y(n_87)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_23),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_54),
.A2(n_26),
.B(n_37),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_40),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_56),
.A2(n_60),
.B1(n_61),
.B2(n_36),
.Y(n_66)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_28),
.B1(n_34),
.B2(n_18),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_64),
.A2(n_65),
.B1(n_68),
.B2(n_71),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_28),
.B1(n_34),
.B2(n_16),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

BUFx24_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_41),
.B1(n_36),
.B2(n_39),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_17),
.B1(n_20),
.B2(n_21),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_74),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_61),
.A2(n_37),
.B1(n_39),
.B2(n_36),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_79),
.A2(n_83),
.B1(n_45),
.B2(n_57),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_81),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_82),
.A2(n_85),
.B1(n_42),
.B2(n_27),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_36),
.B1(n_52),
.B2(n_39),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_30),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_86),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_45),
.A2(n_42),
.B1(n_37),
.B2(n_30),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_19),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_87),
.B(n_24),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_88),
.B(n_21),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_61),
.B(n_29),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_89),
.A2(n_88),
.B(n_100),
.Y(n_126)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_92),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_80),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_93),
.Y(n_117)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_96),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_67),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_97),
.A2(n_111),
.B1(n_74),
.B2(n_72),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_58),
.C(n_37),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_100),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_69),
.B(n_57),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_42),
.Y(n_104)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

NAND2xp33_ASAP7_75t_SL g105 ( 
.A(n_82),
.B(n_1),
.Y(n_105)
);

AO21x1_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_20),
.B(n_24),
.Y(n_120)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_107),
.Y(n_132)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

INVx3_ASAP7_75t_SL g110 ( 
.A(n_72),
.Y(n_110)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_104),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_113),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_102),
.Y(n_113)
);

AO21x2_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_85),
.B(n_78),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_109),
.B1(n_94),
.B2(n_108),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_91),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_115),
.Y(n_139)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_123),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_96),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_118),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_120),
.A2(n_89),
.B(n_29),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_107),
.A2(n_75),
.B1(n_85),
.B2(n_77),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_124),
.B1(n_125),
.B2(n_129),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_95),
.A2(n_85),
.B1(n_77),
.B2(n_70),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_111),
.A2(n_70),
.B1(n_42),
.B2(n_78),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_126),
.A2(n_33),
.B(n_32),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_92),
.A2(n_50),
.B1(n_74),
.B2(n_72),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_101),
.A2(n_103),
.B1(n_99),
.B2(n_106),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_131),
.A2(n_137),
.B1(n_98),
.B2(n_93),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_102),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_135),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_94),
.B1(n_110),
.B2(n_108),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_31),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_103),
.A2(n_74),
.B1(n_16),
.B2(n_17),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_141),
.Y(n_166)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_142),
.A2(n_152),
.B(n_159),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_131),
.A2(n_98),
.B1(n_105),
.B2(n_90),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_143),
.A2(n_145),
.B1(n_113),
.B2(n_32),
.Y(n_188)
);

XNOR2x1_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_114),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_146),
.B(n_33),
.Y(n_186)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_157),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_148),
.A2(n_149),
.B1(n_130),
.B2(n_164),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_114),
.A2(n_110),
.B(n_109),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_31),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_121),
.C(n_124),
.Y(n_171)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_158),
.B(n_19),
.Y(n_175)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_126),
.A2(n_31),
.B(n_32),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_115),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_162),
.B(n_135),
.Y(n_184)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_114),
.A2(n_31),
.B(n_33),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_123),
.B(n_33),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_165),
.A2(n_173),
.B1(n_174),
.B2(n_185),
.Y(n_199)
);

AO21x1_ASAP7_75t_L g167 ( 
.A1(n_163),
.A2(n_120),
.B(n_137),
.Y(n_167)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_125),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_171),
.C(n_177),
.Y(n_192)
);

XOR2x1_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_121),
.Y(n_173)
);

O2A1O1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_152),
.A2(n_136),
.B(n_130),
.C(n_123),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_175),
.B(n_176),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_139),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_133),
.C(n_123),
.Y(n_177)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_182),
.Y(n_206)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_183),
.A2(n_187),
.B1(n_188),
.B2(n_140),
.Y(n_190)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_156),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_147),
.A2(n_113),
.B(n_2),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_193),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_195),
.Y(n_217)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_174),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_143),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_140),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_200),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_185),
.A2(n_161),
.B1(n_142),
.B2(n_159),
.Y(n_197)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_166),
.B(n_153),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_198),
.B(n_182),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_171),
.B(n_151),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_141),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_1),
.Y(n_221)
);

INVxp33_ASAP7_75t_SL g202 ( 
.A(n_178),
.Y(n_202)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_138),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_204),
.C(n_207),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_157),
.C(n_160),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_81),
.C(n_32),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_169),
.B(n_27),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_209),
.C(n_179),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_27),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_202),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_210),
.B(n_221),
.Y(n_229)
);

OAI322xp33_ASAP7_75t_L g211 ( 
.A1(n_206),
.A2(n_167),
.A3(n_183),
.B1(n_172),
.B2(n_188),
.C1(n_187),
.C2(n_170),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_211),
.B(n_4),
.Y(n_235)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_4),
.Y(n_233)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_216),
.A2(n_4),
.B(n_5),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_179),
.C(n_181),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_204),
.C(n_192),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_199),
.A2(n_170),
.B1(n_180),
.B2(n_81),
.Y(n_220)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_3),
.Y(n_222)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_3),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_226),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_27),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_213),
.C(n_225),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_218),
.A2(n_196),
.B1(n_203),
.B2(n_208),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_228),
.A2(n_225),
.B1(n_217),
.B2(n_226),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_224),
.A2(n_191),
.B1(n_209),
.B2(n_19),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_230),
.A2(n_236),
.B1(n_6),
.B2(n_8),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_232),
.A2(n_214),
.B(n_215),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_235),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_223),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_236),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_214),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_240),
.A2(n_247),
.B1(n_238),
.B2(n_229),
.Y(n_251)
);

FAx1_ASAP7_75t_SL g241 ( 
.A(n_228),
.B(n_213),
.CI(n_219),
.CON(n_241),
.SN(n_241)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_233),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_242),
.A2(n_245),
.B(n_249),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_237),
.A2(n_231),
.B1(n_216),
.B2(n_235),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_243),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_244),
.B(n_250),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_217),
.C(n_7),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_11),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_239),
.A2(n_6),
.B(n_8),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_230),
.A2(n_9),
.B(n_10),
.Y(n_250)
);

AOI221xp5_ASAP7_75t_L g260 ( 
.A1(n_251),
.A2(n_244),
.B1(n_246),
.B2(n_241),
.C(n_245),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_241),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_257),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_255),
.B(n_256),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_10),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_259),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_250),
.B(n_246),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_254),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_252),
.B(n_242),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_265),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_13),
.Y(n_265)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_266),
.Y(n_271)
);

AOI21xp33_ASAP7_75t_L g267 ( 
.A1(n_262),
.A2(n_258),
.B(n_14),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_267),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_13),
.C(n_15),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_271),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_269),
.C(n_264),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_270),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_274),
.B(n_268),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_15),
.Y(n_276)
);


endmodule