module fake_ibex_1529_n_4 (n_1, n_0, n_4);

input n_1;
input n_0;

output n_4;



endmodule