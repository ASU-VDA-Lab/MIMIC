module fake_jpeg_14806_n_314 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_314);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx2_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

INVx11_ASAP7_75t_SL g16 ( 
.A(n_9),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

AOI21xp33_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_13),
.B(n_12),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_36),
.Y(n_43)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_34),
.B(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_22),
.Y(n_46)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_29),
.A2(n_25),
.B1(n_17),
.B2(n_22),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_31),
.B1(n_35),
.B2(n_18),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_53),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_22),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_38),
.B(n_16),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_14),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_29),
.B1(n_38),
.B2(n_33),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_69),
.B1(n_72),
.B2(n_75),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_55),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_58),
.B(n_74),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_14),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_64),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_45),
.A2(n_29),
.B1(n_25),
.B2(n_33),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_63),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_29),
.B1(n_25),
.B2(n_33),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_33),
.B1(n_35),
.B2(n_17),
.Y(n_66)
);

O2A1O1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_53),
.B(n_51),
.C(n_49),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_68),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_41),
.A2(n_35),
.B1(n_20),
.B2(n_28),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_39),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_71),
.B(n_76),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_42),
.A2(n_30),
.B1(n_36),
.B2(n_31),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_37),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_45),
.A2(n_28),
.B1(n_14),
.B2(n_26),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_50),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_48),
.A2(n_26),
.B1(n_24),
.B2(n_27),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_77),
.A2(n_18),
.B1(n_15),
.B2(n_19),
.Y(n_97)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_98),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_59),
.B(n_26),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_86),
.B(n_23),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_58),
.A2(n_55),
.B1(n_40),
.B2(n_48),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_93),
.B1(n_70),
.B2(n_73),
.Y(n_114)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_78),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_88),
.A2(n_73),
.B1(n_57),
.B2(n_31),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_58),
.A2(n_19),
.B(n_27),
.C(n_24),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_101),
.Y(n_103)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_74),
.B(n_14),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_59),
.C(n_62),
.Y(n_112)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_61),
.A2(n_40),
.B1(n_30),
.B2(n_50),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_69),
.A2(n_40),
.B1(n_31),
.B2(n_30),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_94),
.A2(n_67),
.B1(n_66),
.B2(n_77),
.Y(n_107)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_75),
.B(n_71),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_76),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_80),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_104),
.B(n_105),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_85),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_107),
.A2(n_114),
.B1(n_101),
.B2(n_79),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_100),
.A2(n_74),
.B1(n_68),
.B2(n_71),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_108),
.A2(n_82),
.B1(n_93),
.B2(n_101),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_109),
.A2(n_121),
.B(n_122),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_68),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_70),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_123),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_116),
.B(n_125),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_97),
.B(n_83),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_86),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_72),
.C(n_50),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_91),
.Y(n_136)
);

OR2x2_ASAP7_75t_SL g121 ( 
.A(n_89),
.B(n_19),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_100),
.A2(n_19),
.B(n_15),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_65),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_84),
.B(n_50),
.Y(n_125)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_96),
.Y(n_129)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_151),
.B(n_122),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_80),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_133),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_115),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_87),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_110),
.B(n_114),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_72),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_81),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_137),
.B(n_139),
.Y(n_178)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_89),
.Y(n_141)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_142),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_143),
.A2(n_125),
.B1(n_105),
.B2(n_118),
.Y(n_165)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_101),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_148),
.Y(n_157)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_124),
.A2(n_79),
.B1(n_82),
.B2(n_83),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_109),
.A2(n_94),
.B1(n_85),
.B2(n_81),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_152),
.A2(n_123),
.B1(n_120),
.B2(n_107),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_156),
.B(n_163),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_158),
.A2(n_161),
.B(n_168),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_128),
.A2(n_122),
.B(n_108),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_162),
.Y(n_183)
);

MAJx2_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_112),
.C(n_121),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_151),
.A2(n_143),
.B1(n_128),
.B2(n_130),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_164),
.A2(n_160),
.B1(n_158),
.B2(n_156),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_165),
.A2(n_180),
.B1(n_144),
.B2(n_149),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_116),
.Y(n_167)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_135),
.A2(n_113),
.B(n_121),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_135),
.A2(n_127),
.B(n_141),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_170),
.A2(n_147),
.B(n_18),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_134),
.A2(n_113),
.B1(n_88),
.B2(n_92),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_171),
.A2(n_176),
.B1(n_15),
.B2(n_21),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_63),
.Y(n_172)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_132),
.C(n_136),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_134),
.A2(n_15),
.B1(n_18),
.B2(n_21),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_129),
.B(n_138),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_179),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_37),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_0),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_169),
.Y(n_217)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_184),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_145),
.C(n_140),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_191),
.C(n_203),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_186),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_146),
.Y(n_188)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_166),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_190),
.B(n_194),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_152),
.C(n_146),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_155),
.Y(n_192)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_192),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_193),
.A2(n_180),
.B(n_23),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_153),
.B(n_147),
.Y(n_194)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_195),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_166),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_196),
.B(n_197),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_154),
.B(n_150),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_154),
.B(n_150),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_202),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_153),
.B(n_13),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_206),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_160),
.A2(n_139),
.B1(n_21),
.B2(n_27),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_201),
.A2(n_172),
.B1(n_157),
.B2(n_24),
.Y(n_213)
);

O2A1O1Ixp33_ASAP7_75t_L g202 ( 
.A1(n_168),
.A2(n_27),
.B(n_24),
.C(n_23),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_139),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_163),
.B(n_14),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_204),
.B(n_159),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_166),
.Y(n_206)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_213),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_192),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_199),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_203),
.A2(n_157),
.B(n_164),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_215),
.A2(n_28),
.B(n_14),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_182),
.B(n_155),
.C(n_162),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_218),
.C(n_221),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_219),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_173),
.C(n_179),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_178),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_173),
.C(n_159),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_28),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_223),
.A2(n_202),
.B(n_23),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_187),
.B(n_184),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_28),
.C(n_52),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_183),
.A2(n_175),
.B1(n_180),
.B2(n_21),
.Y(n_226)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_226),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_220),
.A2(n_208),
.B1(n_205),
.B2(n_225),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_229),
.A2(n_236),
.B1(n_240),
.B2(n_241),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_207),
.B(n_211),
.Y(n_230)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

O2A1O1Ixp33_ASAP7_75t_L g232 ( 
.A1(n_210),
.A2(n_189),
.B(n_205),
.C(n_199),
.Y(n_232)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_232),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_234),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_226),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_224),
.A2(n_187),
.B1(n_189),
.B2(n_186),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_242),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_221),
.A2(n_181),
.B1(n_188),
.B2(n_193),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_198),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_237),
.B(n_239),
.Y(n_260)
);

AO21x1_ASAP7_75t_L g255 ( 
.A1(n_238),
.A2(n_243),
.B(n_227),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_210),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_218),
.A2(n_181),
.B1(n_206),
.B2(n_175),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_212),
.A2(n_201),
.B1(n_1),
.B2(n_2),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_36),
.C(n_30),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_242),
.C(n_212),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_219),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_252),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_232),
.A2(n_215),
.B(n_223),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_251),
.A2(n_263),
.B(n_265),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_217),
.C(n_222),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_259),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_258),
.Y(n_267)
);

A2O1A1O1Ixp25_ASAP7_75t_L g256 ( 
.A1(n_235),
.A2(n_213),
.B(n_13),
.C(n_2),
.D(n_3),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_256),
.A2(n_238),
.B(n_2),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_0),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_0),
.Y(n_259)
);

NAND3xp33_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_0),
.C(n_1),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_1),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_264),
.B(n_1),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_229),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_253),
.A2(n_248),
.B1(n_231),
.B2(n_246),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_266),
.B(n_275),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_265),
.A2(n_262),
.B1(n_250),
.B2(n_257),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_5),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_245),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_52),
.C(n_37),
.Y(n_290)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_271),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_247),
.Y(n_272)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_272),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_245),
.Y(n_274)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_36),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_277),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_36),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_243),
.Y(n_278)
);

AOI322xp5_ASAP7_75t_L g286 ( 
.A1(n_278),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_263),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_289),
.Y(n_295)
);

AOI21x1_ASAP7_75t_SL g301 ( 
.A1(n_286),
.A2(n_6),
.B(n_7),
.Y(n_301)
);

OAI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_270),
.A2(n_44),
.B1(n_30),
.B2(n_5),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_287),
.B(n_291),
.Y(n_298)
);

AOI31xp67_ASAP7_75t_L g288 ( 
.A1(n_267),
.A2(n_3),
.A3(n_4),
.B(n_5),
.Y(n_288)
);

AOI31xp67_ASAP7_75t_L g293 ( 
.A1(n_288),
.A2(n_287),
.A3(n_278),
.B(n_280),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_44),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_290),
.B(n_269),
.Y(n_292)
);

AOI21xp33_ASAP7_75t_L g307 ( 
.A1(n_292),
.A2(n_52),
.B(n_47),
.Y(n_307)
);

OAI321xp33_ASAP7_75t_L g302 ( 
.A1(n_293),
.A2(n_296),
.A3(n_301),
.B1(n_6),
.B2(n_10),
.C(n_11),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_284),
.B(n_268),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_294),
.A2(n_300),
.B(n_298),
.Y(n_304)
);

AOI31xp67_ASAP7_75t_L g296 ( 
.A1(n_281),
.A2(n_272),
.A3(n_273),
.B(n_8),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_37),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_299),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_283),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_290),
.A2(n_47),
.B(n_44),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_302),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_305),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_291),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_294),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_306),
.A2(n_307),
.B(n_10),
.Y(n_310)
);

AOI322xp5_ASAP7_75t_L g312 ( 
.A1(n_310),
.A2(n_10),
.A3(n_37),
.B1(n_47),
.B2(n_52),
.C1(n_288),
.C2(n_296),
.Y(n_312)
);

OAI221xp5_ASAP7_75t_L g311 ( 
.A1(n_308),
.A2(n_303),
.B1(n_47),
.B2(n_10),
.C(n_44),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_311),
.B(n_312),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_309),
.Y(n_314)
);


endmodule