module fake_netlist_6_3051_n_2774 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_695, n_507, n_580, n_762, n_209, n_367, n_465, n_680, n_741, n_760, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_726, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_740, n_578, n_703, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_106, n_725, n_358, n_160, n_751, n_449, n_131, n_749, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_396, n_495, n_350, n_78, n_84, n_585, n_732, n_568, n_392, n_442, n_480, n_142, n_724, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_698, n_255, n_739, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_768, n_38, n_471, n_289, n_421, n_781, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_769, n_202, n_320, n_108, n_639, n_676, n_327, n_727, n_369, n_597, n_685, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_718, n_747, n_667, n_71, n_74, n_229, n_542, n_644, n_682, n_621, n_305, n_72, n_721, n_750, n_532, n_742, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_704, n_748, n_506, n_56, n_763, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_710, n_387, n_452, n_616, n_658, n_744, n_39, n_344, n_73, n_581, n_428, n_761, n_746, n_609, n_765, n_432, n_641, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_720, n_525, n_758, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_772, n_96, n_8, n_666, n_371, n_770, n_567, n_189, n_738, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_752, n_112, n_172, n_713, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_782, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_734, n_708, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_779, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_709, n_366, n_777, n_407, n_450, n_103, n_272, n_526, n_185, n_712, n_348, n_711, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_717, n_46, n_330, n_771, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_686, n_252, n_757, n_228, n_565, n_594, n_719, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_745, n_654, n_323, n_606, n_393, n_411, n_503, n_716, n_152, n_623, n_92, n_599, n_513, n_776, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_731, n_406, n_483, n_735, n_102, n_204, n_482, n_755, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_714, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_767, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_345, n_409, n_231, n_354, n_689, n_40, n_505, n_240, n_756, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_635, n_95, n_311, n_10, n_403, n_723, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_764, n_556, n_159, n_157, n_162, n_692, n_733, n_754, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_560, n_753, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_737, n_318, n_303, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_674, n_775, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_759, n_355, n_426, n_317, n_149, n_632, n_702, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_780, n_773, n_675, n_85, n_99, n_257, n_730, n_655, n_13, n_706, n_670, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_690, n_29, n_75, n_401, n_324, n_743, n_766, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_728, n_681, n_729, n_110, n_151, n_774, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_688, n_722, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_637, n_295, n_385, n_701, n_629, n_388, n_190, n_262, n_484, n_613, n_736, n_187, n_501, n_531, n_60, n_361, n_508, n_663, n_379, n_170, n_778, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_2774);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_695;
input n_507;
input n_580;
input n_762;
input n_209;
input n_367;
input n_465;
input n_680;
input n_741;
input n_760;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_726;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_740;
input n_578;
input n_703;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_106;
input n_725;
input n_358;
input n_160;
input n_751;
input n_449;
input n_131;
input n_749;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_732;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_724;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_255;
input n_739;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_768;
input n_38;
input n_471;
input n_289;
input n_421;
input n_781;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_769;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_727;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_718;
input n_747;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_682;
input n_621;
input n_305;
input n_72;
input n_721;
input n_750;
input n_532;
input n_742;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_704;
input n_748;
input n_506;
input n_56;
input n_763;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_387;
input n_452;
input n_616;
input n_658;
input n_744;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_761;
input n_746;
input n_609;
input n_765;
input n_432;
input n_641;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_720;
input n_525;
input n_758;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_772;
input n_96;
input n_8;
input n_666;
input n_371;
input n_770;
input n_567;
input n_189;
input n_738;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_752;
input n_112;
input n_172;
input n_713;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_782;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_734;
input n_708;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_779;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_709;
input n_366;
input n_777;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_712;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_717;
input n_46;
input n_330;
input n_771;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_686;
input n_252;
input n_757;
input n_228;
input n_565;
input n_594;
input n_719;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_745;
input n_654;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_716;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_776;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_731;
input n_406;
input n_483;
input n_735;
input n_102;
input n_204;
input n_482;
input n_755;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_767;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_505;
input n_240;
input n_756;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_635;
input n_95;
input n_311;
input n_10;
input n_403;
input n_723;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_764;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_733;
input n_754;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_560;
input n_753;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_737;
input n_318;
input n_303;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_674;
input n_775;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_759;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_780;
input n_773;
input n_675;
input n_85;
input n_99;
input n_257;
input n_730;
input n_655;
input n_13;
input n_706;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_690;
input n_29;
input n_75;
input n_401;
input n_324;
input n_743;
input n_766;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_728;
input n_681;
input n_729;
input n_110;
input n_151;
input n_774;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_688;
input n_722;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_637;
input n_295;
input n_385;
input n_701;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_736;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_663;
input n_379;
input n_170;
input n_778;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_2774;

wire n_992;
wire n_2542;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_1027;
wire n_1351;
wire n_1189;
wire n_1212;
wire n_2157;
wire n_2332;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_2291;
wire n_830;
wire n_2299;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_2480;
wire n_2739;
wire n_822;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_2729;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_1591;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_940;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_1467;
wire n_976;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2599;
wire n_1978;
wire n_2085;
wire n_917;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_1986;
wire n_2300;
wire n_2397;
wire n_824;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_2735;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_2059;
wire n_2198;
wire n_2669;
wire n_2073;
wire n_2273;
wire n_2546;
wire n_792;
wire n_2522;
wire n_1328;
wire n_1957;
wire n_2616;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_2674;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_2455;
wire n_2654;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_2355;
wire n_966;
wire n_2751;
wire n_2764;
wire n_1663;
wire n_2009;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1722;
wire n_1664;
wire n_2641;
wire n_1165;
wire n_2008;
wire n_2749;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_835;
wire n_1214;
wire n_928;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_2319;
wire n_2519;
wire n_825;
wire n_1063;
wire n_1588;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_2476;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_2733;
wire n_890;
wire n_2377;
wire n_2178;
wire n_950;
wire n_2644;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_949;
wire n_1630;
wire n_2075;
wire n_2194;
wire n_2619;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2728;
wire n_2349;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_2436;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_794;
wire n_2767;
wire n_894;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_2707;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_851;
wire n_2537;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_2517;
wire n_2713;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_2643;
wire n_2590;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_797;
wire n_2689;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2675;
wire n_1426;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_1049;
wire n_2771;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_919;
wire n_1698;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_1299;
wire n_2718;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_998;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_1475;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_2682;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_931;
wire n_1021;
wire n_811;
wire n_1207;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_1250;
wire n_958;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_889;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_1314;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_1877;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2596;
wire n_2274;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_914;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_1243;
wire n_848;
wire n_2732;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_2159;
wire n_906;
wire n_1390;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2289;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_2627;
wire n_956;
wire n_960;
wire n_2276;
wire n_856;
wire n_2100;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_793;
wire n_1593;
wire n_1202;
wire n_1030;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_999;
wire n_1254;
wire n_2420;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_974;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_1871;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_2302;
wire n_1667;
wire n_1206;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_901;
wire n_1499;
wire n_2755;
wire n_923;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_991;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_785;
wire n_2740;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2401;
wire n_2337;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2716;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2037;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2244;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_962;
wire n_1041;
wire n_2346;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2541;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_1823;
wire n_2479;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_2406;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_2567;
wire n_2322;
wire n_2154;
wire n_2727;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2759;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2668;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_2695;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1949;
wire n_2671;
wire n_2761;
wire n_2715;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_2054;
wire n_876;
wire n_1337;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_853;
wire n_1542;
wire n_2587;
wire n_875;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_1953;
wire n_933;
wire n_978;
wire n_2752;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2186;
wire n_2163;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_1379;
wire n_2528;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_2380;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_814;
wire n_2746;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_1461;
wire n_2076;
wire n_2736;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_2182;
wire n_1283;
wire n_2385;
wire n_918;
wire n_1114;
wire n_1848;
wire n_1147;
wire n_1785;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_971;
wire n_2702;
wire n_946;
wire n_1303;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_2685;
wire n_1083;
wire n_1561;
wire n_2741;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_839;
wire n_2437;
wire n_2743;
wire n_1973;
wire n_2267;
wire n_990;
wire n_1500;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_1584;
wire n_2425;
wire n_924;
wire n_1582;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_1972;
wire n_2592;
wire n_1525;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_2600;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_2033;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_981;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_980;
wire n_2681;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_1996;
wire n_2367;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_849;
wire n_2662;
wire n_1753;
wire n_2471;
wire n_2540;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_1170;
wire n_1629;
wire n_2221;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_2632;
wire n_2579;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_2659;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_1742;
wire n_1612;
wire n_1240;

CKINVDCx16_ASAP7_75t_R g783 ( 
.A(n_96),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_694),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_10),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_261),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_744),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_157),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_382),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_278),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_686),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_152),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_772),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_219),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_242),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_732),
.Y(n_796)
);

CKINVDCx16_ASAP7_75t_R g797 ( 
.A(n_607),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_761),
.Y(n_798)
);

CKINVDCx16_ASAP7_75t_R g799 ( 
.A(n_108),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_531),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_603),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_775),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_737),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_98),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_722),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_681),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_767),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_723),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_779),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_312),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_682),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_170),
.Y(n_812)
);

INVx1_ASAP7_75t_SL g813 ( 
.A(n_236),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_626),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_740),
.Y(n_815)
);

INVxp67_ASAP7_75t_SL g816 ( 
.A(n_660),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_753),
.Y(n_817)
);

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_773),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_746),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_76),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_325),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_571),
.Y(n_822)
);

CKINVDCx20_ASAP7_75t_R g823 ( 
.A(n_762),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_177),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_233),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_217),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_516),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_341),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_66),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_717),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_194),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_120),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_679),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_165),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_194),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_215),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_349),
.Y(n_837)
);

BUFx5_ASAP7_75t_L g838 ( 
.A(n_223),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_755),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_691),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_776),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_754),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_235),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_616),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_536),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_781),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_592),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_483),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_648),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_575),
.Y(n_850)
);

CKINVDCx20_ASAP7_75t_R g851 ( 
.A(n_769),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_680),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_18),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_170),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_711),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_638),
.Y(n_856)
);

INVxp67_ASAP7_75t_L g857 ( 
.A(n_238),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_714),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_710),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_765),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_633),
.Y(n_861)
);

BUFx10_ASAP7_75t_L g862 ( 
.A(n_436),
.Y(n_862)
);

BUFx2_ASAP7_75t_L g863 ( 
.A(n_739),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_742),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_698),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_677),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_573),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_703),
.Y(n_868)
);

CKINVDCx20_ASAP7_75t_R g869 ( 
.A(n_630),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_554),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_696),
.Y(n_871)
);

BUFx2_ASAP7_75t_L g872 ( 
.A(n_759),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_128),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_764),
.Y(n_874)
);

CKINVDCx20_ASAP7_75t_R g875 ( 
.A(n_624),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_414),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_225),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_209),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_184),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_726),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_756),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_297),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_363),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_615),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_191),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_443),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_692),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_768),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_505),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_727),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_628),
.Y(n_891)
);

INVxp33_ASAP7_75t_SL g892 ( 
.A(n_211),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_777),
.Y(n_893)
);

INVx1_ASAP7_75t_SL g894 ( 
.A(n_550),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_704),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_760),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_650),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_405),
.Y(n_898)
);

BUFx8_ASAP7_75t_SL g899 ( 
.A(n_253),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_595),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_152),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_664),
.Y(n_902)
);

CKINVDCx20_ASAP7_75t_R g903 ( 
.A(n_411),
.Y(n_903)
);

INVx1_ASAP7_75t_SL g904 ( 
.A(n_226),
.Y(n_904)
);

BUFx3_ASAP7_75t_L g905 ( 
.A(n_725),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_119),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_663),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_715),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_331),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_454),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_689),
.Y(n_911)
);

INVxp67_ASAP7_75t_L g912 ( 
.A(n_750),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_645),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_588),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_644),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_233),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_523),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_629),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_219),
.Y(n_919)
);

BUFx10_ASAP7_75t_L g920 ( 
.A(n_319),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_465),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_265),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_341),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_74),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_204),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_266),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_225),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_613),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_358),
.Y(n_929)
);

CKINVDCx20_ASAP7_75t_R g930 ( 
.A(n_683),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_366),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_567),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_731),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_138),
.Y(n_934)
);

CKINVDCx20_ASAP7_75t_R g935 ( 
.A(n_8),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_372),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_585),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_749),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_215),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_413),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_335),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_209),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_469),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_459),
.Y(n_944)
);

BUFx10_ASAP7_75t_L g945 ( 
.A(n_734),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_178),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_47),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_702),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_500),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_296),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_738),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_63),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_504),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_701),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_13),
.Y(n_955)
);

INVxp33_ASAP7_75t_R g956 ( 
.A(n_11),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_113),
.Y(n_957)
);

BUFx10_ASAP7_75t_L g958 ( 
.A(n_586),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_88),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_770),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_319),
.Y(n_961)
);

BUFx10_ASAP7_75t_L g962 ( 
.A(n_687),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_61),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_434),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_707),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_133),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_411),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_685),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_688),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_266),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_20),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_673),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_13),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_721),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_539),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_455),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_162),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_733),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_45),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_0),
.Y(n_980)
);

INVx1_ASAP7_75t_SL g981 ( 
.A(n_110),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_184),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_461),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_541),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_61),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_712),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_259),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_709),
.Y(n_988)
);

CKINVDCx20_ASAP7_75t_R g989 ( 
.A(n_574),
.Y(n_989)
);

INVx1_ASAP7_75t_SL g990 ( 
.A(n_171),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_427),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_92),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_741),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_189),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_328),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_26),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_771),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_166),
.Y(n_998)
);

INVx2_ASAP7_75t_SL g999 ( 
.A(n_327),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_126),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_2),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_52),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_598),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_463),
.Y(n_1004)
);

CKINVDCx20_ASAP7_75t_R g1005 ( 
.A(n_315),
.Y(n_1005)
);

INVx1_ASAP7_75t_SL g1006 ( 
.A(n_706),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_255),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_298),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_757),
.Y(n_1009)
);

CKINVDCx20_ASAP7_75t_R g1010 ( 
.A(n_577),
.Y(n_1010)
);

INVx2_ASAP7_75t_SL g1011 ( 
.A(n_395),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_172),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_210),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_275),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_29),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_513),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_724),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_587),
.Y(n_1018)
);

HB1xp67_ASAP7_75t_L g1019 ( 
.A(n_474),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_41),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_404),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_525),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_204),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_735),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_409),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_736),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_240),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_684),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_261),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_700),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_220),
.Y(n_1031)
);

CKINVDCx20_ASAP7_75t_R g1032 ( 
.A(n_758),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_748),
.Y(n_1033)
);

CKINVDCx20_ASAP7_75t_R g1034 ( 
.A(n_752),
.Y(n_1034)
);

INVx2_ASAP7_75t_SL g1035 ( 
.A(n_695),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_665),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_676),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_672),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_443),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_426),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_445),
.Y(n_1041)
);

CKINVDCx20_ASAP7_75t_R g1042 ( 
.A(n_678),
.Y(n_1042)
);

CKINVDCx20_ASAP7_75t_R g1043 ( 
.A(n_417),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_287),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_543),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_747),
.Y(n_1046)
);

INVx1_ASAP7_75t_SL g1047 ( 
.A(n_331),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_471),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_68),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_766),
.Y(n_1050)
);

BUFx2_ASAP7_75t_L g1051 ( 
.A(n_697),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_778),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_36),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_719),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_306),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_50),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_275),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_318),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_169),
.Y(n_1059)
);

CKINVDCx16_ASAP7_75t_R g1060 ( 
.A(n_561),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_67),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_634),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_425),
.Y(n_1063)
);

BUFx3_ASAP7_75t_L g1064 ( 
.A(n_493),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_197),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_693),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_566),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_41),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_332),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_713),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_730),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_708),
.Y(n_1072)
);

CKINVDCx16_ASAP7_75t_R g1073 ( 
.A(n_718),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_279),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_187),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_432),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_431),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_774),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_720),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_67),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_618),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_314),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_468),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_751),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_690),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_729),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_705),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_407),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_303),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_297),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_699),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_362),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_530),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_728),
.Y(n_1094)
);

BUFx10_ASAP7_75t_L g1095 ( 
.A(n_763),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_399),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_557),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_324),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_213),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_393),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_416),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_380),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_716),
.Y(n_1103)
);

INVxp33_ASAP7_75t_L g1104 ( 
.A(n_432),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_780),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_59),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_526),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_743),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_745),
.Y(n_1109)
);

INVxp67_ASAP7_75t_SL g1110 ( 
.A(n_802),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_783),
.Y(n_1111)
);

CKINVDCx20_ASAP7_75t_R g1112 ( 
.A(n_809),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_899),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_863),
.B(n_1),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_838),
.Y(n_1115)
);

INVxp67_ASAP7_75t_SL g1116 ( 
.A(n_1019),
.Y(n_1116)
);

CKINVDCx20_ASAP7_75t_R g1117 ( 
.A(n_818),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_838),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_787),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_923),
.B(n_0),
.Y(n_1120)
);

NOR2xp67_ASAP7_75t_L g1121 ( 
.A(n_849),
.B(n_1),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_838),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_838),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_791),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_800),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_801),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_806),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_872),
.B(n_3),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_838),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_1051),
.B(n_3),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_811),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_792),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_792),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_823),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_792),
.Y(n_1135)
);

INVxp67_ASAP7_75t_SL g1136 ( 
.A(n_849),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_898),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_814),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_898),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_898),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_815),
.Y(n_1141)
);

CKINVDCx16_ASAP7_75t_R g1142 ( 
.A(n_799),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_916),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_916),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_916),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_817),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1044),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_827),
.Y(n_1148)
);

INVxp67_ASAP7_75t_L g1149 ( 
.A(n_999),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1044),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1044),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_830),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_877),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_841),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_980),
.Y(n_1155)
);

INVxp67_ASAP7_75t_L g1156 ( 
.A(n_1011),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1049),
.Y(n_1157)
);

CKINVDCx20_ASAP7_75t_R g1158 ( 
.A(n_851),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_844),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1082),
.Y(n_1160)
);

OR2x2_ASAP7_75t_L g1161 ( 
.A(n_794),
.B(n_2),
.Y(n_1161)
);

NAND2xp33_ASAP7_75t_L g1162 ( 
.A(n_1120),
.B(n_1106),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1132),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1133),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1135),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_1111),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_1136),
.B(n_793),
.Y(n_1167)
);

BUFx3_ASAP7_75t_L g1168 ( 
.A(n_1153),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1137),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1139),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1140),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1143),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1119),
.B(n_805),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_1144),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1145),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_1147),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1110),
.B(n_797),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1124),
.B(n_1060),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1150),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_1116),
.B(n_848),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1151),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1129),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1125),
.B(n_1126),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_1127),
.Y(n_1184)
);

CKINVDCx8_ASAP7_75t_R g1185 ( 
.A(n_1142),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1131),
.B(n_1073),
.Y(n_1186)
);

INVx3_ASAP7_75t_L g1187 ( 
.A(n_1155),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1115),
.A2(n_819),
.B(n_808),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_1114),
.B(n_1095),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1118),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1173),
.B(n_1138),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1190),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_1186),
.B(n_1141),
.Y(n_1193)
);

NAND3xp33_ASAP7_75t_L g1194 ( 
.A(n_1178),
.B(n_1130),
.C(n_1128),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_1168),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1182),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1167),
.B(n_1146),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1176),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1163),
.Y(n_1199)
);

AND2x6_ASAP7_75t_L g1200 ( 
.A(n_1177),
.B(n_864),
.Y(n_1200)
);

INVxp33_ASAP7_75t_L g1201 ( 
.A(n_1166),
.Y(n_1201)
);

INVx2_ASAP7_75t_SL g1202 ( 
.A(n_1180),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1184),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_1183),
.B(n_1148),
.Y(n_1204)
);

INVx2_ASAP7_75t_SL g1205 ( 
.A(n_1180),
.Y(n_1205)
);

INVx2_ASAP7_75t_SL g1206 ( 
.A(n_1166),
.Y(n_1206)
);

INVx2_ASAP7_75t_SL g1207 ( 
.A(n_1167),
.Y(n_1207)
);

NAND2xp33_ASAP7_75t_L g1208 ( 
.A(n_1189),
.B(n_1152),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1162),
.B(n_1154),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_1184),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_1176),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1170),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1187),
.B(n_1159),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1176),
.B(n_1113),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1185),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1171),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_1174),
.Y(n_1217)
);

NOR2x1p5_ASAP7_75t_L g1218 ( 
.A(n_1175),
.B(n_1161),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1164),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_1181),
.B(n_1121),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1188),
.A2(n_1123),
.B1(n_1122),
.B2(n_786),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1165),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_1169),
.B(n_945),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1172),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1179),
.B(n_913),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1182),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1190),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_1166),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1182),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_1186),
.B(n_945),
.Y(n_1230)
);

INVx1_ASAP7_75t_SL g1231 ( 
.A(n_1166),
.Y(n_1231)
);

BUFx10_ASAP7_75t_L g1232 ( 
.A(n_1178),
.Y(n_1232)
);

BUFx10_ASAP7_75t_L g1233 ( 
.A(n_1178),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1167),
.B(n_1035),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1190),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1190),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_1218),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1199),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1194),
.A2(n_892),
.B1(n_860),
.B2(n_887),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1226),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_1202),
.B(n_869),
.Y(n_1241)
);

BUFx5_ASAP7_75t_L g1242 ( 
.A(n_1236),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1229),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_1215),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1204),
.B(n_816),
.Y(n_1245)
);

AO221x1_ASAP7_75t_L g1246 ( 
.A1(n_1217),
.A2(n_857),
.B1(n_912),
.B2(n_884),
.C(n_864),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_SL g1247 ( 
.A(n_1205),
.B(n_875),
.Y(n_1247)
);

NAND2xp33_ASAP7_75t_SL g1248 ( 
.A(n_1230),
.B(n_1112),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1231),
.B(n_1117),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_1207),
.B(n_930),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1212),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1191),
.A2(n_989),
.B1(n_1032),
.B2(n_1010),
.Y(n_1252)
);

A2O1A1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1234),
.A2(n_796),
.B(n_798),
.C(n_784),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_1213),
.B(n_1197),
.Y(n_1254)
);

INVxp67_ASAP7_75t_L g1255 ( 
.A(n_1228),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1192),
.B(n_803),
.Y(n_1256)
);

NOR2xp67_ASAP7_75t_L g1257 ( 
.A(n_1206),
.B(n_1149),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_1209),
.B(n_1034),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1216),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1227),
.B(n_807),
.Y(n_1260)
);

CKINVDCx20_ASAP7_75t_R g1261 ( 
.A(n_1203),
.Y(n_1261)
);

A2O1A1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1235),
.A2(n_822),
.B(n_839),
.C(n_833),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1200),
.B(n_840),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1200),
.A2(n_943),
.B1(n_948),
.B2(n_845),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1200),
.B(n_842),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1200),
.B(n_847),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1196),
.B(n_850),
.Y(n_1267)
);

INVx3_ASAP7_75t_L g1268 ( 
.A(n_1195),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1232),
.B(n_1042),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_SL g1270 ( 
.A(n_1232),
.B(n_1072),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1198),
.B(n_852),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1222),
.B(n_861),
.Y(n_1272)
);

AOI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1208),
.A2(n_1193),
.B1(n_1220),
.B2(n_1158),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1211),
.B(n_867),
.Y(n_1274)
);

INVx3_ASAP7_75t_L g1275 ( 
.A(n_1219),
.Y(n_1275)
);

O2A1O1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1225),
.A2(n_824),
.B(n_828),
.C(n_826),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1224),
.Y(n_1277)
);

INVxp67_ASAP7_75t_L g1278 ( 
.A(n_1210),
.Y(n_1278)
);

HB1xp67_ASAP7_75t_L g1279 ( 
.A(n_1201),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1223),
.Y(n_1280)
);

INVx3_ASAP7_75t_L g1281 ( 
.A(n_1233),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1221),
.B(n_891),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1214),
.B(n_893),
.Y(n_1283)
);

NAND2xp33_ASAP7_75t_L g1284 ( 
.A(n_1233),
.B(n_846),
.Y(n_1284)
);

INVxp67_ASAP7_75t_SL g1285 ( 
.A(n_1211),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1199),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1204),
.B(n_900),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1231),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1204),
.B(n_914),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1204),
.B(n_917),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1204),
.B(n_921),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1199),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1191),
.B(n_1134),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1204),
.B(n_938),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1204),
.B(n_965),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1195),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1191),
.B(n_1104),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_1202),
.B(n_894),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1204),
.B(n_975),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1231),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1226),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1202),
.B(n_1006),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_1195),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1204),
.B(n_983),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1226),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1226),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_SL g1307 ( 
.A(n_1202),
.B(n_1105),
.Y(n_1307)
);

BUFx5_ASAP7_75t_L g1308 ( 
.A(n_1192),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1199),
.Y(n_1309)
);

INVx2_ASAP7_75t_SL g1310 ( 
.A(n_1218),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1204),
.B(n_984),
.Y(n_1311)
);

INVx4_ASAP7_75t_L g1312 ( 
.A(n_1215),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1202),
.B(n_1109),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_L g1314 ( 
.A(n_1191),
.B(n_956),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1204),
.B(n_997),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1199),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1204),
.B(n_1003),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1199),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1204),
.B(n_1022),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1191),
.B(n_813),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1204),
.B(n_1026),
.Y(n_1321)
);

O2A1O1Ixp5_ASAP7_75t_L g1322 ( 
.A1(n_1234),
.A2(n_1016),
.B(n_1045),
.C(n_953),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1199),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1191),
.B(n_904),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_SL g1325 ( 
.A(n_1202),
.B(n_1097),
.Y(n_1325)
);

NOR2x1p5_ASAP7_75t_L g1326 ( 
.A(n_1215),
.B(n_1157),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_SL g1327 ( 
.A(n_1202),
.B(n_855),
.Y(n_1327)
);

NAND2xp33_ASAP7_75t_L g1328 ( 
.A(n_1200),
.B(n_856),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1226),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1204),
.B(n_1033),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1204),
.B(n_1048),
.Y(n_1331)
);

INVxp67_ASAP7_75t_L g1332 ( 
.A(n_1228),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_SL g1333 ( 
.A(n_1202),
.B(n_858),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1204),
.B(n_1054),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1204),
.B(n_1066),
.Y(n_1335)
);

OR2x2_ASAP7_75t_L g1336 ( 
.A(n_1231),
.B(n_1160),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1199),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1202),
.B(n_859),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_SL g1339 ( 
.A(n_1202),
.B(n_865),
.Y(n_1339)
);

AOI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1282),
.A2(n_1085),
.B(n_1084),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1320),
.B(n_1086),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1238),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1324),
.B(n_1149),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1297),
.B(n_1093),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1251),
.Y(n_1345)
);

AOI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1245),
.A2(n_1108),
.B1(n_1103),
.B2(n_868),
.Y(n_1346)
);

BUFx8_ASAP7_75t_L g1347 ( 
.A(n_1249),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1287),
.B(n_866),
.Y(n_1348)
);

AOI22x1_ASAP7_75t_L g1349 ( 
.A1(n_1259),
.A2(n_870),
.B1(n_874),
.B2(n_871),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1289),
.B(n_880),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1288),
.B(n_1156),
.Y(n_1351)
);

OAI321xp33_ASAP7_75t_L g1352 ( 
.A1(n_1239),
.A2(n_1290),
.A3(n_1291),
.B1(n_1299),
.B2(n_1295),
.C(n_1294),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1304),
.B(n_881),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1254),
.A2(n_884),
.B(n_864),
.Y(n_1354)
);

A2O1A1Ixp33_ASAP7_75t_L g1355 ( 
.A1(n_1311),
.A2(n_1030),
.B(n_1064),
.C(n_905),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1315),
.B(n_888),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1317),
.A2(n_1083),
.B(n_884),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1319),
.A2(n_1083),
.B(n_890),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1286),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1240),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1292),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1321),
.B(n_889),
.Y(n_1362)
);

AOI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1271),
.A2(n_835),
.B(n_829),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1330),
.B(n_895),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1331),
.B(n_896),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1334),
.B(n_897),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1335),
.A2(n_1083),
.B(n_907),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1309),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1316),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1243),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1252),
.B(n_902),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1318),
.A2(n_910),
.B(n_908),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1242),
.B(n_911),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1323),
.A2(n_918),
.B(n_915),
.Y(n_1374)
);

A2O1A1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1314),
.A2(n_1107),
.B(n_1070),
.C(n_990),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1301),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1242),
.B(n_1308),
.Y(n_1377)
);

OAI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1322),
.A2(n_932),
.B(n_928),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1242),
.B(n_933),
.Y(n_1379)
);

CKINVDCx11_ASAP7_75t_R g1380 ( 
.A(n_1261),
.Y(n_1380)
);

INVxp67_ASAP7_75t_L g1381 ( 
.A(n_1300),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1337),
.A2(n_944),
.B(n_937),
.Y(n_1382)
);

NOR3xp33_ASAP7_75t_L g1383 ( 
.A(n_1269),
.B(n_1047),
.C(n_981),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_L g1384 ( 
.A(n_1293),
.B(n_832),
.Y(n_1384)
);

OAI21xp33_ASAP7_75t_L g1385 ( 
.A1(n_1336),
.A2(n_1156),
.B(n_788),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1242),
.B(n_949),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1308),
.B(n_951),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_SL g1388 ( 
.A(n_1308),
.B(n_954),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1296),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1285),
.A2(n_968),
.B(n_960),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1258),
.A2(n_972),
.B(n_969),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1308),
.B(n_974),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1283),
.A2(n_978),
.B(n_976),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1307),
.A2(n_988),
.B(n_986),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1305),
.B(n_1306),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1329),
.B(n_993),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1279),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1273),
.A2(n_935),
.B1(n_1005),
.B2(n_903),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1257),
.B(n_862),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1255),
.B(n_1015),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1256),
.B(n_1004),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1313),
.A2(n_1327),
.B(n_1325),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1260),
.A2(n_1017),
.B(n_1009),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1333),
.A2(n_1024),
.B(n_1018),
.Y(n_1404)
);

BUFx3_ASAP7_75t_L g1405 ( 
.A(n_1303),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1277),
.B(n_1028),
.Y(n_1406)
);

AND2x4_ASAP7_75t_L g1407 ( 
.A(n_1268),
.B(n_836),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1272),
.B(n_1036),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1332),
.B(n_1278),
.Y(n_1409)
);

A2O1A1Ixp33_ASAP7_75t_L g1410 ( 
.A1(n_1280),
.A2(n_843),
.B(n_873),
.C(n_854),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_SL g1411 ( 
.A(n_1281),
.B(n_1037),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1275),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1267),
.B(n_1038),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_SL g1414 ( 
.A(n_1312),
.B(n_1041),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1274),
.B(n_1298),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1302),
.B(n_1046),
.Y(n_1416)
);

A2O1A1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1248),
.A2(n_879),
.B(n_931),
.C(n_924),
.Y(n_1417)
);

OAI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1338),
.A2(n_1052),
.B(n_1050),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_L g1419 ( 
.A(n_1241),
.B(n_1043),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1339),
.A2(n_1067),
.B(n_1062),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1263),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1246),
.B(n_1071),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1237),
.A2(n_1310),
.B1(n_1247),
.B2(n_1250),
.Y(n_1423)
);

NOR3xp33_ASAP7_75t_L g1424 ( 
.A(n_1270),
.B(n_789),
.C(n_785),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1265),
.B(n_1078),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1266),
.A2(n_1081),
.B(n_1079),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1253),
.B(n_1087),
.Y(n_1427)
);

INVx3_ASAP7_75t_L g1428 ( 
.A(n_1244),
.Y(n_1428)
);

OAI21xp33_ASAP7_75t_L g1429 ( 
.A1(n_1284),
.A2(n_795),
.B(n_790),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1264),
.B(n_1262),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_1326),
.B(n_934),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1328),
.B(n_862),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_L g1433 ( 
.A(n_1276),
.B(n_810),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1320),
.B(n_1091),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1245),
.A2(n_1094),
.B(n_940),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1320),
.B(n_812),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1320),
.B(n_820),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1245),
.A2(n_947),
.B(n_936),
.Y(n_1438)
);

BUFx12f_ASAP7_75t_L g1439 ( 
.A(n_1244),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1320),
.B(n_821),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1240),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1245),
.A2(n_959),
.B(n_950),
.Y(n_1442)
);

A2O1A1Ixp33_ASAP7_75t_L g1443 ( 
.A1(n_1320),
.A2(n_970),
.B(n_971),
.C(n_966),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_SL g1444 ( 
.A(n_1320),
.B(n_958),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1288),
.Y(n_1445)
);

AOI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1320),
.A2(n_962),
.B1(n_1095),
.B2(n_958),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1320),
.B(n_825),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1245),
.A2(n_1002),
.B(n_1001),
.Y(n_1448)
);

NOR2xp67_ASAP7_75t_L g1449 ( 
.A(n_1312),
.B(n_444),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1240),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1240),
.Y(n_1451)
);

AOI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1282),
.A2(n_1056),
.B(n_1027),
.Y(n_1452)
);

INVx2_ASAP7_75t_SL g1453 ( 
.A(n_1288),
.Y(n_1453)
);

AOI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1282),
.A2(n_1068),
.B(n_1059),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_SL g1455 ( 
.A(n_1320),
.B(n_962),
.Y(n_1455)
);

NOR2xp33_ASAP7_75t_L g1456 ( 
.A(n_1320),
.B(n_831),
.Y(n_1456)
);

AOI21xp33_ASAP7_75t_L g1457 ( 
.A1(n_1320),
.A2(n_837),
.B(n_834),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1238),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1245),
.A2(n_1076),
.B(n_1075),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1320),
.B(n_853),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_1320),
.B(n_876),
.Y(n_1461)
);

AOI21xp33_ASAP7_75t_L g1462 ( 
.A1(n_1320),
.A2(n_882),
.B(n_878),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1245),
.A2(n_883),
.B1(n_886),
.B2(n_885),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_L g1464 ( 
.A(n_1320),
.B(n_901),
.Y(n_1464)
);

OAI21xp33_ASAP7_75t_SL g1465 ( 
.A1(n_1287),
.A2(n_1101),
.B(n_1089),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1245),
.A2(n_1102),
.B(n_922),
.Y(n_1466)
);

INVx2_ASAP7_75t_SL g1467 ( 
.A(n_1288),
.Y(n_1467)
);

A2O1A1Ixp33_ASAP7_75t_L g1468 ( 
.A1(n_1320),
.A2(n_967),
.B(n_979),
.C(n_804),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1320),
.B(n_906),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1320),
.B(n_909),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1245),
.A2(n_1020),
.B(n_1014),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1288),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1320),
.B(n_919),
.Y(n_1473)
);

OAI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1282),
.A2(n_1065),
.B(n_1063),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_1320),
.B(n_925),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1240),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1240),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1282),
.A2(n_1074),
.B(n_1069),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1245),
.A2(n_927),
.B(n_926),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1320),
.B(n_929),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1238),
.Y(n_1481)
);

AOI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1282),
.A2(n_447),
.B(n_446),
.Y(n_1482)
);

O2A1O1Ixp33_ASAP7_75t_L g1483 ( 
.A1(n_1320),
.A2(n_939),
.B(n_942),
.C(n_941),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1320),
.B(n_946),
.Y(n_1484)
);

O2A1O1Ixp33_ASAP7_75t_L g1485 ( 
.A1(n_1320),
.A2(n_952),
.B(n_957),
.C(n_955),
.Y(n_1485)
);

AOI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1245),
.A2(n_963),
.B(n_961),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1320),
.B(n_964),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1288),
.Y(n_1488)
);

OAI21xp33_ASAP7_75t_L g1489 ( 
.A1(n_1320),
.A2(n_977),
.B(n_973),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_SL g1490 ( 
.A(n_1320),
.B(n_982),
.Y(n_1490)
);

AOI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1245),
.A2(n_987),
.B(n_985),
.Y(n_1491)
);

AOI21xp33_ASAP7_75t_L g1492 ( 
.A1(n_1456),
.A2(n_992),
.B(n_991),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1464),
.B(n_994),
.Y(n_1493)
);

BUFx12f_ASAP7_75t_L g1494 ( 
.A(n_1380),
.Y(n_1494)
);

AOI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1473),
.A2(n_995),
.B1(n_998),
.B2(n_996),
.Y(n_1495)
);

O2A1O1Ixp33_ASAP7_75t_L g1496 ( 
.A1(n_1341),
.A2(n_920),
.B(n_1007),
.C(n_1000),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1342),
.Y(n_1497)
);

INVx1_ASAP7_75t_SL g1498 ( 
.A(n_1472),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1345),
.Y(n_1499)
);

BUFx6f_ASAP7_75t_L g1500 ( 
.A(n_1389),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1377),
.A2(n_1012),
.B1(n_1013),
.B2(n_1008),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1343),
.B(n_920),
.Y(n_1502)
);

AO32x2_ASAP7_75t_L g1503 ( 
.A1(n_1423),
.A2(n_6),
.A3(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1384),
.B(n_1487),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1344),
.B(n_1021),
.Y(n_1505)
);

A2O1A1Ixp33_ASAP7_75t_L g1506 ( 
.A1(n_1352),
.A2(n_1025),
.B(n_1029),
.C(n_1023),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1399),
.B(n_1031),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_SL g1508 ( 
.A(n_1453),
.B(n_1467),
.Y(n_1508)
);

NOR2x1_ASAP7_75t_R g1509 ( 
.A(n_1439),
.B(n_1039),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1360),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1436),
.B(n_1437),
.Y(n_1511)
);

O2A1O1Ixp33_ASAP7_75t_SL g1512 ( 
.A1(n_1375),
.A2(n_449),
.B(n_450),
.C(n_448),
.Y(n_1512)
);

AOI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1388),
.A2(n_452),
.B(n_451),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1370),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1359),
.Y(n_1515)
);

INVx1_ASAP7_75t_SL g1516 ( 
.A(n_1488),
.Y(n_1516)
);

AOI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1373),
.A2(n_456),
.B(n_453),
.Y(n_1517)
);

AOI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1379),
.A2(n_458),
.B(n_457),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_R g1519 ( 
.A(n_1428),
.B(n_1389),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1440),
.B(n_1040),
.Y(n_1520)
);

NOR3xp33_ASAP7_75t_SL g1521 ( 
.A(n_1398),
.B(n_1055),
.C(n_1053),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_R g1522 ( 
.A(n_1428),
.B(n_1057),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1376),
.Y(n_1523)
);

CKINVDCx8_ASAP7_75t_R g1524 ( 
.A(n_1389),
.Y(n_1524)
);

AOI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1386),
.A2(n_462),
.B(n_460),
.Y(n_1525)
);

NAND2xp33_ASAP7_75t_SL g1526 ( 
.A(n_1432),
.B(n_1058),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1434),
.A2(n_1077),
.B1(n_1080),
.B2(n_1061),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1361),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1447),
.B(n_1088),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_SL g1530 ( 
.A(n_1381),
.B(n_1090),
.Y(n_1530)
);

INVxp67_ASAP7_75t_SL g1531 ( 
.A(n_1445),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_SL g1532 ( 
.A(n_1460),
.B(n_1092),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1368),
.Y(n_1533)
);

AND2x2_ASAP7_75t_SL g1534 ( 
.A(n_1419),
.B(n_4),
.Y(n_1534)
);

NAND2xp33_ASAP7_75t_SL g1535 ( 
.A(n_1371),
.B(n_1096),
.Y(n_1535)
);

BUFx6f_ASAP7_75t_L g1536 ( 
.A(n_1405),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1441),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1397),
.B(n_464),
.Y(n_1538)
);

AOI21xp5_ASAP7_75t_L g1539 ( 
.A1(n_1387),
.A2(n_467),
.B(n_466),
.Y(n_1539)
);

AND2x2_ASAP7_75t_SL g1540 ( 
.A(n_1383),
.B(n_5),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1469),
.B(n_1098),
.Y(n_1541)
);

O2A1O1Ixp33_ASAP7_75t_L g1542 ( 
.A1(n_1470),
.A2(n_1100),
.B(n_1099),
.C(n_8),
.Y(n_1542)
);

NOR3xp33_ASAP7_75t_L g1543 ( 
.A(n_1457),
.B(n_6),
.C(n_7),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1450),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1347),
.Y(n_1545)
);

AOI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1392),
.A2(n_472),
.B(n_470),
.Y(n_1546)
);

AOI21xp33_ASAP7_75t_L g1547 ( 
.A1(n_1480),
.A2(n_9),
.B(n_10),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1347),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1484),
.B(n_9),
.Y(n_1549)
);

BUFx6f_ASAP7_75t_L g1550 ( 
.A(n_1407),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1451),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1476),
.Y(n_1552)
);

NOR3xp33_ASAP7_75t_L g1553 ( 
.A(n_1462),
.B(n_11),
.C(n_12),
.Y(n_1553)
);

OR2x6_ASAP7_75t_L g1554 ( 
.A(n_1351),
.B(n_1402),
.Y(n_1554)
);

OAI21x1_ASAP7_75t_L g1555 ( 
.A1(n_1482),
.A2(n_475),
.B(n_473),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1369),
.B(n_12),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_1407),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1400),
.B(n_14),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1458),
.B(n_14),
.Y(n_1559)
);

BUFx12f_ASAP7_75t_L g1560 ( 
.A(n_1431),
.Y(n_1560)
);

AOI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1421),
.A2(n_477),
.B(n_476),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1481),
.Y(n_1562)
);

INVx4_ASAP7_75t_L g1563 ( 
.A(n_1431),
.Y(n_1563)
);

O2A1O1Ixp33_ASAP7_75t_L g1564 ( 
.A1(n_1444),
.A2(n_17),
.B(n_15),
.C(n_16),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_SL g1565 ( 
.A(n_1415),
.B(n_478),
.Y(n_1565)
);

AOI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1395),
.A2(n_480),
.B(n_479),
.Y(n_1566)
);

A2O1A1Ixp33_ASAP7_75t_L g1567 ( 
.A1(n_1474),
.A2(n_17),
.B(n_15),
.C(n_16),
.Y(n_1567)
);

INVxp67_ASAP7_75t_L g1568 ( 
.A(n_1409),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1348),
.B(n_18),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_SL g1570 ( 
.A(n_1483),
.B(n_481),
.Y(n_1570)
);

INVx4_ASAP7_75t_L g1571 ( 
.A(n_1412),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1461),
.B(n_19),
.Y(n_1572)
);

AOI21xp5_ASAP7_75t_L g1573 ( 
.A1(n_1350),
.A2(n_1356),
.B(n_1353),
.Y(n_1573)
);

BUFx2_ASAP7_75t_L g1574 ( 
.A(n_1465),
.Y(n_1574)
);

AOI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1362),
.A2(n_484),
.B(n_482),
.Y(n_1575)
);

AO32x1_ASAP7_75t_L g1576 ( 
.A1(n_1463),
.A2(n_21),
.A3(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1477),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1364),
.B(n_21),
.Y(n_1578)
);

AOI21xp5_ASAP7_75t_L g1579 ( 
.A1(n_1365),
.A2(n_486),
.B(n_485),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_SL g1580 ( 
.A(n_1485),
.B(n_487),
.Y(n_1580)
);

NOR2xp33_ASAP7_75t_L g1581 ( 
.A(n_1475),
.B(n_22),
.Y(n_1581)
);

AOI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1366),
.A2(n_489),
.B(n_488),
.Y(n_1582)
);

AOI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1430),
.A2(n_491),
.B(n_490),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1490),
.B(n_23),
.Y(n_1584)
);

AOI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1396),
.A2(n_494),
.B(n_492),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1401),
.A2(n_496),
.B(n_495),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1478),
.B(n_23),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1452),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1425),
.A2(n_498),
.B(n_497),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1454),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1438),
.B(n_24),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1363),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_SL g1593 ( 
.A(n_1424),
.B(n_499),
.Y(n_1593)
);

A2O1A1Ixp33_ASAP7_75t_L g1594 ( 
.A1(n_1346),
.A2(n_1489),
.B(n_1435),
.C(n_1433),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1442),
.B(n_24),
.Y(n_1595)
);

CKINVDCx16_ASAP7_75t_R g1596 ( 
.A(n_1446),
.Y(n_1596)
);

AND2x2_ASAP7_75t_SL g1597 ( 
.A(n_1422),
.B(n_25),
.Y(n_1597)
);

AOI221xp5_ASAP7_75t_L g1598 ( 
.A1(n_1455),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.C(n_28),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_R g1599 ( 
.A(n_1340),
.B(n_501),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1406),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1448),
.B(n_27),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1385),
.B(n_28),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1413),
.A2(n_503),
.B(n_502),
.Y(n_1603)
);

OAI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1479),
.A2(n_507),
.B(n_506),
.Y(n_1604)
);

BUFx12f_ASAP7_75t_L g1605 ( 
.A(n_1449),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_L g1606 ( 
.A1(n_1429),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_1606)
);

INVx3_ASAP7_75t_L g1607 ( 
.A(n_1416),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_1414),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1459),
.B(n_1466),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1417),
.Y(n_1610)
);

AO31x2_ASAP7_75t_L g1611 ( 
.A1(n_1590),
.A2(n_1354),
.A3(n_1355),
.B(n_1468),
.Y(n_1611)
);

AO31x2_ASAP7_75t_L g1612 ( 
.A1(n_1592),
.A2(n_1594),
.A3(n_1573),
.B(n_1567),
.Y(n_1612)
);

INVx1_ASAP7_75t_SL g1613 ( 
.A(n_1498),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1497),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1516),
.B(n_1486),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_1494),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1502),
.B(n_1443),
.Y(n_1617)
);

AOI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1511),
.A2(n_1408),
.B(n_1411),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1504),
.B(n_1491),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1529),
.B(n_1471),
.Y(n_1620)
);

BUFx8_ASAP7_75t_L g1621 ( 
.A(n_1545),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1568),
.B(n_1410),
.Y(n_1622)
);

AO32x2_ASAP7_75t_L g1623 ( 
.A1(n_1501),
.A2(n_1378),
.A3(n_1349),
.B1(n_1418),
.B2(n_1391),
.Y(n_1623)
);

AOI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1609),
.A2(n_1367),
.B(n_1358),
.Y(n_1624)
);

AOI21xp5_ASAP7_75t_L g1625 ( 
.A1(n_1600),
.A2(n_1403),
.B(n_1357),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1493),
.B(n_1372),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1563),
.B(n_1374),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1499),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1519),
.Y(n_1629)
);

AOI21xp5_ASAP7_75t_L g1630 ( 
.A1(n_1604),
.A2(n_1427),
.B(n_1393),
.Y(n_1630)
);

O2A1O1Ixp33_ASAP7_75t_L g1631 ( 
.A1(n_1558),
.A2(n_1492),
.B(n_1587),
.C(n_1584),
.Y(n_1631)
);

BUFx4f_ASAP7_75t_L g1632 ( 
.A(n_1500),
.Y(n_1632)
);

NOR2xp67_ASAP7_75t_L g1633 ( 
.A(n_1605),
.B(n_1390),
.Y(n_1633)
);

OAI21x1_ASAP7_75t_SL g1634 ( 
.A1(n_1583),
.A2(n_1404),
.B(n_1394),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1515),
.Y(n_1635)
);

OAI21x1_ASAP7_75t_L g1636 ( 
.A1(n_1555),
.A2(n_1382),
.B(n_1426),
.Y(n_1636)
);

AOI21xp5_ASAP7_75t_L g1637 ( 
.A1(n_1554),
.A2(n_1420),
.B(n_509),
.Y(n_1637)
);

OAI21x1_ASAP7_75t_SL g1638 ( 
.A1(n_1513),
.A2(n_510),
.B(n_508),
.Y(n_1638)
);

AO32x2_ASAP7_75t_L g1639 ( 
.A1(n_1503),
.A2(n_32),
.A3(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_1639)
);

NOR2x1_ASAP7_75t_SL g1640 ( 
.A(n_1554),
.B(n_511),
.Y(n_1640)
);

OAI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1517),
.A2(n_514),
.B(n_512),
.Y(n_1641)
);

OAI21x1_ASAP7_75t_L g1642 ( 
.A1(n_1518),
.A2(n_517),
.B(n_515),
.Y(n_1642)
);

AOI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1570),
.A2(n_1580),
.B(n_1565),
.Y(n_1643)
);

A2O1A1Ixp33_ASAP7_75t_L g1644 ( 
.A1(n_1581),
.A2(n_34),
.B(n_32),
.C(n_33),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1528),
.Y(n_1645)
);

INVx4_ASAP7_75t_L g1646 ( 
.A(n_1536),
.Y(n_1646)
);

BUFx6f_ASAP7_75t_L g1647 ( 
.A(n_1524),
.Y(n_1647)
);

AOI21x1_ASAP7_75t_L g1648 ( 
.A1(n_1588),
.A2(n_519),
.B(n_518),
.Y(n_1648)
);

AOI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1520),
.A2(n_521),
.B(n_520),
.Y(n_1649)
);

AOI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1541),
.A2(n_524),
.B(n_522),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1593),
.A2(n_528),
.B(n_527),
.Y(n_1651)
);

AOI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1525),
.A2(n_532),
.B(n_529),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1533),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_1653)
);

AOI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1539),
.A2(n_1546),
.B(n_1575),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1562),
.Y(n_1655)
);

OAI221xp5_ASAP7_75t_L g1656 ( 
.A1(n_1495),
.A2(n_1521),
.B1(n_1526),
.B2(n_1606),
.C(n_1496),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1505),
.B(n_35),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1607),
.B(n_37),
.Y(n_1658)
);

A2O1A1Ixp33_ASAP7_75t_L g1659 ( 
.A1(n_1549),
.A2(n_39),
.B(n_37),
.C(n_38),
.Y(n_1659)
);

OAI21x1_ASAP7_75t_L g1660 ( 
.A1(n_1589),
.A2(n_534),
.B(n_533),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1510),
.Y(n_1661)
);

AO31x2_ASAP7_75t_L g1662 ( 
.A1(n_1574),
.A2(n_537),
.A3(n_538),
.B(n_535),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1507),
.B(n_1569),
.Y(n_1663)
);

AO31x2_ASAP7_75t_L g1664 ( 
.A1(n_1506),
.A2(n_542),
.A3(n_544),
.B(n_540),
.Y(n_1664)
);

INVx3_ASAP7_75t_L g1665 ( 
.A(n_1536),
.Y(n_1665)
);

AOI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1579),
.A2(n_546),
.B(n_545),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1578),
.B(n_38),
.Y(n_1667)
);

AOI21x1_ASAP7_75t_L g1668 ( 
.A1(n_1610),
.A2(n_548),
.B(n_547),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1534),
.B(n_39),
.Y(n_1669)
);

NOR2xp67_ASAP7_75t_L g1670 ( 
.A(n_1571),
.B(n_549),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1514),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1572),
.B(n_40),
.Y(n_1672)
);

OAI21x1_ASAP7_75t_L g1673 ( 
.A1(n_1561),
.A2(n_552),
.B(n_551),
.Y(n_1673)
);

INVx3_ASAP7_75t_L g1674 ( 
.A(n_1500),
.Y(n_1674)
);

A2O1A1Ixp33_ASAP7_75t_L g1675 ( 
.A1(n_1535),
.A2(n_43),
.B(n_40),
.C(n_42),
.Y(n_1675)
);

A2O1A1Ixp33_ASAP7_75t_L g1676 ( 
.A1(n_1542),
.A2(n_44),
.B(n_42),
.C(n_43),
.Y(n_1676)
);

AOI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1582),
.A2(n_555),
.B(n_553),
.Y(n_1677)
);

NOR4xp25_ASAP7_75t_L g1678 ( 
.A(n_1564),
.B(n_46),
.C(n_44),
.D(n_45),
.Y(n_1678)
);

AOI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1586),
.A2(n_1603),
.B(n_1532),
.Y(n_1679)
);

BUFx3_ASAP7_75t_L g1680 ( 
.A(n_1560),
.Y(n_1680)
);

OAI21x1_ASAP7_75t_L g1681 ( 
.A1(n_1566),
.A2(n_558),
.B(n_556),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1556),
.B(n_46),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1550),
.B(n_1557),
.Y(n_1683)
);

AOI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1585),
.A2(n_560),
.B(n_559),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1577),
.Y(n_1685)
);

AOI21xp5_ASAP7_75t_L g1686 ( 
.A1(n_1512),
.A2(n_563),
.B(n_562),
.Y(n_1686)
);

AOI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1596),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_1687)
);

OAI21x1_ASAP7_75t_L g1688 ( 
.A1(n_1523),
.A2(n_565),
.B(n_564),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1602),
.B(n_48),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_SL g1690 ( 
.A(n_1550),
.B(n_49),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1531),
.B(n_50),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1508),
.Y(n_1692)
);

BUFx4_ASAP7_75t_SL g1693 ( 
.A(n_1548),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1559),
.B(n_51),
.Y(n_1694)
);

AOI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1591),
.A2(n_569),
.B(n_568),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1557),
.B(n_570),
.Y(n_1696)
);

OAI21x1_ASAP7_75t_L g1697 ( 
.A1(n_1537),
.A2(n_576),
.B(n_572),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1544),
.B(n_51),
.Y(n_1698)
);

AOI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1595),
.A2(n_579),
.B(n_578),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1540),
.B(n_52),
.Y(n_1700)
);

A2O1A1Ixp33_ASAP7_75t_L g1701 ( 
.A1(n_1543),
.A2(n_55),
.B(n_53),
.C(n_54),
.Y(n_1701)
);

O2A1O1Ixp33_ASAP7_75t_L g1702 ( 
.A1(n_1547),
.A2(n_55),
.B(n_53),
.C(n_54),
.Y(n_1702)
);

AO22x1_ASAP7_75t_L g1703 ( 
.A1(n_1553),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_1703)
);

OAI21x1_ASAP7_75t_L g1704 ( 
.A1(n_1551),
.A2(n_581),
.B(n_580),
.Y(n_1704)
);

OA21x2_ASAP7_75t_L g1705 ( 
.A1(n_1601),
.A2(n_583),
.B(n_582),
.Y(n_1705)
);

A2O1A1Ixp33_ASAP7_75t_L g1706 ( 
.A1(n_1598),
.A2(n_58),
.B(n_56),
.C(n_57),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1552),
.A2(n_589),
.B(n_584),
.Y(n_1707)
);

BUFx6f_ASAP7_75t_L g1708 ( 
.A(n_1538),
.Y(n_1708)
);

O2A1O1Ixp33_ASAP7_75t_L g1709 ( 
.A1(n_1527),
.A2(n_62),
.B(n_59),
.C(n_60),
.Y(n_1709)
);

AOI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1608),
.A2(n_591),
.B(n_590),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1503),
.Y(n_1711)
);

OAI21x1_ASAP7_75t_L g1712 ( 
.A1(n_1530),
.A2(n_594),
.B(n_593),
.Y(n_1712)
);

O2A1O1Ixp33_ASAP7_75t_SL g1713 ( 
.A1(n_1576),
.A2(n_1597),
.B(n_1599),
.C(n_1522),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1576),
.A2(n_63),
.B1(n_60),
.B2(n_62),
.Y(n_1714)
);

AND3x2_ASAP7_75t_L g1715 ( 
.A(n_1509),
.B(n_64),
.C(n_65),
.Y(n_1715)
);

AOI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1573),
.A2(n_597),
.B(n_596),
.Y(n_1716)
);

INVxp67_ASAP7_75t_SL g1717 ( 
.A(n_1531),
.Y(n_1717)
);

AOI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1573),
.A2(n_600),
.B(n_599),
.Y(n_1718)
);

HB1xp67_ASAP7_75t_L g1719 ( 
.A(n_1498),
.Y(n_1719)
);

AOI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1504),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1504),
.B(n_68),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1497),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1563),
.B(n_601),
.Y(n_1723)
);

A2O1A1Ixp33_ASAP7_75t_L g1724 ( 
.A1(n_1504),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_1724)
);

OAI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1504),
.A2(n_604),
.B(n_602),
.Y(n_1725)
);

AO31x2_ASAP7_75t_L g1726 ( 
.A1(n_1590),
.A2(n_606),
.A3(n_608),
.B(n_605),
.Y(n_1726)
);

AO31x2_ASAP7_75t_L g1727 ( 
.A1(n_1590),
.A2(n_610),
.A3(n_611),
.B(n_609),
.Y(n_1727)
);

AOI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1504),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_1728)
);

INVxp67_ASAP7_75t_L g1729 ( 
.A(n_1531),
.Y(n_1729)
);

OAI21x1_ASAP7_75t_SL g1730 ( 
.A1(n_1604),
.A2(n_614),
.B(n_612),
.Y(n_1730)
);

OA21x2_ASAP7_75t_L g1731 ( 
.A1(n_1590),
.A2(n_619),
.B(n_617),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1502),
.B(n_72),
.Y(n_1732)
);

AO31x2_ASAP7_75t_L g1733 ( 
.A1(n_1590),
.A2(n_621),
.A3(n_622),
.B(n_620),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1497),
.Y(n_1734)
);

INVx3_ASAP7_75t_L g1735 ( 
.A(n_1524),
.Y(n_1735)
);

OAI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1504),
.A2(n_625),
.B(n_623),
.Y(n_1736)
);

OAI21x1_ASAP7_75t_L g1737 ( 
.A1(n_1555),
.A2(n_631),
.B(n_627),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_L g1738 ( 
.A(n_1504),
.B(n_72),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1504),
.B(n_73),
.Y(n_1739)
);

O2A1O1Ixp33_ASAP7_75t_L g1740 ( 
.A1(n_1504),
.A2(n_75),
.B(n_73),
.C(n_74),
.Y(n_1740)
);

OAI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1596),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_1741)
);

AOI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1573),
.A2(n_635),
.B(n_632),
.Y(n_1742)
);

CKINVDCx11_ASAP7_75t_R g1743 ( 
.A(n_1494),
.Y(n_1743)
);

AOI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1504),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_1744)
);

BUFx6f_ASAP7_75t_L g1745 ( 
.A(n_1524),
.Y(n_1745)
);

NOR2x1_ASAP7_75t_R g1746 ( 
.A(n_1494),
.B(n_636),
.Y(n_1746)
);

AO31x2_ASAP7_75t_L g1747 ( 
.A1(n_1590),
.A2(n_639),
.A3(n_640),
.B(n_637),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1497),
.Y(n_1748)
);

OAI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1721),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_1749)
);

BUFx12f_ASAP7_75t_L g1750 ( 
.A(n_1743),
.Y(n_1750)
);

INVx4_ASAP7_75t_SL g1751 ( 
.A(n_1647),
.Y(n_1751)
);

INVx6_ASAP7_75t_L g1752 ( 
.A(n_1647),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1614),
.Y(n_1753)
);

INVx6_ASAP7_75t_L g1754 ( 
.A(n_1745),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1748),
.Y(n_1755)
);

INVxp67_ASAP7_75t_L g1756 ( 
.A(n_1719),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1628),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1635),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1661),
.Y(n_1759)
);

INVx3_ASAP7_75t_L g1760 ( 
.A(n_1745),
.Y(n_1760)
);

AOI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1738),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_1761)
);

CKINVDCx11_ASAP7_75t_R g1762 ( 
.A(n_1629),
.Y(n_1762)
);

AOI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1656),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1619),
.B(n_83),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1645),
.Y(n_1765)
);

AOI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1739),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_1766)
);

AOI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1669),
.A2(n_1617),
.B1(n_1700),
.B2(n_1667),
.Y(n_1767)
);

OAI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1631),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1655),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1671),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1722),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1657),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_1772)
);

HB1xp67_ASAP7_75t_L g1773 ( 
.A(n_1613),
.Y(n_1773)
);

OAI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1663),
.A2(n_90),
.B1(n_87),
.B2(n_89),
.Y(n_1774)
);

AOI22xp33_ASAP7_75t_L g1775 ( 
.A1(n_1615),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_1775)
);

CKINVDCx5p33_ASAP7_75t_R g1776 ( 
.A(n_1693),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1682),
.B(n_91),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1734),
.Y(n_1778)
);

CKINVDCx5p33_ASAP7_75t_R g1779 ( 
.A(n_1616),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1685),
.Y(n_1780)
);

OR2x2_ASAP7_75t_L g1781 ( 
.A(n_1694),
.B(n_93),
.Y(n_1781)
);

OAI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1687),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_1782)
);

CKINVDCx20_ASAP7_75t_R g1783 ( 
.A(n_1621),
.Y(n_1783)
);

AOI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1732),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_1784)
);

AOI22xp33_ASAP7_75t_L g1785 ( 
.A1(n_1672),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1689),
.B(n_97),
.Y(n_1786)
);

BUFx12f_ASAP7_75t_L g1787 ( 
.A(n_1646),
.Y(n_1787)
);

OAI22xp33_ASAP7_75t_L g1788 ( 
.A1(n_1720),
.A2(n_1728),
.B1(n_1744),
.B2(n_1622),
.Y(n_1788)
);

OAI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1741),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1698),
.Y(n_1790)
);

BUFx3_ASAP7_75t_L g1791 ( 
.A(n_1632),
.Y(n_1791)
);

CKINVDCx5p33_ASAP7_75t_R g1792 ( 
.A(n_1665),
.Y(n_1792)
);

BUFx3_ASAP7_75t_L g1793 ( 
.A(n_1735),
.Y(n_1793)
);

INVx6_ASAP7_75t_L g1794 ( 
.A(n_1708),
.Y(n_1794)
);

AOI22xp33_ASAP7_75t_L g1795 ( 
.A1(n_1725),
.A2(n_102),
.B1(n_100),
.B2(n_101),
.Y(n_1795)
);

BUFx2_ASAP7_75t_L g1796 ( 
.A(n_1674),
.Y(n_1796)
);

AOI22xp33_ASAP7_75t_L g1797 ( 
.A1(n_1736),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_1797)
);

BUFx8_ASAP7_75t_L g1798 ( 
.A(n_1708),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1717),
.Y(n_1799)
);

CKINVDCx12_ASAP7_75t_R g1800 ( 
.A(n_1746),
.Y(n_1800)
);

AOI22xp33_ASAP7_75t_SL g1801 ( 
.A1(n_1730),
.A2(n_111),
.B1(n_119),
.B2(n_103),
.Y(n_1801)
);

OAI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1729),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_1802)
);

OAI22x1_ASAP7_75t_L g1803 ( 
.A1(n_1690),
.A2(n_107),
.B1(n_105),
.B2(n_106),
.Y(n_1803)
);

BUFx2_ASAP7_75t_L g1804 ( 
.A(n_1692),
.Y(n_1804)
);

BUFx6f_ASAP7_75t_L g1805 ( 
.A(n_1683),
.Y(n_1805)
);

AOI22xp33_ASAP7_75t_L g1806 ( 
.A1(n_1626),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1612),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1658),
.Y(n_1808)
);

CKINVDCx11_ASAP7_75t_R g1809 ( 
.A(n_1680),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1620),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_1810)
);

INVx1_ASAP7_75t_SL g1811 ( 
.A(n_1691),
.Y(n_1811)
);

BUFx6f_ASAP7_75t_L g1812 ( 
.A(n_1696),
.Y(n_1812)
);

OAI22xp5_ASAP7_75t_L g1813 ( 
.A1(n_1706),
.A2(n_114),
.B1(n_112),
.B2(n_113),
.Y(n_1813)
);

AOI22xp33_ASAP7_75t_L g1814 ( 
.A1(n_1627),
.A2(n_115),
.B1(n_112),
.B2(n_114),
.Y(n_1814)
);

CKINVDCx20_ASAP7_75t_R g1815 ( 
.A(n_1710),
.Y(n_1815)
);

INVx1_ASAP7_75t_SL g1816 ( 
.A(n_1723),
.Y(n_1816)
);

BUFx10_ASAP7_75t_L g1817 ( 
.A(n_1715),
.Y(n_1817)
);

AOI22xp33_ASAP7_75t_L g1818 ( 
.A1(n_1618),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1639),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1612),
.Y(n_1820)
);

BUFx4f_ASAP7_75t_SL g1821 ( 
.A(n_1633),
.Y(n_1821)
);

INVx2_ASAP7_75t_SL g1822 ( 
.A(n_1712),
.Y(n_1822)
);

BUFx8_ASAP7_75t_L g1823 ( 
.A(n_1639),
.Y(n_1823)
);

BUFx2_ASAP7_75t_L g1824 ( 
.A(n_1611),
.Y(n_1824)
);

OAI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1653),
.A2(n_118),
.B1(n_116),
.B2(n_117),
.Y(n_1825)
);

AND2x4_ASAP7_75t_L g1826 ( 
.A(n_1670),
.B(n_641),
.Y(n_1826)
);

AOI22xp33_ASAP7_75t_SL g1827 ( 
.A1(n_1640),
.A2(n_127),
.B1(n_135),
.B2(n_118),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1611),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1662),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1662),
.Y(n_1830)
);

BUFx4_ASAP7_75t_R g1831 ( 
.A(n_1703),
.Y(n_1831)
);

AOI22xp33_ASAP7_75t_L g1832 ( 
.A1(n_1651),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1726),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1726),
.Y(n_1834)
);

BUFx4f_ASAP7_75t_SL g1835 ( 
.A(n_1711),
.Y(n_1835)
);

BUFx6f_ASAP7_75t_L g1836 ( 
.A(n_1688),
.Y(n_1836)
);

INVx2_ASAP7_75t_SL g1837 ( 
.A(n_1727),
.Y(n_1837)
);

OAI21xp33_ASAP7_75t_L g1838 ( 
.A1(n_1701),
.A2(n_121),
.B(n_122),
.Y(n_1838)
);

NAND2x1p5_ASAP7_75t_L g1839 ( 
.A(n_1673),
.B(n_642),
.Y(n_1839)
);

BUFx3_ASAP7_75t_L g1840 ( 
.A(n_1638),
.Y(n_1840)
);

BUFx3_ASAP7_75t_L g1841 ( 
.A(n_1697),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_SL g1842 ( 
.A1(n_1714),
.A2(n_1630),
.B1(n_1650),
.B2(n_1649),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1727),
.Y(n_1843)
);

CKINVDCx20_ASAP7_75t_R g1844 ( 
.A(n_1705),
.Y(n_1844)
);

INVx6_ASAP7_75t_L g1845 ( 
.A(n_1644),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1733),
.Y(n_1846)
);

CKINVDCx6p67_ASAP7_75t_R g1847 ( 
.A(n_1675),
.Y(n_1847)
);

INVxp33_ASAP7_75t_L g1848 ( 
.A(n_1625),
.Y(n_1848)
);

CKINVDCx6p67_ASAP7_75t_R g1849 ( 
.A(n_1659),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1704),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1733),
.Y(n_1851)
);

AOI22xp33_ASAP7_75t_L g1852 ( 
.A1(n_1643),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1747),
.Y(n_1853)
);

BUFx2_ASAP7_75t_SL g1854 ( 
.A(n_1637),
.Y(n_1854)
);

BUFx3_ASAP7_75t_L g1855 ( 
.A(n_1641),
.Y(n_1855)
);

AOI22xp33_ASAP7_75t_L g1856 ( 
.A1(n_1695),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_1856)
);

OAI22xp5_ASAP7_75t_L g1857 ( 
.A1(n_1676),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1737),
.Y(n_1858)
);

OAI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1724),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1747),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_SL g1861 ( 
.A1(n_1716),
.A2(n_137),
.B1(n_145),
.B2(n_129),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1681),
.Y(n_1862)
);

BUFx12f_ASAP7_75t_L g1863 ( 
.A(n_1678),
.Y(n_1863)
);

AOI22xp5_ASAP7_75t_L g1864 ( 
.A1(n_1679),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.Y(n_1864)
);

CKINVDCx11_ASAP7_75t_R g1865 ( 
.A(n_1709),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1660),
.Y(n_1866)
);

BUFx6f_ASAP7_75t_L g1867 ( 
.A(n_1642),
.Y(n_1867)
);

INVx2_ASAP7_75t_SL g1868 ( 
.A(n_1664),
.Y(n_1868)
);

OAI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1740),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_1869)
);

AOI22xp33_ASAP7_75t_L g1870 ( 
.A1(n_1699),
.A2(n_136),
.B1(n_134),
.B2(n_135),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1664),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1702),
.B(n_136),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1648),
.Y(n_1873)
);

BUFx3_ASAP7_75t_L g1874 ( 
.A(n_1634),
.Y(n_1874)
);

AOI22xp33_ASAP7_75t_L g1875 ( 
.A1(n_1718),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.Y(n_1875)
);

NAND2x1p5_ASAP7_75t_L g1876 ( 
.A(n_1731),
.B(n_643),
.Y(n_1876)
);

AOI22xp33_ASAP7_75t_L g1877 ( 
.A1(n_1742),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.Y(n_1877)
);

AOI22xp33_ASAP7_75t_L g1878 ( 
.A1(n_1666),
.A2(n_1677),
.B1(n_1684),
.B2(n_1652),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1668),
.Y(n_1879)
);

AOI22xp33_ASAP7_75t_L g1880 ( 
.A1(n_1654),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1808),
.B(n_1713),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1804),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1759),
.Y(n_1883)
);

HB1xp67_ASAP7_75t_L g1884 ( 
.A(n_1799),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1767),
.B(n_1623),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1807),
.Y(n_1886)
);

INVx2_ASAP7_75t_SL g1887 ( 
.A(n_1752),
.Y(n_1887)
);

CKINVDCx11_ASAP7_75t_R g1888 ( 
.A(n_1750),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1757),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1770),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1758),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1765),
.Y(n_1892)
);

OAI22xp5_ASAP7_75t_L g1893 ( 
.A1(n_1849),
.A2(n_1686),
.B1(n_1707),
.B2(n_1624),
.Y(n_1893)
);

BUFx3_ASAP7_75t_L g1894 ( 
.A(n_1791),
.Y(n_1894)
);

BUFx3_ASAP7_75t_L g1895 ( 
.A(n_1787),
.Y(n_1895)
);

AOI21xp5_ASAP7_75t_L g1896 ( 
.A1(n_1878),
.A2(n_1636),
.B(n_1623),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1769),
.Y(n_1897)
);

INVx2_ASAP7_75t_SL g1898 ( 
.A(n_1752),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1773),
.B(n_142),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1771),
.Y(n_1900)
);

INVx4_ASAP7_75t_SL g1901 ( 
.A(n_1821),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1753),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1755),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1786),
.B(n_646),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1778),
.Y(n_1905)
);

INVx1_ASAP7_75t_SL g1906 ( 
.A(n_1762),
.Y(n_1906)
);

OAI22xp5_ASAP7_75t_L g1907 ( 
.A1(n_1811),
.A2(n_1845),
.B1(n_1847),
.B2(n_1763),
.Y(n_1907)
);

AOI21x1_ASAP7_75t_L g1908 ( 
.A1(n_1873),
.A2(n_649),
.B(n_647),
.Y(n_1908)
);

NOR2xp33_ASAP7_75t_L g1909 ( 
.A(n_1816),
.B(n_1756),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1780),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1829),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1764),
.B(n_651),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1830),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1833),
.Y(n_1914)
);

OAI21x1_ASAP7_75t_L g1915 ( 
.A1(n_1862),
.A2(n_653),
.B(n_652),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1790),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1834),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1777),
.B(n_654),
.Y(n_1918)
);

BUFx12f_ASAP7_75t_L g1919 ( 
.A(n_1776),
.Y(n_1919)
);

AND2x4_ASAP7_75t_L g1920 ( 
.A(n_1751),
.B(n_655),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1781),
.B(n_656),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1820),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1796),
.Y(n_1923)
);

INVx2_ASAP7_75t_SL g1924 ( 
.A(n_1754),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1843),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1835),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1872),
.B(n_143),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1846),
.Y(n_1928)
);

NOR2x1_ASAP7_75t_R g1929 ( 
.A(n_1809),
.B(n_657),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1851),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1853),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1860),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1823),
.Y(n_1933)
);

INVx3_ASAP7_75t_L g1934 ( 
.A(n_1840),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1819),
.Y(n_1935)
);

BUFx3_ASAP7_75t_L g1936 ( 
.A(n_1754),
.Y(n_1936)
);

CKINVDCx14_ASAP7_75t_R g1937 ( 
.A(n_1783),
.Y(n_1937)
);

INVx1_ASAP7_75t_SL g1938 ( 
.A(n_1792),
.Y(n_1938)
);

OR2x2_ASAP7_75t_L g1939 ( 
.A(n_1760),
.B(n_143),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1874),
.Y(n_1940)
);

INVx3_ASAP7_75t_L g1941 ( 
.A(n_1805),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1837),
.Y(n_1942)
);

INVxp33_ASAP7_75t_L g1943 ( 
.A(n_1805),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1871),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1824),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1879),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1788),
.B(n_144),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1828),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1844),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1845),
.B(n_144),
.Y(n_1950)
);

HB1xp67_ASAP7_75t_L g1951 ( 
.A(n_1863),
.Y(n_1951)
);

OAI21x1_ASAP7_75t_L g1952 ( 
.A1(n_1866),
.A2(n_659),
.B(n_658),
.Y(n_1952)
);

AOI22xp33_ASAP7_75t_L g1953 ( 
.A1(n_1865),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1868),
.Y(n_1954)
);

OR2x2_ASAP7_75t_L g1955 ( 
.A(n_1812),
.B(n_1793),
.Y(n_1955)
);

AO21x2_ASAP7_75t_L g1956 ( 
.A1(n_1850),
.A2(n_146),
.B(n_147),
.Y(n_1956)
);

AND2x4_ASAP7_75t_L g1957 ( 
.A(n_1751),
.B(n_661),
.Y(n_1957)
);

BUFx3_ASAP7_75t_L g1958 ( 
.A(n_1798),
.Y(n_1958)
);

INVx3_ASAP7_75t_L g1959 ( 
.A(n_1812),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1803),
.B(n_1784),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1858),
.Y(n_1961)
);

INVx3_ASAP7_75t_L g1962 ( 
.A(n_1794),
.Y(n_1962)
);

AOI22xp33_ASAP7_75t_L g1963 ( 
.A1(n_1838),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_1963)
);

O2A1O1Ixp33_ASAP7_75t_L g1964 ( 
.A1(n_1947),
.A2(n_1869),
.B(n_1857),
.C(n_1859),
.Y(n_1964)
);

NOR2xp33_ASAP7_75t_L g1965 ( 
.A(n_1938),
.B(n_1800),
.Y(n_1965)
);

NOR2xp33_ASAP7_75t_L g1966 ( 
.A(n_1943),
.B(n_1955),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1949),
.B(n_1848),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1933),
.B(n_1801),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1923),
.B(n_1827),
.Y(n_1969)
);

AOI221xp5_ASAP7_75t_L g1970 ( 
.A1(n_1953),
.A2(n_1782),
.B1(n_1789),
.B2(n_1749),
.C(n_1768),
.Y(n_1970)
);

AOI22xp33_ASAP7_75t_L g1971 ( 
.A1(n_1960),
.A2(n_1815),
.B1(n_1795),
.B2(n_1797),
.Y(n_1971)
);

NOR2xp33_ASAP7_75t_L g1972 ( 
.A(n_1909),
.B(n_1779),
.Y(n_1972)
);

A2O1A1Ixp33_ASAP7_75t_L g1973 ( 
.A1(n_1963),
.A2(n_1864),
.B(n_1813),
.C(n_1761),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1882),
.B(n_1855),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1884),
.B(n_1794),
.Y(n_1975)
);

BUFx12f_ASAP7_75t_L g1976 ( 
.A(n_1888),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1946),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1889),
.B(n_1842),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1891),
.B(n_1822),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1892),
.B(n_1841),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1897),
.Y(n_1981)
);

O2A1O1Ixp33_ASAP7_75t_L g1982 ( 
.A1(n_1907),
.A2(n_1774),
.B(n_1825),
.C(n_1802),
.Y(n_1982)
);

OAI22xp5_ASAP7_75t_L g1983 ( 
.A1(n_1951),
.A2(n_1766),
.B1(n_1772),
.B2(n_1852),
.Y(n_1983)
);

BUFx6f_ASAP7_75t_L g1984 ( 
.A(n_1936),
.Y(n_1984)
);

INVx3_ASAP7_75t_L g1985 ( 
.A(n_1894),
.Y(n_1985)
);

INVx8_ASAP7_75t_L g1986 ( 
.A(n_1919),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1916),
.B(n_1775),
.Y(n_1987)
);

OAI21xp5_ASAP7_75t_L g1988 ( 
.A1(n_1893),
.A2(n_1870),
.B(n_1856),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1902),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1900),
.B(n_1861),
.Y(n_1990)
);

OAI21xp5_ASAP7_75t_L g1991 ( 
.A1(n_1896),
.A2(n_1875),
.B(n_1877),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1905),
.B(n_1880),
.Y(n_1992)
);

AOI211xp5_ASAP7_75t_L g1993 ( 
.A1(n_1927),
.A2(n_1831),
.B(n_1826),
.C(n_1867),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1903),
.B(n_1810),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1910),
.B(n_1814),
.Y(n_1995)
);

O2A1O1Ixp33_ASAP7_75t_L g1996 ( 
.A1(n_1950),
.A2(n_1881),
.B(n_1818),
.C(n_1832),
.Y(n_1996)
);

OR2x6_ASAP7_75t_L g1997 ( 
.A(n_1934),
.B(n_1854),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1883),
.B(n_1806),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1885),
.B(n_1817),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1918),
.B(n_1785),
.Y(n_2000)
);

NOR2x1_ASAP7_75t_SL g2001 ( 
.A(n_1945),
.B(n_1867),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1921),
.B(n_1876),
.Y(n_2002)
);

OR2x6_ASAP7_75t_L g2003 ( 
.A(n_1934),
.B(n_1839),
.Y(n_2003)
);

OR2x2_ASAP7_75t_L g2004 ( 
.A(n_1935),
.B(n_1836),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1890),
.B(n_1836),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1911),
.Y(n_2006)
);

AOI22xp5_ASAP7_75t_L g2007 ( 
.A1(n_1912),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_2007)
);

AOI22xp5_ASAP7_75t_SL g2008 ( 
.A1(n_1926),
.A2(n_154),
.B1(n_151),
.B2(n_153),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1925),
.Y(n_2009)
);

AND2x4_ASAP7_75t_L g2010 ( 
.A(n_1940),
.B(n_662),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1904),
.B(n_151),
.Y(n_2011)
);

OAI21xp5_ASAP7_75t_L g2012 ( 
.A1(n_1915),
.A2(n_1952),
.B(n_1908),
.Y(n_2012)
);

NOR2xp33_ASAP7_75t_L g2013 ( 
.A(n_1906),
.B(n_153),
.Y(n_2013)
);

OAI21xp5_ASAP7_75t_L g2014 ( 
.A1(n_1908),
.A2(n_667),
.B(n_666),
.Y(n_2014)
);

CKINVDCx5p33_ASAP7_75t_R g2015 ( 
.A(n_1937),
.Y(n_2015)
);

A2O1A1Ixp33_ASAP7_75t_L g2016 ( 
.A1(n_1920),
.A2(n_156),
.B(n_154),
.C(n_155),
.Y(n_2016)
);

NOR2x1_ASAP7_75t_SL g2017 ( 
.A(n_1956),
.B(n_668),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1913),
.Y(n_2018)
);

AO22x2_ASAP7_75t_L g2019 ( 
.A1(n_1914),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_2019)
);

OAI22xp5_ASAP7_75t_L g2020 ( 
.A1(n_1959),
.A2(n_160),
.B1(n_158),
.B2(n_159),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1941),
.B(n_158),
.Y(n_2021)
);

AOI21x1_ASAP7_75t_L g2022 ( 
.A1(n_1942),
.A2(n_159),
.B(n_160),
.Y(n_2022)
);

HB1xp67_ASAP7_75t_L g2023 ( 
.A(n_1928),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1930),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1917),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1931),
.Y(n_2026)
);

NOR2x1_ASAP7_75t_SL g2027 ( 
.A(n_1954),
.B(n_669),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1899),
.B(n_161),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1941),
.B(n_161),
.Y(n_2029)
);

AND2x4_ASAP7_75t_L g2030 ( 
.A(n_1959),
.B(n_670),
.Y(n_2030)
);

AND2x4_ASAP7_75t_L g2031 ( 
.A(n_1887),
.B(n_671),
.Y(n_2031)
);

AO21x2_ASAP7_75t_L g2032 ( 
.A1(n_1944),
.A2(n_162),
.B(n_163),
.Y(n_2032)
);

O2A1O1Ixp33_ASAP7_75t_SL g2033 ( 
.A1(n_1939),
.A2(n_172),
.B(n_180),
.C(n_163),
.Y(n_2033)
);

AOI22xp33_ASAP7_75t_L g2034 ( 
.A1(n_1920),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.Y(n_2034)
);

AND2x6_ASAP7_75t_L g2035 ( 
.A(n_1957),
.B(n_674),
.Y(n_2035)
);

AO21x2_ASAP7_75t_L g2036 ( 
.A1(n_1886),
.A2(n_164),
.B(n_167),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1962),
.B(n_167),
.Y(n_2037)
);

BUFx2_ASAP7_75t_R g2038 ( 
.A(n_1958),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1999),
.B(n_1962),
.Y(n_2039)
);

OR2x2_ASAP7_75t_L g2040 ( 
.A(n_2023),
.B(n_1932),
.Y(n_2040)
);

INVxp67_ASAP7_75t_SL g2041 ( 
.A(n_1978),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1981),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1967),
.B(n_1989),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1974),
.B(n_1898),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1977),
.Y(n_2045)
);

OR2x2_ASAP7_75t_L g2046 ( 
.A(n_2006),
.B(n_1886),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_2009),
.Y(n_2047)
);

OR2x6_ASAP7_75t_SL g2048 ( 
.A(n_2015),
.B(n_1901),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_2018),
.Y(n_2049)
);

HB1xp67_ASAP7_75t_L g2050 ( 
.A(n_2004),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_2024),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2025),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_1975),
.B(n_1924),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_2026),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1979),
.Y(n_2055)
);

INVxp67_ASAP7_75t_L g2056 ( 
.A(n_1966),
.Y(n_2056)
);

BUFx6f_ASAP7_75t_L g2057 ( 
.A(n_1984),
.Y(n_2057)
);

HB1xp67_ASAP7_75t_L g2058 ( 
.A(n_1980),
.Y(n_2058)
);

AND2x4_ASAP7_75t_L g2059 ( 
.A(n_1997),
.B(n_1922),
.Y(n_2059)
);

INVxp67_ASAP7_75t_SL g2060 ( 
.A(n_2005),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2036),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2032),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_2022),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_2001),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2019),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_1985),
.B(n_1961),
.Y(n_2066)
);

OR2x2_ASAP7_75t_L g2067 ( 
.A(n_1997),
.B(n_1948),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2019),
.Y(n_2068)
);

NOR2x1p5_ASAP7_75t_L g2069 ( 
.A(n_1976),
.B(n_1895),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1990),
.B(n_1901),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1992),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_2021),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_2002),
.B(n_1957),
.Y(n_2073)
);

HB1xp67_ASAP7_75t_L g2074 ( 
.A(n_1995),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_1969),
.B(n_168),
.Y(n_2075)
);

NOR2xp33_ASAP7_75t_L g2076 ( 
.A(n_1972),
.B(n_1929),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_1968),
.B(n_168),
.Y(n_2077)
);

OAI22xp33_ASAP7_75t_L g2078 ( 
.A1(n_1988),
.A2(n_173),
.B1(n_169),
.B2(n_171),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_2029),
.Y(n_2079)
);

HB1xp67_ASAP7_75t_L g2080 ( 
.A(n_2012),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_1984),
.B(n_173),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_2037),
.B(n_174),
.Y(n_2082)
);

AND2x4_ASAP7_75t_L g2083 ( 
.A(n_2003),
.B(n_174),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_1993),
.B(n_175),
.Y(n_2084)
);

AOI21xp5_ASAP7_75t_L g2085 ( 
.A1(n_1991),
.A2(n_175),
.B(n_176),
.Y(n_2085)
);

BUFx2_ASAP7_75t_L g2086 ( 
.A(n_2003),
.Y(n_2086)
);

HB1xp67_ASAP7_75t_L g2087 ( 
.A(n_1994),
.Y(n_2087)
);

INVx2_ASAP7_75t_SL g2088 ( 
.A(n_1986),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_SL g2089 ( 
.A(n_1996),
.B(n_675),
.Y(n_2089)
);

INVxp67_ASAP7_75t_SL g2090 ( 
.A(n_2017),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_2027),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1987),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_2010),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1998),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2014),
.Y(n_2095)
);

INVx2_ASAP7_75t_SL g2096 ( 
.A(n_1986),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_2028),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_2000),
.B(n_176),
.Y(n_2098)
);

BUFx2_ASAP7_75t_L g2099 ( 
.A(n_2035),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_2011),
.B(n_177),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2033),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_1965),
.B(n_178),
.Y(n_2102)
);

OAI21xp5_ASAP7_75t_L g2103 ( 
.A1(n_1964),
.A2(n_179),
.B(n_180),
.Y(n_2103)
);

INVxp67_ASAP7_75t_SL g2104 ( 
.A(n_1982),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_2013),
.B(n_179),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_2038),
.B(n_181),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2008),
.Y(n_2107)
);

AOI22xp33_ASAP7_75t_L g2108 ( 
.A1(n_1970),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.Y(n_2108)
);

HB1xp67_ASAP7_75t_L g2109 ( 
.A(n_2031),
.Y(n_2109)
);

AOI22xp33_ASAP7_75t_L g2110 ( 
.A1(n_1971),
.A2(n_185),
.B1(n_182),
.B2(n_183),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_2030),
.B(n_185),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2020),
.Y(n_2112)
);

OR2x2_ASAP7_75t_L g2113 ( 
.A(n_1983),
.B(n_186),
.Y(n_2113)
);

INVxp67_ASAP7_75t_SL g2114 ( 
.A(n_2007),
.Y(n_2114)
);

INVxp33_ASAP7_75t_L g2115 ( 
.A(n_2034),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_2035),
.B(n_2016),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2035),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1973),
.Y(n_2118)
);

OR2x2_ASAP7_75t_L g2119 ( 
.A(n_2023),
.B(n_186),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_2074),
.B(n_187),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_2058),
.B(n_188),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2054),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_2050),
.B(n_188),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_2054),
.Y(n_2124)
);

OR2x2_ASAP7_75t_L g2125 ( 
.A(n_2071),
.B(n_189),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2041),
.B(n_190),
.Y(n_2126)
);

OR2x2_ASAP7_75t_L g2127 ( 
.A(n_2055),
.B(n_2040),
.Y(n_2127)
);

BUFx2_ASAP7_75t_L g2128 ( 
.A(n_2086),
.Y(n_2128)
);

AOI21xp5_ASAP7_75t_L g2129 ( 
.A1(n_2089),
.A2(n_2085),
.B(n_2103),
.Y(n_2129)
);

AND2x4_ASAP7_75t_SL g2130 ( 
.A(n_2057),
.B(n_782),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2042),
.Y(n_2131)
);

BUFx2_ASAP7_75t_L g2132 ( 
.A(n_2080),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_2087),
.B(n_190),
.Y(n_2133)
);

OR2x2_ASAP7_75t_SL g2134 ( 
.A(n_2107),
.B(n_191),
.Y(n_2134)
);

NAND5xp2_ASAP7_75t_L g2135 ( 
.A(n_2108),
.B(n_195),
.C(n_192),
.D(n_193),
.E(n_196),
.Y(n_2135)
);

NAND2x1p5_ASAP7_75t_SL g2136 ( 
.A(n_2116),
.B(n_192),
.Y(n_2136)
);

AOI221xp5_ASAP7_75t_L g2137 ( 
.A1(n_2078),
.A2(n_196),
.B1(n_193),
.B2(n_195),
.C(n_197),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_2060),
.B(n_2039),
.Y(n_2138)
);

OAI31xp33_ASAP7_75t_L g2139 ( 
.A1(n_2118),
.A2(n_200),
.A3(n_198),
.B(n_199),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_2045),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_2049),
.Y(n_2141)
);

OAI221xp5_ASAP7_75t_L g2142 ( 
.A1(n_2118),
.A2(n_200),
.B1(n_198),
.B2(n_199),
.C(n_201),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2052),
.Y(n_2143)
);

AOI221xp5_ASAP7_75t_L g2144 ( 
.A1(n_2104),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.C(n_205),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_2047),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_2051),
.Y(n_2146)
);

HB1xp67_ASAP7_75t_L g2147 ( 
.A(n_2043),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2092),
.B(n_202),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2046),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2094),
.B(n_203),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2065),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_2044),
.B(n_205),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_2068),
.B(n_206),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_2097),
.B(n_206),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_2066),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_2072),
.B(n_207),
.Y(n_2156)
);

OAI33xp33_ASAP7_75t_L g2157 ( 
.A1(n_2113),
.A2(n_210),
.A3(n_212),
.B1(n_207),
.B2(n_208),
.B3(n_211),
.Y(n_2157)
);

OR2x2_ASAP7_75t_L g2158 ( 
.A(n_2079),
.B(n_208),
.Y(n_2158)
);

OR2x2_ASAP7_75t_L g2159 ( 
.A(n_2056),
.B(n_212),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2053),
.B(n_213),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_2067),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_2062),
.B(n_214),
.Y(n_2162)
);

AND2x2_ASAP7_75t_L g2163 ( 
.A(n_2099),
.B(n_214),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_L g2164 ( 
.A(n_2095),
.B(n_216),
.Y(n_2164)
);

INVx1_ASAP7_75t_SL g2165 ( 
.A(n_2057),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_2064),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2061),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2063),
.Y(n_2168)
);

NOR2xp33_ASAP7_75t_L g2169 ( 
.A(n_2070),
.B(n_216),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2119),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_2117),
.B(n_217),
.Y(n_2171)
);

HB1xp67_ASAP7_75t_L g2172 ( 
.A(n_2059),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_2073),
.B(n_2059),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_2095),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_2091),
.Y(n_2175)
);

AND2x4_ASAP7_75t_L g2176 ( 
.A(n_2090),
.B(n_218),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_2098),
.B(n_218),
.Y(n_2177)
);

CKINVDCx5p33_ASAP7_75t_R g2178 ( 
.A(n_2048),
.Y(n_2178)
);

NOR3xp33_ASAP7_75t_L g2179 ( 
.A(n_2114),
.B(n_220),
.C(n_221),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_2109),
.B(n_221),
.Y(n_2180)
);

OAI33xp33_ASAP7_75t_L g2181 ( 
.A1(n_2101),
.A2(n_224),
.A3(n_227),
.B1(n_222),
.B2(n_223),
.B3(n_226),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2093),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_2057),
.Y(n_2183)
);

INVx3_ASAP7_75t_L g2184 ( 
.A(n_2088),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_2096),
.B(n_222),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2069),
.B(n_224),
.Y(n_2186)
);

INVxp67_ASAP7_75t_SL g2187 ( 
.A(n_2083),
.Y(n_2187)
);

HB1xp67_ASAP7_75t_L g2188 ( 
.A(n_2083),
.Y(n_2188)
);

OR2x2_ASAP7_75t_L g2189 ( 
.A(n_2112),
.B(n_227),
.Y(n_2189)
);

OAI22xp33_ASAP7_75t_L g2190 ( 
.A1(n_2115),
.A2(n_230),
.B1(n_228),
.B2(n_229),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_2077),
.B(n_228),
.Y(n_2191)
);

AND2x2_ASAP7_75t_L g2192 ( 
.A(n_2102),
.B(n_229),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_2081),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_2082),
.Y(n_2194)
);

AND2x2_ASAP7_75t_L g2195 ( 
.A(n_2075),
.B(n_230),
.Y(n_2195)
);

AND2x4_ASAP7_75t_L g2196 ( 
.A(n_2084),
.B(n_231),
.Y(n_2196)
);

OAI31xp33_ASAP7_75t_L g2197 ( 
.A1(n_2110),
.A2(n_234),
.A3(n_231),
.B(n_232),
.Y(n_2197)
);

OR2x2_ASAP7_75t_L g2198 ( 
.A(n_2100),
.B(n_232),
.Y(n_2198)
);

OAI31xp33_ASAP7_75t_L g2199 ( 
.A1(n_2106),
.A2(n_236),
.A3(n_234),
.B(n_235),
.Y(n_2199)
);

BUFx3_ASAP7_75t_L g2200 ( 
.A(n_2111),
.Y(n_2200)
);

OAI21xp5_ASAP7_75t_SL g2201 ( 
.A1(n_2076),
.A2(n_237),
.B(n_238),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_2105),
.B(n_237),
.Y(n_2202)
);

INVx5_ASAP7_75t_L g2203 ( 
.A(n_2083),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_2087),
.B(n_239),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2054),
.Y(n_2205)
);

AND2x2_ASAP7_75t_L g2206 ( 
.A(n_2074),
.B(n_239),
.Y(n_2206)
);

BUFx2_ASAP7_75t_L g2207 ( 
.A(n_2086),
.Y(n_2207)
);

BUFx3_ASAP7_75t_L g2208 ( 
.A(n_2057),
.Y(n_2208)
);

OR2x2_ASAP7_75t_L g2209 ( 
.A(n_2074),
.B(n_240),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2054),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_2074),
.B(n_241),
.Y(n_2211)
);

OR2x2_ASAP7_75t_L g2212 ( 
.A(n_2074),
.B(n_241),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_2074),
.B(n_242),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_2074),
.B(n_243),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_2074),
.B(n_243),
.Y(n_2215)
);

INVxp67_ASAP7_75t_L g2216 ( 
.A(n_2087),
.Y(n_2216)
);

AOI22xp33_ASAP7_75t_L g2217 ( 
.A1(n_2118),
.A2(n_246),
.B1(n_244),
.B2(n_245),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2054),
.Y(n_2218)
);

INVx2_ASAP7_75t_L g2219 ( 
.A(n_2124),
.Y(n_2219)
);

AND2x4_ASAP7_75t_L g2220 ( 
.A(n_2151),
.B(n_244),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_2216),
.B(n_2174),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_2128),
.B(n_245),
.Y(n_2222)
);

INVx1_ASAP7_75t_SL g2223 ( 
.A(n_2207),
.Y(n_2223)
);

INVx2_ASAP7_75t_SL g2224 ( 
.A(n_2203),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_2175),
.Y(n_2225)
);

HB1xp67_ASAP7_75t_L g2226 ( 
.A(n_2132),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_2122),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_2205),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2168),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2210),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_2218),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_2173),
.B(n_246),
.Y(n_2232)
);

AND2x2_ASAP7_75t_L g2233 ( 
.A(n_2172),
.B(n_247),
.Y(n_2233)
);

INVx3_ASAP7_75t_L g2234 ( 
.A(n_2203),
.Y(n_2234)
);

AND2x2_ASAP7_75t_L g2235 ( 
.A(n_2138),
.B(n_247),
.Y(n_2235)
);

OR2x2_ASAP7_75t_L g2236 ( 
.A(n_2127),
.B(n_248),
.Y(n_2236)
);

AND2x2_ASAP7_75t_SL g2237 ( 
.A(n_2179),
.B(n_248),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_2161),
.B(n_249),
.Y(n_2238)
);

NOR2xp33_ASAP7_75t_SL g2239 ( 
.A(n_2178),
.B(n_249),
.Y(n_2239)
);

AND2x2_ASAP7_75t_L g2240 ( 
.A(n_2147),
.B(n_2155),
.Y(n_2240)
);

NOR2xp67_ASAP7_75t_L g2241 ( 
.A(n_2203),
.B(n_250),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_2132),
.B(n_2166),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_2140),
.Y(n_2243)
);

AND2x2_ASAP7_75t_L g2244 ( 
.A(n_2170),
.B(n_250),
.Y(n_2244)
);

AND2x2_ASAP7_75t_L g2245 ( 
.A(n_2188),
.B(n_251),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_2141),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_2149),
.B(n_251),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_2182),
.B(n_252),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2167),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_2187),
.B(n_252),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_2194),
.B(n_253),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2131),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_2165),
.B(n_254),
.Y(n_2253)
);

OR2x2_ASAP7_75t_L g2254 ( 
.A(n_2145),
.B(n_254),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_2183),
.B(n_2208),
.Y(n_2255)
);

AND2x2_ASAP7_75t_L g2256 ( 
.A(n_2146),
.B(n_255),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2143),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2162),
.Y(n_2258)
);

OR2x2_ASAP7_75t_L g2259 ( 
.A(n_2209),
.B(n_256),
.Y(n_2259)
);

OR2x2_ASAP7_75t_L g2260 ( 
.A(n_2212),
.B(n_256),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_2164),
.B(n_257),
.Y(n_2261)
);

INVx3_ASAP7_75t_L g2262 ( 
.A(n_2176),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2184),
.B(n_257),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_2133),
.B(n_258),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2193),
.B(n_258),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2200),
.B(n_259),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2153),
.Y(n_2267)
);

HB1xp67_ASAP7_75t_L g2268 ( 
.A(n_2125),
.Y(n_2268)
);

INVxp67_ASAP7_75t_SL g2269 ( 
.A(n_2204),
.Y(n_2269)
);

AND2x2_ASAP7_75t_L g2270 ( 
.A(n_2120),
.B(n_260),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_2206),
.B(n_260),
.Y(n_2271)
);

AND2x2_ASAP7_75t_L g2272 ( 
.A(n_2211),
.B(n_262),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_2213),
.B(n_2214),
.Y(n_2273)
);

INVx1_ASAP7_75t_SL g2274 ( 
.A(n_2186),
.Y(n_2274)
);

OR2x2_ASAP7_75t_L g2275 ( 
.A(n_2158),
.B(n_262),
.Y(n_2275)
);

AND2x2_ASAP7_75t_L g2276 ( 
.A(n_2215),
.B(n_263),
.Y(n_2276)
);

HB1xp67_ASAP7_75t_L g2277 ( 
.A(n_2123),
.Y(n_2277)
);

AND2x2_ASAP7_75t_L g2278 ( 
.A(n_2121),
.B(n_263),
.Y(n_2278)
);

AND2x4_ASAP7_75t_L g2279 ( 
.A(n_2176),
.B(n_264),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_2126),
.B(n_264),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2150),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_2189),
.B(n_265),
.Y(n_2282)
);

OAI22xp5_ASAP7_75t_L g2283 ( 
.A1(n_2129),
.A2(n_2142),
.B1(n_2137),
.B2(n_2201),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_2180),
.B(n_267),
.Y(n_2284)
);

HB1xp67_ASAP7_75t_L g2285 ( 
.A(n_2171),
.Y(n_2285)
);

AND2x2_ASAP7_75t_L g2286 ( 
.A(n_2163),
.B(n_267),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_2196),
.B(n_268),
.Y(n_2287)
);

AND2x2_ASAP7_75t_L g2288 ( 
.A(n_2196),
.B(n_268),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_2152),
.B(n_269),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_2148),
.B(n_269),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_2156),
.Y(n_2291)
);

AND2x4_ASAP7_75t_L g2292 ( 
.A(n_2185),
.B(n_270),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_2160),
.B(n_270),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2154),
.B(n_271),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_2191),
.B(n_271),
.Y(n_2295)
);

AND2x2_ASAP7_75t_L g2296 ( 
.A(n_2195),
.B(n_272),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_2159),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2177),
.Y(n_2298)
);

HB1xp67_ASAP7_75t_L g2299 ( 
.A(n_2198),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2136),
.Y(n_2300)
);

AND2x4_ASAP7_75t_SL g2301 ( 
.A(n_2192),
.B(n_272),
.Y(n_2301)
);

NOR2x1_ASAP7_75t_L g2302 ( 
.A(n_2169),
.B(n_273),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2134),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_2202),
.B(n_2130),
.Y(n_2304)
);

NOR2x1p5_ASAP7_75t_L g2305 ( 
.A(n_2199),
.B(n_273),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2190),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2144),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2217),
.Y(n_2308)
);

AND2x2_ASAP7_75t_L g2309 ( 
.A(n_2139),
.B(n_274),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_2197),
.B(n_274),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2157),
.B(n_276),
.Y(n_2311)
);

BUFx2_ASAP7_75t_L g2312 ( 
.A(n_2181),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2135),
.Y(n_2313)
);

AND4x1_ASAP7_75t_L g2314 ( 
.A(n_2129),
.B(n_278),
.C(n_276),
.D(n_277),
.Y(n_2314)
);

NOR2xp33_ASAP7_75t_L g2315 ( 
.A(n_2178),
.B(n_277),
.Y(n_2315)
);

AOI22xp5_ASAP7_75t_L g2316 ( 
.A1(n_2129),
.A2(n_281),
.B1(n_279),
.B2(n_280),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2216),
.B(n_280),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2216),
.B(n_281),
.Y(n_2318)
);

AND2x2_ASAP7_75t_L g2319 ( 
.A(n_2128),
.B(n_282),
.Y(n_2319)
);

INVx1_ASAP7_75t_SL g2320 ( 
.A(n_2128),
.Y(n_2320)
);

AND2x2_ASAP7_75t_L g2321 ( 
.A(n_2128),
.B(n_282),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2216),
.B(n_283),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2168),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_2124),
.Y(n_2324)
);

OAI222xp33_ASAP7_75t_L g2325 ( 
.A1(n_2129),
.A2(n_285),
.B1(n_287),
.B2(n_283),
.C1(n_284),
.C2(n_286),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2168),
.Y(n_2326)
);

OR2x2_ASAP7_75t_L g2327 ( 
.A(n_2216),
.B(n_284),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2128),
.B(n_285),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2168),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2168),
.Y(n_2330)
);

NOR2x1_ASAP7_75t_L g2331 ( 
.A(n_2234),
.B(n_286),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2326),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_2269),
.B(n_288),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2326),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2229),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2323),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2300),
.B(n_288),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_2223),
.B(n_289),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2320),
.B(n_289),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2329),
.Y(n_2340)
);

NOR2xp33_ASAP7_75t_L g2341 ( 
.A(n_2303),
.B(n_290),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2258),
.B(n_290),
.Y(n_2342)
);

AOI21xp33_ASAP7_75t_L g2343 ( 
.A1(n_2283),
.A2(n_291),
.B(n_292),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2330),
.Y(n_2344)
);

INVx1_ASAP7_75t_SL g2345 ( 
.A(n_2274),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2230),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2262),
.B(n_291),
.Y(n_2347)
);

AOI22xp5_ASAP7_75t_L g2348 ( 
.A1(n_2307),
.A2(n_294),
.B1(n_292),
.B2(n_293),
.Y(n_2348)
);

OR2x2_ASAP7_75t_L g2349 ( 
.A(n_2297),
.B(n_293),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_2234),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2252),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2257),
.Y(n_2352)
);

AND2x2_ASAP7_75t_L g2353 ( 
.A(n_2262),
.B(n_294),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2249),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2227),
.Y(n_2355)
);

INVx1_ASAP7_75t_SL g2356 ( 
.A(n_2222),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2281),
.B(n_295),
.Y(n_2357)
);

AND2x4_ASAP7_75t_L g2358 ( 
.A(n_2224),
.B(n_295),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2240),
.B(n_296),
.Y(n_2359)
);

BUFx2_ASAP7_75t_L g2360 ( 
.A(n_2226),
.Y(n_2360)
);

AND2x2_ASAP7_75t_L g2361 ( 
.A(n_2242),
.B(n_298),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_SL g2362 ( 
.A(n_2241),
.B(n_299),
.Y(n_2362)
);

OR2x2_ASAP7_75t_L g2363 ( 
.A(n_2299),
.B(n_2221),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2267),
.B(n_299),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_2298),
.B(n_300),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2228),
.Y(n_2366)
);

INVx3_ASAP7_75t_SL g2367 ( 
.A(n_2301),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2231),
.Y(n_2368)
);

INVx3_ASAP7_75t_L g2369 ( 
.A(n_2255),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2268),
.B(n_2277),
.Y(n_2370)
);

OR2x2_ASAP7_75t_L g2371 ( 
.A(n_2236),
.B(n_300),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2243),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2246),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2219),
.Y(n_2374)
);

NAND2x1_ASAP7_75t_L g2375 ( 
.A(n_2324),
.B(n_301),
.Y(n_2375)
);

INVxp67_ASAP7_75t_L g2376 ( 
.A(n_2302),
.Y(n_2376)
);

INVx2_ASAP7_75t_SL g2377 ( 
.A(n_2285),
.Y(n_2377)
);

OR2x2_ASAP7_75t_L g2378 ( 
.A(n_2291),
.B(n_301),
.Y(n_2378)
);

INVx1_ASAP7_75t_SL g2379 ( 
.A(n_2319),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2247),
.B(n_302),
.Y(n_2380)
);

NAND2x1p5_ASAP7_75t_L g2381 ( 
.A(n_2279),
.B(n_302),
.Y(n_2381)
);

OR2x2_ASAP7_75t_L g2382 ( 
.A(n_2273),
.B(n_303),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2256),
.B(n_304),
.Y(n_2383)
);

NAND2x1_ASAP7_75t_L g2384 ( 
.A(n_2225),
.B(n_304),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_2220),
.Y(n_2385)
);

NOR2xp33_ASAP7_75t_L g2386 ( 
.A(n_2261),
.B(n_305),
.Y(n_2386)
);

AND2x2_ASAP7_75t_L g2387 ( 
.A(n_2235),
.B(n_305),
.Y(n_2387)
);

INVxp67_ASAP7_75t_SL g2388 ( 
.A(n_2254),
.Y(n_2388)
);

INVx3_ASAP7_75t_L g2389 ( 
.A(n_2279),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_2220),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2327),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2238),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2317),
.Y(n_2393)
);

INVx3_ASAP7_75t_L g2394 ( 
.A(n_2292),
.Y(n_2394)
);

NOR2x1p5_ASAP7_75t_SL g2395 ( 
.A(n_2306),
.B(n_306),
.Y(n_2395)
);

NOR4xp25_ASAP7_75t_L g2396 ( 
.A(n_2325),
.B(n_309),
.C(n_307),
.D(n_308),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2248),
.B(n_307),
.Y(n_2397)
);

OR2x2_ASAP7_75t_L g2398 ( 
.A(n_2318),
.B(n_308),
.Y(n_2398)
);

INVxp67_ASAP7_75t_SL g2399 ( 
.A(n_2282),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_2253),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2322),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2233),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2312),
.B(n_309),
.Y(n_2403)
);

INVxp67_ASAP7_75t_L g2404 ( 
.A(n_2239),
.Y(n_2404)
);

AND2x4_ASAP7_75t_L g2405 ( 
.A(n_2245),
.B(n_310),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2251),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_2312),
.B(n_310),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2244),
.Y(n_2408)
);

INVxp67_ASAP7_75t_SL g2409 ( 
.A(n_2321),
.Y(n_2409)
);

AOI32xp33_ASAP7_75t_L g2410 ( 
.A1(n_2310),
.A2(n_313),
.A3(n_311),
.B1(n_312),
.B2(n_314),
.Y(n_2410)
);

AND2x2_ASAP7_75t_L g2411 ( 
.A(n_2232),
.B(n_311),
.Y(n_2411)
);

OR2x2_ASAP7_75t_L g2412 ( 
.A(n_2275),
.B(n_313),
.Y(n_2412)
);

AND2x2_ASAP7_75t_L g2413 ( 
.A(n_2328),
.B(n_315),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_L g2414 ( 
.A(n_2250),
.B(n_316),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_2265),
.B(n_316),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2259),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2260),
.Y(n_2417)
);

INVx3_ASAP7_75t_L g2418 ( 
.A(n_2292),
.Y(n_2418)
);

AND2x2_ASAP7_75t_L g2419 ( 
.A(n_2304),
.B(n_317),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2308),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2263),
.Y(n_2421)
);

INVx2_ASAP7_75t_L g2422 ( 
.A(n_2266),
.Y(n_2422)
);

AND2x2_ASAP7_75t_L g2423 ( 
.A(n_2270),
.B(n_317),
.Y(n_2423)
);

OAI21xp33_ASAP7_75t_L g2424 ( 
.A1(n_2316),
.A2(n_318),
.B(n_320),
.Y(n_2424)
);

OA21x2_ASAP7_75t_L g2425 ( 
.A1(n_2264),
.A2(n_2290),
.B(n_2294),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_2287),
.Y(n_2426)
);

OR2x2_ASAP7_75t_L g2427 ( 
.A(n_2271),
.B(n_320),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_2272),
.B(n_321),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2276),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2278),
.B(n_321),
.Y(n_2430)
);

AND2x2_ASAP7_75t_L g2431 ( 
.A(n_2280),
.B(n_322),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2288),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2311),
.Y(n_2433)
);

INVxp67_ASAP7_75t_SL g2434 ( 
.A(n_2305),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_2237),
.B(n_322),
.Y(n_2435)
);

OA211x2_ASAP7_75t_L g2436 ( 
.A1(n_2315),
.A2(n_325),
.B(n_323),
.C(n_324),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2284),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_2286),
.B(n_323),
.Y(n_2438)
);

HB1xp67_ASAP7_75t_L g2439 ( 
.A(n_2289),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2293),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2295),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_2296),
.Y(n_2442)
);

OAI22xp5_ASAP7_75t_L g2443 ( 
.A1(n_2313),
.A2(n_2309),
.B1(n_2314),
.B2(n_328),
.Y(n_2443)
);

INVx3_ASAP7_75t_L g2444 ( 
.A(n_2234),
.Y(n_2444)
);

INVxp67_ASAP7_75t_L g2445 ( 
.A(n_2300),
.Y(n_2445)
);

NOR2xp33_ASAP7_75t_L g2446 ( 
.A(n_2303),
.B(n_326),
.Y(n_2446)
);

AND2x2_ASAP7_75t_L g2447 ( 
.A(n_2223),
.B(n_326),
.Y(n_2447)
);

OR2x2_ASAP7_75t_L g2448 ( 
.A(n_2269),
.B(n_327),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2326),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2269),
.B(n_329),
.Y(n_2450)
);

NOR2x1_ASAP7_75t_L g2451 ( 
.A(n_2234),
.B(n_329),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_2234),
.Y(n_2452)
);

AND2x2_ASAP7_75t_L g2453 ( 
.A(n_2223),
.B(n_330),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2269),
.B(n_330),
.Y(n_2454)
);

INVx2_ASAP7_75t_L g2455 ( 
.A(n_2234),
.Y(n_2455)
);

INVx2_ASAP7_75t_SL g2456 ( 
.A(n_2234),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_2234),
.Y(n_2457)
);

OAI21xp33_ASAP7_75t_L g2458 ( 
.A1(n_2283),
.A2(n_332),
.B(n_333),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2326),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2326),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_2269),
.B(n_333),
.Y(n_2461)
);

OR2x2_ASAP7_75t_L g2462 ( 
.A(n_2269),
.B(n_334),
.Y(n_2462)
);

OR2x2_ASAP7_75t_L g2463 ( 
.A(n_2269),
.B(n_334),
.Y(n_2463)
);

NOR2x2_ASAP7_75t_L g2464 ( 
.A(n_2297),
.B(n_335),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2234),
.Y(n_2465)
);

AND2x2_ASAP7_75t_L g2466 ( 
.A(n_2223),
.B(n_336),
.Y(n_2466)
);

INVx2_ASAP7_75t_SL g2467 ( 
.A(n_2234),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2326),
.Y(n_2468)
);

INVx3_ASAP7_75t_L g2469 ( 
.A(n_2234),
.Y(n_2469)
);

BUFx3_ASAP7_75t_L g2470 ( 
.A(n_2292),
.Y(n_2470)
);

BUFx2_ASAP7_75t_L g2471 ( 
.A(n_2234),
.Y(n_2471)
);

OR2x2_ASAP7_75t_L g2472 ( 
.A(n_2269),
.B(n_336),
.Y(n_2472)
);

AND2x2_ASAP7_75t_L g2473 ( 
.A(n_2223),
.B(n_337),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_L g2474 ( 
.A(n_2269),
.B(n_337),
.Y(n_2474)
);

AND2x2_ASAP7_75t_L g2475 ( 
.A(n_2223),
.B(n_338),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2326),
.Y(n_2476)
);

BUFx3_ASAP7_75t_L g2477 ( 
.A(n_2292),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2326),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2326),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2326),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2326),
.Y(n_2481)
);

HB1xp67_ASAP7_75t_L g2482 ( 
.A(n_2226),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2269),
.B(n_338),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2326),
.Y(n_2484)
);

AND2x2_ASAP7_75t_L g2485 ( 
.A(n_2223),
.B(n_339),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2326),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2326),
.Y(n_2487)
);

OR2x2_ASAP7_75t_L g2488 ( 
.A(n_2269),
.B(n_339),
.Y(n_2488)
);

AND2x2_ASAP7_75t_L g2489 ( 
.A(n_2223),
.B(n_340),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2269),
.B(n_340),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2269),
.B(n_342),
.Y(n_2491)
);

AND2x2_ASAP7_75t_L g2492 ( 
.A(n_2223),
.B(n_342),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_2269),
.B(n_343),
.Y(n_2493)
);

NAND2xp67_ASAP7_75t_SL g2494 ( 
.A(n_2309),
.B(n_343),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2326),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2326),
.Y(n_2496)
);

NAND2x1_ASAP7_75t_L g2497 ( 
.A(n_2234),
.B(n_344),
.Y(n_2497)
);

AND2x2_ASAP7_75t_L g2498 ( 
.A(n_2369),
.B(n_344),
.Y(n_2498)
);

AND2x2_ASAP7_75t_L g2499 ( 
.A(n_2399),
.B(n_345),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_SL g2500 ( 
.A(n_2376),
.B(n_345),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_2471),
.Y(n_2501)
);

AND2x2_ASAP7_75t_L g2502 ( 
.A(n_2345),
.B(n_346),
.Y(n_2502)
);

OR2x2_ASAP7_75t_L g2503 ( 
.A(n_2370),
.B(n_346),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_SL g2504 ( 
.A(n_2377),
.B(n_347),
.Y(n_2504)
);

INVx2_ASAP7_75t_SL g2505 ( 
.A(n_2470),
.Y(n_2505)
);

INVx1_ASAP7_75t_SL g2506 ( 
.A(n_2367),
.Y(n_2506)
);

INVxp67_ASAP7_75t_L g2507 ( 
.A(n_2434),
.Y(n_2507)
);

AOI21xp5_ASAP7_75t_L g2508 ( 
.A1(n_2403),
.A2(n_347),
.B(n_348),
.Y(n_2508)
);

OR2x2_ASAP7_75t_L g2509 ( 
.A(n_2445),
.B(n_348),
.Y(n_2509)
);

NOR2x1_ASAP7_75t_L g2510 ( 
.A(n_2331),
.B(n_349),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2332),
.Y(n_2511)
);

HB1xp67_ASAP7_75t_L g2512 ( 
.A(n_2360),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_L g2513 ( 
.A(n_2433),
.B(n_2388),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2334),
.Y(n_2514)
);

NOR2xp33_ASAP7_75t_L g2515 ( 
.A(n_2394),
.B(n_350),
.Y(n_2515)
);

NAND4xp25_ASAP7_75t_L g2516 ( 
.A(n_2410),
.B(n_352),
.C(n_350),
.D(n_351),
.Y(n_2516)
);

AND2x2_ASAP7_75t_L g2517 ( 
.A(n_2418),
.B(n_351),
.Y(n_2517)
);

HB1xp67_ASAP7_75t_L g2518 ( 
.A(n_2482),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2416),
.B(n_352),
.Y(n_2519)
);

OR2x2_ASAP7_75t_L g2520 ( 
.A(n_2363),
.B(n_2420),
.Y(n_2520)
);

AND2x2_ASAP7_75t_L g2521 ( 
.A(n_2385),
.B(n_353),
.Y(n_2521)
);

AND2x2_ASAP7_75t_L g2522 ( 
.A(n_2390),
.B(n_353),
.Y(n_2522)
);

AO21x2_ASAP7_75t_L g2523 ( 
.A1(n_2407),
.A2(n_354),
.B(n_355),
.Y(n_2523)
);

AND2x2_ASAP7_75t_L g2524 ( 
.A(n_2389),
.B(n_354),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_L g2525 ( 
.A(n_2417),
.B(n_355),
.Y(n_2525)
);

OR2x2_ASAP7_75t_L g2526 ( 
.A(n_2425),
.B(n_356),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_2391),
.B(n_356),
.Y(n_2527)
);

INVx2_ASAP7_75t_SL g2528 ( 
.A(n_2477),
.Y(n_2528)
);

INVx2_ASAP7_75t_L g2529 ( 
.A(n_2444),
.Y(n_2529)
);

INVx2_ASAP7_75t_L g2530 ( 
.A(n_2469),
.Y(n_2530)
);

AND2x2_ASAP7_75t_L g2531 ( 
.A(n_2439),
.B(n_357),
.Y(n_2531)
);

NOR2xp33_ASAP7_75t_L g2532 ( 
.A(n_2404),
.B(n_2393),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2449),
.Y(n_2533)
);

AOI22xp5_ASAP7_75t_L g2534 ( 
.A1(n_2458),
.A2(n_359),
.B1(n_357),
.B2(n_358),
.Y(n_2534)
);

AOI21xp5_ASAP7_75t_L g2535 ( 
.A1(n_2343),
.A2(n_359),
.B(n_360),
.Y(n_2535)
);

AND2x4_ASAP7_75t_L g2536 ( 
.A(n_2456),
.B(n_360),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2459),
.Y(n_2537)
);

AND2x2_ASAP7_75t_L g2538 ( 
.A(n_2409),
.B(n_361),
.Y(n_2538)
);

AOI21xp33_ASAP7_75t_L g2539 ( 
.A1(n_2467),
.A2(n_361),
.B(n_362),
.Y(n_2539)
);

AND2x2_ASAP7_75t_L g2540 ( 
.A(n_2425),
.B(n_363),
.Y(n_2540)
);

AND2x2_ASAP7_75t_L g2541 ( 
.A(n_2401),
.B(n_364),
.Y(n_2541)
);

OR2x2_ASAP7_75t_L g2542 ( 
.A(n_2356),
.B(n_2379),
.Y(n_2542)
);

AND2x2_ASAP7_75t_L g2543 ( 
.A(n_2426),
.B(n_364),
.Y(n_2543)
);

AND2x2_ASAP7_75t_L g2544 ( 
.A(n_2432),
.B(n_365),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_L g2545 ( 
.A(n_2400),
.B(n_365),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2350),
.Y(n_2546)
);

NAND2xp33_ASAP7_75t_L g2547 ( 
.A(n_2451),
.B(n_366),
.Y(n_2547)
);

AND2x2_ASAP7_75t_L g2548 ( 
.A(n_2452),
.B(n_367),
.Y(n_2548)
);

HB1xp67_ASAP7_75t_L g2549 ( 
.A(n_2460),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2468),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2455),
.Y(n_2551)
);

INVxp67_ASAP7_75t_L g2552 ( 
.A(n_2341),
.Y(n_2552)
);

OR2x2_ASAP7_75t_L g2553 ( 
.A(n_2402),
.B(n_367),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2421),
.B(n_368),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2476),
.Y(n_2555)
);

OR2x2_ASAP7_75t_L g2556 ( 
.A(n_2408),
.B(n_368),
.Y(n_2556)
);

OAI22xp33_ASAP7_75t_L g2557 ( 
.A1(n_2443),
.A2(n_371),
.B1(n_369),
.B2(n_370),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2478),
.Y(n_2558)
);

INVx1_ASAP7_75t_SL g2559 ( 
.A(n_2464),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2479),
.Y(n_2560)
);

AND2x2_ASAP7_75t_L g2561 ( 
.A(n_2457),
.B(n_369),
.Y(n_2561)
);

AOI31xp33_ASAP7_75t_L g2562 ( 
.A1(n_2381),
.A2(n_372),
.A3(n_370),
.B(n_371),
.Y(n_2562)
);

AND2x2_ASAP7_75t_L g2563 ( 
.A(n_2465),
.B(n_373),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2480),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2481),
.Y(n_2565)
);

OR2x2_ASAP7_75t_L g2566 ( 
.A(n_2372),
.B(n_373),
.Y(n_2566)
);

OR2x2_ASAP7_75t_L g2567 ( 
.A(n_2373),
.B(n_374),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2484),
.Y(n_2568)
);

OR2x2_ASAP7_75t_L g2569 ( 
.A(n_2392),
.B(n_374),
.Y(n_2569)
);

INVx1_ASAP7_75t_SL g2570 ( 
.A(n_2497),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2486),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2487),
.Y(n_2572)
);

OR2x2_ASAP7_75t_L g2573 ( 
.A(n_2429),
.B(n_375),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_SL g2574 ( 
.A(n_2396),
.B(n_375),
.Y(n_2574)
);

NAND2x1_ASAP7_75t_L g2575 ( 
.A(n_2335),
.B(n_376),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_L g2576 ( 
.A(n_2395),
.B(n_376),
.Y(n_2576)
);

OAI33xp33_ASAP7_75t_L g2577 ( 
.A1(n_2494),
.A2(n_379),
.A3(n_381),
.B1(n_377),
.B2(n_378),
.B3(n_380),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2347),
.B(n_2353),
.Y(n_2578)
);

HB1xp67_ASAP7_75t_L g2579 ( 
.A(n_2495),
.Y(n_2579)
);

NOR2x1_ASAP7_75t_L g2580 ( 
.A(n_2448),
.B(n_377),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2422),
.B(n_378),
.Y(n_2581)
);

NOR2xp33_ASAP7_75t_L g2582 ( 
.A(n_2337),
.B(n_379),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_L g2583 ( 
.A(n_2406),
.B(n_381),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2496),
.Y(n_2584)
);

NAND4xp25_ASAP7_75t_L g2585 ( 
.A(n_2436),
.B(n_384),
.C(n_382),
.D(n_383),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2346),
.Y(n_2586)
);

OR2x2_ASAP7_75t_L g2587 ( 
.A(n_2437),
.B(n_383),
.Y(n_2587)
);

NOR2xp33_ASAP7_75t_L g2588 ( 
.A(n_2382),
.B(n_384),
.Y(n_2588)
);

NOR2x1_ASAP7_75t_L g2589 ( 
.A(n_2462),
.B(n_385),
.Y(n_2589)
);

OR2x2_ASAP7_75t_L g2590 ( 
.A(n_2440),
.B(n_385),
.Y(n_2590)
);

OR2x2_ASAP7_75t_L g2591 ( 
.A(n_2441),
.B(n_386),
.Y(n_2591)
);

AND2x2_ASAP7_75t_L g2592 ( 
.A(n_2442),
.B(n_386),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2336),
.Y(n_2593)
);

INVx1_ASAP7_75t_SL g2594 ( 
.A(n_2338),
.Y(n_2594)
);

OR2x2_ASAP7_75t_L g2595 ( 
.A(n_2374),
.B(n_387),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2361),
.B(n_387),
.Y(n_2596)
);

AND2x4_ASAP7_75t_L g2597 ( 
.A(n_2358),
.B(n_388),
.Y(n_2597)
);

AND2x2_ASAP7_75t_L g2598 ( 
.A(n_2359),
.B(n_388),
.Y(n_2598)
);

AND2x2_ASAP7_75t_L g2599 ( 
.A(n_2339),
.B(n_389),
.Y(n_2599)
);

AND2x2_ASAP7_75t_L g2600 ( 
.A(n_2447),
.B(n_389),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2333),
.B(n_390),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2340),
.Y(n_2602)
);

OR2x6_ASAP7_75t_L g2603 ( 
.A(n_2384),
.B(n_2375),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2358),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2453),
.B(n_2466),
.Y(n_2605)
);

INVx4_ASAP7_75t_L g2606 ( 
.A(n_2405),
.Y(n_2606)
);

OR2x2_ASAP7_75t_L g2607 ( 
.A(n_2355),
.B(n_390),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2344),
.Y(n_2608)
);

OA21x2_ASAP7_75t_L g2609 ( 
.A1(n_2351),
.A2(n_391),
.B(n_392),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_2450),
.B(n_391),
.Y(n_2610)
);

AND2x2_ASAP7_75t_L g2611 ( 
.A(n_2473),
.B(n_392),
.Y(n_2611)
);

AND2x2_ASAP7_75t_L g2612 ( 
.A(n_2475),
.B(n_393),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2352),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_L g2614 ( 
.A(n_2454),
.B(n_394),
.Y(n_2614)
);

OR2x2_ASAP7_75t_L g2615 ( 
.A(n_2366),
.B(n_394),
.Y(n_2615)
);

INVx1_ASAP7_75t_SL g2616 ( 
.A(n_2485),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2354),
.Y(n_2617)
);

INVx1_ASAP7_75t_SL g2618 ( 
.A(n_2489),
.Y(n_2618)
);

NAND2x1p5_ASAP7_75t_L g2619 ( 
.A(n_2362),
.B(n_2492),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2368),
.Y(n_2620)
);

BUFx2_ASAP7_75t_L g2621 ( 
.A(n_2463),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2549),
.Y(n_2622)
);

INVx1_ASAP7_75t_SL g2623 ( 
.A(n_2506),
.Y(n_2623)
);

AOI221xp5_ASAP7_75t_L g2624 ( 
.A1(n_2574),
.A2(n_2424),
.B1(n_2446),
.B2(n_2435),
.C(n_2386),
.Y(n_2624)
);

OAI21xp33_ASAP7_75t_SL g2625 ( 
.A1(n_2526),
.A2(n_2474),
.B(n_2461),
.Y(n_2625)
);

OAI221xp5_ASAP7_75t_L g2626 ( 
.A1(n_2507),
.A2(n_2348),
.B1(n_2483),
.B2(n_2491),
.C(n_2490),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_2606),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_L g2628 ( 
.A(n_2559),
.B(n_2493),
.Y(n_2628)
);

HB1xp67_ASAP7_75t_L g2629 ( 
.A(n_2512),
.Y(n_2629)
);

O2A1O1Ixp33_ASAP7_75t_L g2630 ( 
.A1(n_2547),
.A2(n_2488),
.B(n_2472),
.C(n_2357),
.Y(n_2630)
);

AOI222xp33_ASAP7_75t_L g2631 ( 
.A1(n_2557),
.A2(n_2380),
.B1(n_2364),
.B2(n_2342),
.C1(n_2365),
.C2(n_2414),
.Y(n_2631)
);

OAI21xp5_ASAP7_75t_L g2632 ( 
.A1(n_2508),
.A2(n_2398),
.B(n_2349),
.Y(n_2632)
);

INVxp67_ASAP7_75t_SL g2633 ( 
.A(n_2510),
.Y(n_2633)
);

A2O1A1Ixp33_ASAP7_75t_L g2634 ( 
.A1(n_2516),
.A2(n_2371),
.B(n_2412),
.C(n_2413),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2579),
.Y(n_2635)
);

OAI211xp5_ASAP7_75t_SL g2636 ( 
.A1(n_2513),
.A2(n_2383),
.B(n_2397),
.C(n_2438),
.Y(n_2636)
);

OAI322xp33_ASAP7_75t_L g2637 ( 
.A1(n_2500),
.A2(n_2378),
.A3(n_2427),
.B1(n_2415),
.B2(n_2430),
.C1(n_2428),
.C2(n_2387),
.Y(n_2637)
);

AO21x1_ASAP7_75t_L g2638 ( 
.A1(n_2540),
.A2(n_2423),
.B(n_2431),
.Y(n_2638)
);

AOI221xp5_ASAP7_75t_L g2639 ( 
.A1(n_2518),
.A2(n_2419),
.B1(n_2411),
.B2(n_397),
.C(n_395),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2511),
.Y(n_2640)
);

A2O1A1Ixp33_ASAP7_75t_L g2641 ( 
.A1(n_2535),
.A2(n_398),
.B(n_396),
.C(n_397),
.Y(n_2641)
);

OR2x2_ASAP7_75t_L g2642 ( 
.A(n_2542),
.B(n_2621),
.Y(n_2642)
);

NAND2x1_ASAP7_75t_L g2643 ( 
.A(n_2603),
.B(n_396),
.Y(n_2643)
);

HB1xp67_ASAP7_75t_L g2644 ( 
.A(n_2594),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2514),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2533),
.Y(n_2646)
);

OR2x6_ASAP7_75t_L g2647 ( 
.A(n_2575),
.B(n_398),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2537),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2550),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2555),
.Y(n_2650)
);

AND2x4_ASAP7_75t_L g2651 ( 
.A(n_2604),
.B(n_399),
.Y(n_2651)
);

AOI22xp5_ASAP7_75t_L g2652 ( 
.A1(n_2505),
.A2(n_402),
.B1(n_400),
.B2(n_401),
.Y(n_2652)
);

AND2x2_ASAP7_75t_L g2653 ( 
.A(n_2570),
.B(n_400),
.Y(n_2653)
);

AND2x2_ASAP7_75t_L g2654 ( 
.A(n_2528),
.B(n_401),
.Y(n_2654)
);

AOI21xp33_ASAP7_75t_SL g2655 ( 
.A1(n_2619),
.A2(n_402),
.B(n_403),
.Y(n_2655)
);

NAND4xp25_ASAP7_75t_L g2656 ( 
.A(n_2532),
.B(n_405),
.C(n_403),
.D(n_404),
.Y(n_2656)
);

NAND2x1p5_ASAP7_75t_L g2657 ( 
.A(n_2504),
.B(n_406),
.Y(n_2657)
);

INVx3_ASAP7_75t_L g2658 ( 
.A(n_2536),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2558),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_L g2660 ( 
.A(n_2616),
.B(n_406),
.Y(n_2660)
);

AOI22xp5_ASAP7_75t_L g2661 ( 
.A1(n_2529),
.A2(n_409),
.B1(n_407),
.B2(n_408),
.Y(n_2661)
);

OAI221xp5_ASAP7_75t_L g2662 ( 
.A1(n_2534),
.A2(n_412),
.B1(n_408),
.B2(n_410),
.C(n_413),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2501),
.Y(n_2663)
);

A2O1A1Ixp33_ASAP7_75t_L g2664 ( 
.A1(n_2585),
.A2(n_414),
.B(n_410),
.C(n_412),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2560),
.Y(n_2665)
);

AOI22xp5_ASAP7_75t_L g2666 ( 
.A1(n_2530),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.Y(n_2666)
);

OAI211xp5_ASAP7_75t_L g2667 ( 
.A1(n_2580),
.A2(n_419),
.B(n_415),
.C(n_418),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2564),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_L g2669 ( 
.A(n_2618),
.B(n_418),
.Y(n_2669)
);

INVxp67_ASAP7_75t_L g2670 ( 
.A(n_2589),
.Y(n_2670)
);

INVx1_ASAP7_75t_SL g2671 ( 
.A(n_2605),
.Y(n_2671)
);

OAI21xp5_ASAP7_75t_SL g2672 ( 
.A1(n_2562),
.A2(n_419),
.B(n_420),
.Y(n_2672)
);

NOR2x1_ASAP7_75t_L g2673 ( 
.A(n_2523),
.B(n_420),
.Y(n_2673)
);

OR2x2_ASAP7_75t_L g2674 ( 
.A(n_2520),
.B(n_421),
.Y(n_2674)
);

AND2x2_ASAP7_75t_L g2675 ( 
.A(n_2546),
.B(n_421),
.Y(n_2675)
);

AND2x2_ASAP7_75t_L g2676 ( 
.A(n_2551),
.B(n_422),
.Y(n_2676)
);

AND2x2_ASAP7_75t_L g2677 ( 
.A(n_2603),
.B(n_422),
.Y(n_2677)
);

A2O1A1Ixp33_ASAP7_75t_L g2678 ( 
.A1(n_2539),
.A2(n_425),
.B(n_423),
.C(n_424),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2565),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2568),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_SL g2681 ( 
.A(n_2552),
.B(n_2503),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_L g2682 ( 
.A(n_2536),
.B(n_423),
.Y(n_2682)
);

AOI21xp5_ASAP7_75t_L g2683 ( 
.A1(n_2633),
.A2(n_2576),
.B(n_2582),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2644),
.Y(n_2684)
);

AO22x2_ASAP7_75t_L g2685 ( 
.A1(n_2670),
.A2(n_2509),
.B1(n_2593),
.B2(n_2586),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2629),
.Y(n_2686)
);

NOR2x1_ASAP7_75t_L g2687 ( 
.A(n_2643),
.B(n_2609),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2642),
.Y(n_2688)
);

A2O1A1Ixp33_ASAP7_75t_SL g2689 ( 
.A1(n_2662),
.A2(n_2588),
.B(n_2515),
.C(n_2527),
.Y(n_2689)
);

AOI31xp33_ASAP7_75t_L g2690 ( 
.A1(n_2673),
.A2(n_2577),
.A3(n_2499),
.B(n_2531),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2622),
.Y(n_2691)
);

O2A1O1Ixp5_ASAP7_75t_L g2692 ( 
.A1(n_2667),
.A2(n_2620),
.B(n_2608),
.C(n_2613),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2635),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2640),
.Y(n_2694)
);

AOI22xp5_ASAP7_75t_L g2695 ( 
.A1(n_2623),
.A2(n_2609),
.B1(n_2578),
.B2(n_2617),
.Y(n_2695)
);

AOI21xp33_ASAP7_75t_SL g2696 ( 
.A1(n_2657),
.A2(n_2553),
.B(n_2573),
.Y(n_2696)
);

OAI221xp5_ASAP7_75t_SL g2697 ( 
.A1(n_2672),
.A2(n_2614),
.B1(n_2610),
.B2(n_2601),
.C(n_2525),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2645),
.Y(n_2698)
);

OAI22xp5_ASAP7_75t_L g2699 ( 
.A1(n_2664),
.A2(n_2519),
.B1(n_2583),
.B2(n_2554),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2646),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2648),
.Y(n_2701)
);

OAI21xp5_ASAP7_75t_L g2702 ( 
.A1(n_2625),
.A2(n_2545),
.B(n_2581),
.Y(n_2702)
);

NOR3xp33_ASAP7_75t_L g2703 ( 
.A(n_2628),
.B(n_2627),
.C(n_2681),
.Y(n_2703)
);

NOR2xp33_ASAP7_75t_L g2704 ( 
.A(n_2637),
.B(n_2569),
.Y(n_2704)
);

AOI321xp33_ASAP7_75t_L g2705 ( 
.A1(n_2624),
.A2(n_2502),
.A3(n_2602),
.B1(n_2538),
.B2(n_2600),
.C(n_2599),
.Y(n_2705)
);

AOI222xp33_ASAP7_75t_L g2706 ( 
.A1(n_2639),
.A2(n_2541),
.B1(n_2612),
.B2(n_2611),
.C1(n_2596),
.C2(n_2598),
.Y(n_2706)
);

OAI22xp5_ASAP7_75t_L g2707 ( 
.A1(n_2626),
.A2(n_2590),
.B1(n_2591),
.B2(n_2587),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2658),
.B(n_2548),
.Y(n_2708)
);

INVx3_ASAP7_75t_SL g2709 ( 
.A(n_2651),
.Y(n_2709)
);

OAI221xp5_ASAP7_75t_L g2710 ( 
.A1(n_2671),
.A2(n_2572),
.B1(n_2584),
.B2(n_2571),
.C(n_2556),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2649),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_L g2712 ( 
.A(n_2677),
.B(n_2561),
.Y(n_2712)
);

OR2x2_ASAP7_75t_L g2713 ( 
.A(n_2663),
.B(n_2566),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2650),
.Y(n_2714)
);

OAI322xp33_ASAP7_75t_L g2715 ( 
.A1(n_2659),
.A2(n_2615),
.A3(n_2607),
.B1(n_2567),
.B2(n_2595),
.C1(n_2592),
.C2(n_2544),
.Y(n_2715)
);

AOI22xp33_ASAP7_75t_L g2716 ( 
.A1(n_2638),
.A2(n_2522),
.B1(n_2521),
.B2(n_2543),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2709),
.B(n_2653),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2684),
.Y(n_2718)
);

AND2x2_ASAP7_75t_L g2719 ( 
.A(n_2688),
.B(n_2632),
.Y(n_2719)
);

INVx2_ASAP7_75t_L g2720 ( 
.A(n_2686),
.Y(n_2720)
);

NOR2xp67_ASAP7_75t_L g2721 ( 
.A(n_2696),
.B(n_2674),
.Y(n_2721)
);

OAI21xp5_ASAP7_75t_L g2722 ( 
.A1(n_2687),
.A2(n_2641),
.B(n_2655),
.Y(n_2722)
);

OAI22xp5_ASAP7_75t_L g2723 ( 
.A1(n_2690),
.A2(n_2647),
.B1(n_2666),
.B2(n_2661),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2713),
.Y(n_2724)
);

XNOR2xp5_ASAP7_75t_L g2725 ( 
.A(n_2716),
.B(n_2656),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_2703),
.B(n_2704),
.Y(n_2726)
);

O2A1O1Ixp33_ASAP7_75t_L g2727 ( 
.A1(n_2683),
.A2(n_2689),
.B(n_2692),
.C(n_2702),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2691),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2693),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2685),
.Y(n_2730)
);

XNOR2xp5_ASAP7_75t_L g2731 ( 
.A(n_2707),
.B(n_2699),
.Y(n_2731)
);

OAI22xp5_ASAP7_75t_L g2732 ( 
.A1(n_2695),
.A2(n_2647),
.B1(n_2678),
.B2(n_2652),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_2706),
.B(n_2634),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2685),
.B(n_2631),
.Y(n_2734)
);

NOR2xp67_ASAP7_75t_L g2735 ( 
.A(n_2710),
.B(n_2665),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2724),
.Y(n_2736)
);

AOI21xp5_ASAP7_75t_L g2737 ( 
.A1(n_2727),
.A2(n_2726),
.B(n_2734),
.Y(n_2737)
);

AOI22xp5_ASAP7_75t_L g2738 ( 
.A1(n_2723),
.A2(n_2708),
.B1(n_2712),
.B2(n_2636),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_2721),
.B(n_2654),
.Y(n_2739)
);

OAI21x1_ASAP7_75t_L g2740 ( 
.A1(n_2730),
.A2(n_2722),
.B(n_2717),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2719),
.B(n_2630),
.Y(n_2741)
);

NOR4xp25_ASAP7_75t_L g2742 ( 
.A(n_2733),
.B(n_2705),
.C(n_2698),
.D(n_2700),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_SL g2743 ( 
.A(n_2732),
.B(n_2597),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2718),
.Y(n_2744)
);

AOI221xp5_ASAP7_75t_L g2745 ( 
.A1(n_2742),
.A2(n_2731),
.B1(n_2725),
.B2(n_2720),
.C(n_2729),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2737),
.B(n_2735),
.Y(n_2746)
);

AOI21xp33_ASAP7_75t_L g2747 ( 
.A1(n_2739),
.A2(n_2728),
.B(n_2701),
.Y(n_2747)
);

AOI211xp5_ASAP7_75t_SL g2748 ( 
.A1(n_2741),
.A2(n_2711),
.B(n_2714),
.C(n_2694),
.Y(n_2748)
);

AOI22xp5_ASAP7_75t_L g2749 ( 
.A1(n_2743),
.A2(n_2679),
.B1(n_2680),
.B2(n_2668),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2736),
.Y(n_2750)
);

A2O1A1Ixp33_ASAP7_75t_L g2751 ( 
.A1(n_2740),
.A2(n_2697),
.B(n_2669),
.C(n_2660),
.Y(n_2751)
);

AOI211xp5_ASAP7_75t_L g2752 ( 
.A1(n_2738),
.A2(n_2744),
.B(n_2715),
.C(n_2682),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2750),
.Y(n_2753)
);

NAND4xp75_ASAP7_75t_L g2754 ( 
.A(n_2746),
.B(n_2676),
.C(n_2675),
.D(n_2563),
.Y(n_2754)
);

AOI222xp33_ASAP7_75t_L g2755 ( 
.A1(n_2745),
.A2(n_2524),
.B1(n_2517),
.B2(n_2498),
.C1(n_428),
.C2(n_429),
.Y(n_2755)
);

OAI211xp5_ASAP7_75t_L g2756 ( 
.A1(n_2752),
.A2(n_427),
.B(n_424),
.C(n_426),
.Y(n_2756)
);

OAI211xp5_ASAP7_75t_SL g2757 ( 
.A1(n_2751),
.A2(n_430),
.B(n_428),
.C(n_429),
.Y(n_2757)
);

XNOR2xp5_ASAP7_75t_L g2758 ( 
.A(n_2754),
.B(n_2749),
.Y(n_2758)
);

HB1xp67_ASAP7_75t_L g2759 ( 
.A(n_2753),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2759),
.B(n_2755),
.Y(n_2760)
);

AOI22xp5_ASAP7_75t_L g2761 ( 
.A1(n_2760),
.A2(n_2756),
.B1(n_2757),
.B2(n_2758),
.Y(n_2761)
);

HB1xp67_ASAP7_75t_L g2762 ( 
.A(n_2761),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2762),
.Y(n_2763)
);

AOI21xp5_ASAP7_75t_SL g2764 ( 
.A1(n_2762),
.A2(n_2748),
.B(n_2747),
.Y(n_2764)
);

HB1xp67_ASAP7_75t_L g2765 ( 
.A(n_2763),
.Y(n_2765)
);

AOI22xp33_ASAP7_75t_L g2766 ( 
.A1(n_2764),
.A2(n_433),
.B1(n_430),
.B2(n_431),
.Y(n_2766)
);

INVxp67_ASAP7_75t_L g2767 ( 
.A(n_2765),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_L g2768 ( 
.A(n_2767),
.B(n_2766),
.Y(n_2768)
);

OAI222xp33_ASAP7_75t_SL g2769 ( 
.A1(n_2768),
.A2(n_433),
.B1(n_434),
.B2(n_435),
.C1(n_436),
.C2(n_437),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_SL g2770 ( 
.A(n_2768),
.B(n_435),
.Y(n_2770)
);

OAI22xp33_ASAP7_75t_L g2771 ( 
.A1(n_2770),
.A2(n_439),
.B1(n_437),
.B2(n_438),
.Y(n_2771)
);

XNOR2xp5_ASAP7_75t_L g2772 ( 
.A(n_2769),
.B(n_438),
.Y(n_2772)
);

AOI221xp5_ASAP7_75t_L g2773 ( 
.A1(n_2772),
.A2(n_441),
.B1(n_439),
.B2(n_440),
.C(n_442),
.Y(n_2773)
);

AOI211xp5_ASAP7_75t_L g2774 ( 
.A1(n_2773),
.A2(n_2771),
.B(n_442),
.C(n_440),
.Y(n_2774)
);


endmodule