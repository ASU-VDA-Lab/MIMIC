module real_jpeg_25431_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_2),
.B(n_47),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_2),
.B(n_67),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_2),
.B(n_49),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_2),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_2),
.B(n_33),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_2),
.B(n_27),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx8_ASAP7_75t_SL g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_5),
.B(n_43),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_5),
.B(n_47),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_5),
.B(n_67),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_5),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_5),
.B(n_33),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_5),
.B(n_52),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_5),
.B(n_49),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_6),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_6),
.B(n_27),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_6),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_6),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_6),
.B(n_33),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_6),
.B(n_52),
.Y(n_277)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVxp33_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_8),
.B(n_43),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_8),
.B(n_33),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_8),
.B(n_52),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_8),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_8),
.B(n_49),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_8),
.B(n_47),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_8),
.B(n_67),
.Y(n_292)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_10),
.B(n_47),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_10),
.B(n_67),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_10),
.B(n_17),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_10),
.B(n_33),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_10),
.B(n_52),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_11),
.B(n_43),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_11),
.B(n_49),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_11),
.B(n_47),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_11),
.B(n_52),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_11),
.B(n_33),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_11),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_11),
.B(n_67),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_11),
.B(n_27),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_12),
.B(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_12),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_12),
.B(n_49),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_12),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_12),
.B(n_47),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_13),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_13),
.B(n_47),
.Y(n_86)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_13),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_13),
.B(n_52),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_13),
.B(n_67),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_13),
.B(n_269),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_15),
.B(n_52),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_16),
.B(n_27),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_16),
.B(n_52),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_16),
.B(n_49),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_16),
.B(n_33),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_16),
.B(n_17),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_16),
.B(n_47),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_16),
.B(n_67),
.Y(n_270)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_17),
.Y(n_112)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_17),
.Y(n_172)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_17),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_146),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_116),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_77),
.C(n_89),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_21),
.B(n_77),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_54),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_22),
.B(n_55),
.C(n_71),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.C(n_45),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_23),
.B(n_322),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_24),
.B(n_30),
.C(n_37),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_26),
.B(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_26),
.B(n_61),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_30),
.A2(n_38),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_SL g130 ( 
.A(n_30),
.B(n_79),
.C(n_82),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_31),
.B(n_62),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_32),
.B(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_35),
.A2(n_37),
.B1(n_40),
.B2(n_101),
.Y(n_100)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_36),
.Y(n_181)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_36),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_40),
.C(n_41),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_39),
.B(n_45),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_40),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_41),
.A2(n_42),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g274 ( 
.A(n_43),
.Y(n_274)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_44),
.Y(n_140)
);

BUFx24_ASAP7_75t_SL g330 ( 
.A(n_45),
.Y(n_330)
);

FAx1_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_48),
.CI(n_51),
.CON(n_45),
.SN(n_45)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_48),
.C(n_51),
.Y(n_84)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx13_ASAP7_75t_L g213 ( 
.A(n_52),
.Y(n_213)
);

BUFx24_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_71),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_66),
.C(n_70),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_56),
.A2(n_57),
.B1(n_103),
.B2(n_105),
.Y(n_102)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_60),
.C(n_63),
.Y(n_57)
);

FAx1_ASAP7_75t_SL g91 ( 
.A(n_58),
.B(n_60),
.CI(n_63),
.CON(n_91),
.SN(n_91)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_64),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_66),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_66),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_66),
.A2(n_70),
.B1(n_75),
.B2(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_66),
.B(n_74),
.C(n_76),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_70),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_76),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_73),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_83),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_78),
.B(n_84),
.C(n_85),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_81),
.A2(n_82),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_85),
.Y(n_328)
);

FAx1_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_87),
.CI(n_88),
.CON(n_85),
.SN(n_85)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_86),
.B(n_87),
.C(n_88),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_89),
.B(n_327),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_102),
.C(n_106),
.Y(n_89)
);

FAx1_ASAP7_75t_SL g323 ( 
.A(n_90),
.B(n_102),
.CI(n_106),
.CON(n_323),
.SN(n_323)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.C(n_98),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_91),
.B(n_307),
.Y(n_306)
);

BUFx24_ASAP7_75t_SL g331 ( 
.A(n_91),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_92),
.B(n_98),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.C(n_96),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_95),
.B(n_287),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_103),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_114),
.C(n_115),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_107),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_107),
.B(n_313),
.Y(n_312)
);

FAx1_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_110),
.CI(n_113),
.CON(n_107),
.SN(n_107)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_114),
.B(n_115),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_131),
.B2(n_132),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_127),
.B2(n_128),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_125),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_144),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_325),
.C(n_326),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_316),
.C(n_317),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_302),
.C(n_303),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_280),
.C(n_281),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_248),
.C(n_249),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_223),
.C(n_224),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_183),
.C(n_195),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_167),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_162),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_155),
.B(n_162),
.C(n_167),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_160),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_156),
.A2(n_157),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_186)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_163),
.B(n_165),
.C(n_166),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_175),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_168),
.B(n_176),
.C(n_177),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_173),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_169),
.A2(n_170),
.B1(n_173),
.B2(n_174),
.Y(n_194)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_172),
.Y(n_269)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_182),
.Y(n_177)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_178),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_179),
.B(n_182),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.C(n_194),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_187),
.A2(n_188),
.B1(n_194),
.B2(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_199)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_194),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_219),
.C(n_220),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_204),
.C(n_209),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_202),
.C(n_203),
.Y(n_219)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_205),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.C(n_214),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_212),
.B(n_274),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_237),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_238),
.C(n_247),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_233),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_232),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_232),
.C(n_233),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_228),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_231),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx24_ASAP7_75t_SL g332 ( 
.A(n_233),
.Y(n_332)
);

FAx1_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_235),
.CI(n_236),
.CON(n_233),
.SN(n_233)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_235),
.C(n_236),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_247),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_245),
.B2(n_246),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_241),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_244),
.C(n_246),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_245),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_264),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_252),
.B(n_253),
.C(n_264),
.Y(n_280)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_259),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_260),
.C(n_263),
.Y(n_284)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_255),
.Y(n_333)
);

FAx1_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_257),
.CI(n_258),
.CON(n_255),
.SN(n_255)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_256),
.B(n_257),
.C(n_258),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_265),
.B(n_272),
.C(n_278),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_272),
.B1(n_278),
.B2(n_279),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_267),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_270),
.B(n_271),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_268),
.B(n_270),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_271),
.B(n_299),
.C(n_300),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_272),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_275),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_276),
.C(n_277),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_295),
.B2(n_301),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_296),
.C(n_297),
.Y(n_302)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_286),
.C(n_288),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_288),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_294),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_290),
.B(n_293),
.C(n_294),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_292),
.Y(n_293)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_295),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_300),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_314),
.B2(n_315),
.Y(n_303)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_304),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_305),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_308),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_308),
.C(n_314),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_311),
.C(n_312),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_320),
.C(n_324),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_321),
.B1(n_323),
.B2(n_324),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_323),
.Y(n_324)
);

BUFx24_ASAP7_75t_SL g334 ( 
.A(n_323),
.Y(n_334)
);


endmodule