module fake_jpeg_9260_n_46 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_46);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_46;

wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_40;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_37;
wire n_29;
wire n_43;
wire n_32;

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_20),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_8),
.B(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_34),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_26),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_35),
.B(n_37),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_0),
.B(n_22),
.Y(n_36)
);

MAJx2_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_38),
.C(n_3),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_31),
.A2(n_32),
.B1(n_23),
.B2(n_29),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_1),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_41),
.A2(n_37),
.B(n_25),
.Y(n_42)
);

OAI322xp33_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_39),
.A3(n_40),
.B1(n_10),
.B2(n_11),
.C1(n_13),
.C2(n_6),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_21),
.B1(n_16),
.B2(n_18),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

NAND3xp33_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_7),
.C(n_19),
.Y(n_46)
);


endmodule