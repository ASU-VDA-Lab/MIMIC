module fake_aes_4038_n_43 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_10, n_8, n_0, n_43);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_10;
input n_8;
input n_0;
output n_43;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_25;
wire n_30;
wire n_26;
wire n_16;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
INVx1_ASAP7_75t_L g15 ( .A(n_4), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_6), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_10), .Y(n_17) );
CKINVDCx16_ASAP7_75t_R g18 ( .A(n_11), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_8), .Y(n_19) );
HB1xp67_ASAP7_75t_L g20 ( .A(n_0), .Y(n_20) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_8), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_12), .B(n_7), .Y(n_22) );
HB1xp67_ASAP7_75t_L g23 ( .A(n_20), .Y(n_23) );
HB1xp67_ASAP7_75t_L g24 ( .A(n_21), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_19), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_18), .B(n_0), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
OAI22xp5_ASAP7_75t_L g28 ( .A1(n_23), .A2(n_18), .B1(n_15), .B2(n_19), .Y(n_28) );
AND2x2_ASAP7_75t_L g29 ( .A(n_28), .B(n_24), .Y(n_29) );
NAND2xp5_ASAP7_75t_L g30 ( .A(n_27), .B(n_26), .Y(n_30) );
OR2x2_ASAP7_75t_L g31 ( .A(n_29), .B(n_15), .Y(n_31) );
OR2x2_ASAP7_75t_L g32 ( .A(n_30), .B(n_19), .Y(n_32) );
INVxp67_ASAP7_75t_L g33 ( .A(n_32), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_31), .Y(n_34) );
OAI22xp5_ASAP7_75t_L g35 ( .A1(n_33), .A2(n_16), .B1(n_22), .B2(n_17), .Y(n_35) );
AOI322xp5_ASAP7_75t_L g36 ( .A1(n_34), .A2(n_22), .A3(n_2), .B1(n_3), .B2(n_4), .C1(n_5), .C2(n_1), .Y(n_36) );
AOI221xp5_ASAP7_75t_L g37 ( .A1(n_34), .A2(n_1), .B1(n_2), .B2(n_3), .C(n_5), .Y(n_37) );
OAI221xp5_ASAP7_75t_L g38 ( .A1(n_35), .A2(n_6), .B1(n_7), .B2(n_9), .C(n_13), .Y(n_38) );
INVx1_ASAP7_75t_L g39 ( .A(n_37), .Y(n_39) );
NOR2x1p5_ASAP7_75t_L g40 ( .A(n_36), .B(n_14), .Y(n_40) );
HB1xp67_ASAP7_75t_L g41 ( .A(n_40), .Y(n_41) );
INVx1_ASAP7_75t_SL g42 ( .A(n_39), .Y(n_42) );
AOI22xp33_ASAP7_75t_L g43 ( .A1(n_41), .A2(n_38), .B1(n_39), .B2(n_42), .Y(n_43) );
endmodule