module fake_jpeg_17129_n_294 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_294);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_294;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_SL g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_0),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_24),
.Y(n_40)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_22),
.B(n_29),
.C(n_28),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_42),
.A2(n_27),
.B(n_21),
.Y(n_85)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_18),
.B1(n_19),
.B2(n_22),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_54),
.B1(n_18),
.B2(n_19),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_18),
.B1(n_19),
.B2(n_22),
.Y(n_54)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_15),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_64),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_33),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_83),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_70),
.Y(n_90)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_15),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_65),
.A2(n_40),
.B1(n_16),
.B2(n_21),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_68),
.B(n_69),
.Y(n_106)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_33),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_49),
.A2(n_34),
.B1(n_22),
.B2(n_39),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_71),
.A2(n_37),
.B1(n_36),
.B2(n_21),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_75),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_42),
.B(n_35),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_74),
.B(n_81),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_29),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_76),
.B(n_78),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_49),
.A2(n_40),
.B1(n_39),
.B2(n_41),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_77),
.A2(n_44),
.B1(n_43),
.B2(n_56),
.Y(n_94)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_28),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_84),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_50),
.B(n_35),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_17),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_82),
.B(n_88),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_32),
.C(n_40),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_53),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_16),
.Y(n_98)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_87),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_52),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_59),
.A2(n_52),
.B1(n_56),
.B2(n_44),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_93),
.A2(n_111),
.B1(n_77),
.B2(n_84),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_103),
.B1(n_105),
.B2(n_107),
.Y(n_125)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_99),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_0),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_96),
.A2(n_27),
.B(n_31),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_98),
.B(n_82),
.Y(n_126)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_70),
.A2(n_44),
.B1(n_40),
.B2(n_41),
.Y(n_103)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_110),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_59),
.B(n_32),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_112),
.Y(n_119)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_65),
.A2(n_41),
.B1(n_39),
.B2(n_37),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_32),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_62),
.B(n_24),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_114),
.B(n_106),
.Y(n_130)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_73),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_83),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_118),
.A2(n_123),
.B(n_140),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_136),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_122),
.A2(n_95),
.B1(n_99),
.B2(n_104),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_112),
.A2(n_63),
.B(n_69),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_126),
.B(n_129),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_103),
.A2(n_63),
.B1(n_68),
.B2(n_76),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_134),
.B1(n_97),
.B2(n_109),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_92),
.B(n_31),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_141),
.Y(n_146)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_90),
.B(n_71),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_132),
.B(n_133),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_97),
.A2(n_80),
.B1(n_86),
.B2(n_72),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_80),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_135),
.B(n_37),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_102),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_139),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_138),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_102),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_113),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_92),
.B(n_88),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_108),
.A2(n_78),
.B(n_24),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_144),
.A2(n_36),
.B(n_27),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_147),
.A2(n_167),
.B1(n_122),
.B2(n_137),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_98),
.B(n_90),
.C(n_96),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_148),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_114),
.C(n_111),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_150),
.B(n_151),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_132),
.C(n_119),
.Y(n_151)
);

OAI21x1_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_113),
.B(n_96),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_153),
.A2(n_164),
.B(n_165),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_89),
.C(n_94),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_162),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_107),
.Y(n_155)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_120),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_156),
.B(n_158),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_120),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_161),
.B(n_139),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_24),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_123),
.B(n_30),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_140),
.A2(n_131),
.B(n_124),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_169),
.A2(n_170),
.B(n_173),
.Y(n_190)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_126),
.A2(n_20),
.B(n_23),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_166),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_176),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_157),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_127),
.Y(n_178)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_180),
.A2(n_189),
.B1(n_195),
.B2(n_200),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_163),
.B(n_129),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_181),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_128),
.Y(n_182)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

A2O1A1Ixp33_ASAP7_75t_SL g185 ( 
.A1(n_167),
.A2(n_125),
.B(n_115),
.C(n_110),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_185),
.A2(n_198),
.B1(n_179),
.B2(n_184),
.Y(n_206)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_186),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_133),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_188),
.B(n_199),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_160),
.A2(n_125),
.B1(n_101),
.B2(n_67),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_173),
.B(n_146),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_193),
.A2(n_197),
.B1(n_201),
.B2(n_188),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_194),
.A2(n_162),
.B1(n_145),
.B2(n_0),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_154),
.A2(n_101),
.B1(n_23),
.B2(n_17),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_101),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_152),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_26),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_159),
.A2(n_20),
.B1(n_26),
.B2(n_30),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_159),
.B(n_8),
.Y(n_201)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_151),
.C(n_164),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_210),
.C(n_219),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_150),
.C(n_149),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_196),
.B(n_145),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_221),
.Y(n_227)
);

OR2x6_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_165),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_198),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_180),
.A2(n_155),
.B1(n_149),
.B2(n_148),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_214),
.A2(n_216),
.B1(n_190),
.B2(n_199),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_194),
.A2(n_30),
.B1(n_2),
.B2(n_3),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_218),
.A2(n_200),
.B(n_190),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_1),
.C(n_2),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_220),
.B(n_195),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_1),
.C(n_2),
.Y(n_221)
);

BUFx24_ASAP7_75t_SL g222 ( 
.A(n_202),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_224),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_204),
.A2(n_174),
.B1(n_192),
.B2(n_185),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_223),
.A2(n_225),
.B1(n_226),
.B2(n_234),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_212),
.Y(n_224)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_196),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_211),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_175),
.Y(n_232)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_215),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_236),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_213),
.A2(n_174),
.B1(n_185),
.B2(n_179),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_235),
.A2(n_218),
.B1(n_185),
.B2(n_189),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_209),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_206),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_205),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_221),
.B(n_177),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_238),
.B(n_239),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_219),
.B(n_186),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_235),
.A2(n_217),
.B(n_213),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_240),
.A2(n_3),
.B(n_4),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_210),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_242),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_208),
.Y(n_242)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_247),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_248),
.B(n_14),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_229),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_208),
.C(n_213),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_254),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_213),
.Y(n_253)
);

BUFx24_ASAP7_75t_SL g259 ( 
.A(n_253),
.Y(n_259)
);

INVxp33_ASAP7_75t_L g256 ( 
.A(n_245),
.Y(n_256)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_244),
.A2(n_225),
.B1(n_223),
.B2(n_234),
.Y(n_257)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_257),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_261),
.Y(n_269)
);

NAND3xp33_ASAP7_75t_SL g262 ( 
.A(n_249),
.B(n_3),
.C(n_5),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_263),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_7),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_252),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_255),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_10),
.Y(n_279)
);

BUFx24_ASAP7_75t_SL g267 ( 
.A(n_265),
.Y(n_267)
);

BUFx24_ASAP7_75t_SL g282 ( 
.A(n_267),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_272),
.B(n_253),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_260),
.C(n_251),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_242),
.C(n_248),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_243),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_11),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_275),
.A2(n_276),
.B1(n_280),
.B2(n_281),
.Y(n_283)
);

NOR2xp67_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_241),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_278),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_8),
.C(n_9),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_279),
.A2(n_268),
.B1(n_12),
.B2(n_13),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_10),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_285),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_282),
.A2(n_270),
.B(n_12),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_11),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_286),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_13),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_289),
.A2(n_13),
.B(n_14),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_292),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_287),
.C(n_286),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_290),
.Y(n_294)
);


endmodule