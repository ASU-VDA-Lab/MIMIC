module fake_jpeg_27168_n_198 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_198);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_198;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_15),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_40),
.Y(n_49)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_1),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_42),
.B(n_30),
.Y(n_69)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_53),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_21),
.B1(n_28),
.B2(n_25),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_48),
.A2(n_31),
.B1(n_35),
.B2(n_34),
.Y(n_61)
);

AND2x2_ASAP7_75t_SL g50 ( 
.A(n_33),
.B(n_28),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_36),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_19),
.B1(n_20),
.B2(n_27),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_32),
.A2(n_20),
.B1(n_22),
.B2(n_27),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_52),
.A2(n_23),
.B1(n_30),
.B2(n_29),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_22),
.B1(n_23),
.B2(n_26),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_56),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_58),
.B(n_65),
.Y(n_80)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_66),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_32),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_70),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_79),
.B1(n_41),
.B2(n_54),
.Y(n_82)
);

AOI211xp5_ASAP7_75t_SL g64 ( 
.A1(n_50),
.A2(n_38),
.B(n_40),
.C(n_24),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_64),
.A2(n_45),
.B1(n_55),
.B2(n_18),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_26),
.Y(n_66)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_76),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_49),
.B(n_30),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_71),
.B(n_74),
.Y(n_101)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_75),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_25),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_25),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_47),
.B(n_29),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_77),
.Y(n_94)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_54),
.A2(n_31),
.B1(n_35),
.B2(n_34),
.Y(n_79)
);

MAJx2_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_35),
.C(n_36),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_71),
.C(n_64),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_82),
.A2(n_83),
.B1(n_92),
.B2(n_95),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_46),
.B1(n_55),
.B2(n_41),
.Y(n_83)
);

NAND3xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_14),
.C(n_2),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_87),
.B(n_91),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_88),
.B(n_24),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_67),
.A2(n_45),
.B1(n_28),
.B2(n_25),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_93),
.B(n_100),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_73),
.A2(n_45),
.B1(n_43),
.B2(n_36),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_74),
.A2(n_43),
.B1(n_18),
.B2(n_24),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_61),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_78),
.B(n_43),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_75),
.B(n_79),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_24),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_58),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_110),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_107),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_105),
.A2(n_113),
.B(n_82),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_106),
.B(n_108),
.Y(n_122)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_80),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_115),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_116),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_70),
.C(n_62),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_99),
.B(n_94),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_118),
.B(n_121),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_62),
.Y(n_119)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_72),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_120),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_99),
.B(n_28),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_105),
.A2(n_88),
.B(n_101),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_128),
.Y(n_140)
);

NOR2x1_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_99),
.Y(n_128)
);

NOR4xp25_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_119),
.C(n_101),
.D(n_110),
.Y(n_129)
);

NAND3xp33_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_132),
.C(n_115),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_133),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_86),
.B(n_81),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_116),
.B(n_94),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_139),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_114),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_124),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_108),
.A2(n_98),
.B(n_86),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_138),
.A2(n_98),
.B(n_96),
.Y(n_150)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_125),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_141),
.B(n_148),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_135),
.A2(n_107),
.B1(n_95),
.B2(n_68),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_145),
.B1(n_151),
.B2(n_154),
.Y(n_162)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_153),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_106),
.B1(n_111),
.B2(n_112),
.Y(n_145)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_146),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_126),
.A2(n_111),
.B1(n_98),
.B2(n_109),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_149),
.A2(n_139),
.B1(n_136),
.B2(n_17),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_150),
.A2(n_103),
.B(n_53),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_17),
.B1(n_68),
.B2(n_102),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_137),
.B(n_17),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_127),
.Y(n_157)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_126),
.B1(n_130),
.B2(n_131),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_160),
.Y(n_173)
);

NOR2x1_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_130),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_163),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_143),
.B(n_123),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_159),
.B(n_153),
.Y(n_172)
);

AOI221xp5_ASAP7_75t_L g160 ( 
.A1(n_140),
.A2(n_137),
.B1(n_129),
.B2(n_136),
.C(n_133),
.Y(n_160)
);

BUFx12_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_164),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_165),
.A2(n_150),
.B(n_144),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_1),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_149),
.C(n_147),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_169),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_147),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_171),
.B(n_172),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_161),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_174),
.A2(n_156),
.B(n_155),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_2),
.C(n_3),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_166),
.C(n_163),
.Y(n_176)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_176),
.Y(n_184)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_177),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_167),
.A2(n_158),
.B1(n_162),
.B2(n_164),
.Y(n_178)
);

AOI322xp5_ASAP7_75t_L g187 ( 
.A1(n_178),
.A2(n_181),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_157),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_170),
.A2(n_165),
.B1(n_164),
.B2(n_4),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_182),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_186)
);

AOI31xp67_ASAP7_75t_SL g185 ( 
.A1(n_180),
.A2(n_175),
.A3(n_168),
.B(n_173),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_185),
.B(n_186),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_187),
.A2(n_5),
.B(n_7),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_188),
.A2(n_10),
.B(n_11),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_183),
.A2(n_176),
.B(n_179),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_189),
.A2(n_8),
.B(n_10),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_182),
.Y(n_190)
);

AOI31xp33_ASAP7_75t_L g192 ( 
.A1(n_190),
.A2(n_184),
.A3(n_181),
.B(n_11),
.Y(n_192)
);

NAND2xp33_ASAP7_75t_R g195 ( 
.A(n_192),
.B(n_191),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_194),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_195),
.B(n_10),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_196),
.Y(n_198)
);


endmodule