module fake_jpeg_24798_n_299 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_299);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_299;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_282;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_1),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_8),
.B(n_2),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_32),
.Y(n_49)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_42),
.B(n_46),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_39),
.B(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_44),
.B(n_50),
.Y(n_71)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_55),
.Y(n_75)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_33),
.A2(n_31),
.B1(n_32),
.B2(n_23),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_34),
.B1(n_35),
.B2(n_39),
.Y(n_70)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_34),
.Y(n_80)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_61),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx24_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_33),
.B1(n_35),
.B2(n_31),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_62),
.A2(n_23),
.B1(n_17),
.B2(n_30),
.Y(n_100)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_69),
.Y(n_99)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_65),
.B(n_66),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_47),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_33),
.B1(n_35),
.B2(n_40),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_67),
.A2(n_34),
.B1(n_39),
.B2(n_37),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_18),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_73),
.Y(n_91)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_70),
.A2(n_16),
.B1(n_29),
.B2(n_24),
.Y(n_110)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_74),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_40),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_76),
.Y(n_105)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_78),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_56),
.A2(n_28),
.B1(n_23),
.B2(n_32),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_40),
.Y(n_82)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_40),
.Y(n_83)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_84),
.Y(n_112)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_86),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_44),
.B(n_25),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_90),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_61),
.A2(n_32),
.B(n_23),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_93),
.A2(n_111),
.B(n_27),
.Y(n_136)
);

FAx1_ASAP7_75t_SL g96 ( 
.A(n_68),
.B(n_71),
.CI(n_73),
.CON(n_96),
.SN(n_96)
);

MAJx2_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_64),
.C(n_38),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_32),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_79),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_100),
.A2(n_101),
.B1(n_108),
.B2(n_81),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_66),
.A2(n_17),
.B1(n_30),
.B2(n_39),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_65),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_59),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_67),
.A2(n_30),
.B1(n_17),
.B2(n_38),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_110),
.A2(n_29),
.B1(n_25),
.B2(n_21),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_16),
.B(n_24),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_75),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_113),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_115),
.B(n_122),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_59),
.C(n_60),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_128),
.C(n_88),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_101),
.Y(n_149)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_123),
.B(n_125),
.Y(n_165)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_126),
.A2(n_133),
.B(n_21),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_95),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_127),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_77),
.C(n_69),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_74),
.Y(n_129)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_106),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_130),
.B(n_131),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

NAND3xp33_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_8),
.C(n_1),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_134),
.A2(n_137),
.B(n_140),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_95),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_135),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_139),
.B1(n_27),
.B2(n_101),
.Y(n_146)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_111),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_96),
.B(n_97),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_141),
.A2(n_90),
.B1(n_102),
.B2(n_108),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_143),
.A2(n_154),
.B1(n_161),
.B2(n_26),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_102),
.B(n_96),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_144),
.A2(n_145),
.B(n_164),
.Y(n_176)
);

AO22x1_ASAP7_75t_L g145 ( 
.A1(n_118),
.A2(n_100),
.B1(n_101),
.B2(n_36),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_146),
.A2(n_157),
.B(n_162),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_151),
.C(n_168),
.Y(n_175)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_121),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_141),
.A2(n_88),
.B1(n_114),
.B2(n_107),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_116),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_156),
.Y(n_201)
);

NOR2x1_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_114),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_122),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_107),
.B1(n_57),
.B2(n_63),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_115),
.A2(n_87),
.B(n_89),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_126),
.A2(n_87),
.B(n_89),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_120),
.A2(n_112),
.B(n_105),
.C(n_0),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_167),
.A2(n_84),
.B1(n_26),
.B2(n_22),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_117),
.B(n_38),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_129),
.A2(n_85),
.B(n_0),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_172),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_125),
.B(n_38),
.C(n_36),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_38),
.C(n_36),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_105),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_136),
.A2(n_28),
.B1(n_105),
.B2(n_63),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_174),
.Y(n_180)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_177),
.B(n_182),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_178),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_161),
.B(n_123),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_179),
.B(n_185),
.Y(n_220)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_142),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_138),
.Y(n_183)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_148),
.B(n_72),
.Y(n_186)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_78),
.Y(n_187)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_188),
.A2(n_193),
.B1(n_197),
.B2(n_199),
.Y(n_210)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_145),
.A2(n_164),
.A3(n_147),
.B1(n_149),
.B2(n_167),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_189),
.A2(n_191),
.B(n_150),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_144),
.B(n_36),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_192),
.C(n_172),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_36),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_158),
.B(n_10),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_194),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_170),
.Y(n_195)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_195),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_166),
.B(n_10),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_196),
.Y(n_216)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_153),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_154),
.B(n_173),
.Y(n_198)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_200),
.A2(n_26),
.B1(n_22),
.B2(n_20),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_203),
.A2(n_200),
.B(n_202),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_206),
.C(n_208),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_151),
.C(n_147),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_143),
.C(n_167),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_191),
.A2(n_150),
.B1(n_145),
.B2(n_174),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_209),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_180),
.A2(n_167),
.B1(n_160),
.B2(n_138),
.Y(n_212)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_214),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_180),
.A2(n_76),
.B1(n_22),
.B2(n_0),
.Y(n_217)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_199),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_201),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_220),
.B(n_189),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_224),
.B(n_232),
.Y(n_247)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_211),
.B(n_185),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_231),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_192),
.Y(n_231)
);

MAJx2_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_176),
.C(n_190),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_176),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_239),
.C(n_240),
.Y(n_250)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_235),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_197),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_236),
.A2(n_223),
.B1(n_205),
.B2(n_221),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_215),
.Y(n_237)
);

INVxp33_ASAP7_75t_L g244 ( 
.A(n_237),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_238),
.A2(n_222),
.B1(n_205),
.B2(n_214),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_179),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_184),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_178),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_251),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_240),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_241),
.A2(n_221),
.B(n_222),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_246),
.B(n_231),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_248),
.A2(n_252),
.B1(n_255),
.B2(n_4),
.Y(n_265)
);

NOR3xp33_ASAP7_75t_SL g251 ( 
.A(n_224),
.B(n_218),
.C(n_184),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_226),
.A2(n_217),
.B1(n_213),
.B2(n_211),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_207),
.C(n_213),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_229),
.C(n_233),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_238),
.A2(n_76),
.B1(n_1),
.B2(n_2),
.Y(n_255)
);

OAI321xp33_ASAP7_75t_L g256 ( 
.A1(n_227),
.A2(n_7),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_4),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_262),
.C(n_247),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_259),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_239),
.Y(n_260)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_260),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_265),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_232),
.C(n_0),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_3),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_264),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_3),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_268),
.Y(n_277)
);

FAx1_ASAP7_75t_SL g267 ( 
.A(n_251),
.B(n_5),
.CI(n_6),
.CON(n_267),
.SN(n_267)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_242),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_249),
.A2(n_6),
.B(n_8),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_264),
.B(n_244),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_271),
.B(n_275),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_247),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_274),
.C(n_262),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_267),
.Y(n_281)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_263),
.Y(n_275)
);

INVxp33_ASAP7_75t_L g280 ( 
.A(n_270),
.Y(n_280)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_280),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_281),
.A2(n_279),
.B1(n_273),
.B2(n_269),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_283),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_278),
.Y(n_283)
);

OAI21x1_ASAP7_75t_L g284 ( 
.A1(n_275),
.A2(n_244),
.B(n_258),
.Y(n_284)
);

AOI31xp67_ASAP7_75t_L g291 ( 
.A1(n_284),
.A2(n_286),
.A3(n_269),
.B(n_12),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_277),
.B(n_246),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_285),
.A2(n_276),
.B(n_243),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_245),
.Y(n_286)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_289),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_291),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_286),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_287),
.C(n_12),
.Y(n_295)
);

AO21x1_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_292),
.B(n_293),
.Y(n_296)
);

NAND2xp33_ASAP7_75t_R g297 ( 
.A(n_296),
.B(n_11),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_13),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_13),
.B(n_15),
.Y(n_299)
);


endmodule