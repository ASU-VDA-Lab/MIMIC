module real_aes_2952_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_0), .B(n_490), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_1), .A2(n_492), .B(n_493), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_2), .B(n_797), .Y(n_796) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_3), .Y(n_779) );
AOI21xp5_ASAP7_75t_L g780 ( .A1(n_3), .A2(n_781), .B(n_785), .Y(n_780) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_4), .Y(n_786) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_5), .B(n_201), .Y(n_527) );
INVx1_ASAP7_75t_L g133 ( .A(n_6), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_7), .B(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_8), .B(n_201), .Y(n_576) );
INVx1_ASAP7_75t_L g171 ( .A(n_9), .Y(n_171) );
CKINVDCx16_ASAP7_75t_R g797 ( .A(n_10), .Y(n_797) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_11), .Y(n_139) );
NAND2xp33_ASAP7_75t_L g568 ( .A(n_12), .B(n_198), .Y(n_568) );
INVx2_ASAP7_75t_L g115 ( .A(n_13), .Y(n_115) );
AOI221x1_ASAP7_75t_L g512 ( .A1(n_14), .A2(n_26), .B1(n_490), .B2(n_492), .C(n_513), .Y(n_512) );
CKINVDCx16_ASAP7_75t_R g473 ( .A(n_15), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_16), .B(n_490), .Y(n_564) );
INVx1_ASAP7_75t_L g199 ( .A(n_17), .Y(n_199) );
AO21x2_ASAP7_75t_L g562 ( .A1(n_18), .A2(n_168), .B(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_19), .B(n_163), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_20), .B(n_201), .Y(n_501) );
AO21x1_ASAP7_75t_L g522 ( .A1(n_21), .A2(n_490), .B(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g477 ( .A(n_22), .Y(n_477) );
INVx1_ASAP7_75t_L g196 ( .A(n_23), .Y(n_196) );
INVx1_ASAP7_75t_SL g183 ( .A(n_24), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_25), .B(n_126), .Y(n_241) );
AOI33xp33_ASAP7_75t_L g221 ( .A1(n_27), .A2(n_52), .A3(n_119), .B1(n_144), .B2(n_222), .B3(n_223), .Y(n_221) );
NAND2x1_ASAP7_75t_L g543 ( .A(n_28), .B(n_201), .Y(n_543) );
NAND2x1_ASAP7_75t_L g575 ( .A(n_29), .B(n_198), .Y(n_575) );
INVx1_ASAP7_75t_L g124 ( .A(n_30), .Y(n_124) );
OA21x2_ASAP7_75t_L g114 ( .A1(n_31), .A2(n_85), .B(n_115), .Y(n_114) );
OR2x2_ASAP7_75t_L g165 ( .A(n_31), .B(n_85), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_32), .B(n_148), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_33), .B(n_198), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_34), .B(n_201), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_35), .B(n_198), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_36), .A2(n_492), .B(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g132 ( .A(n_37), .B(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g143 ( .A(n_37), .Y(n_143) );
AND2x2_ASAP7_75t_L g152 ( .A(n_37), .B(n_122), .Y(n_152) );
OR2x6_ASAP7_75t_L g475 ( .A(n_38), .B(n_476), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_39), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_40), .B(n_490), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_41), .B(n_148), .Y(n_156) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_42), .A2(n_113), .B1(n_190), .B2(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_43), .B(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_44), .B(n_126), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_45), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_46), .B(n_198), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_47), .B(n_168), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_48), .B(n_126), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_49), .A2(n_492), .B(n_574), .Y(n_573) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_50), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_51), .B(n_198), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_53), .B(n_126), .Y(n_160) );
INVx1_ASAP7_75t_L g120 ( .A(n_54), .Y(n_120) );
INVx1_ASAP7_75t_L g128 ( .A(n_54), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_55), .Y(n_804) );
AND2x2_ASAP7_75t_L g162 ( .A(n_56), .B(n_163), .Y(n_162) );
AOI221xp5_ASAP7_75t_L g169 ( .A1(n_57), .A2(n_73), .B1(n_141), .B2(n_148), .C(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_58), .B(n_148), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_59), .B(n_201), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_60), .B(n_113), .Y(n_146) );
AOI21xp5_ASAP7_75t_SL g208 ( .A1(n_61), .A2(n_141), .B(n_209), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_62), .A2(n_492), .B(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g193 ( .A(n_63), .Y(n_193) );
AO21x1_ASAP7_75t_L g524 ( .A1(n_64), .A2(n_492), .B(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_65), .B(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g159 ( .A(n_66), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_67), .B(n_490), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_68), .A2(n_141), .B(n_158), .Y(n_157) );
AND2x2_ASAP7_75t_L g537 ( .A(n_69), .B(n_164), .Y(n_537) );
INVx1_ASAP7_75t_L g122 ( .A(n_70), .Y(n_122) );
INVx1_ASAP7_75t_L g130 ( .A(n_70), .Y(n_130) );
AND2x2_ASAP7_75t_L g578 ( .A(n_71), .B(n_112), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_72), .B(n_148), .Y(n_224) );
AND2x2_ASAP7_75t_L g185 ( .A(n_74), .B(n_112), .Y(n_185) );
INVx1_ASAP7_75t_L g194 ( .A(n_75), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_76), .A2(n_141), .B(n_182), .Y(n_181) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_77), .A2(n_141), .B(n_216), .C(n_240), .Y(n_239) );
OAI22xp33_ASAP7_75t_SL g808 ( .A1(n_78), .A2(n_479), .B1(n_783), .B2(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_78), .Y(n_809) );
INVx1_ASAP7_75t_L g478 ( .A(n_79), .Y(n_478) );
AND2x2_ASAP7_75t_L g487 ( .A(n_80), .B(n_112), .Y(n_487) );
AND2x2_ASAP7_75t_SL g206 ( .A(n_81), .B(n_112), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_82), .B(n_490), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_83), .A2(n_141), .B1(n_219), .B2(n_220), .Y(n_218) );
AND2x2_ASAP7_75t_L g523 ( .A(n_84), .B(n_190), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_86), .B(n_198), .Y(n_502) );
AND2x2_ASAP7_75t_L g546 ( .A(n_87), .B(n_112), .Y(n_546) );
INVx1_ASAP7_75t_L g210 ( .A(n_88), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_89), .B(n_201), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_90), .A2(n_492), .B(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_91), .B(n_198), .Y(n_514) );
AND2x2_ASAP7_75t_L g225 ( .A(n_92), .B(n_112), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_93), .B(n_201), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g116 ( .A1(n_94), .A2(n_117), .B(n_123), .C(n_131), .Y(n_116) );
BUFx2_ASAP7_75t_L g798 ( .A(n_95), .Y(n_798) );
BUFx2_ASAP7_75t_SL g816 ( .A(n_95), .Y(n_816) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_96), .A2(n_492), .B(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_97), .B(n_126), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g98 ( .A1(n_99), .A2(n_790), .B(n_801), .Y(n_98) );
OAI21xp5_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_778), .B(n_780), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
OAI22x1_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_470), .B1(n_479), .B2(n_774), .Y(n_101) );
INVxp67_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
OAI22xp5_ASAP7_75t_SL g781 ( .A1(n_103), .A2(n_782), .B1(n_783), .B2(n_784), .Y(n_781) );
NAND3x1_ASAP7_75t_L g103 ( .A(n_104), .B(n_349), .C(n_416), .Y(n_103) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_309), .Y(n_104) );
NOR3x1_ASAP7_75t_L g105 ( .A(n_106), .B(n_260), .C(n_289), .Y(n_105) );
OAI221xp5_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_174), .B1(n_213), .B2(n_228), .C(n_245), .Y(n_106) );
A2O1A1Ixp33_ASAP7_75t_SL g423 ( .A1(n_107), .A2(n_187), .B(n_424), .C(n_425), .Y(n_423) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_108), .A2(n_395), .B1(n_398), .B2(n_400), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_108), .B(n_214), .Y(n_469) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_153), .Y(n_108) );
BUFx2_ASAP7_75t_L g388 ( .A(n_109), .Y(n_388) );
INVx1_ASAP7_75t_SL g401 ( .A(n_109), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_109), .B(n_256), .Y(n_443) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x4_ASAP7_75t_L g226 ( .A(n_110), .B(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g271 ( .A(n_110), .B(n_167), .Y(n_271) );
INVx1_ASAP7_75t_L g282 ( .A(n_110), .Y(n_282) );
INVx2_ASAP7_75t_L g286 ( .A(n_110), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_110), .B(n_257), .Y(n_413) );
OR2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_136), .Y(n_110) );
OAI22xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_116), .B1(n_134), .B2(n_135), .Y(n_111) );
INVx3_ASAP7_75t_L g135 ( .A(n_112), .Y(n_135) );
INVx4_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_113), .B(n_138), .Y(n_137) );
INVx3_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
BUFx4f_ASAP7_75t_L g168 ( .A(n_114), .Y(n_168) );
AND2x2_ASAP7_75t_SL g164 ( .A(n_115), .B(n_165), .Y(n_164) );
AND2x4_ASAP7_75t_L g190 ( .A(n_115), .B(n_165), .Y(n_190) );
INVxp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
O2A1O1Ixp33_ASAP7_75t_L g158 ( .A1(n_118), .A2(n_159), .B(n_160), .C(n_161), .Y(n_158) );
O2A1O1Ixp33_ASAP7_75t_SL g170 ( .A1(n_118), .A2(n_161), .B(n_171), .C(n_172), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_SL g182 ( .A1(n_118), .A2(n_161), .B(n_183), .C(n_184), .Y(n_182) );
OAI22xp5_ASAP7_75t_L g192 ( .A1(n_118), .A2(n_125), .B1(n_193), .B2(n_194), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g209 ( .A1(n_118), .A2(n_161), .B(n_210), .C(n_211), .Y(n_209) );
INVx2_ASAP7_75t_L g243 ( .A(n_118), .Y(n_243) );
OR2x6_ASAP7_75t_L g118 ( .A(n_119), .B(n_121), .Y(n_118) );
AND2x2_ASAP7_75t_L g149 ( .A(n_119), .B(n_150), .Y(n_149) );
INVxp33_ASAP7_75t_L g222 ( .A(n_119), .Y(n_222) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g145 ( .A(n_120), .B(n_133), .Y(n_145) );
AND2x4_ASAP7_75t_L g201 ( .A(n_120), .B(n_129), .Y(n_201) );
INVx3_ASAP7_75t_L g144 ( .A(n_121), .Y(n_144) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x6_ASAP7_75t_L g198 ( .A(n_122), .B(n_127), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x4_ASAP7_75t_L g490 ( .A(n_126), .B(n_132), .Y(n_490) );
AND2x4_ASAP7_75t_L g126 ( .A(n_127), .B(n_129), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx5_ASAP7_75t_L g161 ( .A(n_132), .Y(n_161) );
HB1xp67_ASAP7_75t_L g150 ( .A(n_133), .Y(n_150) );
AO21x2_ASAP7_75t_L g154 ( .A1(n_135), .A2(n_155), .B(n_162), .Y(n_154) );
AO21x2_ASAP7_75t_L g257 ( .A1(n_135), .A2(n_155), .B(n_162), .Y(n_257) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_135), .A2(n_531), .B(n_537), .Y(n_530) );
AO21x2_ASAP7_75t_L g539 ( .A1(n_135), .A2(n_540), .B(n_546), .Y(n_539) );
AO21x2_ASAP7_75t_L g552 ( .A1(n_135), .A2(n_540), .B(n_546), .Y(n_552) );
AO21x2_ASAP7_75t_L g555 ( .A1(n_135), .A2(n_531), .B(n_537), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_140), .B1(n_146), .B2(n_147), .Y(n_136) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVxp67_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_145), .Y(n_141) );
NOR2x1p5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
INVx1_ASAP7_75t_L g223 ( .A(n_144), .Y(n_223) );
AND2x6_ASAP7_75t_L g492 ( .A(n_145), .B(n_152), .Y(n_492) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
INVx1_ASAP7_75t_L g236 ( .A(n_149), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_151), .Y(n_237) );
BUFx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AND2x2_ASAP7_75t_L g362 ( .A(n_153), .B(n_363), .Y(n_362) );
NOR2x1_ASAP7_75t_L g153 ( .A(n_154), .B(n_166), .Y(n_153) );
INVx2_ASAP7_75t_L g265 ( .A(n_154), .Y(n_265) );
AND2x2_ASAP7_75t_L g285 ( .A(n_154), .B(n_286), .Y(n_285) );
NOR2xp67_ASAP7_75t_L g410 ( .A(n_154), .B(n_286), .Y(n_410) );
AND2x2_ASAP7_75t_L g435 ( .A(n_154), .B(n_278), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_161), .B(n_190), .Y(n_202) );
INVx1_ASAP7_75t_L g219 ( .A(n_161), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_161), .A2(n_241), .B(n_242), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_161), .A2(n_494), .B(n_495), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_161), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_161), .A2(n_514), .B(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_161), .A2(n_526), .B(n_527), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_161), .A2(n_534), .B(n_535), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_161), .A2(n_543), .B(n_544), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_161), .A2(n_567), .B(n_568), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_161), .A2(n_575), .B(n_576), .Y(n_574) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_163), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_163), .A2(n_489), .B(n_491), .Y(n_488) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_163), .A2(n_512), .B(n_516), .Y(n_511) );
OA21x2_ASAP7_75t_L g582 ( .A1(n_163), .A2(n_512), .B(n_516), .Y(n_582) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g227 ( .A(n_167), .Y(n_227) );
INVx1_ASAP7_75t_L g249 ( .A(n_167), .Y(n_249) );
INVxp67_ASAP7_75t_L g288 ( .A(n_167), .Y(n_288) );
AND2x4_ASAP7_75t_L g328 ( .A(n_167), .B(n_329), .Y(n_328) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_167), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_167), .B(n_279), .Y(n_414) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_173), .Y(n_167) );
INVx2_ASAP7_75t_SL g216 ( .A(n_168), .Y(n_216) );
INVx1_ASAP7_75t_SL g174 ( .A(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_186), .Y(n_175) );
AND2x2_ASAP7_75t_L g302 ( .A(n_176), .B(n_274), .Y(n_302) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_177), .Y(n_230) );
AND2x2_ASAP7_75t_L g258 ( .A(n_177), .B(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g269 ( .A(n_177), .Y(n_269) );
INVx1_ASAP7_75t_L g293 ( .A(n_177), .Y(n_293) );
AND2x2_ASAP7_75t_L g296 ( .A(n_177), .B(n_188), .Y(n_296) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_177), .Y(n_318) );
AO21x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_185), .Y(n_177) );
AO21x2_ASAP7_75t_L g571 ( .A1(n_178), .A2(n_572), .B(n_578), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
NOR2x1_ASAP7_75t_L g186 ( .A(n_187), .B(n_203), .Y(n_186) );
AND2x2_ASAP7_75t_L g283 ( .A(n_187), .B(n_205), .Y(n_283) );
NAND2x1_ASAP7_75t_L g316 ( .A(n_187), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g419 ( .A(n_187), .Y(n_419) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx3_ASAP7_75t_L g259 ( .A(n_188), .Y(n_259) );
AND2x2_ASAP7_75t_L g274 ( .A(n_188), .B(n_233), .Y(n_274) );
NOR2x1_ASAP7_75t_SL g343 ( .A(n_188), .B(n_205), .Y(n_343) );
AND2x4_ASAP7_75t_L g188 ( .A(n_189), .B(n_191), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_190), .A2(n_208), .B(n_212), .Y(n_207) );
INVx1_ASAP7_75t_SL g497 ( .A(n_190), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_190), .B(n_529), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_190), .A2(n_564), .B(n_565), .Y(n_563) );
OAI21xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_195), .B(n_202), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B1(n_199), .B2(n_200), .Y(n_195) );
INVxp67_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVxp67_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NOR2x1_ASAP7_75t_L g380 ( .A(n_203), .B(n_367), .Y(n_380) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g305 ( .A(n_204), .B(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx4_ASAP7_75t_L g244 ( .A(n_205), .Y(n_244) );
AND2x4_ASAP7_75t_L g251 ( .A(n_205), .B(n_252), .Y(n_251) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_205), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_205), .B(n_268), .Y(n_368) );
AND2x2_ASAP7_75t_L g396 ( .A(n_205), .B(n_233), .Y(n_396) );
OR2x6_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
NAND2x1_ASAP7_75t_SL g213 ( .A(n_214), .B(n_226), .Y(n_213) );
OR2x2_ASAP7_75t_L g424 ( .A(n_214), .B(n_336), .Y(n_424) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x4_ASAP7_75t_L g264 ( .A(n_215), .B(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g329 ( .A(n_215), .Y(n_329) );
AND2x2_ASAP7_75t_L g363 ( .A(n_215), .B(n_286), .Y(n_363) );
AO21x2_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B(n_225), .Y(n_215) );
AO21x2_ASAP7_75t_L g279 ( .A1(n_216), .A2(n_217), .B(n_225), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_218), .B(n_224), .Y(n_217) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx3_ASAP7_75t_L g336 ( .A(n_226), .Y(n_336) );
AND2x2_ASAP7_75t_L g344 ( .A(n_226), .B(n_277), .Y(n_344) );
AND2x2_ASAP7_75t_L g461 ( .A(n_226), .B(n_264), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_229), .B(n_231), .Y(n_228) );
BUFx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g415 ( .A(n_230), .B(n_356), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_230), .B(n_255), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_231), .A2(n_292), .B(n_295), .Y(n_291) );
AND2x2_ASAP7_75t_L g361 ( .A(n_231), .B(n_267), .Y(n_361) );
INVx2_ASAP7_75t_SL g448 ( .A(n_231), .Y(n_448) );
AND2x4_ASAP7_75t_SL g231 ( .A(n_232), .B(n_244), .Y(n_231) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g252 ( .A(n_233), .Y(n_252) );
INVx2_ASAP7_75t_L g299 ( .A(n_233), .Y(n_299) );
AND2x4_ASAP7_75t_L g306 ( .A(n_233), .B(n_259), .Y(n_306) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_239), .Y(n_233) );
NOR3xp33_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .C(n_238), .Y(n_235) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_244), .Y(n_262) );
AND2x4_ASAP7_75t_L g338 ( .A(n_244), .B(n_252), .Y(n_338) );
OR2x2_ASAP7_75t_L g464 ( .A(n_244), .B(n_465), .Y(n_464) );
NAND4xp25_ASAP7_75t_L g245 ( .A(n_246), .B(n_250), .C(n_253), .D(n_258), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g311 ( .A(n_247), .B(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g408 ( .A(n_247), .Y(n_408) );
INVx3_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
NAND2x1p5_ASAP7_75t_L g308 ( .A(n_248), .B(n_256), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_248), .B(n_313), .Y(n_442) );
BUFx3_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_251), .B(n_267), .Y(n_320) );
INVx2_ASAP7_75t_L g422 ( .A(n_251), .Y(n_422) );
AND2x2_ASAP7_75t_SL g432 ( .A(n_251), .B(n_292), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_251), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g324 ( .A(n_255), .B(n_271), .Y(n_324) );
AND2x2_ASAP7_75t_L g392 ( .A(n_255), .B(n_328), .Y(n_392) );
INVx3_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x4_ASAP7_75t_L g277 ( .A(n_256), .B(n_278), .Y(n_277) );
INVx3_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_257), .Y(n_331) );
AND2x2_ASAP7_75t_L g382 ( .A(n_257), .B(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_257), .B(n_279), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_258), .B(n_422), .Y(n_429) );
INVx1_ASAP7_75t_SL g465 ( .A(n_258), .Y(n_465) );
INVx1_ASAP7_75t_L g294 ( .A(n_259), .Y(n_294) );
AND2x2_ASAP7_75t_L g356 ( .A(n_259), .B(n_299), .Y(n_356) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_270), .B(n_272), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
AND2x2_ASAP7_75t_L g322 ( .A(n_264), .B(n_271), .Y(n_322) );
AND2x2_ASAP7_75t_L g430 ( .A(n_264), .B(n_281), .Y(n_430) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g304 ( .A(n_267), .Y(n_304) );
AND2x2_ASAP7_75t_L g337 ( .A(n_267), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g342 ( .A(n_267), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_267), .B(n_306), .Y(n_391) );
NOR3xp33_ASAP7_75t_L g441 ( .A(n_267), .B(n_442), .C(n_443), .Y(n_441) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVxp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_276), .B1(n_283), .B2(n_284), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx2_ASAP7_75t_L g367 ( .A(n_274), .Y(n_367) );
AND2x2_ASAP7_75t_L g301 ( .A(n_275), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g323 ( .A(n_275), .B(n_296), .Y(n_323) );
AND2x2_ASAP7_75t_SL g355 ( .A(n_275), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_280), .Y(n_276) );
INVx1_ASAP7_75t_L g334 ( .A(n_277), .Y(n_334) );
AND2x2_ASAP7_75t_L g287 ( .A(n_278), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g313 ( .A(n_278), .Y(n_313) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g376 ( .A(n_282), .B(n_328), .Y(n_376) );
INVx1_ASAP7_75t_L g434 ( .A(n_282), .Y(n_434) );
INVx1_ASAP7_75t_L g290 ( .A(n_284), .Y(n_290) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
NAND2x1p5_ASAP7_75t_L g312 ( .A(n_285), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g421 ( .A(n_285), .B(n_328), .Y(n_421) );
AND2x2_ASAP7_75t_L g387 ( .A(n_287), .B(n_388), .Y(n_387) );
NAND2x1p5_ASAP7_75t_L g455 ( .A(n_287), .B(n_456), .Y(n_455) );
OAI21xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_291), .B(n_300), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_292), .B(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g348 ( .A(n_292), .B(n_297), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_292), .B(n_338), .Y(n_399) );
AND2x4_ASAP7_75t_SL g292 ( .A(n_293), .B(n_294), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_293), .B(n_356), .Y(n_386) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_293), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g321 ( .A1(n_295), .A2(n_322), .B1(n_323), .B2(n_324), .Y(n_321) );
AND2x2_ASAP7_75t_SL g295 ( .A(n_296), .B(n_297), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_296), .B(n_338), .Y(n_357) );
INVx1_ASAP7_75t_L g458 ( .A(n_296), .Y(n_458) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OAI21xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_303), .B(n_307), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_302), .B(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_L g439 ( .A(n_305), .Y(n_439) );
INVx4_ASAP7_75t_L g341 ( .A(n_306), .Y(n_341) );
INVxp33_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g369 ( .A(n_308), .B(n_370), .Y(n_369) );
NOR2x1_ASAP7_75t_L g309 ( .A(n_310), .B(n_325), .Y(n_309) );
OAI21xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_314), .B(n_321), .Y(n_310) );
INVx1_ASAP7_75t_L g359 ( .A(n_312), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_315), .B(n_319), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g364 ( .A(n_316), .Y(n_364) );
INVx1_ASAP7_75t_L g397 ( .A(n_317), .Y(n_397) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_322), .A2(n_361), .B1(n_362), .B2(n_364), .Y(n_360) );
INVx1_ASAP7_75t_L g374 ( .A(n_323), .Y(n_374) );
NAND4xp25_ASAP7_75t_SL g325 ( .A(n_326), .B(n_332), .C(n_339), .D(n_345), .Y(n_325) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
INVx1_ASAP7_75t_L g347 ( .A(n_328), .Y(n_347) );
AND2x2_ASAP7_75t_L g459 ( .A(n_328), .B(n_456), .Y(n_459) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_337), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g466 ( .A(n_336), .B(n_403), .Y(n_466) );
INVx1_ASAP7_75t_L g463 ( .A(n_337), .Y(n_463) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_338), .Y(n_372) );
OAI21xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_342), .B(n_344), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_377), .Y(n_349) );
NOR3xp33_ASAP7_75t_L g350 ( .A(n_351), .B(n_365), .C(n_373), .Y(n_350) );
OAI21xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_358), .B(n_360), .Y(n_351) );
INVxp67_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_357), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_355), .A2(n_387), .B1(n_390), .B2(n_392), .Y(n_389) );
OAI22xp33_ASAP7_75t_L g365 ( .A1(n_358), .A2(n_366), .B1(n_369), .B2(n_371), .Y(n_365) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g370 ( .A(n_363), .Y(n_370) );
AND2x4_ASAP7_75t_L g381 ( .A(n_363), .B(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_368), .Y(n_468) );
AOI31xp33_ASAP7_75t_L g467 ( .A1(n_371), .A2(n_444), .A3(n_468), .B(n_469), .Y(n_467) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_378), .B(n_393), .Y(n_377) );
NAND2xp5_ASAP7_75t_SL g378 ( .A(n_379), .B(n_389), .Y(n_378) );
AOI22xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_381), .B1(n_384), .B2(n_387), .Y(n_379) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_383), .Y(n_447) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_391), .B(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_394), .B(n_404), .Y(n_393) );
AND2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
AND2x2_ASAP7_75t_L g405 ( .A(n_396), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g444 ( .A(n_396), .Y(n_444) );
AOI22xp33_ASAP7_75t_SL g453 ( .A1(n_396), .A2(n_454), .B1(n_457), .B2(n_459), .Y(n_453) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_401), .B(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_407), .B1(n_411), .B2(n_415), .Y(n_404) );
NOR2xp33_ASAP7_75t_SL g407 ( .A(n_408), .B(n_409), .Y(n_407) );
INVxp67_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
INVx2_ASAP7_75t_SL g456 ( .A(n_413), .Y(n_456) );
INVx2_ASAP7_75t_L g437 ( .A(n_414), .Y(n_437) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_451), .Y(n_416) );
AOI211xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_423), .B(n_426), .C(n_440), .Y(n_417) );
OAI21xp33_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_420), .B(n_422), .Y(n_418) );
INVx1_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g425 ( .A(n_422), .Y(n_425) );
NAND2xp5_ASAP7_75t_SL g426 ( .A(n_427), .B(n_431), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_430), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_433), .B1(n_436), .B2(n_438), .Y(n_431) );
AND2x2_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
AND2x2_ASAP7_75t_L g436 ( .A(n_434), .B(n_437), .Y(n_436) );
AO22x1_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_444), .B1(n_445), .B2(n_449), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_446), .B(n_448), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
NOR3xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_462), .C(n_467), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_453), .B(n_460), .Y(n_452) );
INVx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AOI21xp33_ASAP7_75t_R g462 ( .A1(n_463), .A2(n_464), .B(n_466), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g470 ( .A(n_471), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_471), .Y(n_782) );
CKINVDCx11_ASAP7_75t_R g471 ( .A(n_472), .Y(n_471) );
OR2x6_ASAP7_75t_SL g472 ( .A(n_473), .B(n_474), .Y(n_472) );
AND2x6_ASAP7_75t_SL g777 ( .A(n_473), .B(n_475), .Y(n_777) );
OR2x2_ASAP7_75t_L g789 ( .A(n_473), .B(n_475), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_473), .B(n_474), .Y(n_800) );
CKINVDCx5p33_ASAP7_75t_R g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
BUFx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx3_ASAP7_75t_SL g783 ( .A(n_480), .Y(n_783) );
NOR2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_661), .Y(n_480) );
AO211x2_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_506), .B(n_556), .C(n_629), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVxp67_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
AND3x2_ASAP7_75t_L g710 ( .A(n_484), .B(n_591), .C(n_607), .Y(n_710) );
AND2x4_ASAP7_75t_L g713 ( .A(n_484), .B(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_496), .Y(n_484) );
NAND2x1p5_ASAP7_75t_L g569 ( .A(n_485), .B(n_570), .Y(n_569) );
INVx4_ASAP7_75t_L g622 ( .A(n_485), .Y(n_622) );
AND2x2_ASAP7_75t_SL g707 ( .A(n_485), .B(n_616), .Y(n_707) );
AND2x2_ASAP7_75t_L g750 ( .A(n_485), .B(n_571), .Y(n_750) );
INVx5_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx2_ASAP7_75t_L g599 ( .A(n_486), .Y(n_599) );
AND2x2_ASAP7_75t_L g618 ( .A(n_486), .B(n_562), .Y(n_618) );
AND2x2_ASAP7_75t_L g636 ( .A(n_486), .B(n_571), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_486), .B(n_570), .Y(n_696) );
NOR2x1_ASAP7_75t_SL g723 ( .A(n_486), .B(n_496), .Y(n_723) );
OR2x6_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_496), .B(n_562), .Y(n_561) );
AO21x2_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B(n_504), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_497), .B(n_505), .Y(n_504) );
AO21x2_ASAP7_75t_L g595 ( .A1(n_497), .A2(n_498), .B(n_504), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_499), .B(n_503), .Y(n_498) );
AO21x1_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_538), .B(n_547), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
OAI22xp33_ASAP7_75t_L g604 ( .A1(n_508), .A2(n_605), .B1(n_609), .B2(n_610), .Y(n_604) );
OR2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_517), .Y(n_508) );
AND2x2_ASAP7_75t_L g665 ( .A(n_509), .B(n_553), .Y(n_665) );
BUFx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x4_ASAP7_75t_L g598 ( .A(n_510), .B(n_581), .Y(n_598) );
AND2x2_ASAP7_75t_L g670 ( .A(n_510), .B(n_555), .Y(n_670) );
AND2x2_ASAP7_75t_L g689 ( .A(n_510), .B(n_655), .Y(n_689) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g548 ( .A(n_511), .Y(n_548) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_511), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_517), .B(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g649 ( .A(n_518), .B(n_550), .Y(n_649) );
AND2x4_ASAP7_75t_L g518 ( .A(n_519), .B(n_530), .Y(n_518) );
AND2x2_ASAP7_75t_L g553 ( .A(n_519), .B(n_554), .Y(n_553) );
OR2x2_ASAP7_75t_L g586 ( .A(n_519), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_SL g646 ( .A(n_519), .B(n_582), .Y(n_646) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx2_ASAP7_75t_L g739 ( .A(n_520), .Y(n_739) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g581 ( .A(n_521), .Y(n_581) );
OAI21x1_ASAP7_75t_SL g521 ( .A1(n_522), .A2(n_524), .B(n_528), .Y(n_521) );
INVx1_ASAP7_75t_L g529 ( .A(n_523), .Y(n_529) );
INVx2_ASAP7_75t_L g587 ( .A(n_530), .Y(n_587) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_530), .Y(n_687) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_532), .B(n_536), .Y(n_531) );
INVx2_ASAP7_75t_L g583 ( .A(n_538), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_538), .B(n_715), .Y(n_741) );
AND2x2_ASAP7_75t_L g760 ( .A(n_538), .B(n_750), .Y(n_760) );
BUFx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x4_ASAP7_75t_SL g628 ( .A(n_539), .B(n_587), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_545), .Y(n_540) );
AND2x2_ASAP7_75t_SL g547 ( .A(n_548), .B(n_549), .Y(n_547) );
AND2x2_ASAP7_75t_L g627 ( .A(n_548), .B(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_548), .B(n_597), .Y(n_632) );
INVx1_ASAP7_75t_SL g759 ( .A(n_548), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_549), .B(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_553), .Y(n_549) );
INVx1_ASAP7_75t_L g585 ( .A(n_550), .Y(n_585) );
AND2x2_ASAP7_75t_L g771 ( .A(n_550), .B(n_772), .Y(n_771) );
BUFx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g647 ( .A(n_551), .B(n_554), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_551), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g701 ( .A(n_551), .B(n_555), .Y(n_701) );
AND2x2_ASAP7_75t_L g732 ( .A(n_551), .B(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g597 ( .A(n_552), .B(n_555), .Y(n_597) );
INVxp67_ASAP7_75t_L g614 ( .A(n_552), .Y(n_614) );
BUFx3_ASAP7_75t_L g655 ( .A(n_552), .Y(n_655) );
AND2x2_ASAP7_75t_L g675 ( .A(n_553), .B(n_676), .Y(n_675) );
NAND2xp33_ASAP7_75t_L g688 ( .A(n_553), .B(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_554), .B(n_581), .Y(n_644) );
AND2x2_ASAP7_75t_L g733 ( .A(n_554), .B(n_582), .Y(n_733) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g660 ( .A(n_555), .B(n_582), .Y(n_660) );
OR3x1_ASAP7_75t_L g556 ( .A(n_557), .B(n_604), .C(n_619), .Y(n_556) );
OAI321xp33_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_569), .A3(n_579), .B1(n_584), .B2(n_588), .C(n_596), .Y(n_557) );
INVx1_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVxp67_ASAP7_75t_SL g635 ( .A(n_561), .Y(n_635) );
INVxp67_ASAP7_75t_SL g653 ( .A(n_561), .Y(n_653) );
OR2x2_ASAP7_75t_L g657 ( .A(n_561), .B(n_569), .Y(n_657) );
BUFx3_ASAP7_75t_L g591 ( .A(n_562), .Y(n_591) );
AND2x2_ASAP7_75t_L g608 ( .A(n_562), .B(n_594), .Y(n_608) );
INVx1_ASAP7_75t_L g625 ( .A(n_562), .Y(n_625) );
INVx2_ASAP7_75t_L g641 ( .A(n_562), .Y(n_641) );
OR2x2_ASAP7_75t_L g680 ( .A(n_562), .B(n_570), .Y(n_680) );
INVx2_ASAP7_75t_L g668 ( .A(n_569), .Y(n_668) );
AND2x2_ASAP7_75t_L g592 ( .A(n_570), .B(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g607 ( .A(n_570), .Y(n_607) );
AND2x4_ASAP7_75t_L g616 ( .A(n_570), .B(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_570), .B(n_593), .Y(n_639) );
AND2x2_ASAP7_75t_L g746 ( .A(n_570), .B(n_641), .Y(n_746) );
INVx4_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_571), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_577), .Y(n_572) );
INVx1_ASAP7_75t_L g633 ( .A(n_579), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_580), .B(n_583), .Y(n_579) );
AND2x2_ASAP7_75t_L g720 ( .A(n_580), .B(n_647), .Y(n_720) );
INVx1_ASAP7_75t_SL g737 ( .A(n_580), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_580), .B(n_713), .Y(n_766) );
AND2x4_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
OR2x2_ASAP7_75t_L g609 ( .A(n_581), .B(n_582), .Y(n_609) );
AND2x2_ASAP7_75t_L g702 ( .A(n_583), .B(n_598), .Y(n_702) );
OR2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g725 ( .A(n_587), .B(n_598), .Y(n_725) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_589), .A2(n_738), .B1(n_743), .B2(n_745), .Y(n_742) );
AND2x4_ASAP7_75t_L g589 ( .A(n_590), .B(n_592), .Y(n_589) );
AND2x2_ASAP7_75t_L g667 ( .A(n_590), .B(n_668), .Y(n_667) );
OR2x2_ASAP7_75t_L g762 ( .A(n_590), .B(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g718 ( .A(n_591), .B(n_636), .Y(n_718) );
AND2x4_ASAP7_75t_L g672 ( .A(n_592), .B(n_618), .Y(n_672) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
HB1xp67_ASAP7_75t_L g770 ( .A(n_594), .Y(n_770) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g603 ( .A(n_595), .Y(n_603) );
INVx1_ASAP7_75t_L g617 ( .A(n_595), .Y(n_617) );
NAND4xp25_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .C(n_599), .D(n_600), .Y(n_596) );
AND2x2_ASAP7_75t_L g754 ( .A(n_597), .B(n_739), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_597), .B(n_765), .Y(n_764) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_598), .B(n_674), .Y(n_673) );
OAI322xp33_ASAP7_75t_L g681 ( .A1(n_598), .A2(n_682), .A3(n_686), .B1(n_688), .B2(n_690), .C1(n_692), .C2(n_697), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_598), .B(n_647), .Y(n_697) );
INVx1_ASAP7_75t_L g765 ( .A(n_598), .Y(n_765) );
INVx2_ASAP7_75t_L g611 ( .A(n_599), .Y(n_611) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_602), .B(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_603), .B(n_622), .Y(n_679) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_606), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
INVx1_ASAP7_75t_L g652 ( .A(n_607), .Y(n_652) );
AND2x2_ASAP7_75t_L g724 ( .A(n_607), .B(n_635), .Y(n_724) );
AOI31xp33_ASAP7_75t_L g610 ( .A1(n_608), .A2(n_611), .A3(n_612), .B(n_615), .Y(n_610) );
AND2x2_ASAP7_75t_L g621 ( .A(n_608), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g749 ( .A(n_608), .B(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_SL g756 ( .A(n_608), .B(n_636), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_608), .Y(n_757) );
INVx1_ASAP7_75t_SL g715 ( .A(n_609), .Y(n_715) );
NAND3xp33_ASAP7_75t_SL g743 ( .A(n_609), .B(n_737), .C(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g643 ( .A(n_614), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
AND2x2_ASAP7_75t_L g624 ( .A(n_616), .B(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g685 ( .A(n_616), .Y(n_685) );
AOI322xp5_ASAP7_75t_L g767 ( .A1(n_616), .A2(n_646), .A3(n_649), .B1(n_768), .B2(n_769), .C1(n_771), .C2(n_773), .Y(n_767) );
AND2x2_ASAP7_75t_L g773 ( .A(n_616), .B(n_622), .Y(n_773) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_623), .B(n_626), .Y(n_619) );
INVx1_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_622), .B(n_641), .Y(n_640) );
AND2x4_ASAP7_75t_L g768 ( .A(n_622), .B(n_655), .Y(n_768) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g694 ( .A(n_625), .Y(n_694) );
AND2x2_ASAP7_75t_L g722 ( .A(n_625), .B(n_723), .Y(n_722) );
AND2x2_ASAP7_75t_L g769 ( .A(n_625), .B(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g674 ( .A(n_628), .Y(n_674) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
O2A1O1Ixp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_633), .B(n_634), .C(n_637), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
AND2x2_ASAP7_75t_L g691 ( .A(n_636), .B(n_641), .Y(n_691) );
OAI211xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_642), .B(n_648), .C(n_650), .Y(n_637) );
OAI221xp5_ASAP7_75t_L g663 ( .A1(n_638), .A2(n_664), .B1(n_666), .B2(n_669), .C(n_671), .Y(n_663) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
INVx1_ASAP7_75t_L g683 ( .A(n_640), .Y(n_683) );
OR2x2_ASAP7_75t_L g703 ( .A(n_640), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
INVx1_ASAP7_75t_L g748 ( .A(n_643), .Y(n_748) );
INVx1_ASAP7_75t_L g772 ( .A(n_644), .Y(n_772) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_646), .B(n_647), .Y(n_645) );
AND2x2_ASAP7_75t_L g654 ( .A(n_646), .B(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_646), .B(n_716), .Y(n_728) );
INVx1_ASAP7_75t_L g708 ( .A(n_647), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_654), .B1(n_656), .B2(n_658), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx1_ASAP7_75t_SL g716 ( .A(n_655), .Y(n_716) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NAND4xp75_ASAP7_75t_L g661 ( .A(n_662), .B(n_698), .C(n_726), .D(n_751), .Y(n_661) );
NOR2xp67_ASAP7_75t_L g662 ( .A(n_663), .B(n_681), .Y(n_662) );
INVx1_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_SL g738 ( .A(n_670), .B(n_739), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_673), .B1(n_675), .B2(n_677), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_674), .B(n_737), .Y(n_736) );
INVx2_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
OR2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
INVx2_ASAP7_75t_L g714 ( .A(n_680), .Y(n_714) );
OR2x2_ASAP7_75t_L g729 ( .A(n_680), .B(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_SL g682 ( .A(n_683), .B(n_684), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g744 ( .A(n_689), .Y(n_744) );
INVx1_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
OAI21xp5_ASAP7_75t_SL g735 ( .A1(n_691), .A2(n_736), .B(n_738), .Y(n_735) );
INVxp67_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NOR2x1_ASAP7_75t_L g698 ( .A(n_699), .B(n_711), .Y(n_698) );
OAI221xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_703), .B1(n_706), .B2(n_708), .C(n_709), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
OAI21xp33_ASAP7_75t_L g747 ( .A1(n_701), .A2(n_748), .B(n_749), .Y(n_747) );
INVx3_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
OAI322xp33_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_715), .A3(n_716), .B1(n_717), .B2(n_719), .C1(n_721), .C2(n_725), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
NOR2x1_ASAP7_75t_L g721 ( .A(n_722), .B(n_724), .Y(n_721) );
INVx1_ASAP7_75t_L g734 ( .A(n_722), .Y(n_734) );
INVx1_ASAP7_75t_L g730 ( .A(n_723), .Y(n_730) );
AND2x2_ASAP7_75t_L g745 ( .A(n_723), .B(n_746), .Y(n_745) );
NOR2x1_ASAP7_75t_L g726 ( .A(n_727), .B(n_740), .Y(n_726) );
OAI221xp5_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_729), .B1(n_731), .B2(n_734), .C(n_735), .Y(n_727) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
OAI211xp5_ASAP7_75t_SL g740 ( .A1(n_734), .A2(n_741), .B(n_742), .C(n_747), .Y(n_740) );
INVx2_ASAP7_75t_SL g763 ( .A(n_750), .Y(n_763) );
NOR2x1_ASAP7_75t_L g751 ( .A(n_752), .B(n_761), .Y(n_751) );
OAI22xp33_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_755), .B1(n_757), .B2(n_758), .Y(n_752) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
OAI211xp5_ASAP7_75t_SL g761 ( .A1(n_762), .A2(n_764), .B(n_766), .C(n_767), .Y(n_761) );
CKINVDCx11_ASAP7_75t_R g774 ( .A(n_775), .Y(n_774) );
INVx3_ASAP7_75t_SL g775 ( .A(n_776), .Y(n_775) );
CKINVDCx5p33_ASAP7_75t_R g776 ( .A(n_777), .Y(n_776) );
CKINVDCx11_ASAP7_75t_R g784 ( .A(n_777), .Y(n_784) );
CKINVDCx5p33_ASAP7_75t_R g778 ( .A(n_779), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g785 ( .A(n_786), .B(n_787), .Y(n_785) );
CKINVDCx5p33_ASAP7_75t_R g787 ( .A(n_788), .Y(n_787) );
INVx3_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_791), .Y(n_790) );
INVx2_ASAP7_75t_SL g791 ( .A(n_792), .Y(n_791) );
AND2x2_ASAP7_75t_L g792 ( .A(n_793), .B(n_799), .Y(n_792) );
INVxp67_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
NAND2xp5_ASAP7_75t_SL g794 ( .A(n_795), .B(n_798), .Y(n_794) );
INVx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
OR2x2_ASAP7_75t_SL g812 ( .A(n_796), .B(n_798), .Y(n_812) );
AOI21xp5_ASAP7_75t_L g813 ( .A1(n_796), .A2(n_814), .B(n_817), .Y(n_813) );
BUFx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
BUFx3_ASAP7_75t_L g805 ( .A(n_800), .Y(n_805) );
BUFx2_ASAP7_75t_L g818 ( .A(n_800), .Y(n_818) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_809), .B1(n_810), .B2(n_813), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g802 ( .A(n_803), .B(n_806), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_805), .B(n_808), .Y(n_807) );
INVxp67_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
CKINVDCx11_ASAP7_75t_R g814 ( .A(n_815), .Y(n_814) );
CKINVDCx8_ASAP7_75t_R g815 ( .A(n_816), .Y(n_815) );
INVx2_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
endmodule