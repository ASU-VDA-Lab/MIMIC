module fake_netlist_6_505_n_1692 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1692);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1692;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_32),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_30),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_94),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_128),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_27),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_41),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_41),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_85),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_135),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_111),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_88),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_26),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_10),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_24),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_51),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_59),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_98),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_22),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_14),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_54),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_26),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_97),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_62),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_24),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_147),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_3),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_84),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_45),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_80),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_82),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_32),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_38),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_48),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_75),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_21),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_60),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_140),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_3),
.Y(n_195)
);

BUFx10_ASAP7_75t_L g196 ( 
.A(n_76),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_70),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_13),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_114),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_83),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_138),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_96),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_107),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_123),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_137),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_7),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_92),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_51),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_142),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_63),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_73),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_46),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_109),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_115),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_72),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_125),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_74),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_101),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_113),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_22),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_7),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_49),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_40),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_90),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_14),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_10),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_2),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_86),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_42),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_25),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_48),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_67),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_118),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_6),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_16),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_57),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_4),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_4),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_2),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_117),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_49),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_17),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_65),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_30),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_27),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_52),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_81),
.Y(n_247)
);

BUFx10_ASAP7_75t_L g248 ( 
.A(n_77),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_99),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_102),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_104),
.Y(n_251)
);

BUFx10_ASAP7_75t_L g252 ( 
.A(n_9),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_47),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_116),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_146),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_47),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_58),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_11),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_139),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_121),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_21),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_34),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_64),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_79),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_132),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_148),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_42),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_150),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_55),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_38),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_87),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_25),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_95),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_46),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_5),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_56),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_133),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_103),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_52),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_29),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_6),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_15),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_0),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_106),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_129),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_18),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_1),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_120),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_89),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_122),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_5),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_11),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_91),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_126),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_16),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_29),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_36),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_19),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_1),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_78),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_13),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_20),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_33),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_130),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_159),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_154),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_170),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_157),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_202),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_159),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_161),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_162),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_209),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_159),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_159),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_164),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_172),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_175),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_177),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_159),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_178),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_159),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_288),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_155),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_153),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_171),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_180),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_166),
.Y(n_328)
);

INVxp33_ASAP7_75t_SL g329 ( 
.A(n_152),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_166),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_171),
.B(n_0),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_281),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_281),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_277),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_296),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_193),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_163),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_277),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_194),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_296),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_223),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_223),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_223),
.Y(n_343)
);

INVxp33_ASAP7_75t_SL g344 ( 
.A(n_158),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_197),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_163),
.Y(n_346)
);

INVxp33_ASAP7_75t_SL g347 ( 
.A(n_165),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_199),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_197),
.B(n_8),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_240),
.B(n_8),
.Y(n_350)
);

NOR2xp67_ASAP7_75t_L g351 ( 
.A(n_163),
.B(n_9),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_153),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_160),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_169),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_160),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_211),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_155),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_167),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_156),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_167),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_240),
.B(n_12),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_265),
.B(n_12),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_200),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_201),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_190),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_204),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_207),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_213),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_190),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_215),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_217),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_198),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_218),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_219),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_305),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_305),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_354),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_341),
.B(n_265),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_310),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_310),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_341),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_314),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_314),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_315),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_337),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_315),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_342),
.B(n_186),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_320),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_342),
.B(n_186),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_337),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_320),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_343),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_334),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_337),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_322),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_337),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_322),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_337),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_346),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_346),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_346),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_343),
.B(n_163),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_357),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_351),
.B(n_214),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_357),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_359),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_346),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_331),
.B(n_196),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_359),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_346),
.B(n_214),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_355),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_364),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_324),
.B(n_214),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_355),
.B(n_214),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_328),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_328),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_330),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_330),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_332),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_358),
.B(n_224),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_332),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_358),
.B(n_228),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_333),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_333),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_326),
.B(n_189),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_338),
.B(n_239),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_335),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_345),
.B(n_189),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_335),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_360),
.B(n_184),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_340),
.B(n_230),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_353),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_325),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_340),
.Y(n_434)
);

OR2x6_ASAP7_75t_L g435 ( 
.A(n_349),
.B(n_208),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_352),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_360),
.B(n_233),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_356),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_365),
.B(n_184),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_376),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_394),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_381),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_402),
.B(n_156),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_375),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_402),
.B(n_365),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_394),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_381),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_392),
.Y(n_448)
);

INVxp33_ASAP7_75t_L g449 ( 
.A(n_426),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_412),
.Y(n_450)
);

NOR2x1p5_ASAP7_75t_L g451 ( 
.A(n_378),
.B(n_230),
.Y(n_451)
);

OR2x6_ASAP7_75t_L g452 ( 
.A(n_435),
.B(n_350),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_408),
.B(n_329),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_385),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_375),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_375),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_392),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g458 ( 
.A(n_426),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_408),
.B(n_344),
.Y(n_459)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_394),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_433),
.Y(n_461)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_394),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_394),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_L g464 ( 
.A1(n_435),
.A2(n_361),
.B1(n_362),
.B2(n_208),
.Y(n_464)
);

AND3x2_ASAP7_75t_L g465 ( 
.A(n_433),
.B(n_264),
.C(n_260),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_411),
.Y(n_466)
);

BUFx4f_ASAP7_75t_L g467 ( 
.A(n_404),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_436),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_425),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_425),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_375),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_432),
.B(n_306),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_425),
.A2(n_374),
.B1(n_366),
.B2(n_367),
.Y(n_473)
);

INVx2_ASAP7_75t_SL g474 ( 
.A(n_428),
.Y(n_474)
);

AND2x6_ASAP7_75t_L g475 ( 
.A(n_410),
.B(n_260),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_410),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_376),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_420),
.B(n_347),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_391),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_391),
.Y(n_480)
);

AND2x6_ASAP7_75t_L g481 ( 
.A(n_410),
.B(n_264),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_385),
.B(n_308),
.Y(n_482)
);

AND2x2_ASAP7_75t_SL g483 ( 
.A(n_404),
.B(n_269),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_411),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_410),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_420),
.B(n_311),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_378),
.B(n_422),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_379),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_422),
.B(n_312),
.Y(n_489)
);

BUFx4f_ASAP7_75t_L g490 ( 
.A(n_404),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_394),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_379),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_432),
.B(n_316),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_379),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_385),
.Y(n_495)
);

BUFx6f_ASAP7_75t_SL g496 ( 
.A(n_435),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_390),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_379),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_390),
.B(n_317),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g500 ( 
.A1(n_435),
.A2(n_279),
.B1(n_198),
.B2(n_235),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_383),
.Y(n_501)
);

AO22x2_ASAP7_75t_L g502 ( 
.A1(n_404),
.A2(n_291),
.B1(n_235),
.B2(n_238),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_410),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_428),
.B(n_318),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_412),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_383),
.Y(n_506)
);

INVx5_ASAP7_75t_L g507 ( 
.A(n_394),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_410),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_390),
.B(n_319),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_380),
.Y(n_510)
);

INVx4_ASAP7_75t_L g511 ( 
.A(n_394),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_398),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_383),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_383),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_428),
.Y(n_515)
);

NAND3xp33_ASAP7_75t_L g516 ( 
.A(n_437),
.B(n_327),
.C(n_321),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_377),
.B(n_336),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_380),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_377),
.B(n_339),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_380),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_437),
.B(n_348),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_388),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_402),
.B(n_369),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_382),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_431),
.B(n_369),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_404),
.Y(n_526)
);

AND3x2_ASAP7_75t_L g527 ( 
.A(n_436),
.B(n_271),
.C(n_269),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_388),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_390),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_388),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_404),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_390),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_435),
.B(n_363),
.Y(n_533)
);

AND2x6_ASAP7_75t_L g534 ( 
.A(n_413),
.B(n_271),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_396),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_398),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_388),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_435),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_398),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_398),
.Y(n_540)
);

NAND2xp33_ASAP7_75t_L g541 ( 
.A(n_398),
.B(n_294),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_396),
.B(n_368),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_382),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_396),
.B(n_370),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_435),
.A2(n_256),
.B1(n_238),
.B2(n_246),
.Y(n_545)
);

OAI21xp33_ASAP7_75t_SL g546 ( 
.A1(n_387),
.A2(n_182),
.B(n_168),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g547 ( 
.A(n_438),
.B(n_307),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_382),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_431),
.B(n_372),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_397),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_398),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_397),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_397),
.Y(n_553)
);

AND2x6_ASAP7_75t_L g554 ( 
.A(n_413),
.B(n_294),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_384),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_398),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_438),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_397),
.Y(n_558)
);

NAND3xp33_ASAP7_75t_L g559 ( 
.A(n_387),
.B(n_373),
.C(n_371),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_396),
.Y(n_560)
);

OR2x2_ASAP7_75t_L g561 ( 
.A(n_389),
.B(n_431),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_396),
.B(n_236),
.Y(n_562)
);

NAND3xp33_ASAP7_75t_L g563 ( 
.A(n_389),
.B(n_174),
.C(n_173),
.Y(n_563)
);

NAND2xp33_ASAP7_75t_SL g564 ( 
.A(n_414),
.B(n_261),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_415),
.B(n_309),
.Y(n_565)
);

OR2x6_ASAP7_75t_L g566 ( 
.A(n_438),
.B(n_246),
.Y(n_566)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_398),
.Y(n_567)
);

NAND3xp33_ASAP7_75t_L g568 ( 
.A(n_413),
.B(n_226),
.C(n_303),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_399),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_384),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_384),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_399),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_386),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_415),
.B(n_416),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_386),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_413),
.B(n_196),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_386),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_395),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_395),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_413),
.B(n_196),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_395),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_430),
.Y(n_582)
);

OR2x6_ASAP7_75t_L g583 ( 
.A(n_393),
.B(n_256),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_419),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_415),
.B(n_372),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_503),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_486),
.B(n_489),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_483),
.B(n_469),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_503),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_487),
.B(n_393),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_483),
.B(n_413),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_469),
.B(n_313),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_L g593 ( 
.A1(n_508),
.A2(n_401),
.B(n_400),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_487),
.B(n_400),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_478),
.B(n_400),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_470),
.B(n_399),
.Y(n_596)
);

INVx2_ASAP7_75t_SL g597 ( 
.A(n_451),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_444),
.Y(n_598)
);

AND2x2_ASAP7_75t_SL g599 ( 
.A(n_453),
.B(n_168),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_470),
.B(n_399),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_474),
.B(n_399),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_474),
.B(n_399),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_515),
.B(n_399),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_515),
.B(n_400),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_508),
.Y(n_605)
);

O2A1O1Ixp5_ASAP7_75t_L g606 ( 
.A1(n_582),
.A2(n_414),
.B(n_430),
.C(n_439),
.Y(n_606)
);

OR2x6_ASAP7_75t_L g607 ( 
.A(n_461),
.B(n_393),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_476),
.Y(n_608)
);

CKINVDCx11_ASAP7_75t_R g609 ( 
.A(n_458),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_461),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_SL g611 ( 
.A(n_459),
.B(n_323),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_526),
.B(n_401),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_526),
.B(n_401),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_504),
.B(n_176),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_531),
.B(n_401),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_468),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_476),
.Y(n_617)
);

OAI22xp33_ASAP7_75t_L g618 ( 
.A1(n_561),
.A2(n_291),
.B1(n_292),
.B2(n_262),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_531),
.B(n_399),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_445),
.B(n_407),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_467),
.B(n_407),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_467),
.B(n_407),
.Y(n_622)
);

BUFx5_ASAP7_75t_L g623 ( 
.A(n_534),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_485),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_445),
.B(n_407),
.Y(n_625)
);

OR2x6_ASAP7_75t_L g626 ( 
.A(n_566),
.B(n_262),
.Y(n_626)
);

A2O1A1Ixp33_ASAP7_75t_L g627 ( 
.A1(n_561),
.A2(n_292),
.B(n_279),
.C(n_280),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_523),
.B(n_414),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_444),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_525),
.Y(n_630)
);

OR2x2_ASAP7_75t_L g631 ( 
.A(n_442),
.B(n_426),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_525),
.B(n_414),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_549),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_447),
.B(n_179),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_523),
.B(n_466),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_585),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_484),
.B(n_414),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_585),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_443),
.B(n_414),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_549),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_443),
.B(n_454),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_467),
.B(n_430),
.Y(n_642)
);

O2A1O1Ixp33_ASAP7_75t_L g643 ( 
.A1(n_538),
.A2(n_439),
.B(n_430),
.C(n_280),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_443),
.B(n_430),
.Y(n_644)
);

NOR2xp67_ASAP7_75t_L g645 ( 
.A(n_559),
.B(n_416),
.Y(n_645)
);

AND2x4_ASAP7_75t_L g646 ( 
.A(n_448),
.B(n_430),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_490),
.B(n_439),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_490),
.B(n_439),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_455),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_565),
.B(n_473),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_582),
.B(n_439),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_457),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_502),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_490),
.B(n_538),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_533),
.B(n_439),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_500),
.B(n_243),
.Y(n_656)
);

OAI21xp33_ASAP7_75t_L g657 ( 
.A1(n_464),
.A2(n_283),
.B(n_297),
.Y(n_657)
);

INVxp67_ASAP7_75t_SL g658 ( 
.A(n_512),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_SL g659 ( 
.A1(n_496),
.A2(n_298),
.B1(n_196),
.B2(n_248),
.Y(n_659)
);

INVx8_ASAP7_75t_L g660 ( 
.A(n_496),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_455),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_472),
.B(n_493),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_583),
.B(n_252),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_571),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_571),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_440),
.B(n_477),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_456),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_SL g668 ( 
.A(n_450),
.B(n_248),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_583),
.B(n_252),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_440),
.B(n_403),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_456),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_477),
.B(n_403),
.Y(n_672)
);

AND2x4_ASAP7_75t_L g673 ( 
.A(n_568),
.B(n_182),
.Y(n_673)
);

OAI22xp5_ASAP7_75t_L g674 ( 
.A1(n_452),
.A2(n_255),
.B1(n_232),
.B2(n_216),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_479),
.B(n_405),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_479),
.B(n_405),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_471),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_521),
.B(n_181),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_480),
.B(n_405),
.Y(n_679)
);

A2O1A1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_545),
.A2(n_283),
.B(n_297),
.C(n_301),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_480),
.B(n_406),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_471),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_502),
.A2(n_301),
.B1(n_185),
.B2(n_273),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_510),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_574),
.B(n_406),
.Y(n_685)
);

NAND2xp33_ASAP7_75t_L g686 ( 
.A(n_475),
.B(n_247),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_488),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_510),
.Y(n_688)
);

OAI221xp5_ASAP7_75t_L g689 ( 
.A1(n_546),
.A2(n_452),
.B1(n_564),
.B2(n_563),
.C(n_516),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_575),
.B(n_406),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_518),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_517),
.B(n_183),
.Y(n_692)
);

OAI221xp5_ASAP7_75t_L g693 ( 
.A1(n_452),
.A2(n_255),
.B1(n_187),
.B2(n_191),
.C(n_203),
.Y(n_693)
);

OAI22xp5_ASAP7_75t_SL g694 ( 
.A1(n_449),
.A2(n_227),
.B1(n_231),
.B2(n_302),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_577),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_578),
.B(n_409),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_495),
.B(n_249),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_583),
.B(n_252),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_518),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_482),
.A2(n_429),
.B(n_419),
.Y(n_700)
);

A2O1A1Ixp33_ASAP7_75t_L g701 ( 
.A1(n_564),
.A2(n_304),
.B(n_185),
.C(n_187),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_497),
.B(n_250),
.Y(n_702)
);

INVxp67_ASAP7_75t_L g703 ( 
.A(n_547),
.Y(n_703)
);

AOI21xp5_ASAP7_75t_L g704 ( 
.A1(n_499),
.A2(n_429),
.B(n_419),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_488),
.Y(n_705)
);

AND2x4_ASAP7_75t_L g706 ( 
.A(n_509),
.B(n_191),
.Y(n_706)
);

AND2x6_ASAP7_75t_L g707 ( 
.A(n_520),
.B(n_203),
.Y(n_707)
);

HB1xp67_ASAP7_75t_L g708 ( 
.A(n_502),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_520),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_519),
.B(n_188),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_583),
.B(n_252),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_579),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_529),
.B(n_251),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_532),
.B(n_254),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_566),
.B(n_192),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_465),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_524),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_535),
.B(n_257),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_566),
.B(n_195),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_524),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_560),
.B(n_259),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_542),
.B(n_417),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_SL g723 ( 
.A(n_450),
.B(n_505),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_496),
.A2(n_289),
.B1(n_263),
.B2(n_266),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_544),
.B(n_417),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_543),
.B(n_417),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_543),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_502),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_475),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_452),
.B(n_206),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_548),
.Y(n_731)
);

NAND2xp33_ASAP7_75t_L g732 ( 
.A(n_475),
.B(n_268),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_548),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_576),
.A2(n_293),
.B1(n_278),
.B2(n_285),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_555),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_555),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_570),
.B(n_290),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_570),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_573),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_492),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_566),
.B(n_434),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_492),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_SL g743 ( 
.A(n_505),
.B(n_248),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_580),
.A2(n_304),
.B1(n_210),
.B2(n_216),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_557),
.B(n_434),
.Y(n_745)
);

BUFx10_ASAP7_75t_L g746 ( 
.A(n_527),
.Y(n_746)
);

A2O1A1Ixp33_ASAP7_75t_L g747 ( 
.A1(n_573),
.A2(n_210),
.B(n_300),
.C(n_284),
.Y(n_747)
);

OR2x6_ASAP7_75t_L g748 ( 
.A(n_562),
.B(n_205),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_579),
.B(n_212),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_581),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_441),
.B(n_417),
.Y(n_751)
);

INVxp67_ASAP7_75t_L g752 ( 
.A(n_557),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_587),
.B(n_534),
.Y(n_753)
);

NOR3xp33_ASAP7_75t_L g754 ( 
.A(n_752),
.B(n_273),
.C(n_232),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_642),
.A2(n_511),
.B(n_460),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_586),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_599),
.A2(n_554),
.B1(n_534),
.B2(n_475),
.Y(n_757)
);

AO21x1_ASAP7_75t_L g758 ( 
.A1(n_674),
.A2(n_205),
.B(n_300),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_599),
.B(n_534),
.Y(n_759)
);

A2O1A1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_657),
.A2(n_284),
.B(n_276),
.C(n_421),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_594),
.B(n_534),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_630),
.B(n_534),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_642),
.A2(n_511),
.B(n_460),
.Y(n_763)
);

OAI21xp5_ASAP7_75t_L g764 ( 
.A1(n_606),
.A2(n_628),
.B(n_591),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_595),
.B(n_554),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_589),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_590),
.B(n_441),
.Y(n_767)
);

O2A1O1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_588),
.A2(n_541),
.B(n_276),
.C(n_584),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_647),
.A2(n_511),
.B(n_460),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_623),
.B(n_441),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_647),
.A2(n_567),
.B(n_462),
.Y(n_771)
);

AOI21x1_ASAP7_75t_L g772 ( 
.A1(n_621),
.A2(n_552),
.B(n_528),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_609),
.Y(n_773)
);

OAI21xp5_ASAP7_75t_L g774 ( 
.A1(n_639),
.A2(n_491),
.B(n_463),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_623),
.B(n_446),
.Y(n_775)
);

BUFx4f_ASAP7_75t_L g776 ( 
.A(n_607),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_623),
.B(n_446),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_706),
.B(n_554),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_706),
.B(n_554),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_648),
.A2(n_567),
.B(n_462),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_605),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_683),
.A2(n_554),
.B1(n_475),
.B2(n_481),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_R g783 ( 
.A(n_723),
.B(n_554),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_695),
.Y(n_784)
);

BUFx3_ASAP7_75t_L g785 ( 
.A(n_652),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_648),
.A2(n_567),
.B(n_462),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_695),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_722),
.A2(n_539),
.B(n_572),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_632),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_632),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_725),
.A2(n_539),
.B(n_572),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_636),
.B(n_475),
.Y(n_792)
);

OAI21xp5_ASAP7_75t_L g793 ( 
.A1(n_593),
.A2(n_463),
.B(n_491),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_650),
.B(n_446),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_623),
.B(n_463),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_616),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_638),
.B(n_481),
.Y(n_797)
);

BUFx4f_ASAP7_75t_L g798 ( 
.A(n_607),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_655),
.A2(n_512),
.B(n_572),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_684),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_635),
.B(n_481),
.Y(n_801)
);

A2O1A1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_627),
.A2(n_416),
.B(n_418),
.C(n_421),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_655),
.A2(n_512),
.B(n_572),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_641),
.A2(n_658),
.B(n_644),
.Y(n_804)
);

OAI21xp5_ASAP7_75t_L g805 ( 
.A1(n_588),
.A2(n_651),
.B(n_625),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_633),
.B(n_481),
.Y(n_806)
);

AO21x1_ASAP7_75t_L g807 ( 
.A1(n_654),
.A2(n_541),
.B(n_584),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_621),
.A2(n_572),
.B(n_569),
.Y(n_808)
);

AOI21xp33_ASAP7_75t_L g809 ( 
.A1(n_678),
.A2(n_244),
.B(n_220),
.Y(n_809)
);

INVx1_ASAP7_75t_SL g810 ( 
.A(n_592),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_623),
.B(n_491),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_729),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_617),
.A2(n_481),
.B1(n_536),
.B2(n_540),
.Y(n_813)
);

INVx3_ASAP7_75t_L g814 ( 
.A(n_608),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_712),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_622),
.A2(n_569),
.B(n_512),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_688),
.Y(n_817)
);

AO21x1_ASAP7_75t_L g818 ( 
.A1(n_654),
.A2(n_513),
.B(n_553),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_622),
.A2(n_569),
.B(n_512),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_619),
.A2(n_569),
.B(n_556),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_640),
.B(n_481),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_624),
.A2(n_536),
.B1(n_540),
.B2(n_551),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_623),
.B(n_536),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_691),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_666),
.B(n_540),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_620),
.A2(n_551),
.B(n_553),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_699),
.B(n_709),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_646),
.B(n_418),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_619),
.A2(n_556),
.B(n_539),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_SL g830 ( 
.A(n_611),
.B(n_248),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_612),
.A2(n_556),
.B(n_539),
.Y(n_831)
);

BUFx2_ASAP7_75t_L g832 ( 
.A(n_607),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_717),
.B(n_551),
.Y(n_833)
);

AOI21x1_ASAP7_75t_L g834 ( 
.A1(n_596),
.A2(n_558),
.B(n_494),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_720),
.B(n_539),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_613),
.A2(n_556),
.B(n_507),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_727),
.B(n_558),
.Y(n_837)
);

AO21x1_ASAP7_75t_L g838 ( 
.A1(n_678),
.A2(n_552),
.B(n_550),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_637),
.A2(n_550),
.B(n_537),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_700),
.A2(n_537),
.B(n_530),
.Y(n_840)
);

NOR2x1_ASAP7_75t_L g841 ( 
.A(n_652),
.B(n_530),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_731),
.B(n_494),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_608),
.B(n_498),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_729),
.A2(n_528),
.B1(n_522),
.B2(n_514),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_662),
.B(n_498),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_733),
.B(n_522),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_615),
.A2(n_507),
.B(n_513),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_645),
.B(n_501),
.Y(n_848)
);

HB1xp67_ASAP7_75t_L g849 ( 
.A(n_610),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_735),
.Y(n_850)
);

NAND3xp33_ASAP7_75t_L g851 ( 
.A(n_692),
.B(n_275),
.C(n_222),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_703),
.B(n_221),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_604),
.A2(n_507),
.B(n_506),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_745),
.B(n_225),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_736),
.Y(n_855)
);

A2O1A1Ixp33_ASAP7_75t_L g856 ( 
.A1(n_627),
.A2(n_434),
.B(n_421),
.C(n_418),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_L g857 ( 
.A1(n_683),
.A2(n_274),
.B1(n_234),
.B2(n_237),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_664),
.Y(n_858)
);

AO21x1_ASAP7_75t_L g859 ( 
.A1(n_737),
.A2(n_419),
.B(n_429),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_738),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_634),
.B(n_229),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_596),
.A2(n_507),
.B(n_429),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_600),
.A2(n_507),
.B(n_427),
.Y(n_863)
);

INVxp67_ASAP7_75t_L g864 ( 
.A(n_634),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_653),
.B(n_708),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_739),
.Y(n_866)
);

INVxp33_ASAP7_75t_SL g867 ( 
.A(n_668),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_653),
.B(n_241),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_744),
.B(n_427),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_750),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_749),
.B(n_427),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_600),
.A2(n_427),
.B(n_424),
.Y(n_872)
);

A2O1A1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_701),
.A2(n_282),
.B(n_245),
.C(n_253),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_601),
.A2(n_427),
.B(n_424),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_749),
.B(n_427),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_664),
.Y(n_876)
);

AOI21x1_ASAP7_75t_L g877 ( 
.A1(n_601),
.A2(n_602),
.B(n_603),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_741),
.B(n_287),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_665),
.B(n_427),
.Y(n_879)
);

INVx11_ASAP7_75t_L g880 ( 
.A(n_707),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_602),
.A2(n_427),
.B(n_424),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_685),
.B(n_673),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_665),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_603),
.A2(n_424),
.B(n_423),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_663),
.B(n_286),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_669),
.B(n_272),
.Y(n_886)
);

A2O1A1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_701),
.A2(n_295),
.B(n_258),
.C(n_267),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_598),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_673),
.B(n_424),
.Y(n_889)
);

AOI22x1_ASAP7_75t_SL g890 ( 
.A1(n_659),
.A2(n_242),
.B1(n_270),
.B2(n_299),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_646),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_751),
.A2(n_424),
.B(n_423),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_660),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_686),
.A2(n_424),
.B(n_423),
.Y(n_894)
);

NOR3xp33_ASAP7_75t_L g895 ( 
.A(n_692),
.B(n_15),
.C(n_17),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_708),
.A2(n_424),
.B1(n_423),
.B2(n_417),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_732),
.A2(n_423),
.B(n_417),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_698),
.B(n_423),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_629),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_737),
.B(n_423),
.Y(n_900)
);

OAI21xp5_ASAP7_75t_L g901 ( 
.A1(n_704),
.A2(n_423),
.B(n_417),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_670),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_614),
.B(n_18),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_614),
.B(n_19),
.Y(n_904)
);

BUFx3_ASAP7_75t_L g905 ( 
.A(n_660),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_748),
.B(n_20),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_730),
.B(n_68),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_689),
.A2(n_66),
.B1(n_145),
.B2(n_144),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_649),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_726),
.A2(n_61),
.B(n_143),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_730),
.B(n_149),
.Y(n_911)
);

INVxp67_ASAP7_75t_L g912 ( 
.A(n_597),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_SL g913 ( 
.A1(n_631),
.A2(n_23),
.B1(n_28),
.B2(n_31),
.Y(n_913)
);

NOR3xp33_ASAP7_75t_L g914 ( 
.A(n_710),
.B(n_23),
.C(n_28),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_697),
.A2(n_141),
.B(n_127),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_672),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_661),
.Y(n_917)
);

O2A1O1Ixp5_ASAP7_75t_L g918 ( 
.A1(n_697),
.A2(n_119),
.B(n_112),
.C(n_110),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_711),
.B(n_31),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_748),
.B(n_33),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_728),
.B(n_34),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_675),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_702),
.A2(n_108),
.B(n_100),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_728),
.B(n_93),
.Y(n_924)
);

OAI21xp5_ASAP7_75t_L g925 ( 
.A1(n_643),
.A2(n_71),
.B(n_69),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_748),
.B(n_35),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_693),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_713),
.A2(n_37),
.B(n_39),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_676),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_667),
.A2(n_39),
.B(n_40),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_710),
.B(n_43),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_671),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_677),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_715),
.B(n_43),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_787),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_804),
.A2(n_714),
.B(n_713),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_864),
.B(n_743),
.Y(n_937)
);

AO22x1_ASAP7_75t_L g938 ( 
.A1(n_931),
.A2(n_716),
.B1(n_707),
.B2(n_618),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_902),
.B(n_681),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_796),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_916),
.B(n_679),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_867),
.B(n_719),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_922),
.B(n_690),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_753),
.A2(n_761),
.B(n_764),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_849),
.Y(n_945)
);

NAND2xp33_ASAP7_75t_SL g946 ( 
.A(n_783),
.B(n_656),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_929),
.B(n_696),
.Y(n_947)
);

CKINVDCx11_ASAP7_75t_R g948 ( 
.A(n_832),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_756),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_810),
.B(n_626),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_854),
.B(n_626),
.Y(n_951)
);

OAI22x1_ASAP7_75t_L g952 ( 
.A1(n_931),
.A2(n_724),
.B1(n_626),
.B2(n_656),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_903),
.A2(n_714),
.B(n_718),
.C(n_721),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_882),
.B(n_707),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_785),
.B(n_660),
.Y(n_955)
);

NOR3xp33_ASAP7_75t_SL g956 ( 
.A(n_913),
.B(n_773),
.C(n_694),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_854),
.B(n_618),
.Y(n_957)
);

AOI21x1_ASAP7_75t_L g958 ( 
.A1(n_871),
.A2(n_718),
.B(n_742),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_765),
.A2(n_687),
.B(n_740),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_778),
.A2(n_682),
.B(n_705),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_893),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_794),
.B(n_707),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_794),
.B(n_707),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_785),
.B(n_734),
.Y(n_964)
);

NAND2x1p5_ASAP7_75t_L g965 ( 
.A(n_812),
.B(n_747),
.Y(n_965)
);

O2A1O1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_904),
.A2(n_680),
.B(n_747),
.C(n_746),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_878),
.B(n_746),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_809),
.A2(n_680),
.B(n_45),
.C(n_50),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_779),
.A2(n_44),
.B(n_50),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_766),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_801),
.A2(n_44),
.B(n_53),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_875),
.A2(n_53),
.B(n_805),
.Y(n_972)
);

AOI22xp33_ASAP7_75t_L g973 ( 
.A1(n_934),
.A2(n_907),
.B1(n_911),
.B2(n_924),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_SL g974 ( 
.A(n_830),
.B(n_776),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_850),
.B(n_855),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_SL g976 ( 
.A1(n_934),
.A2(n_925),
.B(n_852),
.C(n_767),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_781),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_905),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_755),
.A2(n_769),
.B(n_763),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_776),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_850),
.B(n_855),
.Y(n_981)
);

NOR2x1_ASAP7_75t_L g982 ( 
.A(n_905),
.B(n_851),
.Y(n_982)
);

BUFx8_ASAP7_75t_L g983 ( 
.A(n_919),
.Y(n_983)
);

AOI22xp5_ASAP7_75t_L g984 ( 
.A1(n_861),
.A2(n_891),
.B1(n_789),
.B2(n_790),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_860),
.B(n_866),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_852),
.A2(n_759),
.B(n_866),
.C(n_860),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_812),
.Y(n_987)
);

BUFx2_ASAP7_75t_L g988 ( 
.A(n_798),
.Y(n_988)
);

OR2x6_ASAP7_75t_L g989 ( 
.A(n_812),
.B(n_762),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_812),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_800),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_891),
.B(n_783),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_885),
.B(n_886),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_817),
.Y(n_994)
);

OAI21xp33_ASAP7_75t_L g995 ( 
.A1(n_868),
.A2(n_857),
.B(n_906),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_771),
.A2(n_780),
.B(n_786),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_828),
.B(n_762),
.Y(n_997)
);

NOR3xp33_ASAP7_75t_L g998 ( 
.A(n_920),
.B(n_926),
.C(n_912),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_L g999 ( 
.A1(n_782),
.A2(n_757),
.B1(n_827),
.B2(n_814),
.Y(n_999)
);

NAND3xp33_ASAP7_75t_SL g1000 ( 
.A(n_895),
.B(n_914),
.C(n_754),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_798),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_814),
.Y(n_1002)
);

AOI22xp33_ASAP7_75t_L g1003 ( 
.A1(n_907),
.A2(n_911),
.B1(n_924),
.B2(n_828),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_782),
.A2(n_896),
.B1(n_767),
.B2(n_824),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_898),
.B(n_841),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_774),
.A2(n_797),
.B(n_792),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_784),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_896),
.A2(n_865),
.B1(n_813),
.B2(n_821),
.Y(n_1008)
);

OAI21xp33_ASAP7_75t_L g1009 ( 
.A1(n_868),
.A2(n_930),
.B(n_865),
.Y(n_1009)
);

INVx6_ASAP7_75t_L g1010 ( 
.A(n_845),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_788),
.A2(n_791),
.B(n_826),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_845),
.B(n_825),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_921),
.B(n_890),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_806),
.A2(n_858),
.B1(n_870),
.B2(n_835),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_908),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_815),
.Y(n_1016)
);

NOR2xp67_ASAP7_75t_SL g1017 ( 
.A(n_910),
.B(n_858),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_799),
.A2(n_803),
.B(n_811),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_876),
.B(n_883),
.Y(n_1019)
);

AOI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_921),
.A2(n_889),
.B1(n_848),
.B2(n_917),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_888),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_770),
.A2(n_775),
.B(n_823),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_889),
.B(n_909),
.Y(n_1023)
);

AO32x1_ASAP7_75t_L g1024 ( 
.A1(n_927),
.A2(n_844),
.A3(n_838),
.B1(n_888),
.B2(n_932),
.Y(n_1024)
);

O2A1O1Ixp33_ASAP7_75t_SL g1025 ( 
.A1(n_873),
.A2(n_887),
.B(n_856),
.C(n_802),
.Y(n_1025)
);

AO31x2_ASAP7_75t_L g1026 ( 
.A1(n_807),
.A2(n_859),
.A3(n_818),
.B(n_758),
.Y(n_1026)
);

AOI22xp33_ASAP7_75t_L g1027 ( 
.A1(n_928),
.A2(n_933),
.B1(n_899),
.B2(n_932),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_899),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_933),
.B(n_848),
.Y(n_1029)
);

AOI21x1_ASAP7_75t_L g1030 ( 
.A1(n_772),
.A2(n_900),
.B(n_877),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_837),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_770),
.A2(n_823),
.B(n_795),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_873),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_SL g1034 ( 
.A1(n_833),
.A2(n_842),
.B1(n_846),
.B2(n_822),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_887),
.B(n_760),
.Y(n_1035)
);

INVx3_ASAP7_75t_SL g1036 ( 
.A(n_869),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_775),
.A2(n_811),
.B(n_777),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_880),
.A2(n_793),
.B1(n_777),
.B2(n_795),
.Y(n_1038)
);

AO21x2_ASAP7_75t_L g1039 ( 
.A1(n_901),
.A2(n_840),
.B(n_839),
.Y(n_1039)
);

BUFx8_ASAP7_75t_SL g1040 ( 
.A(n_834),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_768),
.A2(n_918),
.B(n_915),
.C(n_923),
.Y(n_1041)
);

AOI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_843),
.A2(n_879),
.B1(n_869),
.B2(n_808),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_802),
.B(n_856),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_831),
.A2(n_816),
.B(n_819),
.Y(n_1044)
);

CKINVDCx16_ASAP7_75t_R g1045 ( 
.A(n_760),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_879),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_820),
.B(n_829),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_872),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_853),
.B(n_847),
.Y(n_1049)
);

BUFx2_ASAP7_75t_L g1050 ( 
.A(n_874),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_881),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_884),
.A2(n_862),
.B(n_836),
.C(n_892),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_863),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_894),
.B(n_897),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_931),
.A2(n_599),
.B1(n_587),
.B2(n_903),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_902),
.B(n_587),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_785),
.B(n_905),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_931),
.A2(n_587),
.B(n_599),
.C(n_453),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_SL g1059 ( 
.A(n_773),
.B(n_450),
.Y(n_1059)
);

INVx4_ASAP7_75t_L g1060 ( 
.A(n_812),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_804),
.A2(n_490),
.B(n_467),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_902),
.B(n_587),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_787),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_756),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_864),
.B(n_587),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_854),
.B(n_650),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_902),
.B(n_587),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_882),
.A2(n_587),
.B1(n_599),
.B2(n_864),
.Y(n_1068)
);

OAI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_764),
.A2(n_587),
.B(n_805),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_864),
.B(n_587),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_854),
.B(n_650),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_854),
.B(n_650),
.Y(n_1072)
);

NOR2xp67_ASAP7_75t_SL g1073 ( 
.A(n_785),
.B(n_587),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_902),
.B(n_587),
.Y(n_1074)
);

INVx3_ASAP7_75t_SL g1075 ( 
.A(n_773),
.Y(n_1075)
);

INVx4_ASAP7_75t_L g1076 ( 
.A(n_987),
.Y(n_1076)
);

INVx2_ASAP7_75t_SL g1077 ( 
.A(n_940),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1056),
.B(n_1062),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_1060),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_979),
.A2(n_996),
.B(n_1018),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1061),
.A2(n_1069),
.B(n_944),
.Y(n_1081)
);

NOR2x1_ASAP7_75t_SL g1082 ( 
.A(n_989),
.B(n_992),
.Y(n_1082)
);

O2A1O1Ixp33_ASAP7_75t_SL g1083 ( 
.A1(n_1058),
.A2(n_976),
.B(n_953),
.C(n_986),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_SL g1084 ( 
.A(n_957),
.B(n_974),
.Y(n_1084)
);

AOI22x1_ASAP7_75t_L g1085 ( 
.A1(n_952),
.A2(n_972),
.B1(n_936),
.B2(n_1033),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_1055),
.A2(n_1056),
.B1(n_1074),
.B2(n_1062),
.Y(n_1086)
);

AO31x2_ASAP7_75t_L g1087 ( 
.A1(n_972),
.A2(n_1011),
.A3(n_1044),
.B(n_1041),
.Y(n_1087)
);

O2A1O1Ixp5_ASAP7_75t_L g1088 ( 
.A1(n_1073),
.A2(n_1017),
.B(n_1049),
.C(n_937),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_1066),
.B(n_1071),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_949),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_1011),
.A2(n_1039),
.B(n_1047),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1039),
.A2(n_1047),
.B(n_1067),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_1072),
.B(n_1067),
.Y(n_1093)
);

OR2x2_ASAP7_75t_L g1094 ( 
.A(n_1074),
.B(n_945),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_973),
.A2(n_1068),
.B(n_962),
.Y(n_1095)
);

NAND2x1_ASAP7_75t_L g1096 ( 
.A(n_1060),
.B(n_989),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_1044),
.A2(n_1030),
.B(n_959),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_950),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_993),
.B(n_942),
.Y(n_1099)
);

OR2x2_ASAP7_75t_L g1100 ( 
.A(n_1065),
.B(n_1070),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_961),
.Y(n_1101)
);

AO21x1_ASAP7_75t_L g1102 ( 
.A1(n_946),
.A2(n_962),
.B(n_963),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_1075),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_963),
.A2(n_1006),
.B(n_999),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_939),
.A2(n_941),
.B(n_943),
.Y(n_1105)
);

NAND3x1_ASAP7_75t_L g1106 ( 
.A(n_1013),
.B(n_982),
.C(n_998),
.Y(n_1106)
);

NAND2x1p5_ASAP7_75t_L g1107 ( 
.A(n_1057),
.B(n_987),
.Y(n_1107)
);

AOI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_1015),
.A2(n_995),
.B1(n_1000),
.B2(n_1009),
.Y(n_1108)
);

OAI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_1059),
.A2(n_1045),
.B1(n_984),
.B2(n_951),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_SL g1110 ( 
.A1(n_1043),
.A2(n_1003),
.B(n_971),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1043),
.A2(n_1042),
.B(n_954),
.Y(n_1111)
);

AO22x2_ASAP7_75t_L g1112 ( 
.A1(n_1004),
.A2(n_1035),
.B1(n_1008),
.B2(n_1038),
.Y(n_1112)
);

AO31x2_ASAP7_75t_L g1113 ( 
.A1(n_1014),
.A2(n_1050),
.A3(n_1048),
.B(n_1032),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_943),
.B(n_947),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_939),
.A2(n_941),
.B(n_947),
.Y(n_1115)
);

AO31x2_ASAP7_75t_L g1116 ( 
.A1(n_1022),
.A2(n_1037),
.A3(n_954),
.B(n_1053),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_1057),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_1052),
.A2(n_958),
.B(n_960),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_978),
.Y(n_1119)
);

OR2x6_ASAP7_75t_L g1120 ( 
.A(n_989),
.B(n_988),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_965),
.A2(n_1012),
.B(n_975),
.Y(n_1121)
);

CKINVDCx11_ASAP7_75t_R g1122 ( 
.A(n_948),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_968),
.A2(n_964),
.B(n_966),
.C(n_956),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_987),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_965),
.A2(n_1012),
.B(n_985),
.Y(n_1125)
);

NOR2x1_ASAP7_75t_SL g1126 ( 
.A(n_975),
.B(n_985),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_1020),
.A2(n_981),
.B1(n_1031),
.B2(n_994),
.Y(n_1127)
);

BUFx3_ASAP7_75t_L g1128 ( 
.A(n_978),
.Y(n_1128)
);

AOI222xp33_ASAP7_75t_L g1129 ( 
.A1(n_938),
.A2(n_1064),
.B1(n_991),
.B2(n_977),
.C1(n_970),
.C2(n_967),
.Y(n_1129)
);

INVx5_ASAP7_75t_L g1130 ( 
.A(n_990),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1063),
.Y(n_1131)
);

INVx2_ASAP7_75t_SL g1132 ( 
.A(n_978),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1005),
.B(n_1023),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1034),
.A2(n_1051),
.B(n_1025),
.Y(n_1134)
);

AOI221x1_ASAP7_75t_L g1135 ( 
.A1(n_969),
.A2(n_1005),
.B1(n_1029),
.B2(n_1046),
.C(n_1024),
.Y(n_1135)
);

OAI22x1_ASAP7_75t_L g1136 ( 
.A1(n_1036),
.A2(n_980),
.B1(n_1001),
.B2(n_955),
.Y(n_1136)
);

OAI22x1_ASAP7_75t_L g1137 ( 
.A1(n_1029),
.A2(n_1016),
.B1(n_1007),
.B2(n_997),
.Y(n_1137)
);

AO32x2_ASAP7_75t_L g1138 ( 
.A1(n_1024),
.A2(n_1026),
.A3(n_1040),
.B1(n_1010),
.B2(n_1027),
.Y(n_1138)
);

BUFx4f_ASAP7_75t_L g1139 ( 
.A(n_990),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_990),
.B(n_1028),
.Y(n_1140)
);

BUFx2_ASAP7_75t_R g1141 ( 
.A(n_1002),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1028),
.B(n_1021),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1024),
.A2(n_1019),
.B(n_1002),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_983),
.B(n_1010),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_983),
.B(n_1026),
.Y(n_1145)
);

AO21x1_ASAP7_75t_L g1146 ( 
.A1(n_957),
.A2(n_931),
.B(n_587),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1061),
.A2(n_587),
.B(n_1069),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1061),
.A2(n_587),
.B(n_1069),
.Y(n_1148)
);

AO31x2_ASAP7_75t_L g1149 ( 
.A1(n_972),
.A2(n_838),
.A3(n_1058),
.B(n_1011),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1056),
.B(n_587),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1056),
.B(n_587),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_961),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_979),
.A2(n_996),
.B(n_1018),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_978),
.Y(n_1154)
);

INVx2_ASAP7_75t_SL g1155 ( 
.A(n_940),
.Y(n_1155)
);

INVxp67_ASAP7_75t_SL g1156 ( 
.A(n_945),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_1058),
.A2(n_587),
.B(n_957),
.C(n_931),
.Y(n_1157)
);

AO31x2_ASAP7_75t_L g1158 ( 
.A1(n_972),
.A2(n_838),
.A3(n_1058),
.B(n_1011),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1061),
.A2(n_587),
.B(n_1069),
.Y(n_1159)
);

OA21x2_ASAP7_75t_L g1160 ( 
.A1(n_972),
.A2(n_944),
.B(n_1011),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1056),
.B(n_587),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_945),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1058),
.A2(n_587),
.B1(n_1055),
.B2(n_957),
.Y(n_1163)
);

AOI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_957),
.A2(n_587),
.B1(n_931),
.B2(n_599),
.Y(n_1164)
);

AOI221x1_ASAP7_75t_L g1165 ( 
.A1(n_1058),
.A2(n_931),
.B1(n_587),
.B2(n_1009),
.C(n_957),
.Y(n_1165)
);

AOI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1017),
.A2(n_1054),
.B(n_963),
.Y(n_1166)
);

OAI22x1_ASAP7_75t_L g1167 ( 
.A1(n_957),
.A2(n_931),
.B1(n_1013),
.B2(n_951),
.Y(n_1167)
);

AO31x2_ASAP7_75t_L g1168 ( 
.A1(n_972),
.A2(n_838),
.A3(n_1058),
.B(n_1011),
.Y(n_1168)
);

CKINVDCx11_ASAP7_75t_R g1169 ( 
.A(n_1075),
.Y(n_1169)
);

AO31x2_ASAP7_75t_L g1170 ( 
.A1(n_972),
.A2(n_838),
.A3(n_1058),
.B(n_1011),
.Y(n_1170)
);

OAI22x1_ASAP7_75t_L g1171 ( 
.A1(n_957),
.A2(n_931),
.B1(n_1013),
.B2(n_951),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1058),
.A2(n_587),
.B(n_957),
.C(n_931),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_949),
.Y(n_1173)
);

INVx2_ASAP7_75t_SL g1174 ( 
.A(n_940),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1061),
.A2(n_587),
.B(n_1069),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1061),
.A2(n_587),
.B(n_1069),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1058),
.A2(n_587),
.B1(n_1055),
.B2(n_957),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1056),
.B(n_587),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_978),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_1058),
.A2(n_587),
.B(n_957),
.C(n_931),
.Y(n_1180)
);

INVx1_ASAP7_75t_SL g1181 ( 
.A(n_945),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_949),
.Y(n_1182)
);

INVx3_ASAP7_75t_L g1183 ( 
.A(n_1060),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_979),
.A2(n_996),
.B(n_1018),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1061),
.A2(n_587),
.B(n_1069),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1058),
.A2(n_587),
.B(n_957),
.C(n_931),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_1066),
.B(n_587),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_979),
.A2(n_996),
.B(n_1018),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_979),
.A2(n_996),
.B(n_1018),
.Y(n_1189)
);

NAND3xp33_ASAP7_75t_L g1190 ( 
.A(n_1058),
.B(n_587),
.C(n_1055),
.Y(n_1190)
);

INVx6_ASAP7_75t_L g1191 ( 
.A(n_978),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1061),
.A2(n_587),
.B(n_1069),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1058),
.A2(n_1069),
.B(n_1055),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1066),
.B(n_1071),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_SL g1195 ( 
.A1(n_1058),
.A2(n_976),
.B(n_911),
.C(n_907),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1058),
.A2(n_587),
.B1(n_1055),
.B2(n_957),
.Y(n_1196)
);

A2O1A1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1058),
.A2(n_587),
.B(n_957),
.C(n_931),
.Y(n_1197)
);

OR2x2_ASAP7_75t_L g1198 ( 
.A(n_1056),
.B(n_590),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1061),
.A2(n_587),
.B(n_1069),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_SL g1200 ( 
.A(n_957),
.B(n_599),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_979),
.A2(n_996),
.B(n_1018),
.Y(n_1201)
);

A2O1A1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1058),
.A2(n_587),
.B(n_957),
.C(n_931),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1056),
.B(n_587),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1061),
.A2(n_587),
.B(n_1069),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_945),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1058),
.A2(n_1069),
.B(n_1055),
.Y(n_1206)
);

CKINVDCx11_ASAP7_75t_R g1207 ( 
.A(n_1075),
.Y(n_1207)
);

CKINVDCx14_ASAP7_75t_R g1208 ( 
.A(n_948),
.Y(n_1208)
);

AOI221x1_ASAP7_75t_L g1209 ( 
.A1(n_1058),
.A2(n_931),
.B1(n_587),
.B2(n_1009),
.C(n_957),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1056),
.B(n_587),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_935),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1056),
.B(n_587),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_979),
.A2(n_996),
.B(n_1018),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1056),
.B(n_587),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_SL g1215 ( 
.A1(n_1084),
.A2(n_1200),
.B1(n_1163),
.B2(n_1196),
.Y(n_1215)
);

CKINVDCx11_ASAP7_75t_R g1216 ( 
.A(n_1169),
.Y(n_1216)
);

INVx6_ASAP7_75t_L g1217 ( 
.A(n_1130),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_1191),
.Y(n_1218)
);

BUFx12f_ASAP7_75t_L g1219 ( 
.A(n_1122),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_1128),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_SL g1221 ( 
.A1(n_1084),
.A2(n_1200),
.B1(n_1177),
.B2(n_1190),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1164),
.A2(n_1167),
.B1(n_1171),
.B2(n_1190),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_1207),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_1179),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1164),
.A2(n_1108),
.B1(n_1193),
.B2(n_1206),
.Y(n_1225)
);

INVx6_ASAP7_75t_L g1226 ( 
.A(n_1130),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1108),
.A2(n_1193),
.B1(n_1206),
.B2(n_1146),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1187),
.A2(n_1093),
.B1(n_1089),
.B2(n_1194),
.Y(n_1228)
);

CKINVDCx20_ASAP7_75t_R g1229 ( 
.A(n_1103),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1112),
.A2(n_1086),
.B1(n_1109),
.B2(n_1095),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1150),
.B(n_1151),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1112),
.A2(n_1086),
.B1(n_1095),
.B2(n_1134),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1161),
.A2(n_1214),
.B1(n_1212),
.B2(n_1210),
.Y(n_1233)
);

OAI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1178),
.A2(n_1203),
.B1(n_1165),
.B2(n_1209),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1099),
.B(n_1198),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1110),
.A2(n_1129),
.B1(n_1114),
.B2(n_1115),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1129),
.A2(n_1105),
.B1(n_1078),
.B2(n_1085),
.Y(n_1237)
);

BUFx4_ASAP7_75t_SL g1238 ( 
.A(n_1101),
.Y(n_1238)
);

INVx6_ASAP7_75t_L g1239 ( 
.A(n_1130),
.Y(n_1239)
);

CKINVDCx11_ASAP7_75t_R g1240 ( 
.A(n_1181),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1094),
.B(n_1157),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1173),
.Y(n_1242)
);

INVx6_ASAP7_75t_L g1243 ( 
.A(n_1119),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1182),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1211),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_SL g1246 ( 
.A1(n_1082),
.A2(n_1098),
.B1(n_1145),
.B2(n_1156),
.Y(n_1246)
);

BUFx4f_ASAP7_75t_SL g1247 ( 
.A(n_1144),
.Y(n_1247)
);

INVx1_ASAP7_75t_SL g1248 ( 
.A(n_1181),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1131),
.Y(n_1249)
);

AOI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1106),
.A2(n_1180),
.B1(n_1172),
.B2(n_1197),
.Y(n_1250)
);

CKINVDCx11_ASAP7_75t_R g1251 ( 
.A(n_1119),
.Y(n_1251)
);

CKINVDCx11_ASAP7_75t_R g1252 ( 
.A(n_1119),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1142),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1104),
.A2(n_1100),
.B1(n_1111),
.B2(n_1127),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1104),
.A2(n_1111),
.B1(n_1127),
.B2(n_1102),
.Y(n_1255)
);

HB1xp67_ASAP7_75t_L g1256 ( 
.A(n_1162),
.Y(n_1256)
);

OAI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1120),
.A2(n_1133),
.B1(n_1136),
.B2(n_1174),
.Y(n_1257)
);

BUFx8_ASAP7_75t_L g1258 ( 
.A(n_1117),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1140),
.Y(n_1259)
);

BUFx3_ASAP7_75t_L g1260 ( 
.A(n_1191),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1147),
.A2(n_1199),
.B1(n_1185),
.B2(n_1176),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1148),
.A2(n_1159),
.B1(n_1175),
.B2(n_1204),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1202),
.B(n_1186),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1123),
.B(n_1077),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1155),
.B(n_1205),
.Y(n_1265)
);

INVx4_ASAP7_75t_L g1266 ( 
.A(n_1154),
.Y(n_1266)
);

INVx6_ASAP7_75t_L g1267 ( 
.A(n_1154),
.Y(n_1267)
);

AOI21xp33_ASAP7_75t_L g1268 ( 
.A1(n_1088),
.A2(n_1137),
.B(n_1192),
.Y(n_1268)
);

CKINVDCx20_ASAP7_75t_R g1269 ( 
.A(n_1152),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_SL g1270 ( 
.A1(n_1208),
.A2(n_1126),
.B1(n_1120),
.B2(n_1141),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1120),
.A2(n_1107),
.B1(n_1139),
.B2(n_1096),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1121),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1139),
.A2(n_1092),
.B1(n_1132),
.B2(n_1079),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1160),
.A2(n_1091),
.B1(n_1081),
.B2(n_1125),
.Y(n_1274)
);

CKINVDCx6p67_ASAP7_75t_R g1275 ( 
.A(n_1076),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1140),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1124),
.Y(n_1277)
);

CKINVDCx20_ASAP7_75t_R g1278 ( 
.A(n_1076),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_1183),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1183),
.Y(n_1280)
);

CKINVDCx20_ASAP7_75t_R g1281 ( 
.A(n_1143),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_SL g1282 ( 
.A1(n_1160),
.A2(n_1195),
.B1(n_1083),
.B2(n_1138),
.Y(n_1282)
);

BUFx8_ASAP7_75t_L g1283 ( 
.A(n_1138),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1080),
.A2(n_1213),
.B1(n_1184),
.B2(n_1201),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1087),
.Y(n_1285)
);

AOI21xp33_ASAP7_75t_L g1286 ( 
.A1(n_1153),
.A2(n_1189),
.B(n_1188),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1113),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1097),
.A2(n_1118),
.B1(n_1138),
.B2(n_1170),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1113),
.Y(n_1289)
);

OAI21xp33_ASAP7_75t_L g1290 ( 
.A1(n_1166),
.A2(n_1135),
.B(n_1170),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1149),
.B(n_1158),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_SL g1292 ( 
.A1(n_1149),
.A2(n_1158),
.B1(n_1168),
.B2(n_1170),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1149),
.B(n_1158),
.Y(n_1293)
);

BUFx3_ASAP7_75t_L g1294 ( 
.A(n_1116),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1168),
.A2(n_1116),
.B1(n_957),
.B2(n_1200),
.Y(n_1295)
);

BUFx12f_ASAP7_75t_L g1296 ( 
.A(n_1168),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1090),
.Y(n_1297)
);

INVx6_ASAP7_75t_L g1298 ( 
.A(n_1130),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_SL g1299 ( 
.A1(n_1084),
.A2(n_611),
.B1(n_1200),
.B2(n_830),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1187),
.B(n_1093),
.Y(n_1300)
);

BUFx12f_ASAP7_75t_L g1301 ( 
.A(n_1122),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_SL g1302 ( 
.A1(n_1084),
.A2(n_611),
.B1(n_1200),
.B2(n_830),
.Y(n_1302)
);

INVx6_ASAP7_75t_L g1303 ( 
.A(n_1130),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1200),
.A2(n_957),
.B1(n_599),
.B2(n_1164),
.Y(n_1304)
);

BUFx8_ASAP7_75t_L g1305 ( 
.A(n_1117),
.Y(n_1305)
);

CKINVDCx11_ASAP7_75t_R g1306 ( 
.A(n_1169),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_SL g1307 ( 
.A1(n_1084),
.A2(n_611),
.B1(n_1200),
.B2(n_830),
.Y(n_1307)
);

BUFx12f_ASAP7_75t_L g1308 ( 
.A(n_1169),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1187),
.B(n_1093),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1164),
.A2(n_587),
.B1(n_1058),
.B2(n_957),
.Y(n_1310)
);

INVxp67_ASAP7_75t_L g1311 ( 
.A(n_1162),
.Y(n_1311)
);

INVx3_ASAP7_75t_L g1312 ( 
.A(n_1140),
.Y(n_1312)
);

CKINVDCx11_ASAP7_75t_R g1313 ( 
.A(n_1169),
.Y(n_1313)
);

AOI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1084),
.A2(n_611),
.B1(n_957),
.B2(n_1200),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1090),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_SL g1316 ( 
.A1(n_1167),
.A2(n_867),
.B1(n_913),
.B2(n_599),
.Y(n_1316)
);

BUFx3_ASAP7_75t_L g1317 ( 
.A(n_1128),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1128),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1090),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1164),
.A2(n_587),
.B1(n_1058),
.B2(n_957),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1200),
.A2(n_957),
.B1(n_599),
.B2(n_1164),
.Y(n_1321)
);

OAI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1164),
.A2(n_587),
.B(n_1058),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_SL g1323 ( 
.A1(n_1084),
.A2(n_611),
.B1(n_1200),
.B2(n_830),
.Y(n_1323)
);

INVx4_ASAP7_75t_L g1324 ( 
.A(n_1130),
.Y(n_1324)
);

CKINVDCx20_ASAP7_75t_R g1325 ( 
.A(n_1169),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1164),
.A2(n_587),
.B1(n_1058),
.B2(n_957),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_1128),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1187),
.B(n_1093),
.Y(n_1328)
);

OAI21xp33_ASAP7_75t_L g1329 ( 
.A1(n_1164),
.A2(n_957),
.B(n_587),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1200),
.A2(n_957),
.B1(n_599),
.B2(n_1164),
.Y(n_1330)
);

BUFx2_ASAP7_75t_SL g1331 ( 
.A(n_1278),
.Y(n_1331)
);

INVxp67_ASAP7_75t_L g1332 ( 
.A(n_1256),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1300),
.B(n_1309),
.Y(n_1333)
);

INVxp33_ASAP7_75t_SL g1334 ( 
.A(n_1238),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1310),
.A2(n_1326),
.B(n_1320),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1272),
.B(n_1285),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1328),
.B(n_1233),
.Y(n_1337)
);

INVx2_ASAP7_75t_SL g1338 ( 
.A(n_1217),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1233),
.B(n_1231),
.Y(n_1339)
);

INVx2_ASAP7_75t_SL g1340 ( 
.A(n_1217),
.Y(n_1340)
);

INVxp67_ASAP7_75t_L g1341 ( 
.A(n_1265),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1287),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1235),
.B(n_1228),
.Y(n_1343)
);

OAI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1314),
.A2(n_1250),
.B1(n_1322),
.B2(n_1247),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1296),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_SL g1346 ( 
.A1(n_1316),
.A2(n_1283),
.B1(n_1263),
.B2(n_1281),
.Y(n_1346)
);

BUFx2_ASAP7_75t_SL g1347 ( 
.A(n_1324),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1261),
.A2(n_1262),
.B(n_1329),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1289),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1228),
.B(n_1241),
.Y(n_1350)
);

BUFx6f_ASAP7_75t_L g1351 ( 
.A(n_1294),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1291),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_1283),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1264),
.B(n_1253),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1284),
.A2(n_1274),
.B(n_1261),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1293),
.Y(n_1356)
);

INVx6_ASAP7_75t_L g1357 ( 
.A(n_1258),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1284),
.A2(n_1274),
.B(n_1262),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1249),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1248),
.B(n_1299),
.Y(n_1360)
);

INVxp67_ASAP7_75t_L g1361 ( 
.A(n_1311),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1276),
.Y(n_1362)
);

OAI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1302),
.A2(n_1323),
.B(n_1307),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1295),
.B(n_1230),
.Y(n_1364)
);

INVx2_ASAP7_75t_SL g1365 ( 
.A(n_1217),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1249),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1290),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1292),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1295),
.B(n_1230),
.Y(n_1369)
);

INVx2_ASAP7_75t_SL g1370 ( 
.A(n_1226),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1288),
.A2(n_1273),
.B(n_1255),
.Y(n_1371)
);

AO21x2_ASAP7_75t_L g1372 ( 
.A1(n_1268),
.A2(n_1286),
.B(n_1234),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1242),
.Y(n_1373)
);

INVx2_ASAP7_75t_SL g1374 ( 
.A(n_1226),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1244),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1297),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1315),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1319),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1254),
.B(n_1236),
.Y(n_1379)
);

BUFx6f_ASAP7_75t_L g1380 ( 
.A(n_1226),
.Y(n_1380)
);

OR2x2_ASAP7_75t_L g1381 ( 
.A(n_1232),
.B(n_1254),
.Y(n_1381)
);

AO21x2_ASAP7_75t_L g1382 ( 
.A1(n_1257),
.A2(n_1280),
.B(n_1277),
.Y(n_1382)
);

INVxp67_ASAP7_75t_SL g1383 ( 
.A(n_1245),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1282),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1225),
.B(n_1227),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1288),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1304),
.A2(n_1330),
.B(n_1321),
.Y(n_1387)
);

NOR2xp67_ASAP7_75t_L g1388 ( 
.A(n_1237),
.B(n_1236),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1259),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1259),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1255),
.Y(n_1391)
);

BUFx3_ASAP7_75t_L g1392 ( 
.A(n_1258),
.Y(n_1392)
);

BUFx3_ASAP7_75t_L g1393 ( 
.A(n_1305),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1225),
.B(n_1227),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1232),
.Y(n_1395)
);

BUFx2_ASAP7_75t_L g1396 ( 
.A(n_1312),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_SL g1397 ( 
.A(n_1304),
.B(n_1330),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1305),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1237),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1239),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1221),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1222),
.A2(n_1271),
.B(n_1321),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1353),
.B(n_1222),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_1357),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1353),
.B(n_1215),
.Y(n_1405)
);

AO21x2_ASAP7_75t_L g1406 ( 
.A1(n_1372),
.A2(n_1246),
.B(n_1270),
.Y(n_1406)
);

O2A1O1Ixp33_ASAP7_75t_SL g1407 ( 
.A1(n_1344),
.A2(n_1397),
.B(n_1363),
.C(n_1379),
.Y(n_1407)
);

OA21x2_ASAP7_75t_L g1408 ( 
.A1(n_1355),
.A2(n_1279),
.B(n_1218),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1346),
.A2(n_1247),
.B1(n_1317),
.B2(n_1220),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1335),
.A2(n_1229),
.B(n_1269),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1339),
.B(n_1240),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1343),
.B(n_1224),
.Y(n_1412)
);

A2O1A1Ixp33_ASAP7_75t_L g1413 ( 
.A1(n_1388),
.A2(n_1327),
.B(n_1317),
.C(n_1220),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1366),
.B(n_1318),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1345),
.B(n_1318),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1341),
.B(n_1337),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1350),
.B(n_1266),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1334),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_1357),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1354),
.B(n_1327),
.Y(n_1420)
);

A2O1A1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1388),
.A2(n_1224),
.B(n_1260),
.C(n_1298),
.Y(n_1421)
);

AOI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1385),
.A2(n_1325),
.B1(n_1223),
.B2(n_1219),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1387),
.A2(n_1275),
.B1(n_1298),
.B2(n_1239),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1389),
.B(n_1251),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1359),
.B(n_1252),
.Y(n_1425)
);

NAND2x1p5_ASAP7_75t_L g1426 ( 
.A(n_1402),
.B(n_1298),
.Y(n_1426)
);

AO32x2_ASAP7_75t_L g1427 ( 
.A1(n_1338),
.A2(n_1243),
.A3(n_1267),
.B1(n_1239),
.B2(n_1303),
.Y(n_1427)
);

AND2x4_ASAP7_75t_SL g1428 ( 
.A(n_1380),
.B(n_1216),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1331),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1342),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1401),
.B(n_1303),
.Y(n_1431)
);

AO32x2_ASAP7_75t_L g1432 ( 
.A1(n_1338),
.A2(n_1370),
.A3(n_1374),
.B1(n_1365),
.B2(n_1340),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1396),
.B(n_1373),
.Y(n_1433)
);

AOI221xp5_ASAP7_75t_L g1434 ( 
.A1(n_1401),
.A2(n_1306),
.B1(n_1313),
.B2(n_1301),
.C(n_1219),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1375),
.B(n_1308),
.Y(n_1435)
);

O2A1O1Ixp33_ASAP7_75t_SL g1436 ( 
.A1(n_1381),
.A2(n_1267),
.B(n_1301),
.C(n_1399),
.Y(n_1436)
);

INVxp67_ASAP7_75t_L g1437 ( 
.A(n_1362),
.Y(n_1437)
);

A2O1A1Ixp33_ASAP7_75t_L g1438 ( 
.A1(n_1348),
.A2(n_1394),
.B(n_1385),
.C(n_1402),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1333),
.B(n_1332),
.Y(n_1439)
);

A2O1A1Ixp33_ASAP7_75t_L g1440 ( 
.A1(n_1394),
.A2(n_1381),
.B(n_1399),
.C(n_1369),
.Y(n_1440)
);

O2A1O1Ixp33_ASAP7_75t_SL g1441 ( 
.A1(n_1391),
.A2(n_1395),
.B(n_1384),
.C(n_1360),
.Y(n_1441)
);

NOR2x1_ASAP7_75t_SL g1442 ( 
.A(n_1382),
.B(n_1347),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1364),
.B(n_1369),
.Y(n_1443)
);

AOI221xp5_ASAP7_75t_SL g1444 ( 
.A1(n_1384),
.A2(n_1368),
.B1(n_1361),
.B2(n_1367),
.C(n_1386),
.Y(n_1444)
);

A2O1A1Ixp33_ASAP7_75t_L g1445 ( 
.A1(n_1371),
.A2(n_1395),
.B(n_1368),
.C(n_1355),
.Y(n_1445)
);

NOR2x1_ASAP7_75t_SL g1446 ( 
.A(n_1382),
.B(n_1347),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1382),
.B(n_1390),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1383),
.B(n_1376),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1357),
.A2(n_1398),
.B1(n_1393),
.B2(n_1392),
.Y(n_1449)
);

OAI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1371),
.A2(n_1358),
.B(n_1400),
.Y(n_1450)
);

O2A1O1Ixp33_ASAP7_75t_L g1451 ( 
.A1(n_1372),
.A2(n_1367),
.B(n_1393),
.C(n_1392),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1430),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1416),
.B(n_1331),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1443),
.B(n_1352),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1411),
.B(n_1357),
.Y(n_1455)
);

NAND3xp33_ASAP7_75t_L g1456 ( 
.A(n_1407),
.B(n_1377),
.C(n_1378),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1450),
.B(n_1386),
.Y(n_1457)
);

INVxp67_ASAP7_75t_L g1458 ( 
.A(n_1447),
.Y(n_1458)
);

NOR2xp67_ASAP7_75t_L g1459 ( 
.A(n_1447),
.B(n_1378),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1418),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1445),
.B(n_1356),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1445),
.B(n_1358),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1408),
.B(n_1336),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1408),
.B(n_1336),
.Y(n_1464)
);

INVx1_ASAP7_75t_SL g1465 ( 
.A(n_1414),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1429),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1432),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1448),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1440),
.A2(n_1398),
.B1(n_1393),
.B2(n_1392),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1432),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1432),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1438),
.B(n_1352),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1433),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1438),
.B(n_1349),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1467),
.B(n_1372),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1463),
.B(n_1442),
.Y(n_1476)
);

OAI221xp5_ASAP7_75t_SL g1477 ( 
.A1(n_1456),
.A2(n_1440),
.B1(n_1434),
.B2(n_1444),
.C(n_1407),
.Y(n_1477)
);

OAI33xp33_ASAP7_75t_L g1478 ( 
.A1(n_1456),
.A2(n_1437),
.A3(n_1439),
.B1(n_1420),
.B2(n_1451),
.B3(n_1449),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1463),
.B(n_1446),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1467),
.B(n_1427),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1467),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1462),
.B(n_1427),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1463),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1462),
.B(n_1427),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1462),
.B(n_1427),
.Y(n_1485)
);

NAND2x1_ASAP7_75t_L g1486 ( 
.A(n_1464),
.B(n_1351),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1470),
.B(n_1342),
.Y(n_1487)
);

AOI221xp5_ASAP7_75t_L g1488 ( 
.A1(n_1469),
.A2(n_1441),
.B1(n_1409),
.B2(n_1410),
.C(n_1436),
.Y(n_1488)
);

AOI33xp33_ASAP7_75t_L g1489 ( 
.A1(n_1457),
.A2(n_1441),
.A3(n_1403),
.B1(n_1405),
.B2(n_1412),
.B3(n_1422),
.Y(n_1489)
);

AO21x2_ASAP7_75t_L g1490 ( 
.A1(n_1459),
.A2(n_1474),
.B(n_1472),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1471),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1452),
.Y(n_1492)
);

INVxp67_ASAP7_75t_L g1493 ( 
.A(n_1457),
.Y(n_1493)
);

OAI221xp5_ASAP7_75t_L g1494 ( 
.A1(n_1469),
.A2(n_1413),
.B1(n_1421),
.B2(n_1423),
.C(n_1426),
.Y(n_1494)
);

OAI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1474),
.A2(n_1413),
.B(n_1421),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1483),
.B(n_1458),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1483),
.B(n_1458),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1481),
.B(n_1461),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1493),
.B(n_1468),
.Y(n_1499)
);

INVxp67_ASAP7_75t_L g1500 ( 
.A(n_1492),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1493),
.B(n_1468),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1492),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1478),
.A2(n_1406),
.B1(n_1453),
.B2(n_1472),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1482),
.B(n_1473),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1482),
.B(n_1465),
.Y(n_1505)
);

BUFx3_ASAP7_75t_L g1506 ( 
.A(n_1490),
.Y(n_1506)
);

BUFx2_ASAP7_75t_SL g1507 ( 
.A(n_1476),
.Y(n_1507)
);

INVx2_ASAP7_75t_SL g1508 ( 
.A(n_1486),
.Y(n_1508)
);

AND2x4_ASAP7_75t_SL g1509 ( 
.A(n_1482),
.B(n_1425),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1490),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1487),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1482),
.B(n_1465),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1480),
.B(n_1454),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1487),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1481),
.B(n_1461),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1484),
.B(n_1485),
.Y(n_1516)
);

INVx3_ASAP7_75t_L g1517 ( 
.A(n_1486),
.Y(n_1517)
);

BUFx2_ASAP7_75t_L g1518 ( 
.A(n_1490),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1487),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1511),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1511),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1514),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1502),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1516),
.B(n_1484),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1516),
.B(n_1484),
.Y(n_1525)
);

NAND2xp33_ASAP7_75t_SL g1526 ( 
.A(n_1503),
.B(n_1489),
.Y(n_1526)
);

BUFx2_ASAP7_75t_L g1527 ( 
.A(n_1502),
.Y(n_1527)
);

O2A1O1Ixp33_ASAP7_75t_L g1528 ( 
.A1(n_1503),
.A2(n_1477),
.B(n_1478),
.C(n_1495),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1506),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1513),
.B(n_1490),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1516),
.B(n_1504),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1506),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1506),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1514),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1519),
.Y(n_1535)
);

INVx3_ASAP7_75t_L g1536 ( 
.A(n_1506),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1500),
.B(n_1480),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1519),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1498),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1500),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_SL g1541 ( 
.A(n_1509),
.B(n_1489),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1513),
.B(n_1490),
.Y(n_1542)
);

O2A1O1Ixp33_ASAP7_75t_L g1543 ( 
.A1(n_1510),
.A2(n_1477),
.B(n_1495),
.C(n_1488),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1510),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1510),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1504),
.B(n_1484),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1499),
.B(n_1480),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1498),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1499),
.B(n_1490),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1501),
.B(n_1480),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1518),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1501),
.B(n_1481),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1498),
.B(n_1475),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1497),
.B(n_1491),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1504),
.B(n_1485),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1507),
.B(n_1485),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1508),
.B(n_1476),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1515),
.Y(n_1558)
);

NAND2xp33_ASAP7_75t_L g1559 ( 
.A(n_1508),
.B(n_1488),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1497),
.B(n_1491),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1515),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1528),
.B(n_1509),
.Y(n_1562)
);

OR2x6_ASAP7_75t_L g1563 ( 
.A(n_1543),
.B(n_1404),
.Y(n_1563)
);

NOR3xp33_ASAP7_75t_L g1564 ( 
.A(n_1526),
.B(n_1477),
.C(n_1488),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1527),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1531),
.B(n_1527),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1523),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1531),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1541),
.B(n_1509),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1524),
.B(n_1509),
.Y(n_1570)
);

NAND2x1p5_ASAP7_75t_L g1571 ( 
.A(n_1536),
.B(n_1486),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1524),
.B(n_1507),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1525),
.B(n_1507),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1543),
.B(n_1505),
.Y(n_1574)
);

AOI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1559),
.A2(n_1494),
.B1(n_1495),
.B2(n_1406),
.Y(n_1575)
);

AOI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1540),
.A2(n_1494),
.B1(n_1479),
.B2(n_1476),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1554),
.B(n_1454),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1520),
.Y(n_1578)
);

INVx3_ASAP7_75t_L g1579 ( 
.A(n_1557),
.Y(n_1579)
);

NAND4xp25_ASAP7_75t_L g1580 ( 
.A(n_1554),
.B(n_1494),
.C(n_1417),
.D(n_1431),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1557),
.Y(n_1581)
);

INVx1_ASAP7_75t_SL g1582 ( 
.A(n_1560),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1560),
.B(n_1497),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1539),
.B(n_1505),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1525),
.B(n_1508),
.Y(n_1585)
);

NOR2x1_ASAP7_75t_L g1586 ( 
.A(n_1536),
.B(n_1517),
.Y(n_1586)
);

INVx3_ASAP7_75t_L g1587 ( 
.A(n_1557),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1520),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1539),
.B(n_1505),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1521),
.Y(n_1590)
);

AOI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1537),
.A2(n_1518),
.B(n_1436),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1547),
.B(n_1475),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1548),
.B(n_1512),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1546),
.B(n_1496),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1546),
.B(n_1496),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1521),
.Y(n_1596)
);

NAND2x1_ASAP7_75t_SL g1597 ( 
.A(n_1566),
.B(n_1556),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1569),
.B(n_1555),
.Y(n_1598)
);

NAND2x1p5_ASAP7_75t_L g1599 ( 
.A(n_1575),
.B(n_1398),
.Y(n_1599)
);

OAI21xp5_ASAP7_75t_SL g1600 ( 
.A1(n_1564),
.A2(n_1428),
.B(n_1556),
.Y(n_1600)
);

OAI221xp5_ASAP7_75t_L g1601 ( 
.A1(n_1574),
.A2(n_1518),
.B1(n_1537),
.B2(n_1558),
.C(n_1548),
.Y(n_1601)
);

INVx1_ASAP7_75t_SL g1602 ( 
.A(n_1563),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1582),
.B(n_1558),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1562),
.A2(n_1529),
.B1(n_1532),
.B2(n_1533),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1588),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1588),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1583),
.B(n_1561),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1567),
.B(n_1561),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1596),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1566),
.B(n_1557),
.Y(n_1610)
);

XNOR2x1_ASAP7_75t_L g1611 ( 
.A(n_1563),
.B(n_1435),
.Y(n_1611)
);

OAI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1563),
.A2(n_1536),
.B1(n_1549),
.B2(n_1530),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1565),
.B(n_1555),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1566),
.B(n_1547),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1596),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1578),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1580),
.B(n_1590),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1568),
.Y(n_1618)
);

BUFx2_ASAP7_75t_L g1619 ( 
.A(n_1570),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1568),
.B(n_1550),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1594),
.B(n_1550),
.Y(n_1621)
);

AOI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1617),
.A2(n_1591),
.B(n_1586),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1597),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1604),
.B(n_1594),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1616),
.Y(n_1625)
);

OAI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1604),
.A2(n_1576),
.B1(n_1570),
.B2(n_1581),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1602),
.B(n_1595),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1619),
.B(n_1595),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1616),
.Y(n_1629)
);

O2A1O1Ixp33_ASAP7_75t_L g1630 ( 
.A1(n_1612),
.A2(n_1536),
.B(n_1529),
.C(n_1533),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1610),
.B(n_1581),
.Y(n_1631)
);

NAND3xp33_ASAP7_75t_SL g1632 ( 
.A(n_1599),
.B(n_1571),
.C(n_1584),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1610),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1598),
.B(n_1570),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1605),
.B(n_1577),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1606),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1609),
.Y(n_1637)
);

INVx2_ASAP7_75t_SL g1638 ( 
.A(n_1615),
.Y(n_1638)
);

NOR3xp33_ASAP7_75t_SL g1639 ( 
.A(n_1600),
.B(n_1460),
.C(n_1589),
.Y(n_1639)
);

OAI322xp33_ASAP7_75t_L g1640 ( 
.A1(n_1601),
.A2(n_1549),
.A3(n_1530),
.B1(n_1542),
.B2(n_1593),
.C1(n_1522),
.C2(n_1538),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1638),
.B(n_1618),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1634),
.B(n_1633),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1625),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1629),
.Y(n_1644)
);

O2A1O1Ixp5_ASAP7_75t_L g1645 ( 
.A1(n_1640),
.A2(n_1612),
.B(n_1608),
.C(n_1613),
.Y(n_1645)
);

OAI221xp5_ASAP7_75t_L g1646 ( 
.A1(n_1622),
.A2(n_1623),
.B1(n_1639),
.B2(n_1626),
.C(n_1624),
.Y(n_1646)
);

NOR2x1_ASAP7_75t_L g1647 ( 
.A(n_1636),
.B(n_1611),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1633),
.B(n_1611),
.Y(n_1648)
);

AO22x1_ASAP7_75t_L g1649 ( 
.A1(n_1631),
.A2(n_1579),
.B1(n_1587),
.B2(n_1585),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1638),
.Y(n_1650)
);

INVxp67_ASAP7_75t_L g1651 ( 
.A(n_1631),
.Y(n_1651)
);

NAND4xp25_ASAP7_75t_L g1652 ( 
.A(n_1647),
.B(n_1637),
.C(n_1636),
.D(n_1630),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1642),
.B(n_1634),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1650),
.Y(n_1654)
);

NOR2x1_ASAP7_75t_L g1655 ( 
.A(n_1641),
.B(n_1643),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1641),
.Y(n_1656)
);

NAND4xp25_ASAP7_75t_SL g1657 ( 
.A(n_1646),
.B(n_1628),
.C(n_1627),
.D(n_1635),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1651),
.B(n_1599),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1648),
.B(n_1614),
.Y(n_1659)
);

NAND4xp25_ASAP7_75t_L g1660 ( 
.A(n_1645),
.B(n_1632),
.C(n_1603),
.D(n_1607),
.Y(n_1660)
);

NOR2xp67_ASAP7_75t_L g1661 ( 
.A(n_1652),
.B(n_1644),
.Y(n_1661)
);

AOI211x1_ASAP7_75t_SL g1662 ( 
.A1(n_1660),
.A2(n_1620),
.B(n_1649),
.C(n_1533),
.Y(n_1662)
);

OAI211xp5_ASAP7_75t_L g1663 ( 
.A1(n_1652),
.A2(n_1621),
.B(n_1579),
.C(n_1587),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1655),
.Y(n_1664)
);

AOI211xp5_ASAP7_75t_SL g1665 ( 
.A1(n_1654),
.A2(n_1656),
.B(n_1653),
.C(n_1659),
.Y(n_1665)
);

AOI221x1_ASAP7_75t_SL g1666 ( 
.A1(n_1661),
.A2(n_1664),
.B1(n_1662),
.B2(n_1665),
.C(n_1657),
.Y(n_1666)
);

NAND3xp33_ASAP7_75t_L g1667 ( 
.A(n_1663),
.B(n_1658),
.C(n_1532),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1661),
.A2(n_1587),
.B1(n_1579),
.B2(n_1529),
.Y(n_1668)
);

O2A1O1Ixp5_ASAP7_75t_L g1669 ( 
.A1(n_1664),
.A2(n_1532),
.B(n_1551),
.C(n_1545),
.Y(n_1669)
);

OAI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1661),
.A2(n_1571),
.B(n_1572),
.Y(n_1670)
);

INVx1_ASAP7_75t_SL g1671 ( 
.A(n_1664),
.Y(n_1671)
);

XNOR2xp5_ASAP7_75t_L g1672 ( 
.A(n_1666),
.B(n_1428),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_1671),
.B(n_1466),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1667),
.Y(n_1674)
);

NAND4xp75_ASAP7_75t_L g1675 ( 
.A(n_1669),
.B(n_1573),
.C(n_1572),
.D(n_1545),
.Y(n_1675)
);

NOR2x1p5_ASAP7_75t_L g1676 ( 
.A(n_1670),
.B(n_1404),
.Y(n_1676)
);

NAND4xp75_ASAP7_75t_L g1677 ( 
.A(n_1674),
.B(n_1668),
.C(n_1544),
.D(n_1545),
.Y(n_1677)
);

AND3x4_ASAP7_75t_L g1678 ( 
.A(n_1672),
.B(n_1585),
.C(n_1419),
.Y(n_1678)
);

NOR3xp33_ASAP7_75t_L g1679 ( 
.A(n_1673),
.B(n_1675),
.C(n_1676),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1678),
.A2(n_1538),
.B1(n_1535),
.B2(n_1534),
.Y(n_1680)
);

AO22x2_ASAP7_75t_L g1681 ( 
.A1(n_1680),
.A2(n_1677),
.B1(n_1679),
.B2(n_1551),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1681),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1682),
.B(n_1522),
.Y(n_1683)
);

AOI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1683),
.A2(n_1551),
.B(n_1544),
.Y(n_1684)
);

AOI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1684),
.A2(n_1544),
.B1(n_1585),
.B2(n_1573),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_SL g1686 ( 
.A1(n_1684),
.A2(n_1535),
.B1(n_1534),
.B2(n_1517),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1686),
.B(n_1592),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1685),
.B(n_1542),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1687),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1688),
.Y(n_1690)
);

OAI221xp5_ASAP7_75t_R g1691 ( 
.A1(n_1690),
.A2(n_1553),
.B1(n_1508),
.B2(n_1552),
.C(n_1455),
.Y(n_1691)
);

AOI31xp33_ASAP7_75t_L g1692 ( 
.A1(n_1691),
.A2(n_1689),
.A3(n_1424),
.B(n_1415),
.Y(n_1692)
);


endmodule