module fake_jpeg_8087_n_253 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_253);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_253;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_96;

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_16),
.B(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_17),
.B(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_23),
.Y(n_38)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_21),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_46),
.Y(n_55)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_45),
.Y(n_57)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

NAND2x1_ASAP7_75t_SL g46 ( 
.A(n_24),
.B(n_35),
.Y(n_46)
);

CKINVDCx6p67_ASAP7_75t_R g47 ( 
.A(n_23),
.Y(n_47)
);

INVxp67_ASAP7_75t_SL g61 ( 
.A(n_47),
.Y(n_61)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_33),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_43),
.A2(n_21),
.B1(n_20),
.B2(n_34),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_50),
.A2(n_52),
.B1(n_38),
.B2(n_42),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_35),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_20),
.B1(n_34),
.B2(n_33),
.Y(n_52)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_64),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_20),
.B1(n_34),
.B2(n_33),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_59),
.A2(n_32),
.B1(n_45),
.B2(n_44),
.Y(n_85)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_38),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_32),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_42),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_29),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_69),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_29),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g90 ( 
.A(n_70),
.Y(n_90)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_72),
.Y(n_105)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_1),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_39),
.A2(n_18),
.B1(n_22),
.B2(n_30),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_75),
.A2(n_49),
.B1(n_68),
.B2(n_25),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_76),
.A2(n_81),
.B1(n_85),
.B2(n_93),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_77),
.B(n_87),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_51),
.B(n_39),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_91),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_83),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_46),
.B1(n_48),
.B2(n_45),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_66),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_65),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_40),
.Y(n_88)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_49),
.A2(n_32),
.B1(n_45),
.B2(n_44),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_55),
.A2(n_46),
.B1(n_44),
.B2(n_48),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_66),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_94),
.B(n_74),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_57),
.B(n_27),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_26),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_65),
.A2(n_46),
.B1(n_48),
.B2(n_41),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_97),
.B1(n_100),
.B2(n_102),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_59),
.A2(n_18),
.B1(n_22),
.B2(n_30),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_23),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_73),
.Y(n_124)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_103),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_63),
.A2(n_53),
.B1(n_71),
.B2(n_54),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_31),
.C(n_27),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_35),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_53),
.A2(n_31),
.B1(n_28),
.B2(n_24),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_63),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_106),
.Y(n_133)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_111),
.B(n_116),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_124),
.Y(n_144)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_117),
.A2(n_86),
.B1(n_90),
.B2(n_108),
.Y(n_149)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_127),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_91),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_125),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_35),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_106),
.Y(n_141)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_86),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_129),
.Y(n_143)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_83),
.B(n_28),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_130),
.B(n_98),
.Y(n_157)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_132),
.Y(n_148)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_81),
.A2(n_70),
.B(n_28),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_134),
.A2(n_98),
.B(n_89),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_129),
.A2(n_120),
.B1(n_118),
.B2(n_131),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_135),
.A2(n_137),
.B1(n_147),
.B2(n_153),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_93),
.B1(n_87),
.B2(n_80),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_136),
.A2(n_140),
.B1(n_149),
.B2(n_117),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_118),
.A2(n_96),
.B1(n_77),
.B2(n_80),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_139),
.Y(n_166)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_99),
.B1(n_82),
.B2(n_56),
.Y(n_140)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_151),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_121),
.A2(n_82),
.B1(n_108),
.B2(n_103),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_101),
.Y(n_150)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_111),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_158),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_121),
.A2(n_134),
.B1(n_110),
.B2(n_125),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_154),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_84),
.Y(n_155)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_109),
.B(n_88),
.C(n_95),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_130),
.C(n_109),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_157),
.A2(n_160),
.B(n_143),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_84),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_122),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_165),
.C(n_172),
.Y(n_188)
);

AOI21xp33_ASAP7_75t_L g163 ( 
.A1(n_144),
.A2(n_112),
.B(n_159),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_171),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_155),
.B(n_114),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_112),
.C(n_115),
.Y(n_172)
);

XNOR2x1_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_112),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_173),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_175),
.B(n_177),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_160),
.A2(n_146),
.B(n_143),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_176),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_97),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_179),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_137),
.B(n_114),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_144),
.B(n_132),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_183),
.Y(n_194)
);

AOI32xp33_ASAP7_75t_L g181 ( 
.A1(n_153),
.A2(n_86),
.A3(n_89),
.B1(n_3),
.B2(n_4),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_4),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_135),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_182),
.A2(n_145),
.B1(n_151),
.B2(n_140),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_136),
.B(n_3),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_185),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_186),
.A2(n_190),
.B1(n_195),
.B2(n_178),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_169),
.A2(n_148),
.B1(n_147),
.B2(n_145),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_168),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_191),
.A2(n_193),
.B(n_197),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_169),
.A2(n_148),
.B1(n_156),
.B2(n_138),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_152),
.Y(n_196)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_166),
.Y(n_197)
);

OAI32xp33_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_158),
.A3(n_142),
.B1(n_8),
.B2(n_9),
.Y(n_198)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_198),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_161),
.B(n_142),
.Y(n_199)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_199),
.Y(n_211)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_170),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_172),
.C(n_183),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_204),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_208),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_187),
.A2(n_182),
.B1(n_173),
.B2(n_167),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_206),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_215),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_176),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_210),
.B(n_201),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_212),
.A2(n_184),
.B1(n_202),
.B2(n_214),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_180),
.C(n_165),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_188),
.C(n_192),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_175),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_215),
.B(n_192),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_220),
.C(n_225),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_212),
.A2(n_184),
.B1(n_200),
.B2(n_198),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_218),
.A2(n_222),
.B1(n_189),
.B2(n_211),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_221),
.A2(n_208),
.B(n_209),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_202),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_194),
.C(n_195),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_210),
.C(n_206),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_224),
.B(n_162),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_230),
.Y(n_240)
);

MAJx2_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_207),
.C(n_194),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_229),
.A2(n_231),
.B(n_232),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_223),
.B(n_205),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_233),
.A2(n_226),
.B(n_220),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_216),
.A2(n_186),
.B1(n_211),
.B2(n_203),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_5),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_235),
.A2(n_237),
.B(n_10),
.Y(n_245)
);

OAI221xp5_ASAP7_75t_L g236 ( 
.A1(n_229),
.A2(n_219),
.B1(n_199),
.B2(n_203),
.C(n_221),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_236),
.B(n_10),
.Y(n_244)
);

NAND4xp25_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_222),
.C(n_223),
.D(n_9),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_239),
.B(n_6),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_238),
.A2(n_228),
.B1(n_233),
.B2(n_11),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_241),
.B(n_243),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_244),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_6),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_245),
.B(n_11),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_247),
.B(n_12),
.C(n_13),
.Y(n_249)
);

AOI31xp33_ASAP7_75t_L g251 ( 
.A1(n_249),
.A2(n_250),
.A3(n_248),
.B(n_12),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_241),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_12),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_14),
.Y(n_253)
);


endmodule