module real_jpeg_18578_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_470),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_0),
.B(n_471),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_1),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_78)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_1),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_1),
.A2(n_172),
.B1(n_175),
.B2(n_176),
.Y(n_171)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_1),
.Y(n_202)
);

OAI32xp33_ASAP7_75t_L g285 ( 
.A1(n_1),
.A2(n_103),
.A3(n_286),
.B1(n_287),
.B2(n_290),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_1),
.A2(n_202),
.B1(n_295),
.B2(n_297),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_1),
.B(n_132),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_1),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_1),
.B(n_377),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_2),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_2),
.A2(n_77),
.B1(n_96),
.B2(n_194),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_L g238 ( 
.A1(n_2),
.A2(n_77),
.B1(n_239),
.B2(n_242),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_2),
.A2(n_77),
.B1(n_308),
.B2(n_311),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_3),
.Y(n_106)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_3),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_3),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_4),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_4),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_4),
.Y(n_154)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_4),
.Y(n_329)
);

BUFx5_ASAP7_75t_L g332 ( 
.A(n_4),
.Y(n_332)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_5),
.A2(n_89),
.B1(n_90),
.B2(n_95),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g222 ( 
.A(n_6),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_6),
.Y(n_228)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_6),
.Y(n_257)
);

BUFx5_ASAP7_75t_L g316 ( 
.A(n_6),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_7),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_7),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_7),
.Y(n_149)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_7),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_7),
.Y(n_188)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_7),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_8),
.A2(n_54),
.B1(n_57),
.B2(n_58),
.Y(n_53)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_8),
.A2(n_58),
.B1(n_124),
.B2(n_126),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_L g156 ( 
.A1(n_8),
.A2(n_58),
.B1(n_157),
.B2(n_160),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_8),
.A2(n_58),
.B1(n_213),
.B2(n_217),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_9),
.Y(n_471)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_11),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_12),
.Y(n_139)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_12),
.Y(n_142)
);

BUFx4f_ASAP7_75t_L g216 ( 
.A(n_12),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g218 ( 
.A(n_12),
.Y(n_218)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_13),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_63),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_62),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_59),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_18),
.B(n_59),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_18),
.B(n_276),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_18),
.B(n_276),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_33),
.B1(n_41),
.B2(n_53),
.Y(n_18)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_19),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_20),
.B(n_33),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_20),
.A2(n_33),
.B1(n_74),
.B2(n_78),
.Y(n_73)
);

OA22x2_ASAP7_75t_L g165 ( 
.A1(n_20),
.A2(n_33),
.B1(n_74),
.B2(n_78),
.Y(n_165)
);

OAI21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_28),
.B(n_33),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_21),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_30),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g408 ( 
.A(n_32),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_33),
.A2(n_41),
.B(n_272),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_33),
.Y(n_377)
);

OA22x2_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_39),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_46),
.B1(n_48),
.B2(n_52),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_46),
.A2(n_47),
.B1(n_246),
.B2(n_250),
.Y(n_245)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_52),
.A2(n_185),
.B1(n_186),
.B2(n_189),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_53),
.Y(n_60)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_61),
.B(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_277),
.B(n_464),
.Y(n_64)
);

NAND3xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_265),
.C(n_275),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_232),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_67),
.A2(n_466),
.B(n_467),
.Y(n_465)
);

NOR2xp67_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_177),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_68),
.B(n_177),
.Y(n_467)
);

XOR2x2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_167),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_165),
.B2(n_166),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_70),
.B(n_166),
.C(n_167),
.Y(n_266)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_85),
.B2(n_86),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_72),
.A2(n_73),
.B1(n_235),
.B2(n_302),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_72),
.A2(n_73),
.B1(n_192),
.B2(n_378),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_73),
.B(n_235),
.C(n_236),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_73),
.B(n_87),
.C(n_133),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_73),
.B(n_192),
.C(n_438),
.Y(n_437)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_78),
.Y(n_231)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_81),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_81),
.B(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_81),
.B(n_291),
.Y(n_290)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_133),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_100),
.B1(n_123),
.B2(n_132),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_88),
.A2(n_100),
.B1(n_132),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_89),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_90),
.A2(n_396),
.B1(n_405),
.B2(n_409),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g404 ( 
.A(n_94),
.Y(n_404)
);

BUFx2_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx8_ASAP7_75t_L g289 ( 
.A(n_98),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g192 ( 
.A1(n_101),
.A2(n_113),
.B1(n_171),
.B2(n_193),
.Y(n_192)
);

OA22x2_ASAP7_75t_L g235 ( 
.A1(n_101),
.A2(n_113),
.B1(n_171),
.B2(n_193),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_101),
.Y(n_270)
);

AO21x1_ASAP7_75t_L g430 ( 
.A1(n_101),
.A2(n_113),
.B(n_171),
.Y(n_430)
);

NAND2x1p5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_113),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_108),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_107),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_113),
.B(n_270),
.Y(n_269)
);

OA22x2_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_116),
.B1(n_119),
.B2(n_121),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_118),
.Y(n_325)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_123),
.B(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_131),
.Y(n_174)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_133),
.B(n_169),
.Y(n_179)
);

AND2x2_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_156),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_144),
.Y(n_134)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_135),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_135),
.A2(n_184),
.B(n_200),
.Y(n_199)
);

AOI21x1_ASAP7_75t_SL g388 ( 
.A1(n_135),
.A2(n_389),
.B(n_390),
.Y(n_388)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NOR2x1_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_146),
.Y(n_145)
);

AO22x1_ASAP7_75t_L g237 ( 
.A1(n_136),
.A2(n_145),
.B1(n_201),
.B2(n_238),
.Y(n_237)
);

AO22x2_ASAP7_75t_L g301 ( 
.A1(n_136),
.A2(n_145),
.B1(n_201),
.B2(n_238),
.Y(n_301)
);

AO22x2_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_140),
.B2(n_143),
.Y(n_136)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_138),
.Y(n_223)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_139),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_140),
.Y(n_251)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_142),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_144),
.Y(n_190)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_145),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_150),
.B1(n_152),
.B2(n_155),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_148),
.Y(n_243)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_149),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_155),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_156),
.A2(n_183),
.B1(n_190),
.B2(n_191),
.Y(n_182)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_164),
.Y(n_241)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_165),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_179),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_165),
.B(n_430),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_168),
.C(n_169),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_166),
.B(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_166),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_166),
.B(n_302),
.C(n_388),
.Y(n_452)
);

INVxp33_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_175),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_175),
.B(n_406),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.C(n_196),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_178),
.A2(n_180),
.B1(n_181),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_178),
.Y(n_264)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_181),
.A2(n_182),
.B(n_192),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_192),
.Y(n_181)
);

INVxp67_ASAP7_75t_SL g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_189),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_191),
.B(n_357),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_192),
.A2(n_373),
.B1(n_374),
.B2(n_378),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_192),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_192),
.B(n_351),
.C(n_376),
.Y(n_392)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_196),
.B(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_211),
.B(n_229),
.Y(n_196)
);

INVxp33_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_198),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_210),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_199),
.A2(n_210),
.B1(n_211),
.B2(n_421),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_199),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_209),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_201),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B(n_207),
.Y(n_201)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OAI32xp33_ASAP7_75t_L g321 ( 
.A1(n_207),
.A2(n_223),
.A3(n_322),
.B1(n_326),
.B2(n_330),
.Y(n_321)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_209),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_210),
.A2(n_211),
.B1(n_229),
.B2(n_230),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_211),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_219),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_212),
.A2(n_245),
.B1(n_252),
.B2(n_253),
.Y(n_244)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_218),
.Y(n_296)
);

INVx5_ASAP7_75t_L g299 ( 
.A(n_218),
.Y(n_299)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_218),
.Y(n_310)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_218),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_219),
.B(n_293),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_224),
.Y(n_219)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_220),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_220),
.B(n_294),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g350 ( 
.A(n_225),
.Y(n_350)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_231),
.B(n_273),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_262),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_233),
.B(n_262),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_258),
.C(n_259),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_234),
.B(n_415),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_235),
.A2(n_301),
.B1(n_302),
.B2(n_303),
.Y(n_300)
);

INVx3_ASAP7_75t_SL g302 ( 
.A(n_235),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_235),
.A2(n_302),
.B1(n_387),
.B2(n_388),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_236),
.B(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_244),
.Y(n_236)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_237),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_237),
.B(n_317),
.Y(n_339)
);

OAI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_237),
.A2(n_305),
.B1(n_369),
.B2(n_370),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_237),
.A2(n_244),
.B1(n_305),
.B2(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_244),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_245),
.A2(n_354),
.B(n_425),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_249),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OA22x2_ASAP7_75t_L g306 ( 
.A1(n_252),
.A2(n_293),
.B1(n_307),
.B2(n_313),
.Y(n_306)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_257),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_258),
.B(n_260),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

A2O1A1O1Ixp25_ASAP7_75t_L g464 ( 
.A1(n_265),
.A2(n_275),
.B(n_465),
.C(n_468),
.D(n_469),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_266),
.B(n_267),
.Y(n_468)
);

BUFx24_ASAP7_75t_SL g472 ( 
.A(n_267),
.Y(n_472)
);

FAx1_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_271),
.CI(n_274),
.CON(n_267),
.SN(n_267)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_271),
.C(n_274),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_278),
.Y(n_277)
);

AO221x1_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_411),
.B1(n_413),
.B2(n_457),
.C(n_463),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_382),
.B(n_410),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_366),
.B(n_381),
.Y(n_280)
);

OAI21x1_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_318),
.B(n_365),
.Y(n_281)
);

NOR2xp67_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_304),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_283),
.B(n_304),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_300),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_284),
.B(n_301),
.C(n_302),
.Y(n_380)
);

XOR2x2_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_292),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_285),
.B(n_292),
.Y(n_369)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_301),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_301),
.B(n_321),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_301),
.A2(n_303),
.B1(n_321),
.B2(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_301),
.B(n_424),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_301),
.A2(n_303),
.B1(n_424),
.B2(n_450),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.C(n_317),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_305),
.B(n_369),
.C(n_371),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_306),
.A2(n_337),
.B1(n_338),
.B2(n_339),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_306),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_306),
.B(n_356),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_306),
.B(n_356),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_306),
.A2(n_337),
.B1(n_394),
.B2(n_395),
.Y(n_393)
);

OA21x2_ASAP7_75t_L g351 ( 
.A1(n_307),
.A2(n_352),
.B(n_354),
.Y(n_351)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_316),
.Y(n_353)
);

AOI21x1_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_340),
.B(n_364),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_336),
.Y(n_319)
);

NOR2xp67_ASAP7_75t_SL g364 ( 
.A(n_320),
.B(n_336),
.Y(n_364)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_321),
.Y(n_362)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_333),
.Y(n_330)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_337),
.B(n_395),
.Y(n_438)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_359),
.B(n_363),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_342),
.A2(n_355),
.B(n_358),
.Y(n_341)
);

NOR2x1_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_351),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_349),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_351),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_351),
.A2(n_360),
.B1(n_375),
.B2(n_376),
.Y(n_374)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

NAND2xp33_ASAP7_75t_SL g363 ( 
.A(n_360),
.B(n_361),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_367),
.B(n_380),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_367),
.B(n_380),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_371),
.B1(n_372),
.B2(n_379),
.Y(n_367)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_368),
.Y(n_379)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_369),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_383),
.B(n_384),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_391),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_385),
.B(n_392),
.C(n_393),
.Y(n_443)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_393),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_401),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx2_ASAP7_75t_SL g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_441),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_431),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_414),
.B(n_416),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_R g463 ( 
.A(n_414),
.B(n_416),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_420),
.C(n_422),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_418),
.B(n_420),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_422),
.B(n_440),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_428),
.C(n_429),
.Y(n_422)
);

XNOR2x1_ASAP7_75t_L g433 ( 
.A(n_423),
.B(n_434),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_424),
.Y(n_450)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_431),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_439),
.Y(n_431)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_432),
.B(n_439),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_435),
.C(n_437),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_433),
.B(n_435),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_437),
.B(n_455),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_438),
.B(n_446),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_453),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_444),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_443),
.B(n_444),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_447),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_445),
.B(n_449),
.C(n_451),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_448),
.A2(n_449),
.B1(n_451),
.B2(n_452),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_453),
.B(n_460),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_456),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g458 ( 
.A(n_454),
.B(n_456),
.Y(n_458)
);

A2O1A1Ixp33_ASAP7_75t_L g457 ( 
.A1(n_458),
.A2(n_459),
.B(n_461),
.C(n_462),
.Y(n_457)
);


endmodule