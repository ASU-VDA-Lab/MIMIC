module fake_jpeg_14557_n_157 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_157);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_157;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_SL g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_10),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_9),
.B(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_2),
.B(n_3),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_8),
.B(n_12),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_1),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_34),
.A2(n_18),
.B1(n_25),
.B2(n_17),
.Y(n_65)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_23),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_39),
.A2(n_51),
.B1(n_31),
.B2(n_15),
.Y(n_62)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_45),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_50),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_24),
.B(n_7),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_48),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_30),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_28),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_28),
.A2(n_8),
.B1(n_31),
.B2(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_22),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_57),
.B(n_58),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_22),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_27),
.Y(n_59)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_27),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_64),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_57),
.B1(n_58),
.B2(n_55),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_25),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_65),
.A2(n_75),
.B1(n_59),
.B2(n_73),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_28),
.B(n_13),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_68),
.A2(n_76),
.B(n_69),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_17),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_72),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_38),
.B(n_21),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_21),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_64),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_49),
.A2(n_18),
.B1(n_20),
.B2(n_8),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_20),
.C(n_16),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_16),
.B1(n_36),
.B2(n_37),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_77),
.A2(n_53),
.B1(n_55),
.B2(n_78),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_33),
.B(n_47),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_79),
.B(n_52),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_81),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_53),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_84),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_85),
.A2(n_88),
.B1(n_91),
.B2(n_96),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_56),
.B(n_54),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_93),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_63),
.B1(n_78),
.B2(n_54),
.Y(n_91)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

HAxp5_ASAP7_75t_SL g94 ( 
.A(n_68),
.B(n_76),
.CON(n_94),
.SN(n_94)
);

AND2x4_ASAP7_75t_SL g113 ( 
.A(n_94),
.B(n_97),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_63),
.A2(n_61),
.B1(n_60),
.B2(n_71),
.Y(n_96)
);

AO21x2_ASAP7_75t_SL g97 ( 
.A1(n_74),
.A2(n_70),
.B(n_71),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_97),
.A2(n_101),
.B1(n_74),
.B2(n_52),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_101),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_60),
.A2(n_57),
.B1(n_58),
.B2(n_65),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_114),
.B1(n_103),
.B2(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_74),
.C(n_86),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_92),
.C(n_111),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_99),
.Y(n_106)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_99),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_111),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_95),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_116),
.Y(n_124)
);

OAI22x1_ASAP7_75t_L g118 ( 
.A1(n_113),
.A2(n_97),
.B1(n_114),
.B2(n_102),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_97),
.A2(n_90),
.B1(n_88),
.B2(n_91),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_90),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_128),
.B(n_120),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_112),
.B(n_89),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_125),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_122),
.A2(n_110),
.B1(n_107),
.B2(n_115),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_113),
.A2(n_93),
.B1(n_82),
.B2(n_96),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_123),
.A2(n_126),
.B1(n_127),
.B2(n_108),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_109),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_113),
.A2(n_82),
.B1(n_87),
.B2(n_81),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_110),
.A2(n_83),
.B1(n_92),
.B2(n_117),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_107),
.C(n_116),
.Y(n_131)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_123),
.C(n_126),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_121),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_134),
.Y(n_144)
);

BUFx24_ASAP7_75t_SL g134 ( 
.A(n_129),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_135),
.A2(n_138),
.B1(n_127),
.B2(n_120),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_137),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_106),
.B(n_104),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_142),
.C(n_131),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_141),
.B(n_143),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_138),
.B(n_120),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_133),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_148),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_145),
.A2(n_135),
.B(n_137),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_149),
.B(n_150),
.C(n_139),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_145),
.B(n_129),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_151),
.Y(n_154)
);

NAND3xp33_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_124),
.C(n_144),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_152),
.B(n_136),
.Y(n_155)
);

AOI21x1_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_141),
.B(n_153),
.Y(n_156)
);

FAx1_ASAP7_75t_SL g157 ( 
.A(n_156),
.B(n_142),
.CI(n_154),
.CON(n_157),
.SN(n_157)
);


endmodule