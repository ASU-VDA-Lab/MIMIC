module real_jpeg_23740_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_70;
wire n_41;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_1),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx8_ASAP7_75t_SL g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_4),
.B(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_4),
.B(n_36),
.C(n_94),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_4),
.A2(n_28),
.B1(n_69),
.B2(n_70),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_4),
.B(n_87),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_4),
.A2(n_119),
.B1(n_158),
.B2(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_5),
.A2(n_35),
.B1(n_36),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_6),
.A2(n_35),
.B1(n_36),
.B2(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_6),
.A2(n_54),
.B1(n_69),
.B2(n_70),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_7),
.A2(n_25),
.B1(n_32),
.B2(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_62),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_7),
.A2(n_62),
.B1(n_69),
.B2(n_70),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_62),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_9),
.A2(n_35),
.B1(n_36),
.B2(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

NAND3xp33_ASAP7_75t_L g31 ( 
.A(n_10),
.B(n_24),
.C(n_32),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_11),
.A2(n_25),
.B1(n_32),
.B2(n_74),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_11),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_11),
.A2(n_69),
.B1(n_70),
.B2(n_74),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_11),
.A2(n_35),
.B1(n_36),
.B2(n_74),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_12),
.A2(n_25),
.B1(n_32),
.B2(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_12),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_12),
.A2(n_69),
.B1(n_70),
.B2(n_89),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_12),
.A2(n_35),
.B1(n_36),
.B2(n_89),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_13),
.A2(n_69),
.B1(n_70),
.B2(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_13),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_13),
.A2(n_35),
.B1(n_36),
.B2(n_98),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_15),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_124),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_122),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_101),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_19),
.B(n_101),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_75),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_50),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_33),
.B1(n_48),
.B2(n_49),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_22),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_25),
.B(n_27),
.C(n_31),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_32),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_23),
.A2(n_24),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_25),
.A2(n_32),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

HAxp5_ASAP7_75t_SL g116 ( 
.A(n_25),
.B(n_28),
.CON(n_116),
.SN(n_116)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI21xp33_ASAP7_75t_L g77 ( 
.A1(n_27),
.A2(n_28),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_28),
.B(n_96),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_28),
.B(n_165),
.Y(n_164)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

NOR3xp33_ASAP7_75t_L g117 ( 
.A(n_32),
.B(n_66),
.C(n_70),
.Y(n_117)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_39),
.B1(n_42),
.B2(n_46),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_34),
.B(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_34),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_34),
.A2(n_42),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_35),
.A2(n_36),
.B1(n_94),
.B2(n_95),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_35),
.B(n_164),
.Y(n_163)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_38),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_45),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_42),
.B(n_53),
.Y(n_121)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_43),
.A2(n_119),
.B1(n_151),
.B2(n_158),
.Y(n_157)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g139 ( 
.A(n_45),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_55),
.C(n_59),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_51),
.A2(n_55),
.B1(n_56),
.B2(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_77),
.B1(n_79),
.B2(n_83),
.Y(n_76)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_58),
.B(n_80),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_59),
.B(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B1(n_68),
.B2(n_72),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_61),
.A2(n_64),
.B1(n_87),
.B2(n_116),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_64),
.A2(n_73),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_67),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

O2A1O1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_67),
.A2(n_69),
.B(n_115),
.C(n_117),
.Y(n_114)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_69),
.A2(n_70),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_70),
.B(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_85),
.Y(n_75)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_97),
.B(n_99),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_91),
.A2(n_110),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_91),
.A2(n_108),
.B1(n_110),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_92),
.A2(n_107),
.B(n_109),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_92),
.A2(n_96),
.B1(n_134),
.B2(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_96),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_97),
.B(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_106),
.C(n_111),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_102),
.A2(n_103),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_106),
.A2(n_111),
.B1(n_112),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_106),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_118),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_113),
.A2(n_114),
.B1(n_118),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_120),
.B(n_121),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_119),
.A2(n_137),
.B(n_138),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_120),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_179),
.B(n_185),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_169),
.B(n_178),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_147),
.B(n_168),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_135),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_135),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_131),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_141),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_142),
.C(n_145),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_137),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_154),
.B(n_167),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_153),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_153),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_159),
.B(n_166),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_157),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_177),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_177),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_174),
.C(n_175),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_181),
.Y(n_185)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);


endmodule