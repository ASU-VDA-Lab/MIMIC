module fake_jpeg_7912_n_163 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_163);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx11_ASAP7_75t_SL g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

CKINVDCx11_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_24),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_13),
.Y(n_37)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_36),
.A2(n_20),
.B1(n_22),
.B2(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_13),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_22),
.B1(n_25),
.B2(n_20),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_39),
.A2(n_47),
.B1(n_29),
.B2(n_33),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_45),
.A2(n_23),
.B1(n_18),
.B2(n_26),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_25),
.B1(n_17),
.B2(n_24),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_52),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_50),
.B(n_56),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_35),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_0),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_54),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_16),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_17),
.B1(n_16),
.B2(n_21),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_55),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_0),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_32),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_57),
.A2(n_58),
.B(n_69),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_31),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_60),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_21),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_63),
.Y(n_95)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_23),
.B1(n_18),
.B2(n_26),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_27),
.B1(n_30),
.B2(n_28),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_27),
.B1(n_30),
.B2(n_28),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_70),
.B1(n_71),
.B2(n_29),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_48),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_67),
.B(n_73),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_42),
.A2(n_18),
.B1(n_26),
.B2(n_2),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

AOI32xp33_ASAP7_75t_L g69 ( 
.A1(n_42),
.A2(n_33),
.A3(n_26),
.B1(n_29),
.B2(n_14),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_42),
.A2(n_8),
.B1(n_12),
.B2(n_2),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_82),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_76),
.A2(n_59),
.B1(n_63),
.B2(n_67),
.Y(n_112)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_96),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_0),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_1),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_84),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_1),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_1),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_86),
.B(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_2),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_73),
.B1(n_56),
.B2(n_52),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_104),
.B1(n_112),
.B2(n_113),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_94),
.B(n_53),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_100),
.B(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_71),
.Y(n_103)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_79),
.A2(n_58),
.B(n_57),
.Y(n_104)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_108),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_58),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_107),
.B(n_110),
.Y(n_128)
);

A2O1A1O1Ixp25_ASAP7_75t_L g108 ( 
.A1(n_87),
.A2(n_69),
.B(n_4),
.C(n_6),
.D(n_8),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_94),
.B(n_3),
.Y(n_109)
);

XNOR2x1_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_59),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_85),
.A2(n_3),
.B1(n_9),
.B2(n_10),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_12),
.C(n_9),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_84),
.C(n_93),
.Y(n_117)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_115),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_110),
.A2(n_89),
.B1(n_91),
.B2(n_80),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_106),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_108),
.A2(n_104),
.B1(n_107),
.B2(n_112),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_119),
.A2(n_102),
.B(n_109),
.Y(n_134)
);

NOR2x1_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_87),
.Y(n_121)
);

NOR3xp33_ASAP7_75t_SL g136 ( 
.A(n_121),
.B(n_128),
.C(n_125),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_97),
.A2(n_81),
.B1(n_88),
.B2(n_92),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_83),
.C(n_82),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_127),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_98),
.A2(n_90),
.B1(n_86),
.B2(n_75),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_3),
.C(n_9),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_133),
.Y(n_143)
);

OAI31xp33_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_113),
.A3(n_100),
.B(n_101),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_106),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_137),
.C(n_116),
.Y(n_140)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_129),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_10),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_111),
.B(n_115),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_135),
.A2(n_105),
.B1(n_127),
.B2(n_129),
.Y(n_144)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_135),
.A2(n_122),
.B1(n_119),
.B2(n_123),
.Y(n_139)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_142),
.C(n_138),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_117),
.C(n_126),
.Y(n_142)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_144),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_138),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_148),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_151),
.C(n_145),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_143),
.A2(n_134),
.B(n_131),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_139),
.B(n_11),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_155),
.C(n_154),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_149),
.A2(n_141),
.B1(n_140),
.B2(n_142),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_154),
.A2(n_146),
.B1(n_150),
.B2(n_149),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_11),
.Y(n_155)
);

FAx1_ASAP7_75t_SL g156 ( 
.A(n_152),
.B(n_151),
.CI(n_147),
.CON(n_156),
.SN(n_156)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_158),
.Y(n_160)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_158),
.Y(n_159)
);

FAx1_ASAP7_75t_SL g161 ( 
.A(n_160),
.B(n_156),
.CI(n_157),
.CON(n_161),
.SN(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_160),
.C(n_159),
.Y(n_162)
);

BUFx24_ASAP7_75t_SL g163 ( 
.A(n_162),
.Y(n_163)
);


endmodule