module fake_ibex_1739_n_573 (n_85, n_84, n_64, n_3, n_73, n_65, n_55, n_63, n_29, n_2, n_76, n_8, n_67, n_9, n_38, n_37, n_47, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_48, n_57, n_59, n_28, n_39, n_5, n_62, n_71, n_13, n_61, n_14, n_0, n_12, n_42, n_77, n_88, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_22, n_4, n_33, n_30, n_6, n_72, n_26, n_34, n_15, n_24, n_52, n_1, n_25, n_36, n_41, n_45, n_18, n_89, n_83, n_32, n_53, n_50, n_11, n_68, n_79, n_81, n_35, n_31, n_56, n_23, n_54, n_19, n_573);

input n_85;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_55;
input n_63;
input n_29;
input n_2;
input n_76;
input n_8;
input n_67;
input n_9;
input n_38;
input n_37;
input n_47;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_48;
input n_57;
input n_59;
input n_28;
input n_39;
input n_5;
input n_62;
input n_71;
input n_13;
input n_61;
input n_14;
input n_0;
input n_12;
input n_42;
input n_77;
input n_88;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_22;
input n_4;
input n_33;
input n_30;
input n_6;
input n_72;
input n_26;
input n_34;
input n_15;
input n_24;
input n_52;
input n_1;
input n_25;
input n_36;
input n_41;
input n_45;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_50;
input n_11;
input n_68;
input n_79;
input n_81;
input n_35;
input n_31;
input n_56;
input n_23;
input n_54;
input n_19;

output n_573;

wire n_151;
wire n_507;
wire n_540;
wire n_395;
wire n_171;
wire n_103;
wire n_529;
wire n_389;
wire n_204;
wire n_274;
wire n_387;
wire n_130;
wire n_177;
wire n_273;
wire n_330;
wire n_309;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_124;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_446;
wire n_108;
wire n_350;
wire n_165;
wire n_452;
wire n_255;
wire n_175;
wire n_398;
wire n_125;
wire n_304;
wire n_191;
wire n_153;
wire n_545;
wire n_194;
wire n_249;
wire n_334;
wire n_312;
wire n_478;
wire n_239;
wire n_134;
wire n_94;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_449;
wire n_547;
wire n_176;
wire n_216;
wire n_421;
wire n_475;
wire n_166;
wire n_163;
wire n_500;
wire n_542;
wire n_114;
wire n_236;
wire n_376;
wire n_377;
wire n_531;
wire n_556;
wire n_189;
wire n_498;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_105;
wire n_187;
wire n_154;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_144;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_113;
wire n_561;
wire n_117;
wire n_417;
wire n_471;
wire n_265;
wire n_504;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_210;
wire n_348;
wire n_220;
wire n_91;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_228;
wire n_147;
wire n_552;
wire n_251;
wire n_384;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_426;
wire n_323;
wire n_469;
wire n_143;
wire n_106;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_333;
wire n_110;
wire n_306;
wire n_400;
wire n_550;
wire n_169;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_109;
wire n_127;
wire n_121;
wire n_527;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_434;
wire n_296;
wire n_120;
wire n_168;
wire n_526;
wire n_155;
wire n_315;
wire n_441;
wire n_122;
wire n_523;
wire n_116;
wire n_370;
wire n_431;
wire n_289;
wire n_515;
wire n_150;
wire n_286;
wire n_321;
wire n_133;
wire n_569;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_538;
wire n_464;
wire n_136;
wire n_261;
wire n_521;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_437;
wire n_355;
wire n_474;
wire n_407;
wire n_102;
wire n_490;
wire n_568;
wire n_448;
wire n_99;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_126;
wire n_530;
wire n_356;
wire n_104;
wire n_420;
wire n_483;
wire n_543;
wire n_141;
wire n_487;
wire n_222;
wire n_186;
wire n_524;
wire n_349;
wire n_454;
wire n_295;
wire n_331;
wire n_230;
wire n_96;
wire n_185;
wire n_388;
wire n_536;
wire n_352;
wire n_290;
wire n_558;
wire n_174;
wire n_467;
wire n_427;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_146;
wire n_207;
wire n_438;
wire n_167;
wire n_128;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_205;
wire n_488;
wire n_139;
wire n_514;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_98;
wire n_129;
wire n_267;
wire n_245;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_347;
wire n_473;
wire n_445;
wire n_335;
wire n_413;
wire n_263;
wire n_353;
wire n_359;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_137;
wire n_338;
wire n_173;
wire n_477;
wire n_363;
wire n_402;
wire n_180;
wire n_369;
wire n_201;
wire n_351;
wire n_368;
wire n_456;
wire n_257;
wire n_401;
wire n_554;
wire n_553;
wire n_305;
wire n_307;
wire n_192;
wire n_140;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_365;
wire n_539;
wire n_100;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_516;
wire n_548;
wire n_567;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_506;
wire n_562;
wire n_564;
wire n_444;
wire n_546;
wire n_199;
wire n_495;
wire n_410;
wire n_308;
wire n_463;
wire n_411;
wire n_135;
wire n_520;
wire n_512;
wire n_283;
wire n_366;
wire n_397;
wire n_111;
wire n_322;
wire n_227;
wire n_499;
wire n_115;
wire n_248;
wire n_92;
wire n_451;
wire n_101;
wire n_190;
wire n_138;
wire n_409;
wire n_238;
wire n_214;
wire n_332;
wire n_517;
wire n_211;
wire n_218;
wire n_314;
wire n_563;
wire n_132;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_535;
wire n_382;
wire n_502;
wire n_532;
wire n_95;
wire n_405;
wire n_415;
wire n_285;
wire n_288;
wire n_247;
wire n_320;
wire n_379;
wire n_551;
wire n_291;
wire n_318;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_148;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_118;
wire n_378;
wire n_486;
wire n_422;
wire n_264;
wire n_198;
wire n_164;
wire n_217;
wire n_324;
wire n_391;
wire n_537;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_303;
wire n_362;
wire n_93;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_501;
wire n_266;
wire n_294;
wire n_112;
wire n_485;
wire n_284;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_476;
wire n_461;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_119;
wire n_361;
wire n_455;
wire n_419;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_311;
wire n_406;
wire n_97;
wire n_197;
wire n_528;
wire n_181;
wire n_131;
wire n_123;
wire n_260;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_572;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_252;
wire n_396;
wire n_107;
wire n_149;
wire n_489;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_159;
wire n_202;
wire n_231;
wire n_298;
wire n_160;
wire n_184;
wire n_492;
wire n_232;
wire n_380;
wire n_281;
wire n_559;
wire n_425;

INVx2_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_12),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_21),
.Y(n_94)
);

BUFx10_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_39),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_23),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

CKINVDCx5p33_ASAP7_75t_R g102 ( 
.A(n_37),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_22),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_27),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

CKINVDCx5p33_ASAP7_75t_R g108 ( 
.A(n_30),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

CKINVDCx5p33_ASAP7_75t_R g110 ( 
.A(n_90),
.Y(n_110)
);

INVxp67_ASAP7_75t_SL g111 ( 
.A(n_0),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_5),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_10),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_88),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_65),
.Y(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_29),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_33),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_82),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_15),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_47),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_5),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_14),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_59),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_18),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_1),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_32),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_17),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_34),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_7),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_58),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_16),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_50),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_60),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_24),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_9),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_46),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_84),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_53),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_81),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_4),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_51),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_6),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_15),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_2),
.Y(n_147)
);

NOR2xp67_ASAP7_75t_L g148 ( 
.A(n_62),
.B(n_74),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_36),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_45),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_14),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_40),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_52),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_70),
.B(n_4),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_13),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_43),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_9),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g158 ( 
.A(n_41),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_35),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

CKINVDCx11_ASAP7_75t_R g161 ( 
.A(n_120),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_2),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_92),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_92),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_99),
.Y(n_165)
);

AND2x6_ASAP7_75t_L g166 ( 
.A(n_121),
.B(n_48),
.Y(n_166)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_99),
.Y(n_167)
);

CKINVDCx6p67_ASAP7_75t_R g168 ( 
.A(n_134),
.Y(n_168)
);

AND2x6_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_49),
.Y(n_169)
);

AND2x4_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_3),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_99),
.Y(n_172)
);

AND2x4_ASAP7_75t_L g173 ( 
.A(n_128),
.B(n_91),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_144),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_93),
.Y(n_177)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_95),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_98),
.Y(n_179)
);

CKINVDCx6p67_ASAP7_75t_R g180 ( 
.A(n_95),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

OAI22x1_ASAP7_75t_SL g182 ( 
.A1(n_120),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_182)
);

AND2x4_ASAP7_75t_SL g183 ( 
.A(n_95),
.B(n_55),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_91),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_112),
.A2(n_11),
.B1(n_16),
.B2(n_18),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_94),
.Y(n_187)
);

AND2x4_ASAP7_75t_L g188 ( 
.A(n_107),
.B(n_19),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_147),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_113),
.B(n_19),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_100),
.Y(n_191)
);

AND2x6_ASAP7_75t_L g192 ( 
.A(n_107),
.B(n_57),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_147),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_126),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_159),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_99),
.Y(n_197)
);

OAI21x1_ASAP7_75t_L g198 ( 
.A1(n_101),
.A2(n_61),
.B(n_25),
.Y(n_198)
);

AND2x2_ASAP7_75t_SL g199 ( 
.A(n_103),
.B(n_64),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_137),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_104),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g202 ( 
.A(n_96),
.Y(n_202)
);

OAI22x1_ASAP7_75t_L g203 ( 
.A1(n_111),
.A2(n_20),
.B1(n_26),
.B2(n_28),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_105),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_109),
.Y(n_205)
);

AND2x4_ASAP7_75t_L g206 ( 
.A(n_123),
.B(n_20),
.Y(n_206)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_114),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_145),
.Y(n_208)
);

AND2x4_ASAP7_75t_L g209 ( 
.A(n_157),
.B(n_38),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_114),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_114),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_118),
.B(n_42),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_122),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_140),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_125),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_140),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_137),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_130),
.B(n_56),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_137),
.Y(n_219)
);

AND2x6_ASAP7_75t_L g220 ( 
.A(n_132),
.B(n_67),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_136),
.Y(n_221)
);

OAI21x1_ASAP7_75t_L g222 ( 
.A1(n_143),
.A2(n_69),
.B(n_76),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_146),
.Y(n_223)
);

OA21x2_ASAP7_75t_L g224 ( 
.A1(n_153),
.A2(n_156),
.B(n_148),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_168),
.B(n_155),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_178),
.B(n_117),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_178),
.B(n_142),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_170),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_170),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_170),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_174),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_165),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_176),
.Y(n_233)
);

BUFx10_ASAP7_75t_L g234 ( 
.A(n_183),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_176),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_209),
.B(n_110),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_165),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_181),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_181),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_184),
.Y(n_240)
);

NAND2xp33_ASAP7_75t_SL g241 ( 
.A(n_203),
.B(n_119),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_209),
.B(n_173),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_224),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_165),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_168),
.A2(n_119),
.B1(n_138),
.B2(n_131),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_188),
.Y(n_246)
);

INVx8_ASAP7_75t_L g247 ( 
.A(n_166),
.Y(n_247)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_166),
.Y(n_248)
);

AND2x4_ASAP7_75t_L g249 ( 
.A(n_173),
.B(n_137),
.Y(n_249)
);

NAND3xp33_ASAP7_75t_L g250 ( 
.A(n_208),
.B(n_129),
.C(n_151),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_197),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_206),
.Y(n_253)
);

AO22x2_ASAP7_75t_L g254 ( 
.A1(n_175),
.A2(n_186),
.B1(n_206),
.B2(n_199),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_177),
.B(n_116),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_180),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_177),
.B(n_102),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_179),
.B(n_139),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_160),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_224),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_162),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_190),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_179),
.B(n_141),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_191),
.B(n_115),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_191),
.B(n_108),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_195),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_202),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_190),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_185),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_185),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_210),
.Y(n_271)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_166),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_210),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_204),
.B(n_106),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_210),
.Y(n_275)
);

AND2x6_ASAP7_75t_L g276 ( 
.A(n_218),
.B(n_154),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_187),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_161),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_166),
.Y(n_279)
);

AND2x6_ASAP7_75t_L g280 ( 
.A(n_218),
.B(n_154),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_213),
.B(n_215),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_193),
.Y(n_282)
);

CKINVDCx6p67_ASAP7_75t_R g283 ( 
.A(n_202),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_196),
.Y(n_284)
);

AOI21x1_ASAP7_75t_L g285 ( 
.A1(n_212),
.A2(n_97),
.B(n_150),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_215),
.Y(n_286)
);

NAND2xp33_ASAP7_75t_L g287 ( 
.A(n_247),
.B(n_169),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_247),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_258),
.B(n_264),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_253),
.B(n_220),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_259),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_259),
.Y(n_292)
);

A2O1A1Ixp33_ASAP7_75t_L g293 ( 
.A1(n_243),
.A2(n_223),
.B(n_221),
.C(n_205),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_256),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_283),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_248),
.B(n_183),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_270),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_265),
.B(n_221),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_205),
.Y(n_299)
);

A2O1A1Ixp33_ASAP7_75t_L g300 ( 
.A1(n_243),
.A2(n_201),
.B(n_198),
.C(n_222),
.Y(n_300)
);

BUFx6f_ASAP7_75t_SL g301 ( 
.A(n_234),
.Y(n_301)
);

OAI21xp33_ASAP7_75t_L g302 ( 
.A1(n_260),
.A2(n_171),
.B(n_164),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_266),
.Y(n_303)
);

NOR3xp33_ASAP7_75t_L g304 ( 
.A(n_241),
.B(n_194),
.C(n_245),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_270),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_225),
.B(n_124),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_249),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_227),
.B(n_169),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_248),
.B(n_149),
.Y(n_309)
);

INVx8_ASAP7_75t_L g310 ( 
.A(n_247),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_254),
.A2(n_138),
.B1(n_163),
.B2(n_171),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_226),
.B(n_152),
.Y(n_312)
);

OR2x6_ASAP7_75t_L g313 ( 
.A(n_254),
.B(n_203),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_262),
.B(n_169),
.Y(n_314)
);

AND2x4_ASAP7_75t_L g315 ( 
.A(n_268),
.B(n_220),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_253),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_247),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_236),
.B(n_135),
.Y(n_318)
);

BUFx8_ASAP7_75t_L g319 ( 
.A(n_276),
.Y(n_319)
);

O2A1O1Ixp33_ASAP7_75t_L g320 ( 
.A1(n_228),
.A2(n_219),
.B(n_217),
.C(n_200),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_250),
.B(n_255),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_277),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_282),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_257),
.B(n_220),
.Y(n_324)
);

NOR3xp33_ASAP7_75t_L g325 ( 
.A(n_241),
.B(n_161),
.C(n_182),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_282),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_284),
.Y(n_327)
);

OR2x6_ASAP7_75t_L g328 ( 
.A(n_254),
.B(n_189),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_284),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_278),
.B(n_189),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_256),
.B(n_169),
.Y(n_331)
);

BUFx5_ASAP7_75t_L g332 ( 
.A(n_279),
.Y(n_332)
);

AO22x2_ASAP7_75t_L g333 ( 
.A1(n_254),
.A2(n_242),
.B1(n_230),
.B2(n_229),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_263),
.B(n_192),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_276),
.A2(n_192),
.B1(n_217),
.B2(n_200),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_276),
.B(n_192),
.Y(n_336)
);

INVx2_ASAP7_75t_SL g337 ( 
.A(n_234),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_267),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_272),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_276),
.B(n_280),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_269),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_286),
.B(n_280),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_307),
.Y(n_343)
);

OAI21xp33_ASAP7_75t_L g344 ( 
.A1(n_302),
.A2(n_299),
.B(n_293),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_291),
.Y(n_345)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_310),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_287),
.A2(n_272),
.B(n_246),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_290),
.A2(n_272),
.B(n_274),
.Y(n_348)
);

NOR2xp67_ASAP7_75t_L g349 ( 
.A(n_295),
.B(n_285),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_292),
.Y(n_350)
);

OR2x2_ASAP7_75t_L g351 ( 
.A(n_306),
.B(n_238),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_316),
.Y(n_352)
);

BUFx4f_ASAP7_75t_L g353 ( 
.A(n_313),
.Y(n_353)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_307),
.Y(n_354)
);

INVx2_ASAP7_75t_SL g355 ( 
.A(n_338),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_308),
.A2(n_240),
.B(n_239),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_336),
.A2(n_239),
.B(n_238),
.Y(n_357)
);

A2O1A1Ixp33_ASAP7_75t_L g358 ( 
.A1(n_314),
.A2(n_235),
.B(n_233),
.C(n_231),
.Y(n_358)
);

OR2x6_ASAP7_75t_L g359 ( 
.A(n_328),
.B(n_280),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_298),
.B(n_192),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_321),
.B(n_172),
.Y(n_361)
);

O2A1O1Ixp33_ASAP7_75t_L g362 ( 
.A1(n_311),
.A2(n_313),
.B(n_304),
.C(n_340),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_289),
.B(n_172),
.Y(n_363)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_310),
.Y(n_364)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_310),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_341),
.B(n_172),
.Y(n_366)
);

AND2x4_ASAP7_75t_L g367 ( 
.A(n_337),
.B(n_78),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_288),
.B(n_317),
.Y(n_368)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_301),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_301),
.B(n_79),
.Y(n_370)
);

AO21x1_ASAP7_75t_L g371 ( 
.A1(n_335),
.A2(n_244),
.B(n_275),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_288),
.B(n_167),
.Y(n_372)
);

A2O1A1Ixp33_ASAP7_75t_L g373 ( 
.A1(n_324),
.A2(n_216),
.B(n_214),
.C(n_211),
.Y(n_373)
);

A2O1A1Ixp33_ASAP7_75t_L g374 ( 
.A1(n_302),
.A2(n_214),
.B(n_216),
.C(n_271),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_330),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_294),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_322),
.B(n_207),
.Y(n_377)
);

BUFx12f_ASAP7_75t_L g378 ( 
.A(n_328),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_317),
.B(n_319),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_318),
.B(n_80),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_333),
.A2(n_207),
.B1(n_216),
.B2(n_214),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_315),
.A2(n_252),
.B(n_273),
.Y(n_382)
);

NAND3xp33_ASAP7_75t_L g383 ( 
.A(n_320),
.B(n_216),
.C(n_214),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_296),
.A2(n_309),
.B(n_334),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_297),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_312),
.B(n_86),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_331),
.B(n_87),
.Y(n_387)
);

CKINVDCx6p67_ASAP7_75t_R g388 ( 
.A(n_328),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_342),
.A2(n_326),
.B(n_323),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_351),
.Y(n_390)
);

AOI221xp5_ASAP7_75t_L g391 ( 
.A1(n_375),
.A2(n_325),
.B1(n_329),
.B2(n_327),
.C(n_305),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_355),
.B(n_319),
.Y(n_392)
);

INVx4_ASAP7_75t_SL g393 ( 
.A(n_378),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_353),
.A2(n_339),
.B1(n_237),
.B2(n_251),
.Y(n_394)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_376),
.B(n_332),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_346),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g397 ( 
.A(n_369),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_359),
.B(n_232),
.Y(n_398)
);

A2O1A1Ixp33_ASAP7_75t_L g399 ( 
.A1(n_362),
.A2(n_232),
.B(n_237),
.C(n_251),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_356),
.A2(n_232),
.B(n_237),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_357),
.A2(n_251),
.B(n_344),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_359),
.B(n_388),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_344),
.A2(n_358),
.B(n_360),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_352),
.B(n_365),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_347),
.A2(n_348),
.B(n_363),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_364),
.B(n_365),
.Y(n_406)
);

OA21x2_ASAP7_75t_L g407 ( 
.A1(n_374),
.A2(n_381),
.B(n_373),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_367),
.Y(n_408)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_353),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_384),
.A2(n_361),
.B(n_382),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_379),
.A2(n_380),
.B1(n_349),
.B2(n_386),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_343),
.B(n_354),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_385),
.Y(n_413)
);

NAND3xp33_ASAP7_75t_L g414 ( 
.A(n_383),
.B(n_387),
.C(n_370),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_383),
.A2(n_345),
.B1(n_350),
.B2(n_377),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_368),
.A2(n_366),
.B(n_372),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_351),
.B(n_286),
.Y(n_417)
);

OA22x2_ASAP7_75t_L g418 ( 
.A1(n_359),
.A2(n_328),
.B1(n_303),
.B2(n_245),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_346),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_351),
.B(n_286),
.Y(n_420)
);

OA22x2_ASAP7_75t_L g421 ( 
.A1(n_359),
.A2(n_328),
.B1(n_303),
.B2(n_245),
.Y(n_421)
);

OA22x2_ASAP7_75t_L g422 ( 
.A1(n_359),
.A2(n_328),
.B1(n_303),
.B2(n_245),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_351),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_375),
.B(n_303),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_355),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_359),
.A2(n_313),
.B1(n_311),
.B2(n_328),
.Y(n_426)
);

AO31x2_ASAP7_75t_L g427 ( 
.A1(n_371),
.A2(n_300),
.A3(n_374),
.B(n_373),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g428 ( 
.A(n_375),
.B(n_303),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_351),
.B(n_286),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_351),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_375),
.B(n_303),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_351),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_351),
.B(n_286),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_346),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_351),
.B(n_286),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_346),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_355),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_355),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_346),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_359),
.A2(n_313),
.B1(n_311),
.B2(n_328),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_396),
.Y(n_441)
);

NAND2x1p5_ASAP7_75t_L g442 ( 
.A(n_396),
.B(n_409),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_410),
.A2(n_401),
.B(n_405),
.Y(n_443)
);

INVx2_ASAP7_75t_SL g444 ( 
.A(n_396),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_390),
.Y(n_445)
);

AO22x2_ASAP7_75t_L g446 ( 
.A1(n_426),
.A2(n_440),
.B1(n_394),
.B2(n_415),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_401),
.A2(n_403),
.B(n_400),
.Y(n_447)
);

NAND2x1p5_ASAP7_75t_L g448 ( 
.A(n_409),
.B(n_419),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_423),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_403),
.A2(n_400),
.B(n_399),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_418),
.A2(n_422),
.B1(n_421),
.B2(n_440),
.Y(n_451)
);

OAI211xp5_ASAP7_75t_SL g452 ( 
.A1(n_426),
.A2(n_391),
.B(n_428),
.C(n_432),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_437),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_417),
.Y(n_454)
);

NAND3xp33_ASAP7_75t_L g455 ( 
.A(n_414),
.B(n_431),
.C(n_411),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_430),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_419),
.B(n_434),
.Y(n_457)
);

INVx3_ASAP7_75t_SL g458 ( 
.A(n_393),
.Y(n_458)
);

BUFx4f_ASAP7_75t_L g459 ( 
.A(n_436),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_424),
.B(n_435),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_420),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_439),
.B(n_429),
.Y(n_462)
);

AND2x4_ASAP7_75t_L g463 ( 
.A(n_439),
.B(n_433),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_425),
.B(n_438),
.Y(n_464)
);

AND2x6_ASAP7_75t_L g465 ( 
.A(n_402),
.B(n_398),
.Y(n_465)
);

BUFx12f_ASAP7_75t_L g466 ( 
.A(n_397),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_406),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_393),
.B(n_404),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_408),
.A2(n_411),
.B1(n_414),
.B2(n_413),
.Y(n_469)
);

OA21x2_ASAP7_75t_L g470 ( 
.A1(n_389),
.A2(n_416),
.B(n_427),
.Y(n_470)
);

NOR2xp67_ASAP7_75t_L g471 ( 
.A(n_392),
.B(n_395),
.Y(n_471)
);

OA21x2_ASAP7_75t_L g472 ( 
.A1(n_427),
.A2(n_412),
.B(n_407),
.Y(n_472)
);

BUFx12f_ASAP7_75t_L g473 ( 
.A(n_397),
.Y(n_473)
);

AND2x6_ASAP7_75t_L g474 ( 
.A(n_426),
.B(n_440),
.Y(n_474)
);

NOR2x1_ASAP7_75t_L g475 ( 
.A(n_409),
.B(n_369),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_409),
.B(n_439),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_408),
.B(n_353),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_390),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_424),
.B(n_303),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_425),
.Y(n_480)
);

OA21x2_ASAP7_75t_L g481 ( 
.A1(n_443),
.A2(n_450),
.B(n_447),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_467),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_454),
.B(n_460),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_453),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_458),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_453),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_454),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_467),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_474),
.B(n_461),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_441),
.Y(n_490)
);

BUFx12f_ASAP7_75t_L g491 ( 
.A(n_466),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_465),
.B(n_455),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_472),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_451),
.B(n_469),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_487),
.Y(n_495)
);

OR2x2_ASAP7_75t_L g496 ( 
.A(n_483),
.B(n_487),
.Y(n_496)
);

INVx4_ASAP7_75t_L g497 ( 
.A(n_490),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_489),
.B(n_446),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_488),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_489),
.B(n_446),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_483),
.B(n_472),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_493),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_488),
.Y(n_503)
);

INVxp67_ASAP7_75t_R g504 ( 
.A(n_491),
.Y(n_504)
);

BUFx2_ASAP7_75t_L g505 ( 
.A(n_482),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_482),
.B(n_468),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_491),
.B(n_479),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_481),
.B(n_470),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_502),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_495),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_498),
.B(n_481),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_495),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_505),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_496),
.Y(n_514)
);

INVxp33_ASAP7_75t_L g515 ( 
.A(n_506),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_498),
.B(n_481),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_514),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_509),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_510),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_512),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_511),
.B(n_508),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_511),
.B(n_508),
.Y(n_522)
);

NAND2x1p5_ASAP7_75t_L g523 ( 
.A(n_509),
.B(n_497),
.Y(n_523)
);

INVx1_ASAP7_75t_SL g524 ( 
.A(n_515),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_516),
.B(n_501),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_513),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_517),
.B(n_524),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_SL g528 ( 
.A1(n_523),
.A2(n_499),
.B(n_503),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_526),
.B(n_516),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_519),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_521),
.B(n_505),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_521),
.B(n_500),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_521),
.A2(n_492),
.B1(n_494),
.B2(n_515),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_518),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_530),
.B(n_525),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_531),
.B(n_532),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_529),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_527),
.B(n_491),
.Y(n_538)
);

INVxp67_ASAP7_75t_L g539 ( 
.A(n_528),
.Y(n_539)
);

AOI32xp33_ASAP7_75t_L g540 ( 
.A1(n_528),
.A2(n_522),
.A3(n_525),
.B1(n_492),
.B2(n_507),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_534),
.B(n_522),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_536),
.B(n_522),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_538),
.B(n_533),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_537),
.B(n_520),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_539),
.B(n_523),
.Y(n_545)
);

NOR3xp33_ASAP7_75t_L g546 ( 
.A(n_543),
.B(n_540),
.C(n_452),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_SL g547 ( 
.A1(n_543),
.A2(n_535),
.B1(n_541),
.B2(n_492),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_SL g548 ( 
.A1(n_545),
.A2(n_504),
.B(n_494),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_546),
.Y(n_549)
);

NOR2x1_ASAP7_75t_L g550 ( 
.A(n_548),
.B(n_504),
.Y(n_550)
);

NOR3x1_ASAP7_75t_L g551 ( 
.A(n_549),
.B(n_544),
.C(n_535),
.Y(n_551)
);

NAND3x1_ASAP7_75t_L g552 ( 
.A(n_550),
.B(n_475),
.C(n_458),
.Y(n_552)
);

NOR2x1_ASAP7_75t_SL g553 ( 
.A(n_552),
.B(n_473),
.Y(n_553)
);

NOR2xp67_ASAP7_75t_L g554 ( 
.A(n_551),
.B(n_485),
.Y(n_554)
);

OAI211xp5_ASAP7_75t_L g555 ( 
.A1(n_554),
.A2(n_547),
.B(n_480),
.C(n_464),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_553),
.A2(n_480),
.B1(n_542),
.B2(n_492),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_555),
.B(n_468),
.Y(n_557)
);

XOR2x2_ASAP7_75t_L g558 ( 
.A(n_556),
.B(n_442),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_557),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_558),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_558),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_557),
.Y(n_562)
);

A2O1A1Ixp33_ASAP7_75t_L g563 ( 
.A1(n_559),
.A2(n_471),
.B(n_484),
.C(n_486),
.Y(n_563)
);

NOR3xp33_ASAP7_75t_L g564 ( 
.A(n_560),
.B(n_476),
.C(n_452),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_561),
.B(n_459),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_560),
.Y(n_566)
);

OAI21x1_ASAP7_75t_L g567 ( 
.A1(n_566),
.A2(n_562),
.B(n_442),
.Y(n_567)
);

AOI21x1_ASAP7_75t_L g568 ( 
.A1(n_565),
.A2(n_564),
.B(n_563),
.Y(n_568)
);

AOI221xp5_ASAP7_75t_L g569 ( 
.A1(n_568),
.A2(n_478),
.B1(n_445),
.B2(n_449),
.C(n_456),
.Y(n_569)
);

AOI221xp5_ASAP7_75t_L g570 ( 
.A1(n_567),
.A2(n_476),
.B1(n_459),
.B2(n_477),
.C(n_457),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_L g571 ( 
.A1(n_570),
.A2(n_448),
.B(n_477),
.Y(n_571)
);

OAI21x1_ASAP7_75t_L g572 ( 
.A1(n_571),
.A2(n_569),
.B(n_448),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_572),
.A2(n_444),
.B1(n_463),
.B2(n_462),
.Y(n_573)
);


endmodule