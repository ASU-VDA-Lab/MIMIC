module real_aes_8492_n_350 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_350);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_350;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_1004;
wire n_580;
wire n_469;
wire n_987;
wire n_362;
wire n_979;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_841;
wire n_718;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_1014;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_742;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_353;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_666;
wire n_551;
wire n_537;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_856;
wire n_594;
wire n_983;
wire n_767;
wire n_889;
wire n_696;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_932;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1021;
wire n_958;
wire n_677;
wire n_1046;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_994;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_992;
wire n_774;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_1053;
wire n_636;
wire n_559;
wire n_872;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_1025;
wire n_755;
wire n_409;
wire n_748;
wire n_860;
wire n_781;
wire n_523;
wire n_996;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_1049;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_455;
wire n_725;
wire n_973;
wire n_671;
wire n_960;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_1017;
wire n_737;
wire n_1013;
wire n_936;
wire n_581;
wire n_610;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_867;
wire n_745;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_676;
wire n_658;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1037;
wire n_1031;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_999;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_488;
wire n_501;
wire n_1041;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_1028;
wire n_366;
wire n_727;
wire n_649;
wire n_397;
wire n_358;
wire n_385;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_354;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_365;
wire n_899;
wire n_526;
wire n_653;
wire n_637;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_575;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_587;
wire n_546;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_911;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_1045;
wire n_566;
wire n_719;
wire n_837;
wire n_967;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1024;
wire n_842;
wire n_849;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_797;
wire n_668;
wire n_862;
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_0), .A2(n_177), .B1(n_643), .B2(n_986), .Y(n_985) );
INVx1_ASAP7_75t_L g878 ( .A(n_1), .Y(n_878) );
AOI222xp33_ASAP7_75t_L g1028 ( .A1(n_2), .A2(n_169), .B1(n_306), .B2(n_445), .C1(n_469), .C2(n_671), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_3), .A2(n_235), .B1(n_515), .B2(n_572), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_4), .A2(n_102), .B1(n_368), .B2(n_384), .Y(n_367) );
AOI22xp33_ASAP7_75t_SL g552 ( .A1(n_5), .A2(n_154), .B1(n_553), .B2(n_554), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g498 ( .A1(n_6), .A2(n_91), .B1(n_499), .B2(n_502), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_7), .A2(n_75), .B1(n_445), .B2(n_706), .Y(n_726) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_8), .B(n_547), .Y(n_546) );
AO22x2_ASAP7_75t_L g383 ( .A1(n_9), .A2(n_205), .B1(n_374), .B2(n_379), .Y(n_383) );
INVx1_ASAP7_75t_L g1012 ( .A(n_9), .Y(n_1012) );
AOI22xp5_ASAP7_75t_SL g1055 ( .A1(n_10), .A2(n_346), .B1(n_386), .B2(n_418), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_11), .A2(n_163), .B1(n_512), .B2(n_645), .Y(n_1022) );
AOI22xp33_ASAP7_75t_SL g815 ( .A1(n_12), .A2(n_330), .B1(n_466), .B2(n_751), .Y(n_815) );
AOI22xp5_ASAP7_75t_L g967 ( .A1(n_13), .A2(n_150), .B1(n_386), .B2(n_558), .Y(n_967) );
AOI22xp5_ASAP7_75t_SL g1051 ( .A1(n_14), .A2(n_223), .B1(n_528), .B2(n_988), .Y(n_1051) );
CKINVDCx20_ASAP7_75t_R g939 ( .A(n_15), .Y(n_939) );
CKINVDCx20_ASAP7_75t_R g950 ( .A(n_16), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_17), .A2(n_184), .B1(n_424), .B2(n_520), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_18), .A2(n_230), .B1(n_386), .B2(n_528), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_19), .A2(n_296), .B1(n_404), .B2(n_407), .Y(n_403) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_20), .Y(n_786) );
AOI222xp33_ASAP7_75t_L g531 ( .A1(n_21), .A2(n_60), .B1(n_258), .B2(n_466), .C1(n_532), .C2(n_534), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_22), .A2(n_214), .B1(n_492), .B2(n_494), .Y(n_650) );
AOI22xp5_ASAP7_75t_SL g803 ( .A1(n_23), .A2(n_228), .B1(n_558), .B2(n_804), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g957 ( .A(n_24), .Y(n_957) );
AOI22xp33_ASAP7_75t_SL g1049 ( .A1(n_25), .A2(n_182), .B1(n_748), .B2(n_751), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_26), .A2(n_334), .B1(n_530), .B2(n_554), .Y(n_968) );
CKINVDCx20_ASAP7_75t_R g933 ( .A(n_27), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_28), .A2(n_226), .B1(n_502), .B2(n_512), .Y(n_755) );
AO22x2_ASAP7_75t_L g381 ( .A1(n_29), .A2(n_119), .B1(n_374), .B2(n_375), .Y(n_381) );
INVx1_ASAP7_75t_L g618 ( .A(n_30), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_31), .A2(n_166), .B1(n_398), .B2(n_416), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_32), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g973 ( .A1(n_33), .A2(n_974), .B1(n_992), .B2(n_993), .Y(n_973) );
INVx1_ASAP7_75t_L g993 ( .A(n_33), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_34), .A2(n_48), .B1(n_502), .B2(n_636), .Y(n_789) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_35), .Y(n_479) );
AOI22xp33_ASAP7_75t_SL g758 ( .A1(n_36), .A2(n_55), .B1(n_493), .B2(n_645), .Y(n_758) );
INVx1_ASAP7_75t_L g856 ( .A(n_37), .Y(n_856) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_38), .A2(n_269), .B1(n_445), .B2(n_748), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g826 ( .A1(n_39), .A2(n_56), .B1(n_370), .B2(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g592 ( .A(n_40), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_41), .A2(n_158), .B1(n_512), .B2(n_685), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_42), .A2(n_281), .B1(n_368), .B2(n_415), .Y(n_990) );
INVx1_ASAP7_75t_L g915 ( .A(n_43), .Y(n_915) );
AOI22xp5_ASAP7_75t_L g854 ( .A1(n_44), .A2(n_195), .B1(n_434), .B2(n_446), .Y(n_854) );
AOI222xp33_ASAP7_75t_L g437 ( .A1(n_45), .A2(n_276), .B1(n_295), .B2(n_438), .C1(n_440), .C2(n_444), .Y(n_437) );
AOI22xp5_ASAP7_75t_SL g802 ( .A1(n_46), .A2(n_292), .B1(n_515), .B2(n_709), .Y(n_802) );
AOI22xp5_ASAP7_75t_SL g825 ( .A1(n_47), .A2(n_204), .B1(n_386), .B2(n_709), .Y(n_825) );
CKINVDCx20_ASAP7_75t_R g937 ( .A(n_49), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_50), .A2(n_168), .B1(n_494), .B2(n_680), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_51), .A2(n_302), .B1(n_522), .B2(n_523), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_52), .A2(n_279), .B1(n_664), .B2(n_666), .Y(n_663) );
CKINVDCx16_ASAP7_75t_R g929 ( .A(n_53), .Y(n_929) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_54), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_57), .B(n_444), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_58), .Y(n_760) );
AOI22xp33_ASAP7_75t_SL g898 ( .A1(n_59), .A2(n_227), .B1(n_587), .B2(n_899), .Y(n_898) );
AOI22xp5_ASAP7_75t_L g916 ( .A1(n_61), .A2(n_90), .B1(n_445), .B2(n_523), .Y(n_916) );
INVx1_ASAP7_75t_L g625 ( .A(n_62), .Y(n_625) );
AOI22xp33_ASAP7_75t_SL g550 ( .A1(n_63), .A2(n_125), .B1(n_526), .B2(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g1038 ( .A(n_64), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_65), .A2(n_322), .B1(n_643), .B2(n_645), .Y(n_642) );
INVx1_ASAP7_75t_L g876 ( .A(n_66), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_67), .A2(n_140), .B1(n_649), .B2(n_683), .Y(n_795) );
NAND2xp5_ASAP7_75t_SL g865 ( .A(n_68), .B(n_807), .Y(n_865) );
CKINVDCx20_ASAP7_75t_R g977 ( .A(n_69), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_70), .A2(n_89), .B1(n_734), .B2(n_735), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_71), .A2(n_201), .B1(n_424), .B2(n_428), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g965 ( .A(n_72), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_73), .A2(n_211), .B1(n_488), .B2(n_489), .Y(n_487) );
AOI22xp5_ASAP7_75t_SL g1052 ( .A1(n_74), .A2(n_234), .B1(n_393), .B2(n_1053), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_76), .A2(n_95), .B1(n_572), .B2(n_791), .Y(n_790) );
AOI22xp33_ASAP7_75t_SL g902 ( .A1(n_77), .A2(n_209), .B1(n_516), .B2(n_830), .Y(n_902) );
AOI22xp5_ASAP7_75t_SL g829 ( .A1(n_78), .A2(n_96), .B1(n_502), .B2(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g602 ( .A(n_79), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_80), .A2(n_143), .B1(n_497), .B2(n_683), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_81), .A2(n_149), .B1(n_585), .B2(n_587), .Y(n_584) );
AO22x2_ASAP7_75t_L g378 ( .A1(n_82), .A2(n_239), .B1(n_374), .B2(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g1009 ( .A(n_82), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_83), .A2(n_248), .B1(n_398), .B2(n_530), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_84), .A2(n_325), .B1(n_534), .B2(n_596), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_85), .A2(n_323), .B1(n_513), .B2(n_685), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_86), .A2(n_338), .B1(n_680), .B2(n_797), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_87), .A2(n_272), .B1(n_427), .B2(n_519), .Y(n_981) );
AOI22xp5_ASAP7_75t_L g978 ( .A1(n_88), .A2(n_199), .B1(n_444), .B2(n_979), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_92), .A2(n_266), .B1(n_492), .B2(n_494), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_93), .A2(n_288), .B1(n_551), .B2(n_827), .Y(n_969) );
OA22x2_ASAP7_75t_L g363 ( .A1(n_94), .A2(n_364), .B1(n_365), .B2(n_448), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_94), .Y(n_364) );
AOI22xp33_ASAP7_75t_SL g831 ( .A1(n_97), .A2(n_191), .B1(n_415), .B2(n_807), .Y(n_831) );
AOI22xp5_ASAP7_75t_L g920 ( .A1(n_98), .A2(n_115), .B1(n_502), .B2(n_526), .Y(n_920) );
INVx1_ASAP7_75t_L g590 ( .A(n_99), .Y(n_590) );
AOI22xp33_ASAP7_75t_SL g750 ( .A1(n_100), .A2(n_107), .B1(n_440), .B2(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g822 ( .A(n_101), .Y(n_822) );
AOI22xp5_ASAP7_75t_SL g1056 ( .A1(n_103), .A2(n_196), .B1(n_407), .B2(n_516), .Y(n_1056) );
INVx1_ASAP7_75t_L g573 ( .A(n_104), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_105), .A2(n_124), .B1(n_501), .B2(n_988), .Y(n_987) );
AOI22xp33_ASAP7_75t_SL g891 ( .A1(n_106), .A2(n_152), .B1(n_430), .B2(n_666), .Y(n_891) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_108), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g811 ( .A(n_109), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g864 ( .A(n_110), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_111), .B(n_911), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_112), .A2(n_136), .B1(n_404), .B2(n_648), .Y(n_647) );
CKINVDCx20_ASAP7_75t_R g857 ( .A(n_113), .Y(n_857) );
CKINVDCx20_ASAP7_75t_R g662 ( .A(n_114), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_116), .A2(n_257), .B1(n_516), .B2(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g579 ( .A(n_117), .Y(n_579) );
INVx1_ASAP7_75t_L g704 ( .A(n_118), .Y(n_704) );
INVx1_ASAP7_75t_L g1013 ( .A(n_119), .Y(n_1013) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_120), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_121), .A2(n_187), .B1(n_431), .B2(n_702), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_122), .A2(n_128), .B1(n_415), .B2(n_711), .Y(n_923) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_123), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_126), .A2(n_190), .B1(n_488), .B2(n_489), .Y(n_678) );
CKINVDCx20_ASAP7_75t_R g835 ( .A(n_127), .Y(n_835) );
AOI211xp5_ASAP7_75t_L g931 ( .A1(n_129), .A2(n_438), .B(n_932), .C(n_936), .Y(n_931) );
INVx1_ASAP7_75t_L g715 ( .A(n_130), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g861 ( .A(n_131), .Y(n_861) );
CKINVDCx20_ASAP7_75t_R g659 ( .A(n_132), .Y(n_659) );
INVx1_ASAP7_75t_L g924 ( .A(n_133), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_134), .A2(n_308), .B1(n_413), .B2(n_418), .Y(n_412) );
AOI22xp5_ASAP7_75t_L g756 ( .A1(n_135), .A2(n_165), .B1(n_526), .B2(n_713), .Y(n_756) );
AOI22xp5_ASAP7_75t_L g839 ( .A1(n_137), .A2(n_238), .B1(n_600), .B2(n_668), .Y(n_839) );
AOI22xp33_ASAP7_75t_SL g635 ( .A1(n_138), .A2(n_221), .B1(n_636), .B2(n_639), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_139), .A2(n_332), .B1(n_466), .B2(n_751), .Y(n_913) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_141), .A2(n_568), .B1(n_606), .B2(n_607), .Y(n_567) );
CKINVDCx16_ASAP7_75t_R g606 ( .A(n_141), .Y(n_606) );
AOI22xp33_ASAP7_75t_SL g1045 ( .A1(n_142), .A2(n_321), .B1(n_445), .B2(n_624), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_144), .A2(n_244), .B1(n_407), .B2(n_497), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g1020 ( .A1(n_145), .A2(n_174), .B1(n_398), .B2(n_493), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_146), .A2(n_331), .B1(n_430), .B2(n_666), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_147), .A2(n_251), .B1(n_430), .B2(n_434), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_148), .A2(n_216), .B1(n_492), .B2(n_587), .Y(n_991) );
AND2x6_ASAP7_75t_L g353 ( .A(n_151), .B(n_354), .Y(n_353) );
HB1xp67_ASAP7_75t_L g1006 ( .A(n_151), .Y(n_1006) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_153), .A2(n_283), .B1(n_415), .B2(n_577), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g859 ( .A(n_155), .Y(n_859) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_156), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g841 ( .A(n_157), .Y(n_841) );
AOI22xp33_ASAP7_75t_SL g922 ( .A1(n_159), .A2(n_327), .B1(n_493), .B2(n_793), .Y(n_922) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_160), .A2(n_220), .B1(n_434), .B2(n_445), .Y(n_813) );
AOI22xp33_ASAP7_75t_SL g556 ( .A1(n_161), .A2(n_339), .B1(n_502), .B2(n_512), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g559 ( .A(n_162), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_164), .A2(n_246), .B1(n_393), .B2(n_397), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_167), .A2(n_347), .B1(n_472), .B2(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g597 ( .A(n_170), .Y(n_597) );
AOI22xp33_ASAP7_75t_SL g710 ( .A1(n_171), .A2(n_175), .B1(n_649), .B2(n_711), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_172), .Y(n_784) );
AO22x2_ASAP7_75t_L g373 ( .A1(n_173), .A2(n_229), .B1(n_374), .B2(n_375), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g1010 ( .A(n_173), .B(n_1011), .Y(n_1010) );
CKINVDCx20_ASAP7_75t_R g958 ( .A(n_176), .Y(n_958) );
AOI22xp33_ASAP7_75t_SL g557 ( .A1(n_178), .A2(n_245), .B1(n_515), .B2(n_558), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_179), .A2(n_286), .B1(n_600), .B2(n_889), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_180), .A2(n_231), .B1(n_713), .B2(n_827), .Y(n_1019) );
AOI22xp33_ASAP7_75t_SL g712 ( .A1(n_181), .A2(n_318), .B1(n_386), .B2(n_713), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_183), .Y(n_473) );
AOI22xp5_ASAP7_75t_SL g806 ( .A1(n_185), .A2(n_253), .B1(n_577), .B2(n_807), .Y(n_806) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_186), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_188), .A2(n_218), .B1(n_512), .B2(n_513), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_189), .Y(n_775) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_192), .A2(n_314), .B1(n_398), .B2(n_413), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_193), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g1026 ( .A(n_194), .B(n_699), .Y(n_1026) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_197), .Y(n_780) );
AOI22xp33_ASAP7_75t_SL g738 ( .A1(n_198), .A2(n_342), .B1(n_368), .B2(n_709), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g946 ( .A(n_200), .Y(n_946) );
INVx1_ASAP7_75t_L g622 ( .A(n_202), .Y(n_622) );
CKINVDCx20_ASAP7_75t_R g960 ( .A(n_203), .Y(n_960) );
NAND2xp5_ASAP7_75t_SL g1048 ( .A(n_206), .B(n_423), .Y(n_1048) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_207), .A2(n_453), .B1(n_503), .B2(n_504), .Y(n_452) );
INVx1_ASAP7_75t_L g503 ( .A(n_207), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_208), .A2(n_328), .B1(n_413), .B2(n_418), .Y(n_943) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_210), .B(n_520), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_212), .A2(n_274), .B1(n_664), .B2(n_666), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_213), .A2(n_337), .B1(n_513), .B2(n_649), .Y(n_1023) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_215), .Y(n_817) );
AOI22xp33_ASAP7_75t_SL g896 ( .A1(n_217), .A2(n_249), .B1(n_577), .B2(n_897), .Y(n_896) );
AOI22xp5_ASAP7_75t_SL g612 ( .A1(n_219), .A2(n_613), .B1(n_651), .B2(n_652), .Y(n_612) );
INVx1_ASAP7_75t_L g652 ( .A(n_219), .Y(n_652) );
CKINVDCx20_ASAP7_75t_R g1044 ( .A(n_222), .Y(n_1044) );
INVx2_ASAP7_75t_L g358 ( .A(n_224), .Y(n_358) );
AOI22xp33_ASAP7_75t_SL g543 ( .A1(n_225), .A2(n_301), .B1(n_446), .B2(n_466), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_232), .A2(n_243), .B1(n_515), .B2(n_516), .Y(n_514) );
INVx1_ASAP7_75t_L g616 ( .A(n_233), .Y(n_616) );
INVx1_ASAP7_75t_L g631 ( .A(n_236), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_237), .A2(n_291), .B1(n_526), .B2(n_528), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_240), .A2(n_290), .B1(n_553), .B2(n_587), .Y(n_944) );
INVx1_ASAP7_75t_L g853 ( .A(n_241), .Y(n_853) );
CKINVDCx20_ASAP7_75t_R g887 ( .A(n_242), .Y(n_887) );
CKINVDCx20_ASAP7_75t_R g781 ( .A(n_247), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_250), .A2(n_294), .B1(n_423), .B2(n_427), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_252), .B(n_520), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g873 ( .A(n_254), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_255), .A2(n_304), .B1(n_636), .B2(n_687), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_256), .A2(n_335), .B1(n_519), .B2(n_520), .Y(n_518) );
AOI22xp33_ASAP7_75t_SL g903 ( .A1(n_259), .A2(n_349), .B1(n_572), .B2(n_734), .Y(n_903) );
CKINVDCx20_ASAP7_75t_R g836 ( .A(n_260), .Y(n_836) );
INVx1_ASAP7_75t_L g374 ( .A(n_261), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_261), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_262), .A2(n_268), .B1(n_423), .B2(n_893), .Y(n_892) );
INVx1_ASAP7_75t_L g723 ( .A(n_263), .Y(n_723) );
INVx1_ASAP7_75t_L g594 ( .A(n_264), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_265), .A2(n_656), .B1(n_688), .B2(n_689), .Y(n_655) );
CKINVDCx20_ASAP7_75t_R g688 ( .A(n_265), .Y(n_688) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_267), .Y(n_777) );
CKINVDCx20_ASAP7_75t_R g867 ( .A(n_270), .Y(n_867) );
CKINVDCx20_ASAP7_75t_R g871 ( .A(n_271), .Y(n_871) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_273), .A2(n_311), .B1(n_418), .B2(n_526), .Y(n_714) );
INVx1_ASAP7_75t_L g722 ( .A(n_275), .Y(n_722) );
INVx1_ASAP7_75t_L g583 ( .A(n_277), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g843 ( .A(n_278), .Y(n_843) );
AOI211xp5_ASAP7_75t_L g350 ( .A1(n_280), .A2(n_351), .B(n_359), .C(n_1014), .Y(n_350) );
AOI22xp33_ASAP7_75t_SL g548 ( .A1(n_282), .A2(n_320), .B1(n_431), .B2(n_523), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_284), .B(n_627), .Y(n_626) );
CKINVDCx20_ASAP7_75t_R g672 ( .A(n_285), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g964 ( .A(n_287), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_289), .A2(n_312), .B1(n_668), .B2(n_751), .Y(n_1027) );
AO22x2_ASAP7_75t_L g953 ( .A1(n_293), .A2(n_954), .B1(n_971), .B2(n_972), .Y(n_953) );
CKINVDCx20_ASAP7_75t_R g972 ( .A(n_293), .Y(n_972) );
CKINVDCx20_ASAP7_75t_R g882 ( .A(n_297), .Y(n_882) );
AND2x2_ASAP7_75t_L g357 ( .A(n_298), .B(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_299), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g354 ( .A(n_300), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_303), .B(n_699), .Y(n_912) );
INVx1_ASAP7_75t_L g605 ( .A(n_305), .Y(n_605) );
INVx1_ASAP7_75t_L g879 ( .A(n_307), .Y(n_879) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_309), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_310), .B(n_519), .Y(n_934) );
AOI22xp5_ASAP7_75t_L g1015 ( .A1(n_313), .A2(n_1016), .B1(n_1017), .B2(n_1029), .Y(n_1015) );
CKINVDCx20_ASAP7_75t_R g1029 ( .A(n_313), .Y(n_1029) );
CKINVDCx20_ASAP7_75t_R g868 ( .A(n_315), .Y(n_868) );
CKINVDCx20_ASAP7_75t_R g838 ( .A(n_316), .Y(n_838) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_317), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g1025 ( .A(n_319), .Y(n_1025) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_324), .Y(n_730) );
INVx1_ASAP7_75t_L g951 ( .A(n_326), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_329), .B(n_699), .Y(n_698) );
CKINVDCx20_ASAP7_75t_R g948 ( .A(n_333), .Y(n_948) );
INVx1_ASAP7_75t_L g629 ( .A(n_336), .Y(n_629) );
INVx1_ASAP7_75t_L g575 ( .A(n_340), .Y(n_575) );
CKINVDCx20_ASAP7_75t_R g675 ( .A(n_341), .Y(n_675) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_343), .Y(n_725) );
OA22x2_ASAP7_75t_L g770 ( .A1(n_344), .A2(n_771), .B1(n_772), .B2(n_798), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_344), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_345), .B(n_893), .Y(n_1047) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_348), .Y(n_746) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
HB1xp67_ASAP7_75t_L g1005 ( .A(n_354), .Y(n_1005) );
OAI21xp5_ASAP7_75t_L g1036 ( .A1(n_355), .A2(n_1004), .B(n_1037), .Y(n_1036) );
CKINVDCx20_ASAP7_75t_R g355 ( .A(n_356), .Y(n_355) );
INVxp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AOI221xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_763), .B1(n_999), .B2(n_1000), .C(n_1001), .Y(n_359) );
INVx1_ASAP7_75t_L g1000 ( .A(n_360), .Y(n_1000) );
XNOR2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_563), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_449), .B1(n_561), .B2(n_562), .Y(n_362) );
INVx1_ASAP7_75t_L g561 ( .A(n_363), .Y(n_561) );
INVx1_ASAP7_75t_SL g448 ( .A(n_365), .Y(n_448) );
NAND4xp75_ASAP7_75t_L g365 ( .A(n_366), .B(n_402), .C(n_421), .D(n_437), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_392), .Y(n_366) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g497 ( .A(n_369), .Y(n_497) );
INVx2_ASAP7_75t_L g516 ( .A(n_369), .Y(n_516) );
OAI221xp5_ASAP7_75t_SL g578 ( .A1(n_369), .A2(n_579), .B1(n_580), .B2(n_583), .C(n_584), .Y(n_578) );
INVx3_ASAP7_75t_L g645 ( .A(n_369), .Y(n_645) );
OAI22xp5_ASAP7_75t_SL g866 ( .A1(n_369), .A2(n_527), .B1(n_867), .B2(n_868), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g945 ( .A1(n_369), .A2(n_946), .B1(n_947), .B2(n_948), .Y(n_945) );
INVx6_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx3_ASAP7_75t_L g558 ( .A(n_370), .Y(n_558) );
BUFx3_ASAP7_75t_L g793 ( .A(n_370), .Y(n_793) );
AND2x4_ASAP7_75t_L g370 ( .A(n_371), .B(n_380), .Y(n_370) );
AND2x2_ASAP7_75t_L g406 ( .A(n_371), .B(n_390), .Y(n_406) );
AND2x6_ASAP7_75t_L g409 ( .A(n_371), .B(n_410), .Y(n_409) );
AND2x6_ASAP7_75t_L g439 ( .A(n_371), .B(n_436), .Y(n_439) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_377), .Y(n_371) );
AND2x2_ASAP7_75t_L g417 ( .A(n_372), .B(n_378), .Y(n_417) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g388 ( .A(n_373), .B(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_373), .B(n_378), .Y(n_401) );
AND2x2_ASAP7_75t_L g433 ( .A(n_373), .B(n_383), .Y(n_433) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g379 ( .A(n_376), .Y(n_379) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g389 ( .A(n_378), .Y(n_389) );
INVx1_ASAP7_75t_L g443 ( .A(n_378), .Y(n_443) );
AND2x2_ASAP7_75t_L g396 ( .A(n_380), .B(n_388), .Y(n_396) );
AND2x6_ASAP7_75t_L g428 ( .A(n_380), .B(n_417), .Y(n_428) );
NAND2x1p5_ASAP7_75t_L g463 ( .A(n_380), .B(n_417), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g874 ( .A(n_380), .B(n_388), .Y(n_874) );
AND2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
INVx2_ASAP7_75t_L g391 ( .A(n_381), .Y(n_391) );
INVx1_ASAP7_75t_L g400 ( .A(n_381), .Y(n_400) );
OR2x2_ASAP7_75t_L g411 ( .A(n_381), .B(n_382), .Y(n_411) );
AND2x2_ASAP7_75t_L g436 ( .A(n_381), .B(n_383), .Y(n_436) );
AND2x2_ASAP7_75t_L g390 ( .A(n_382), .B(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx3_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx3_ASAP7_75t_L g501 ( .A(n_387), .Y(n_501) );
BUFx3_ASAP7_75t_L g512 ( .A(n_387), .Y(n_512) );
BUFx3_ASAP7_75t_L g638 ( .A(n_387), .Y(n_638) );
AND2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_388), .B(n_390), .Y(n_582) );
INVx1_ASAP7_75t_L g435 ( .A(n_389), .Y(n_435) );
AND2x4_ASAP7_75t_L g416 ( .A(n_390), .B(n_417), .Y(n_416) );
AND2x4_ASAP7_75t_L g419 ( .A(n_390), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g442 ( .A(n_391), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g478 ( .A(n_391), .Y(n_478) );
BUFx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g900 ( .A(n_394), .Y(n_900) );
INVx4_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx5_ASAP7_75t_L g493 ( .A(n_395), .Y(n_493) );
INVx2_ASAP7_75t_L g530 ( .A(n_395), .Y(n_530) );
INVx1_ASAP7_75t_L g553 ( .A(n_395), .Y(n_553) );
BUFx3_ASAP7_75t_L g586 ( .A(n_395), .Y(n_586) );
INVx3_ASAP7_75t_L g709 ( .A(n_395), .Y(n_709) );
INVx8_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
BUFx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx4f_ASAP7_75t_SL g494 ( .A(n_398), .Y(n_494) );
BUFx2_ASAP7_75t_L g554 ( .A(n_398), .Y(n_554) );
BUFx2_ASAP7_75t_L g1053 ( .A(n_398), .Y(n_1053) );
INVx6_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_SL g587 ( .A(n_399), .Y(n_587) );
INVx1_ASAP7_75t_SL g711 ( .A(n_399), .Y(n_711) );
INVx1_ASAP7_75t_L g797 ( .A(n_399), .Y(n_797) );
OR2x6_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
INVx1_ASAP7_75t_L g432 ( .A(n_400), .Y(n_432) );
INVx1_ASAP7_75t_L g420 ( .A(n_401), .Y(n_420) );
AND2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_412), .Y(n_402) );
BUFx3_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
BUFx3_ASAP7_75t_L g488 ( .A(n_405), .Y(n_488) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_405), .Y(n_572) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g527 ( .A(n_406), .Y(n_527) );
BUFx2_ASAP7_75t_SL g804 ( .A(n_406), .Y(n_804) );
BUFx2_ASAP7_75t_SL g988 ( .A(n_406), .Y(n_988) );
INVx1_ASAP7_75t_L g574 ( .A(n_407), .Y(n_574) );
INVx2_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
INVx3_ASAP7_75t_L g515 ( .A(n_408), .Y(n_515) );
INVx4_ASAP7_75t_L g830 ( .A(n_408), .Y(n_830) );
INVx11_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx11_ASAP7_75t_L g644 ( .A(n_409), .Y(n_644) );
AND2x4_ASAP7_75t_L g426 ( .A(n_410), .B(n_417), .Y(n_426) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g459 ( .A(n_411), .B(n_460), .Y(n_459) );
INVx3_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx4_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g490 ( .A(n_416), .Y(n_490) );
BUFx3_ASAP7_75t_L g528 ( .A(n_416), .Y(n_528) );
BUFx3_ASAP7_75t_L g551 ( .A(n_416), .Y(n_551) );
BUFx3_ASAP7_75t_L g649 ( .A(n_416), .Y(n_649) );
INVx1_ASAP7_75t_L g460 ( .A(n_417), .Y(n_460) );
BUFx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx3_ASAP7_75t_L g502 ( .A(n_419), .Y(n_502) );
BUFx3_ASAP7_75t_L g513 ( .A(n_419), .Y(n_513) );
BUFx3_ASAP7_75t_L g577 ( .A(n_419), .Y(n_577) );
BUFx3_ASAP7_75t_L g641 ( .A(n_419), .Y(n_641) );
BUFx2_ASAP7_75t_SL g735 ( .A(n_419), .Y(n_735) );
INVx1_ASAP7_75t_L g872 ( .A(n_419), .Y(n_872) );
BUFx2_ASAP7_75t_SL g986 ( .A(n_419), .Y(n_986) );
AND2x2_ASAP7_75t_L g807 ( .A(n_420), .B(n_478), .Y(n_807) );
AND2x2_ASAP7_75t_SL g421 ( .A(n_422), .B(n_429), .Y(n_421) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx5_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g519 ( .A(n_425), .Y(n_519) );
INVx2_ASAP7_75t_L g547 ( .A(n_425), .Y(n_547) );
INVx2_ASAP7_75t_L g699 ( .A(n_425), .Y(n_699) );
INVx4_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx4f_ASAP7_75t_L g520 ( .A(n_428), .Y(n_520) );
INVx1_ASAP7_75t_SL g894 ( .A(n_428), .Y(n_894) );
BUFx2_ASAP7_75t_L g911 ( .A(n_428), .Y(n_911) );
BUFx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g522 ( .A(n_431), .Y(n_522) );
INVx1_ASAP7_75t_L g665 ( .A(n_431), .Y(n_665) );
BUFx3_ASAP7_75t_L g751 ( .A(n_431), .Y(n_751) );
AND2x4_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
AND2x4_ASAP7_75t_L g441 ( .A(n_433), .B(n_442), .Y(n_441) );
AND2x4_ASAP7_75t_L g446 ( .A(n_433), .B(n_447), .Y(n_446) );
NAND2x1p5_ASAP7_75t_L g477 ( .A(n_433), .B(n_478), .Y(n_477) );
BUFx3_ASAP7_75t_L g523 ( .A(n_434), .Y(n_523) );
BUFx6f_ASAP7_75t_L g668 ( .A(n_434), .Y(n_668) );
BUFx2_ASAP7_75t_SL g706 ( .A(n_434), .Y(n_706) );
BUFx2_ASAP7_75t_SL g748 ( .A(n_434), .Y(n_748) );
AND2x4_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVx1_ASAP7_75t_L g484 ( .A(n_435), .Y(n_484) );
INVx1_ASAP7_75t_L g483 ( .A(n_436), .Y(n_483) );
INVx3_ASAP7_75t_L g961 ( .A(n_438), .Y(n_961) );
BUFx3_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_439), .Y(n_469) );
INVx4_ASAP7_75t_L g533 ( .A(n_439), .Y(n_533) );
INVx2_ASAP7_75t_L g541 ( .A(n_439), .Y(n_541) );
INVx2_ASAP7_75t_L g812 ( .A(n_439), .Y(n_812) );
INVx2_ASAP7_75t_SL g860 ( .A(n_439), .Y(n_860) );
INVx1_ASAP7_75t_L g729 ( .A(n_440), .Y(n_729) );
BUFx4f_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_441), .Y(n_466) );
BUFx2_ASAP7_75t_L g596 ( .A(n_441), .Y(n_596) );
BUFx6f_ASAP7_75t_L g671 ( .A(n_441), .Y(n_671) );
BUFx6f_ASAP7_75t_L g702 ( .A(n_441), .Y(n_702) );
INVx1_ASAP7_75t_L g447 ( .A(n_443), .Y(n_447) );
BUFx4f_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g535 ( .A(n_445), .Y(n_535) );
BUFx12f_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_446), .Y(n_472) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_446), .Y(n_600) );
INVx3_ASAP7_75t_L g562 ( .A(n_449), .Y(n_562) );
BUFx3_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_452), .B1(n_505), .B2(n_506), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g504 ( .A(n_453), .Y(n_504) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_485), .Y(n_453) );
NOR3xp33_ASAP7_75t_L g454 ( .A(n_455), .B(n_464), .C(n_474), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_457), .B1(n_461), .B2(n_462), .Y(n_455) );
OAI221xp5_ASAP7_75t_L g658 ( .A1(n_457), .A2(n_659), .B1(n_660), .B2(n_662), .C(n_663), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g956 ( .A1(n_457), .A2(n_834), .B1(n_957), .B2(n_958), .Y(n_956) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_SL g591 ( .A(n_458), .Y(n_591) );
INVx2_ASAP7_75t_L g776 ( .A(n_458), .Y(n_776) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
BUFx6f_ASAP7_75t_L g617 ( .A(n_459), .Y(n_617) );
OAI21xp5_ASAP7_75t_L g852 ( .A1(n_459), .A2(n_853), .B(n_854), .Y(n_852) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_462), .A2(n_590), .B1(n_591), .B2(n_592), .Y(n_589) );
INVx2_ASAP7_75t_L g661 ( .A(n_462), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_462), .A2(n_591), .B1(n_722), .B2(n_723), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g855 ( .A1(n_462), .A2(n_477), .B1(n_856), .B2(n_857), .Y(n_855) );
OA211x2_ASAP7_75t_L g1024 ( .A1(n_462), .A2(n_1025), .B(n_1026), .C(n_1027), .Y(n_1024) );
BUFx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g620 ( .A(n_463), .Y(n_620) );
OAI222xp33_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_467), .B1(n_468), .B2(n_470), .C1(n_471), .C2(n_473), .Y(n_464) );
INVx3_ASAP7_75t_L g624 ( .A(n_465), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g858 ( .A1(n_465), .A2(n_859), .B1(n_860), .B2(n_861), .Y(n_858) );
INVx4_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g842 ( .A(n_466), .Y(n_842) );
BUFx2_ASAP7_75t_L g889 ( .A(n_466), .Y(n_889) );
OAI221xp5_ASAP7_75t_SL g593 ( .A1(n_468), .A2(n_594), .B1(n_595), .B2(n_597), .C(n_598), .Y(n_593) );
OAI221xp5_ASAP7_75t_L g621 ( .A1(n_468), .A2(n_622), .B1(n_623), .B2(n_625), .C(n_626), .Y(n_621) );
OAI21xp33_ASAP7_75t_L g724 ( .A1(n_468), .A2(n_725), .B(n_726), .Y(n_724) );
INVx2_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g886 ( .A(n_469), .Y(n_886) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx3_ASAP7_75t_L g627 ( .A(n_472), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B1(n_479), .B2(n_480), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_476), .A2(n_728), .B1(n_729), .B2(n_730), .Y(n_727) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx4_ASAP7_75t_L g604 ( .A(n_477), .Y(n_604) );
BUFx3_ASAP7_75t_L g785 ( .A(n_477), .Y(n_785) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_480), .A2(n_602), .B1(n_603), .B2(n_605), .Y(n_601) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
CKINVDCx16_ASAP7_75t_R g481 ( .A(n_482), .Y(n_481) );
BUFx2_ASAP7_75t_L g632 ( .A(n_482), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g963 ( .A1(n_482), .A2(n_603), .B1(n_964), .B2(n_965), .Y(n_963) );
OR2x6_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_486), .B(n_495), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_487), .B(n_491), .Y(n_486) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
OAI21xp5_ASAP7_75t_SL g863 ( .A1(n_490), .A2(n_864), .B(n_865), .Y(n_863) );
INVx2_ASAP7_75t_L g897 ( .A(n_490), .Y(n_897) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
BUFx2_ASAP7_75t_L g680 ( .A(n_493), .Y(n_680) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_496), .B(n_498), .Y(n_495) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx2_ASAP7_75t_L g687 ( .A(n_502), .Y(n_687) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AO22x2_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B1(n_537), .B2(n_560), .Y(n_506) );
INVx2_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
XOR2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_536), .Y(n_508) );
NAND4xp75_ASAP7_75t_L g509 ( .A(n_510), .B(n_517), .C(n_524), .D(n_531), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_514), .Y(n_510) );
INVx1_ASAP7_75t_L g947 ( .A(n_515), .Y(n_947) );
AND2x2_ASAP7_75t_SL g517 ( .A(n_518), .B(n_521), .Y(n_517) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_529), .Y(n_524) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx3_ASAP7_75t_L g827 ( .A(n_527), .Y(n_827) );
INVx4_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
BUFx2_ASAP7_75t_L g779 ( .A(n_533), .Y(n_779) );
OAI22xp5_ASAP7_75t_SL g840 ( .A1(n_533), .A2(n_841), .B1(n_842), .B2(n_843), .Y(n_840) );
OAI21xp5_ASAP7_75t_SL g1043 ( .A1(n_533), .A2(n_1044), .B(n_1045), .Y(n_1043) );
INVx1_ASAP7_75t_L g940 ( .A(n_534), .Y(n_940) );
INVx3_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx4_ASAP7_75t_SL g560 ( .A(n_537), .Y(n_560) );
OA22x2_ASAP7_75t_L g611 ( .A1(n_537), .A2(n_560), .B1(n_612), .B2(n_653), .Y(n_611) );
XOR2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_559), .Y(n_537) );
NAND3x1_ASAP7_75t_L g538 ( .A(n_539), .B(n_549), .C(n_555), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_540), .B(n_544), .Y(n_539) );
OAI21xp5_ASAP7_75t_SL g540 ( .A1(n_541), .A2(n_542), .B(n_543), .Y(n_540) );
OAI222xp33_ASAP7_75t_L g669 ( .A1(n_541), .A2(n_670), .B1(n_672), .B2(n_673), .C1(n_674), .C2(n_675), .Y(n_669) );
OAI21xp5_ASAP7_75t_L g703 ( .A1(n_541), .A2(n_704), .B(n_705), .Y(n_703) );
OAI21xp5_ASAP7_75t_L g745 ( .A1(n_541), .A2(n_746), .B(n_747), .Y(n_745) );
OAI21xp5_ASAP7_75t_SL g914 ( .A1(n_541), .A2(n_915), .B(n_916), .Y(n_914) );
OAI21xp5_ASAP7_75t_SL g976 ( .A1(n_541), .A2(n_977), .B(n_978), .Y(n_976) );
NAND3xp33_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .C(n_548), .Y(n_544) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
AOI22xp5_ASAP7_75t_SL g563 ( .A1(n_564), .A2(n_690), .B1(n_691), .B2(n_762), .Y(n_563) );
INVx1_ASAP7_75t_L g762 ( .A(n_564), .Y(n_762) );
XOR2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_608), .Y(n_564) );
BUFx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g607 ( .A(n_568), .Y(n_607) );
AND2x2_ASAP7_75t_SL g568 ( .A(n_569), .B(n_588), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_578), .Y(n_569) );
OAI221xp5_ASAP7_75t_SL g570 ( .A1(n_571), .A2(n_573), .B1(n_574), .B2(n_575), .C(n_576), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g949 ( .A1(n_571), .A2(n_580), .B1(n_950), .B2(n_951), .Y(n_949) );
INVx1_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g875 ( .A(n_582), .B(n_876), .Y(n_875) );
INVx3_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NOR3xp33_ASAP7_75t_L g588 ( .A(n_589), .B(n_593), .C(n_601), .Y(n_588) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
BUFx4f_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx3_ASAP7_75t_SL g630 ( .A(n_604), .Y(n_630) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OAI22xp5_ASAP7_75t_SL g609 ( .A1(n_610), .A2(n_611), .B1(n_654), .B2(n_655), .Y(n_609) );
INVx2_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g653 ( .A(n_612), .Y(n_653) );
INVx2_ASAP7_75t_SL g651 ( .A(n_613), .Y(n_651) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_633), .Y(n_613) );
NOR3xp33_ASAP7_75t_L g614 ( .A(n_615), .B(n_621), .C(n_628), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_617), .B1(n_618), .B2(n_619), .Y(n_615) );
OAI21xp5_ASAP7_75t_SL g837 ( .A1(n_617), .A2(n_838), .B(n_839), .Y(n_837) );
INVx1_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g834 ( .A(n_620), .Y(n_834) );
OAI221xp5_ASAP7_75t_L g778 ( .A1(n_623), .A2(n_779), .B1(n_780), .B2(n_781), .C(n_782), .Y(n_778) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g674 ( .A(n_627), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_630), .B1(n_631), .B2(n_632), .Y(n_628) );
OAI22xp5_ASAP7_75t_SL g833 ( .A1(n_630), .A2(n_834), .B1(n_835), .B2(n_836), .Y(n_833) );
OAI22xp5_ASAP7_75t_L g783 ( .A1(n_632), .A2(n_784), .B1(n_785), .B2(n_786), .Y(n_783) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_634), .B(n_646), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_642), .Y(n_634) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
BUFx4f_ASAP7_75t_SL g734 ( .A(n_638), .Y(n_734) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_SL g685 ( .A(n_644), .Y(n_685) );
INVx5_ASAP7_75t_SL g713 ( .A(n_644), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g877 ( .A(n_644), .B(n_878), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_650), .Y(n_646) );
BUFx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g689 ( .A(n_656), .Y(n_689) );
AND2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_676), .Y(n_656) );
NOR2xp33_ASAP7_75t_SL g657 ( .A(n_658), .B(n_669), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g774 ( .A1(n_660), .A2(n_775), .B1(n_776), .B2(n_777), .Y(n_774) );
OAI211xp5_ASAP7_75t_L g932 ( .A1(n_660), .A2(n_933), .B(n_934), .C(n_935), .Y(n_932) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g670 ( .A(n_671), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_677), .B(n_681), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g681 ( .A(n_682), .B(n_686), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OA22x2_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_694), .B1(n_716), .B2(n_761), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
XOR2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_715), .Y(n_694) );
NAND4xp75_ASAP7_75t_SL g695 ( .A(n_696), .B(n_707), .C(n_712), .D(n_714), .Y(n_695) );
NOR2xp67_ASAP7_75t_SL g696 ( .A(n_697), .B(n_703), .Y(n_696) );
NAND3xp33_ASAP7_75t_L g697 ( .A(n_698), .B(n_700), .C(n_701), .Y(n_697) );
INVx1_ASAP7_75t_L g938 ( .A(n_702), .Y(n_938) );
BUFx6f_ASAP7_75t_L g979 ( .A(n_702), .Y(n_979) );
AND2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_710), .Y(n_707) );
INVx1_ASAP7_75t_L g761 ( .A(n_716), .Y(n_761) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .B1(n_741), .B2(n_742), .Y(n_716) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
XNOR2x1_ASAP7_75t_L g718 ( .A(n_719), .B(n_740), .Y(n_718) );
AND2x2_ASAP7_75t_L g719 ( .A(n_720), .B(n_731), .Y(n_719) );
NOR3xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_724), .C(n_727), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_732), .B(n_737), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_733), .B(n_736), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
INVx3_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
XOR2x2_ASAP7_75t_L g742 ( .A(n_743), .B(n_760), .Y(n_742) );
NAND2xp5_ASAP7_75t_SL g743 ( .A(n_744), .B(n_753), .Y(n_743) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_745), .B(n_749), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_752), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_754), .B(n_757), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
INVx1_ASAP7_75t_L g999 ( .A(n_763), .Y(n_999) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_765), .B1(n_844), .B2(n_998), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
OAI22xp5_ASAP7_75t_SL g765 ( .A1(n_766), .A2(n_767), .B1(n_819), .B2(n_820), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
HB1xp67_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_799), .B1(n_800), .B2(n_818), .Y(n_769) );
INVx1_ASAP7_75t_L g818 ( .A(n_770), .Y(n_818) );
INVx1_ASAP7_75t_L g798 ( .A(n_772), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_773), .B(n_787), .Y(n_772) );
NOR3xp33_ASAP7_75t_L g773 ( .A(n_774), .B(n_778), .C(n_783), .Y(n_773) );
NOR2xp67_ASAP7_75t_L g787 ( .A(n_788), .B(n_794), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_789), .B(n_790), .Y(n_788) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_795), .B(n_796), .Y(n_794) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
XOR2x2_ASAP7_75t_L g880 ( .A(n_800), .B(n_881), .Y(n_880) );
XOR2x2_ASAP7_75t_L g800 ( .A(n_801), .B(n_817), .Y(n_800) );
NAND4xp75_ASAP7_75t_SL g801 ( .A(n_802), .B(n_803), .C(n_805), .D(n_809), .Y(n_801) );
AND2x2_ASAP7_75t_L g805 ( .A(n_806), .B(n_808), .Y(n_805) );
NOR2xp33_ASAP7_75t_L g809 ( .A(n_810), .B(n_814), .Y(n_809) );
OAI21xp5_ASAP7_75t_L g810 ( .A1(n_811), .A2(n_812), .B(n_813), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .Y(n_814) );
INVx1_ASAP7_75t_SL g819 ( .A(n_820), .Y(n_819) );
HB1xp67_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
XNOR2xp5_ASAP7_75t_L g821 ( .A(n_822), .B(n_823), .Y(n_821) );
NAND3x1_ASAP7_75t_SL g823 ( .A(n_824), .B(n_828), .C(n_832), .Y(n_823) );
AND2x2_ASAP7_75t_L g824 ( .A(n_825), .B(n_826), .Y(n_824) );
AND2x2_ASAP7_75t_L g828 ( .A(n_829), .B(n_831), .Y(n_828) );
NOR3xp33_ASAP7_75t_L g832 ( .A(n_833), .B(n_837), .C(n_840), .Y(n_832) );
INVx1_ASAP7_75t_L g998 ( .A(n_844), .Y(n_998) );
AOI22xp5_ASAP7_75t_L g844 ( .A1(n_845), .A2(n_904), .B1(n_996), .B2(n_997), .Y(n_844) );
INVx1_ASAP7_75t_SL g996 ( .A(n_845), .Y(n_996) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
XNOR2xp5_ASAP7_75t_L g847 ( .A(n_848), .B(n_880), .Y(n_847) );
BUFx2_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
XNOR2x1_ASAP7_75t_L g849 ( .A(n_850), .B(n_879), .Y(n_849) );
AND3x2_ASAP7_75t_L g850 ( .A(n_851), .B(n_862), .C(n_869), .Y(n_850) );
NOR3xp33_ASAP7_75t_L g851 ( .A(n_852), .B(n_855), .C(n_858), .Y(n_851) );
NOR2xp33_ASAP7_75t_L g862 ( .A(n_863), .B(n_866), .Y(n_862) );
NOR3xp33_ASAP7_75t_L g869 ( .A(n_870), .B(n_875), .C(n_877), .Y(n_869) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_872), .B1(n_873), .B2(n_874), .Y(n_870) );
XNOR2xp5_ASAP7_75t_L g881 ( .A(n_882), .B(n_883), .Y(n_881) );
NAND3xp33_ASAP7_75t_L g883 ( .A(n_884), .B(n_895), .C(n_901), .Y(n_883) );
NOR2xp33_ASAP7_75t_L g884 ( .A(n_885), .B(n_890), .Y(n_884) );
OAI21xp5_ASAP7_75t_SL g885 ( .A1(n_886), .A2(n_887), .B(n_888), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_891), .B(n_892), .Y(n_890) );
INVx1_ASAP7_75t_SL g893 ( .A(n_894), .Y(n_893) );
AND2x2_ASAP7_75t_L g895 ( .A(n_896), .B(n_898), .Y(n_895) );
INVx3_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
AND2x2_ASAP7_75t_L g901 ( .A(n_902), .B(n_903), .Y(n_901) );
INVx1_ASAP7_75t_L g997 ( .A(n_904), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_905), .A2(n_906), .B1(n_925), .B2(n_995), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
XOR2x2_ASAP7_75t_SL g906 ( .A(n_907), .B(n_924), .Y(n_906) );
NAND2x1p5_ASAP7_75t_L g907 ( .A(n_908), .B(n_917), .Y(n_907) );
NOR2xp33_ASAP7_75t_L g908 ( .A(n_909), .B(n_914), .Y(n_908) );
NAND3xp33_ASAP7_75t_L g909 ( .A(n_910), .B(n_912), .C(n_913), .Y(n_909) );
NOR2x1_ASAP7_75t_L g917 ( .A(n_918), .B(n_921), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_919), .B(n_920), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_922), .B(n_923), .Y(n_921) );
INVx2_ASAP7_75t_SL g995 ( .A(n_925), .Y(n_995) );
AOI22xp5_ASAP7_75t_L g925 ( .A1(n_926), .A2(n_927), .B1(n_952), .B2(n_994), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
INVx2_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
XNOR2xp5_ASAP7_75t_L g928 ( .A(n_929), .B(n_930), .Y(n_928) );
AND2x2_ASAP7_75t_L g930 ( .A(n_931), .B(n_941), .Y(n_930) );
OAI22xp5_ASAP7_75t_L g936 ( .A1(n_937), .A2(n_938), .B1(n_939), .B2(n_940), .Y(n_936) );
NOR3xp33_ASAP7_75t_L g941 ( .A(n_942), .B(n_945), .C(n_949), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_943), .B(n_944), .Y(n_942) );
INVx2_ASAP7_75t_L g994 ( .A(n_952), .Y(n_994) );
XNOR2x2_ASAP7_75t_L g952 ( .A(n_953), .B(n_973), .Y(n_952) );
INVx1_ASAP7_75t_SL g971 ( .A(n_954), .Y(n_971) );
AND2x2_ASAP7_75t_SL g954 ( .A(n_955), .B(n_966), .Y(n_954) );
NOR3xp33_ASAP7_75t_L g955 ( .A(n_956), .B(n_959), .C(n_963), .Y(n_955) );
OAI21xp33_ASAP7_75t_L g959 ( .A1(n_960), .A2(n_961), .B(n_962), .Y(n_959) );
AND4x1_ASAP7_75t_L g966 ( .A(n_967), .B(n_968), .C(n_969), .D(n_970), .Y(n_966) );
INVx2_ASAP7_75t_SL g992 ( .A(n_974), .Y(n_992) );
AND2x2_ASAP7_75t_L g974 ( .A(n_975), .B(n_983), .Y(n_974) );
NOR2xp33_ASAP7_75t_L g975 ( .A(n_976), .B(n_980), .Y(n_975) );
NAND2xp5_ASAP7_75t_SL g980 ( .A(n_981), .B(n_982), .Y(n_980) );
NOR2xp33_ASAP7_75t_L g983 ( .A(n_984), .B(n_989), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_985), .B(n_987), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_990), .B(n_991), .Y(n_989) );
INVx1_ASAP7_75t_SL g1001 ( .A(n_1002), .Y(n_1001) );
NOR2x1_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1007), .Y(n_1002) );
OR2x2_ASAP7_75t_SL g1059 ( .A(n_1003), .B(n_1008), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1006), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
HB1xp67_ASAP7_75t_L g1030 ( .A(n_1005), .Y(n_1030) );
NAND2xp5_ASAP7_75t_L g1037 ( .A(n_1005), .B(n_1034), .Y(n_1037) );
CKINVDCx16_ASAP7_75t_R g1034 ( .A(n_1006), .Y(n_1034) );
CKINVDCx20_ASAP7_75t_R g1007 ( .A(n_1008), .Y(n_1007) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1010), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1013), .Y(n_1011) );
OAI322xp33_ASAP7_75t_L g1014 ( .A1(n_1015), .A2(n_1030), .A3(n_1031), .B1(n_1035), .B2(n_1038), .C1(n_1039), .C2(n_1057), .Y(n_1014) );
INVx1_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
NAND4xp75_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1021), .C(n_1024), .D(n_1028), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1020), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1021 ( .A(n_1022), .B(n_1023), .Y(n_1021) );
BUFx2_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
HB1xp67_ASAP7_75t_L g1032 ( .A(n_1033), .Y(n_1032) );
INVx1_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
CKINVDCx20_ASAP7_75t_R g1035 ( .A(n_1036), .Y(n_1035) );
XOR2x2_ASAP7_75t_L g1040 ( .A(n_1038), .B(n_1041), .Y(n_1040) );
HB1xp67_ASAP7_75t_L g1039 ( .A(n_1040), .Y(n_1039) );
NAND3x1_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1050), .C(n_1054), .Y(n_1041) );
NOR2x1_ASAP7_75t_L g1042 ( .A(n_1043), .B(n_1046), .Y(n_1042) );
NAND3xp33_ASAP7_75t_L g1046 ( .A(n_1047), .B(n_1048), .C(n_1049), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_1051), .B(n_1052), .Y(n_1050) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1056), .Y(n_1054) );
CKINVDCx20_ASAP7_75t_R g1057 ( .A(n_1058), .Y(n_1057) );
CKINVDCx20_ASAP7_75t_R g1058 ( .A(n_1059), .Y(n_1058) );
endmodule