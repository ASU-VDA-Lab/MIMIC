module fake_jpeg_11653_n_648 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_648);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_648;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_7),
.B(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_3),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_12),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_62),
.Y(n_159)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_63),
.Y(n_150)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_45),
.Y(n_64)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_64),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_65),
.B(n_88),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_66),
.Y(n_176)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_67),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_68),
.Y(n_140)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx11_ASAP7_75t_L g216 ( 
.A(n_69),
.Y(n_216)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx24_ASAP7_75t_L g162 ( 
.A(n_70),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_26),
.B(n_16),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_71),
.B(n_79),
.Y(n_172)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_72),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_73),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_27),
.B(n_16),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_74),
.B(n_81),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_75),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_76),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_77),
.Y(n_152)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_26),
.B(n_16),
.Y(n_79)
);

BUFx24_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

BUFx2_ASAP7_75t_SL g194 ( 
.A(n_80),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_53),
.B(n_0),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_83),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_84),
.Y(n_207)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_85),
.Y(n_165)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g209 ( 
.A(n_86),
.Y(n_209)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_87),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_53),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_89),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_0),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_90),
.B(n_46),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_91),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_92),
.Y(n_210)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_93),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_94),
.Y(n_180)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_23),
.Y(n_95)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_95),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_44),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_96),
.B(n_121),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_97),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_98),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_32),
.Y(n_99)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_99),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_32),
.Y(n_100)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_100),
.Y(n_160)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g154 ( 
.A(n_103),
.Y(n_154)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_104),
.Y(n_177)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_106),
.Y(n_166)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_23),
.Y(n_107)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_107),
.Y(n_198)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_23),
.Y(n_108)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_108),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_27),
.B(n_14),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_109),
.B(n_120),
.Y(n_182)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_30),
.Y(n_110)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_110),
.Y(n_175)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_25),
.Y(n_111)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_28),
.Y(n_112)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_112),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_28),
.Y(n_113)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_113),
.Y(n_196)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_25),
.Y(n_114)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_115),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_51),
.B(n_47),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_116),
.B(n_125),
.Y(n_191)
);

BUFx24_ASAP7_75t_L g117 ( 
.A(n_44),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_117),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g185 ( 
.A(n_118),
.Y(n_185)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_30),
.Y(n_119)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_119),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_38),
.B(n_2),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_25),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_52),
.Y(n_122)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_122),
.Y(n_192)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_34),
.Y(n_123)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_123),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_38),
.B(n_2),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_34),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_126),
.B(n_129),
.Y(n_179)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_56),
.Y(n_127)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_25),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_41),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_130),
.B(n_33),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_117),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_136),
.B(n_164),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_80),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_144),
.A2(n_188),
.B1(n_84),
.B2(n_98),
.Y(n_280)
);

HAxp5_ASAP7_75t_SL g145 ( 
.A(n_80),
.B(n_51),
.CON(n_145),
.SN(n_145)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_145),
.B(n_57),
.Y(n_220)
);

AND2x2_ASAP7_75t_SL g146 ( 
.A(n_117),
.B(n_33),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_146),
.B(n_171),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_61),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_151),
.B(n_183),
.Y(n_234)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_113),
.Y(n_163)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_163),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_90),
.Y(n_164)
);

INVx6_ASAP7_75t_SL g168 ( 
.A(n_64),
.Y(n_168)
);

CKINVDCx9p33_ASAP7_75t_R g269 ( 
.A(n_168),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_70),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_169),
.B(n_195),
.Y(n_268)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_87),
.Y(n_187)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_187),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_66),
.A2(n_31),
.B1(n_36),
.B2(n_22),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_127),
.Y(n_189)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_189),
.Y(n_257)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_68),
.Y(n_190)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_190),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_71),
.B(n_79),
.Y(n_195)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_75),
.Y(n_199)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

INVx6_ASAP7_75t_SL g202 ( 
.A(n_66),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_202),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_76),
.B(n_47),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_204),
.B(n_208),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_L g205 ( 
.A1(n_77),
.A2(n_31),
.B1(n_54),
.B2(n_36),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_205),
.A2(n_211),
.B1(n_214),
.B2(n_146),
.Y(n_224)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_82),
.Y(n_206)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_85),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_83),
.A2(n_36),
.B1(n_22),
.B2(n_54),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_93),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_212),
.B(n_102),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_91),
.A2(n_22),
.B1(n_54),
.B2(n_58),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_92),
.Y(n_215)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_215),
.Y(n_228)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_140),
.Y(n_217)
);

INVx6_ASAP7_75t_L g332 ( 
.A(n_217),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_162),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_218),
.B(n_241),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_220),
.B(n_255),
.Y(n_296)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_165),
.Y(n_222)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_222),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_181),
.B(n_124),
.C(n_122),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_223),
.B(n_248),
.C(n_283),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_224),
.A2(n_235),
.B1(n_261),
.B2(n_286),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_182),
.B(n_57),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_225),
.B(n_278),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_140),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_227),
.Y(n_320)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_148),
.Y(n_229)
);

INVx5_ASAP7_75t_L g295 ( 
.A(n_229),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_141),
.B(n_48),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_230),
.B(n_232),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_191),
.B(n_151),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_231),
.B(n_243),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_171),
.B(n_48),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_148),
.Y(n_233)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_233),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_205),
.A2(n_118),
.B1(n_115),
.B2(n_106),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_196),
.B(n_94),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_236),
.Y(n_342)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_137),
.Y(n_239)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_239),
.Y(n_322)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_173),
.Y(n_240)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_240),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_131),
.Y(n_241)
);

CKINVDCx12_ASAP7_75t_R g242 ( 
.A(n_162),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_242),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_172),
.B(n_59),
.Y(n_243)
);

CKINVDCx12_ASAP7_75t_R g244 ( 
.A(n_162),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_244),
.Y(n_349)
);

INVx6_ASAP7_75t_L g245 ( 
.A(n_152),
.Y(n_245)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_245),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_179),
.B(n_59),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_246),
.B(n_258),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_132),
.B(n_46),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_247),
.B(n_254),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_133),
.B(n_94),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_156),
.Y(n_249)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_249),
.Y(n_293)
);

BUFx24_ASAP7_75t_L g250 ( 
.A(n_134),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_250),
.Y(n_304)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_185),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_251),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_180),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_253),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_142),
.B(n_60),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_176),
.Y(n_255)
);

AND2x4_ASAP7_75t_L g256 ( 
.A(n_145),
.B(n_76),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_256),
.B(n_289),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_201),
.B(n_177),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_185),
.Y(n_259)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_259),
.Y(n_309)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_185),
.Y(n_260)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_260),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_211),
.A2(n_97),
.B1(n_100),
.B2(n_99),
.Y(n_261)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_154),
.Y(n_262)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_262),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_149),
.B(n_58),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_263),
.B(n_270),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_152),
.Y(n_264)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_264),
.Y(n_344)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_143),
.Y(n_266)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_266),
.Y(n_303)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_138),
.Y(n_267)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_267),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_135),
.B(n_35),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_159),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_271),
.B(n_272),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_139),
.B(n_60),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_150),
.B(n_35),
.Y(n_273)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_273),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_176),
.Y(n_274)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_274),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_194),
.Y(n_276)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_276),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_155),
.B(n_61),
.Y(n_277)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_277),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_175),
.B(n_50),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_193),
.Y(n_279)
);

AO21x1_ASAP7_75t_L g331 ( 
.A1(n_279),
.A2(n_280),
.B(n_282),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_175),
.A2(n_84),
.B1(n_50),
.B2(n_43),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_186),
.B(n_102),
.Y(n_283)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_284),
.Y(n_348)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_137),
.Y(n_285)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_285),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_167),
.A2(n_43),
.B1(n_42),
.B2(n_41),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_198),
.A2(n_42),
.B1(n_41),
.B2(n_5),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_287),
.A2(n_218),
.B1(n_250),
.B2(n_207),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_200),
.B(n_3),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_288),
.Y(n_297)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_147),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_186),
.B(n_3),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_290),
.B(n_291),
.Y(n_324)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_200),
.Y(n_291)
);

CKINVDCx12_ASAP7_75t_R g292 ( 
.A(n_193),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_292),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_269),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_301),
.B(n_335),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_221),
.B(n_158),
.C(n_188),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_302),
.B(n_323),
.C(n_347),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_225),
.B(n_221),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_308),
.B(n_325),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_256),
.A2(n_161),
.B1(n_213),
.B2(n_184),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_311),
.A2(n_316),
.B1(n_317),
.B2(n_319),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_256),
.A2(n_161),
.B1(n_213),
.B2(n_184),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_256),
.A2(n_192),
.B1(n_178),
.B2(n_197),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_221),
.A2(n_192),
.B1(n_178),
.B2(n_197),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_223),
.B(n_144),
.C(n_216),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_234),
.B(n_220),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_265),
.A2(n_216),
.B(n_159),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_329),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_269),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_250),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_338),
.B(n_341),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_339),
.B(n_207),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_236),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_267),
.B(n_166),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_343),
.B(n_217),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_237),
.B(n_210),
.C(n_203),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_236),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_352),
.B(n_268),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_353),
.B(n_371),
.Y(n_405)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_326),
.Y(n_354)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_354),
.Y(n_410)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_343),
.Y(n_355)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_355),
.Y(n_417)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_326),
.Y(n_356)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_356),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_312),
.A2(n_224),
.B1(n_261),
.B2(n_166),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g428 ( 
.A1(n_357),
.A2(n_390),
.B1(n_283),
.B2(n_245),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_359),
.B(n_363),
.Y(n_409)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_293),
.Y(n_360)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_360),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_298),
.B(n_281),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_294),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_364),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_298),
.B(n_257),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_365),
.B(n_373),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_366),
.B(n_367),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_327),
.B(n_252),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_321),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_368),
.B(n_384),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_328),
.B(n_238),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_369),
.B(n_377),
.Y(n_406)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_314),
.Y(n_371)
);

OA22x2_ASAP7_75t_L g372 ( 
.A1(n_317),
.A2(n_222),
.B1(n_240),
.B2(n_160),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_372),
.B(n_379),
.Y(n_411)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_293),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_308),
.B(n_324),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_374),
.B(n_381),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_336),
.B(n_266),
.Y(n_377)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_325),
.B(n_262),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_378),
.A2(n_389),
.B(n_396),
.Y(n_420)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_303),
.Y(n_379)
);

INVx13_ASAP7_75t_L g380 ( 
.A(n_299),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_380),
.Y(n_429)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_294),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_306),
.B(n_249),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_382),
.B(n_383),
.Y(n_436)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_350),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_350),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_305),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_385),
.B(n_394),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_324),
.B(n_275),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_386),
.B(n_388),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_302),
.A2(n_157),
.B1(n_153),
.B2(n_203),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_387),
.A2(n_393),
.B1(n_315),
.B2(n_304),
.Y(n_401)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_351),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_342),
.A2(n_291),
.B1(n_274),
.B2(n_253),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g390 ( 
.A1(n_342),
.A2(n_160),
.B1(n_248),
.B2(n_153),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_334),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_391),
.B(n_392),
.Y(n_408)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_322),
.Y(n_392)
);

OAI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_311),
.A2(n_233),
.B1(n_264),
.B2(n_227),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_337),
.B(n_239),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_344),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_395),
.B(n_304),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_331),
.A2(n_248),
.B(n_255),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_324),
.B(n_289),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_397),
.B(n_399),
.Y(n_431)
);

INVx13_ASAP7_75t_L g398 ( 
.A(n_346),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_398),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_310),
.B(n_228),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_401),
.A2(n_407),
.B1(n_414),
.B2(n_427),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_370),
.A2(n_355),
.B1(n_375),
.B2(n_374),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_402),
.B(n_412),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_376),
.A2(n_307),
.B1(n_323),
.B2(n_300),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_370),
.A2(n_331),
.B1(n_316),
.B2(n_300),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_375),
.B(n_307),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_413),
.B(n_419),
.C(n_435),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_376),
.A2(n_307),
.B1(n_296),
.B2(n_348),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_365),
.A2(n_359),
.B1(n_396),
.B2(n_358),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_418),
.B(n_437),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_358),
.B(n_296),
.C(n_347),
.Y(n_419)
);

BUFx24_ASAP7_75t_SL g421 ( 
.A(n_368),
.Y(n_421)
);

BUFx24_ASAP7_75t_SL g440 ( 
.A(n_421),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_378),
.A2(n_329),
.B(n_296),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_422),
.Y(n_456)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_425),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_387),
.A2(n_297),
.B1(n_332),
.B2(n_295),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_428),
.A2(n_430),
.B1(n_392),
.B2(n_354),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_353),
.A2(n_332),
.B1(n_295),
.B2(n_344),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_L g434 ( 
.A1(n_353),
.A2(n_385),
.B1(n_362),
.B2(n_372),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_434),
.Y(n_474)
);

MAJx2_ASAP7_75t_L g435 ( 
.A(n_378),
.B(n_318),
.C(n_283),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_363),
.A2(n_319),
.B1(n_157),
.B2(n_210),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_397),
.A2(n_229),
.B1(n_340),
.B2(n_320),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_438),
.B(n_395),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_404),
.B(n_361),
.Y(n_439)
);

NAND3xp33_ASAP7_75t_L g504 ( 
.A(n_439),
.B(n_441),
.C(n_450),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_404),
.B(n_382),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_420),
.A2(n_386),
.B(n_372),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_442),
.B(n_445),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_405),
.B(n_372),
.Y(n_443)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_443),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_402),
.B(n_391),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_444),
.B(n_448),
.C(n_449),
.Y(n_486)
);

AND2x6_ASAP7_75t_L g445 ( 
.A(n_407),
.B(n_380),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_413),
.B(n_379),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_419),
.B(n_388),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_416),
.B(n_349),
.Y(n_450)
);

INVx13_ASAP7_75t_L g452 ( 
.A(n_432),
.Y(n_452)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_452),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_406),
.B(n_330),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_453),
.B(n_462),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_454),
.A2(n_430),
.B1(n_426),
.B2(n_383),
.Y(n_508)
);

INVx5_ASAP7_75t_L g455 ( 
.A(n_432),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_455),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_409),
.B(n_380),
.Y(n_457)
);

NOR3xp33_ASAP7_75t_L g497 ( 
.A(n_457),
.B(n_398),
.C(n_423),
.Y(n_497)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_459),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_408),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_460),
.B(n_463),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_409),
.B(n_371),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_461),
.B(n_469),
.C(n_426),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_406),
.B(n_345),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_408),
.Y(n_463)
);

CKINVDCx12_ASAP7_75t_R g464 ( 
.A(n_429),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_464),
.B(n_471),
.Y(n_484)
);

CKINVDCx10_ASAP7_75t_R g465 ( 
.A(n_429),
.Y(n_465)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_465),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_415),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_467),
.B(n_470),
.Y(n_475)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_410),
.Y(n_468)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_468),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_435),
.B(n_418),
.C(n_433),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_424),
.B(n_384),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_414),
.B(n_345),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_431),
.B(n_322),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_472),
.B(n_403),
.Y(n_492)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_433),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_473),
.B(n_424),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_474),
.A2(n_427),
.B1(n_401),
.B2(n_417),
.Y(n_477)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_477),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_466),
.B(n_412),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_478),
.B(n_490),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_483),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_474),
.A2(n_417),
.B1(n_431),
.B2(n_420),
.Y(n_485)
);

CKINVDCx14_ASAP7_75t_R g509 ( 
.A(n_485),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_451),
.A2(n_411),
.B1(n_437),
.B2(n_405),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_487),
.A2(n_489),
.B1(n_502),
.B2(n_508),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_446),
.A2(n_436),
.B1(n_422),
.B2(n_400),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_488),
.A2(n_443),
.B1(n_454),
.B2(n_455),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_458),
.A2(n_411),
.B1(n_405),
.B2(n_436),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_466),
.B(n_400),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_449),
.B(n_435),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_491),
.B(n_456),
.C(n_460),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_492),
.B(n_494),
.Y(n_514)
);

A2O1A1O1Ixp25_ASAP7_75t_L g493 ( 
.A1(n_469),
.A2(n_411),
.B(n_346),
.C(n_349),
.D(n_398),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g532 ( 
.A1(n_493),
.A2(n_465),
.B(n_443),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_467),
.B(n_403),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_497),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_447),
.B(n_381),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_498),
.B(n_499),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_447),
.B(n_356),
.Y(n_499)
);

MAJx2_ASAP7_75t_L g500 ( 
.A(n_448),
.B(n_446),
.C(n_461),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_500),
.B(n_507),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_457),
.B(n_360),
.Y(n_501)
);

CKINVDCx16_ASAP7_75t_R g515 ( 
.A(n_501),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_458),
.A2(n_438),
.B1(n_423),
.B2(n_410),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_444),
.B(n_373),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g527 ( 
.A(n_503),
.Y(n_527)
);

XOR2x2_ASAP7_75t_L g511 ( 
.A(n_478),
.B(n_491),
.Y(n_511)
);

OAI21xp33_ASAP7_75t_L g560 ( 
.A1(n_511),
.A2(n_495),
.B(n_505),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_506),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_513),
.B(n_488),
.Y(n_543)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_506),
.Y(n_518)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_518),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_476),
.A2(n_481),
.B(n_456),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g558 ( 
.A1(n_520),
.A2(n_535),
.B(n_508),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_475),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_521),
.B(n_539),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_524),
.B(n_532),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_484),
.B(n_463),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g550 ( 
.A(n_525),
.B(n_533),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_490),
.B(n_473),
.C(n_442),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_526),
.B(n_536),
.C(n_537),
.Y(n_542)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_480),
.Y(n_528)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_528),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_487),
.A2(n_445),
.B1(n_459),
.B2(n_470),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_529),
.A2(n_538),
.B1(n_482),
.B2(n_496),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_530),
.A2(n_534),
.B1(n_532),
.B2(n_535),
.Y(n_551)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_480),
.Y(n_531)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_531),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_479),
.B(n_440),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_476),
.A2(n_468),
.B1(n_452),
.B2(n_333),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_481),
.A2(n_333),
.B(n_315),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_507),
.B(n_309),
.C(n_315),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_486),
.B(n_309),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_489),
.A2(n_320),
.B1(n_340),
.B2(n_313),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_504),
.Y(n_539)
);

XNOR2x1_ASAP7_75t_L g540 ( 
.A(n_526),
.B(n_486),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_540),
.B(n_560),
.Y(n_586)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_543),
.Y(n_567)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_518),
.Y(n_546)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_546),
.Y(n_574)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_528),
.Y(n_548)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_548),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_549),
.A2(n_154),
.B1(n_174),
.B2(n_170),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_551),
.A2(n_510),
.B1(n_529),
.B2(n_519),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_514),
.B(n_493),
.Y(n_552)
);

NAND3xp33_ASAP7_75t_L g578 ( 
.A(n_552),
.B(n_547),
.C(n_550),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_523),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_553),
.B(n_554),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_521),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_517),
.B(n_482),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_SL g571 ( 
.A1(n_556),
.A2(n_558),
.B(n_541),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_536),
.B(n_500),
.C(n_496),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_557),
.B(n_564),
.Y(n_577)
);

XNOR2x1_ASAP7_75t_SL g559 ( 
.A(n_524),
.B(n_502),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_559),
.B(n_530),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_539),
.A2(n_505),
.B1(n_313),
.B2(n_219),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_561),
.Y(n_579)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_531),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g581 ( 
.A1(n_562),
.A2(n_226),
.B1(n_251),
.B2(n_259),
.Y(n_581)
);

FAx1_ASAP7_75t_SL g563 ( 
.A(n_511),
.B(n_41),
.CI(n_285),
.CON(n_563),
.SN(n_563)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_563),
.B(n_515),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_512),
.A2(n_509),
.B1(n_517),
.B2(n_519),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_516),
.B(n_537),
.C(n_522),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_565),
.B(n_516),
.C(n_522),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_555),
.A2(n_520),
.B(n_534),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_566),
.A2(n_558),
.B(n_556),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_568),
.B(n_583),
.Y(n_592)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_569),
.Y(n_588)
);

XOR2xp5_ASAP7_75t_L g598 ( 
.A(n_570),
.B(n_549),
.Y(n_598)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_571),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_572),
.B(n_580),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_551),
.A2(n_510),
.B1(n_512),
.B2(n_538),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_573),
.Y(n_596)
);

BUFx12f_ASAP7_75t_SL g576 ( 
.A(n_555),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_SL g589 ( 
.A(n_576),
.B(n_557),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_578),
.B(n_563),
.Y(n_601)
);

AOI322xp5_ASAP7_75t_L g580 ( 
.A1(n_541),
.A2(n_527),
.A3(n_228),
.B1(n_226),
.B2(n_219),
.C1(n_260),
.C2(n_154),
.Y(n_580)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_581),
.Y(n_595)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_582),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_542),
.B(n_174),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_542),
.B(n_209),
.C(n_5),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_585),
.B(n_4),
.Y(n_597)
);

XOR2xp5_ASAP7_75t_L g617 ( 
.A(n_587),
.B(n_582),
.Y(n_617)
);

OR2x2_ASAP7_75t_L g614 ( 
.A(n_589),
.B(n_590),
.Y(n_614)
);

OAI21xp5_ASAP7_75t_SL g590 ( 
.A1(n_571),
.A2(n_547),
.B(n_546),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_577),
.B(n_565),
.C(n_540),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_594),
.B(n_597),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_598),
.A2(n_544),
.B1(n_563),
.B2(n_8),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_572),
.B(n_559),
.C(n_562),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_599),
.B(n_602),
.Y(n_607)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_601),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_584),
.B(n_548),
.Y(n_602)
);

XOR2xp5_ASAP7_75t_L g603 ( 
.A(n_568),
.B(n_586),
.Y(n_603)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_603),
.B(n_586),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_583),
.B(n_545),
.C(n_544),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_604),
.B(n_545),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_SL g605 ( 
.A(n_588),
.B(n_576),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_605),
.B(n_618),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_593),
.B(n_567),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_608),
.B(n_611),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_609),
.B(n_617),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_599),
.B(n_573),
.Y(n_611)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_612),
.Y(n_620)
);

MAJx2_ASAP7_75t_L g613 ( 
.A(n_591),
.B(n_590),
.C(n_594),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_613),
.B(n_603),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_596),
.A2(n_570),
.B1(n_574),
.B2(n_575),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_615),
.B(n_616),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_604),
.B(n_579),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_L g618 ( 
.A(n_587),
.B(n_585),
.Y(n_618)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_619),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_L g621 ( 
.A1(n_614),
.A2(n_600),
.B(n_595),
.Y(n_621)
);

AO21x1_ASAP7_75t_L g631 ( 
.A1(n_621),
.A2(n_625),
.B(n_610),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_622),
.B(n_618),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_607),
.B(n_598),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_614),
.A2(n_592),
.B(n_7),
.Y(n_626)
);

OAI21x1_ASAP7_75t_L g634 ( 
.A1(n_626),
.A2(n_613),
.B(n_9),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_606),
.B(n_592),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_SL g633 ( 
.A(n_630),
.B(n_609),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g638 ( 
.A(n_631),
.B(n_633),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_632),
.B(n_634),
.Y(n_641)
);

NAND2xp33_ASAP7_75t_L g635 ( 
.A(n_620),
.B(n_617),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_SL g639 ( 
.A1(n_635),
.A2(n_629),
.B(n_623),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_SL g636 ( 
.A(n_628),
.B(n_5),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_636),
.B(n_637),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_624),
.B(n_5),
.Y(n_637)
);

XOR2xp5_ASAP7_75t_L g643 ( 
.A(n_639),
.B(n_9),
.Y(n_643)
);

AOI322xp5_ASAP7_75t_L g642 ( 
.A1(n_638),
.A2(n_627),
.A3(n_625),
.B1(n_623),
.B2(n_12),
.C1(n_11),
.C2(n_10),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_642),
.Y(n_644)
);

XOR2xp5_ASAP7_75t_L g645 ( 
.A(n_644),
.B(n_641),
.Y(n_645)
);

OAI31xp33_ASAP7_75t_L g646 ( 
.A1(n_645),
.A2(n_643),
.A3(n_640),
.B(n_12),
.Y(n_646)
);

OAI321xp33_ASAP7_75t_L g647 ( 
.A1(n_646),
.A2(n_9),
.A3(n_11),
.B1(n_12),
.B2(n_641),
.C(n_547),
.Y(n_647)
);

BUFx24_ASAP7_75t_SL g648 ( 
.A(n_647),
.Y(n_648)
);


endmodule