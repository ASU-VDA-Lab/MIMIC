module real_jpeg_10237_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_4),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_4),
.A2(n_22),
.B(n_29),
.C(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_4),
.B(n_29),
.Y(n_36)
);

AOI21xp33_ASAP7_75t_L g194 ( 
.A1(n_4),
.A2(n_5),
.B(n_23),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_5),
.A2(n_23),
.B1(n_26),
.B2(n_31),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_5),
.A2(n_68),
.B(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_5),
.B(n_68),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_5),
.A2(n_31),
.B1(n_39),
.B2(n_40),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_5),
.B(n_99),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_5),
.B(n_142),
.Y(n_215)
);

O2A1O1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_5),
.A2(n_7),
.B(n_39),
.C(n_226),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_7),
.A2(n_39),
.B(n_42),
.C(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_7),
.B(n_39),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_8),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_41),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_8),
.A2(n_23),
.B1(n_26),
.B2(n_41),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_9),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_9),
.A2(n_10),
.B1(n_68),
.B2(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_9),
.A2(n_11),
.B1(n_34),
.B2(n_68),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_10),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_10),
.A2(n_39),
.B1(n_40),
.B2(n_104),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_10),
.A2(n_23),
.B1(n_26),
.B2(n_104),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_104),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_11),
.A2(n_34),
.B1(n_39),
.B2(n_40),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_11),
.A2(n_23),
.B1(n_26),
.B2(n_34),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_127),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_126),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_106),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_16),
.B(n_106),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_78),
.B2(n_105),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_51),
.B1(n_76),
.B2(n_77),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_19),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_37),
.B(n_50),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_20),
.B(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_32),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_21),
.B(n_218),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_27),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_22),
.B(n_33),
.Y(n_61)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_22),
.B(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_23),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_23),
.B(n_55),
.Y(n_54)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_25),
.A2(n_28),
.B(n_31),
.C(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_26),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_27),
.B(n_35),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_27),
.Y(n_138)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp33_ASAP7_75t_L g226 ( 
.A1(n_29),
.A2(n_31),
.B(n_43),
.Y(n_226)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_31),
.B(n_88),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_31),
.B(n_55),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_32),
.A2(n_60),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_32),
.B(n_197),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_35),
.B(n_198),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_42),
.B(n_44),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_39),
.A2(n_40),
.B1(n_67),
.B2(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_39),
.B(n_71),
.Y(n_162)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_40),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_42),
.B(n_49),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_42),
.A2(n_46),
.B(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_42),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_44),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_48),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_45),
.B(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_46),
.B(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_62),
.B1(n_74),
.B2(n_75),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_52),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_58),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_53),
.A2(n_58),
.B1(n_63),
.B2(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_53),
.A2(n_63),
.B1(n_225),
.B2(n_227),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_53),
.B(n_225),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B(n_57),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_54),
.B(n_85),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_54),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_54),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_55),
.A2(n_83),
.B(n_115),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_56),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_56),
.B(n_86),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_56),
.B(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_58),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_60),
.B(n_61),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_59),
.A2(n_88),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_61),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_61),
.B(n_218),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_62),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_70),
.B(n_72),
.Y(n_65)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_66),
.B(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_66),
.B(n_72),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B(n_69),
.C(n_70),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_68),
.Y(n_69)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_69),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_70),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_70),
.B(n_103),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_73),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_78),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_89),
.C(n_95),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_87),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_80),
.B(n_87),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_83),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_81),
.B(n_203),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_82),
.B(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_84),
.B(n_188),
.Y(n_187)
);

INVxp33_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_90),
.B1(n_95),
.B2(n_96),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_93),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_92),
.B(n_153),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_93),
.B(n_141),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_94),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_94),
.B(n_142),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_99),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_100),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.C(n_112),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_107),
.A2(n_108),
.B1(n_110),
.B2(n_273),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_110),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_112),
.B(n_272),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_119),
.C(n_122),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_113),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_117),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_116),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_116),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_118),
.B(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_119),
.A2(n_120),
.B1(n_122),
.B2(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_122),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_125),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_269),
.B(n_274),
.Y(n_127)
);

O2A1O1Ixp33_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_180),
.B(n_257),
.C(n_268),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_166),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_130),
.B(n_166),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_144),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_132),
.B(n_133),
.C(n_144),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.C(n_139),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_134),
.B(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_136),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_156),
.B1(n_157),
.B2(n_165),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_145),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_150),
.B2(n_155),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_146),
.B(n_155),
.C(n_156),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_150),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.C(n_172),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_167),
.A2(n_168),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_253)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.C(n_176),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_174),
.B(n_241),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_175),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_189),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_190),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_256),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_250),
.B(n_255),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_236),
.B(n_249),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_221),
.B(n_235),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_210),
.B(n_220),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_199),
.B(n_209),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_191),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_191),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_195),
.B2(n_196),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_193),
.B(n_195),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_204),
.B(n_208),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_202),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_212),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_219),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_217),
.C(n_219),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_223),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_228),
.B1(n_229),
.B2(n_234),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_224),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_225),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_230),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_233),
.C(n_234),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_237),
.B(n_238),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_243),
.B2(n_244),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_245),
.C(n_248),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_247),
.B2(n_248),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_245),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_246),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_251),
.B(n_252),
.Y(n_255)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_253),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_258),
.B(n_259),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_266),
.B2(n_267),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_263),
.C(n_267),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_266),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_270),
.B(n_271),
.Y(n_274)
);


endmodule