module real_jpeg_19777_n_12 (n_5, n_4, n_8, n_0, n_278, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_278;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_271;
wire n_47;
wire n_131;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_240;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_216;
wire n_179;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_274;
wire n_256;
wire n_101;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;
wire n_16;

INVx13_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_1),
.A2(n_3),
.B1(n_18),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_54),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_1),
.A2(n_39),
.B1(n_42),
.B2(n_54),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_1),
.A2(n_5),
.B1(n_54),
.B2(n_65),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_L g21 ( 
.A1(n_2),
.A2(n_18),
.B(n_22),
.C(n_25),
.Y(n_21)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_2),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_3),
.A2(n_8),
.B1(n_18),
.B2(n_19),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_3),
.A2(n_9),
.B1(n_18),
.B2(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_3),
.A2(n_7),
.B1(n_18),
.B2(n_50),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_3),
.A2(n_24),
.B(n_50),
.C(n_158),
.Y(n_157)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_4),
.Y(n_78)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_4),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_5),
.A2(n_10),
.B1(n_63),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_5),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_5),
.B(n_78),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_5),
.A2(n_9),
.B1(n_30),
.B2(n_65),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_5),
.A2(n_8),
.B1(n_19),
.B2(n_65),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_5),
.A2(n_7),
.B1(n_50),
.B2(n_65),
.Y(n_148)
);

AOI21xp33_ASAP7_75t_L g185 ( 
.A1(n_5),
.A2(n_7),
.B(n_10),
.Y(n_185)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_7),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_7),
.A2(n_39),
.B1(n_42),
.B2(n_50),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_50),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_SL g158 ( 
.A1(n_7),
.A2(n_23),
.B(n_27),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_7),
.B(n_28),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_SL g209 ( 
.A1(n_7),
.A2(n_40),
.B(n_42),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_8),
.A2(n_19),
.B1(n_26),
.B2(n_27),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_8),
.A2(n_19),
.B1(n_39),
.B2(n_42),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_9),
.A2(n_30),
.B1(n_39),
.B2(n_42),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_10),
.A2(n_39),
.B1(n_42),
.B2(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_10),
.Y(n_63)
);

INVx11_ASAP7_75t_SL g39 ( 
.A(n_11),
.Y(n_39)
);

AO21x1_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_271),
.B(n_274),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_67),
.B(n_270),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_31),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_15),
.B(n_31),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_15),
.B(n_272),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_15),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_20),
.B1(n_28),
.B2(n_29),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_17),
.A2(n_25),
.B(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_20),
.A2(n_28),
.B1(n_53),
.B2(n_55),
.Y(n_52)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_21),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_21),
.B(n_25),
.Y(n_81)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_26),
.A2(n_38),
.B(n_40),
.C(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_40),
.Y(n_45)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_27),
.A2(n_41),
.B(n_50),
.C(n_209),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_28),
.A2(n_48),
.B(n_53),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_29),
.B(n_81),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_32),
.B(n_268),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_32),
.B(n_268),
.Y(n_269)
);

FAx1_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_46),
.CI(n_51),
.CON(n_32),
.SN(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_34),
.A2(n_37),
.B1(n_43),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_36),
.B(n_93),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_43),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_37),
.A2(n_92),
.B(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_38),
.A2(n_44),
.B1(n_91),
.B2(n_93),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_38),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_38),
.B(n_50),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_38)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_42),
.A2(n_50),
.B(n_63),
.C(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_44),
.B(n_93),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_50),
.B(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_50),
.B(n_64),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_56),
.C(n_58),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_52),
.B(n_98),
.C(n_105),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_52),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_52),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_52),
.A2(n_90),
.B1(n_127),
.B2(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_52),
.B(n_154),
.C(n_155),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_52),
.A2(n_105),
.B1(n_127),
.B2(n_165),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_56),
.A2(n_58),
.B1(n_113),
.B2(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_56),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_57),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_58),
.A2(n_113),
.B1(n_114),
.B2(n_117),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_58),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_66),
.Y(n_58)
);

INVxp33_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_60),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_61),
.A2(n_64),
.B1(n_66),
.B2(n_85),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_61),
.A2(n_64),
.B1(n_88),
.B2(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_64),
.A2(n_85),
.B(n_86),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_65),
.B(n_189),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_267),
.B(n_269),
.Y(n_67)
);

OAI321xp33_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_122),
.A3(n_133),
.B1(n_265),
.B2(n_266),
.C(n_278),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_107),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_70),
.B(n_107),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_89),
.C(n_96),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_71),
.B(n_89),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_83),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_80),
.B2(n_82),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_73),
.A2(n_74),
.B1(n_84),
.B2(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_84),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_74),
.A2(n_80),
.B(n_83),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

INVxp33_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_76),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_77),
.A2(n_79),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_77),
.B(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_77),
.A2(n_78),
.B1(n_148),
.B2(n_160),
.Y(n_159)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_80),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_84),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_87),
.A2(n_142),
.B(n_143),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_88),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_94),
.B(n_95),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_94),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_90),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_90),
.B(n_170),
.C(n_172),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_90),
.A2(n_154),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_109),
.C(n_119),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_96),
.A2(n_97),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_98),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_99),
.A2(n_103),
.B1(n_201),
.B2(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_99),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_100),
.A2(n_101),
.B(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_102),
.A2(n_147),
.B(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_103),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_103),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_103),
.B(n_159),
.C(n_200),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_103),
.A2(n_201),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_103),
.B(n_219),
.C(n_224),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_110),
.C(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_105),
.A2(n_150),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_105),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_105),
.A2(n_140),
.B1(n_141),
.B2(n_165),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_105),
.B(n_141),
.C(n_207),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_107)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_118),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_110),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_110),
.A2(n_118),
.B1(n_126),
.B2(n_131),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_110),
.A2(n_118),
.B1(n_163),
.B2(n_166),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_110),
.A2(n_118),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_110),
.B(n_240),
.C(n_242),
.Y(n_257)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_117),
.C(n_118),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_114),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_118),
.B(n_131),
.C(n_132),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_123),
.B(n_124),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_132),
.Y(n_124)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_259),
.B(n_264),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_247),
.B(n_258),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_175),
.B(n_232),
.C(n_246),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_161),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_137),
.B(n_161),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_152),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_149),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_139),
.B(n_149),
.C(n_152),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_144),
.B2(n_145),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_140),
.A2(n_141),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_140),
.B(n_145),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_141),
.B(n_184),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_148),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_150),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_156),
.A2(n_157),
.B1(n_159),
.B2(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

NOR2x1_ASAP7_75t_R g191 ( 
.A(n_159),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_192),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_159),
.A2(n_168),
.B1(n_198),
.B2(n_202),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_160),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_167),
.C(n_169),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_162),
.B(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_163),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_167),
.B(n_169),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_182),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_231),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_226),
.B(n_230),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_216),
.B(n_225),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_204),
.B(n_215),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_195),
.B(n_203),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_186),
.B(n_194),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_191),
.B(n_193),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_197),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_198),
.Y(n_202)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_206),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_214),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_210),
.B1(n_211),
.B2(n_213),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_208),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_213),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_217),
.B(n_218),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_222),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_223),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_228),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_233),
.B(n_234),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_244),
.B2(n_245),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_239),
.C(n_245),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_244),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_248),
.B(n_249),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_257),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_255),
.C(n_257),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_261),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_276),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);


endmodule