module real_jpeg_11815_n_17 (n_5, n_4, n_8, n_0, n_12, n_324, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_324;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx10_ASAP7_75t_L g98 ( 
.A(n_0),
.Y(n_98)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_3),
.A2(n_40),
.B1(n_41),
.B2(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_3),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_110),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_3),
.A2(n_58),
.B1(n_62),
.B2(n_110),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_3),
.A2(n_27),
.B1(n_29),
.B2(n_110),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_4),
.A2(n_40),
.B1(n_41),
.B2(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_4),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_4),
.A2(n_58),
.B1(n_62),
.B2(n_143),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_143),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_4),
.A2(n_27),
.B1(n_29),
.B2(n_143),
.Y(n_253)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_7),
.A2(n_40),
.B1(n_41),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_7),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_7),
.A2(n_27),
.B1(n_29),
.B2(n_81),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_7),
.A2(n_58),
.B1(n_62),
.B2(n_81),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_81),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_8),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_39)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_8),
.A2(n_27),
.B1(n_29),
.B2(n_43),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_43),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_8),
.A2(n_43),
.B1(n_58),
.B2(n_62),
.Y(n_267)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_10),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_10),
.B(n_58),
.C(n_61),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_10),
.B(n_30),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_L g195 ( 
.A1(n_10),
.A2(n_134),
.B(n_179),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_L g205 ( 
.A1(n_10),
.A2(n_28),
.B(n_29),
.C(n_206),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_10),
.A2(n_27),
.B1(n_29),
.B2(n_163),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_10),
.B(n_51),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_10),
.B(n_40),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_11),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_11),
.A2(n_58),
.B1(n_62),
.B2(n_175),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_11),
.A2(n_27),
.B1(n_29),
.B2(n_175),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_11),
.A2(n_40),
.B1(n_41),
.B2(n_175),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_12),
.A2(n_40),
.B1(n_41),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_12),
.A2(n_27),
.B1(n_29),
.B2(n_50),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_50),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_12),
.A2(n_50),
.B1(n_58),
.B2(n_62),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_13),
.A2(n_27),
.B1(n_29),
.B2(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_13),
.A2(n_40),
.B1(n_41),
.B2(n_47),
.Y(n_48)
);

NAND2xp33_ASAP7_75t_SL g263 ( 
.A(n_13),
.B(n_27),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_14),
.A2(n_27),
.B1(n_29),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_14),
.A2(n_36),
.B1(n_58),
.B2(n_62),
.Y(n_100)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_16),
.A2(n_40),
.B1(n_41),
.B2(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_16),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_16),
.A2(n_27),
.B1(n_29),
.B2(n_73),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_16),
.A2(n_31),
.B1(n_32),
.B2(n_73),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_16),
.A2(n_58),
.B1(n_62),
.B2(n_73),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_88),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_87),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_74),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_21),
.B(n_74),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_54),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_37),
.B1(n_52),
.B2(n_53),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_23),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_34),
.Y(n_23)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_24),
.A2(n_30),
.B1(n_84),
.B2(n_86),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_24),
.B(n_213),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_25)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

AO22x1_ASAP7_75t_SL g30 ( 
.A1(n_26),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

OAI21xp33_ASAP7_75t_L g206 ( 
.A1(n_26),
.A2(n_31),
.B(n_163),
.Y(n_206)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

AOI32xp33_ASAP7_75t_L g262 ( 
.A1(n_29),
.A2(n_41),
.A3(n_47),
.B1(n_250),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_30),
.B(n_213),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_31),
.A2(n_32),
.B1(n_60),
.B2(n_61),
.Y(n_64)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_32),
.B(n_167),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_35),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_67)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_44),
.B1(n_49),
.B2(n_51),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_39),
.A2(n_45),
.B1(n_46),
.B2(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

O2A1O1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_41),
.A2(n_45),
.B(n_163),
.C(n_249),
.Y(n_248)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_44),
.B(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_45),
.A2(n_46),
.B1(n_72),
.B2(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_45),
.A2(n_142),
.B(n_144),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_45),
.A2(n_46),
.B1(n_142),
.B2(n_277),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_48),
.Y(n_45)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_46),
.A2(n_80),
.B(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_46),
.B(n_109),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_46),
.A2(n_107),
.B(n_277),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_67),
.C(n_71),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_67),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_55),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_SL g82 ( 
.A(n_55),
.B(n_79),
.C(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_55),
.A2(n_78),
.B1(n_83),
.B2(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_63),
.B(n_65),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_56),
.A2(n_63),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_56),
.A2(n_63),
.B1(n_103),
.B2(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_56),
.B(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_56),
.A2(n_63),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_56),
.A2(n_63),
.B1(n_138),
.B2(n_256),
.Y(n_282)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_57),
.A2(n_66),
.B1(n_105),
.B2(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_57),
.A2(n_174),
.B(n_176),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_57),
.B(n_163),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_57),
.A2(n_176),
.B(n_255),
.Y(n_254)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_57)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_62),
.B(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_62),
.B(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_63),
.B(n_165),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_68),
.A2(n_70),
.B1(n_85),
.B2(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_68),
.A2(n_70),
.B1(n_113),
.B2(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_68),
.A2(n_211),
.B(n_212),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_68),
.A2(n_70),
.B1(n_226),
.B2(n_253),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_68),
.A2(n_212),
.B(n_253),
.Y(n_275)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_70),
.A2(n_226),
.B(n_227),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_70),
.A2(n_140),
.B(n_227),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.C(n_82),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_75),
.A2(n_79),
.B1(n_119),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_75),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_79),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_79),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_82),
.B(n_148),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_83),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AO21x1_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_151),
.B(n_319),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_146),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_121),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_91),
.B(n_121),
.Y(n_320)
);

BUFx24_ASAP7_75t_SL g323 ( 
.A(n_91),
.Y(n_323)
);

FAx1_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_111),
.CI(n_116),
.CON(n_91),
.SN(n_91)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_92),
.B(n_111),
.C(n_116),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_96),
.B(n_106),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_93),
.A2(n_94),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_101),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_96),
.B1(n_106),
.B2(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_95),
.A2(n_96),
.B1(n_101),
.B2(n_102),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_98),
.B(n_99),
.Y(n_96)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_97),
.A2(n_98),
.B1(n_184),
.B2(n_186),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_97),
.B(n_180),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_97),
.A2(n_98),
.B1(n_133),
.B2(n_267),
.Y(n_281)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_98),
.B(n_180),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_100),
.A2(n_132),
.B1(n_134),
.B2(n_135),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_111),
.A2(n_112),
.B(n_114),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_115),
.A2(n_162),
.B(n_164),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_115),
.A2(n_164),
.B(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_127),
.C(n_128),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_122),
.A2(n_123),
.B1(n_127),
.B2(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_127),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_128),
.B(n_316),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_139),
.C(n_141),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_129),
.A2(n_130),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_136),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_131),
.A2(n_136),
.B1(n_137),
.B2(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_131),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_134),
.A2(n_178),
.B(n_179),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_134),
.A2(n_135),
.B1(n_208),
.B2(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_134),
.A2(n_135),
.B1(n_233),
.B2(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_135),
.A2(n_185),
.B(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_135),
.B(n_163),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_135),
.A2(n_193),
.B(n_208),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_139),
.B(n_141),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_145),
.B(n_248),
.Y(n_247)
);

OAI21xp33_ASAP7_75t_L g319 ( 
.A1(n_146),
.A2(n_320),
.B(n_321),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_150),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_147),
.B(n_150),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_313),
.B(n_318),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_301),
.B(n_312),
.Y(n_152)
);

OAI321xp33_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_269),
.A3(n_294),
.B1(n_299),
.B2(n_300),
.C(n_324),
.Y(n_153)
);

AOI21x1_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_242),
.B(n_268),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_220),
.B(n_241),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_201),
.B(n_219),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_181),
.B(n_200),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_168),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_159),
.B(n_168),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_166),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_160),
.A2(n_161),
.B1(n_166),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_166),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_177),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_173),
.C(n_177),
.Y(n_202)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_174),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_178),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_189),
.B(n_199),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_187),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_183),
.B(n_187),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_194),
.B(n_198),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_191),
.B(n_192),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_202),
.B(n_203),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_209),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_214),
.C(n_218),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_207),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_214),
.B1(n_217),
.B2(n_218),
.Y(n_209)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_210),
.Y(n_218)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_214),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_216),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_221),
.B(n_222),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_234),
.B2(n_235),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_237),
.C(n_239),
.Y(n_243)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_228),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_229),
.C(n_232),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_239),
.B2(n_240),
.Y(n_235)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_236),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_237),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_244),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_258),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_245),
.B(n_259),
.C(n_260),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_251),
.B2(n_257),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_246),
.B(n_252),
.C(n_254),
.Y(n_283)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_251),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_264),
.B2(n_265),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_265),
.Y(n_279)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_284),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_284),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_280),
.C(n_283),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_271),
.A2(n_272),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_279),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_276),
.B2(n_278),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_278),
.C(n_279),
.Y(n_293)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_276),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_280),
.B(n_283),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_282),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_293),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_288),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_286),
.B(n_288),
.C(n_293),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_292),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_291),
.C(n_292),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_295),
.B(n_296),
.Y(n_299)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_311),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_311),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_306),
.C(n_307),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_315),
.Y(n_318)
);


endmodule