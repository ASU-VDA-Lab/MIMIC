module fake_jpeg_2776_n_514 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_514);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_514;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_8),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_10),
.B(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_53),
.Y(n_153)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_55),
.B(n_56),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_1),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_57),
.B(n_58),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_23),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_60),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_24),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_61),
.B(n_62),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_21),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_65),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_66),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_30),
.B(n_1),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_83),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_34),
.Y(n_71)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_21),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_73),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_25),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_19),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_75),
.B(n_90),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_80),
.Y(n_137)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_82),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_30),
.B(n_1),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_85),
.Y(n_152)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_86),
.Y(n_148)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

BUFx4f_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

BUFx12_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_88),
.Y(n_154)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_19),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_31),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_91),
.A2(n_2),
.B1(n_5),
.B2(n_7),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_92),
.Y(n_147)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_93),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_18),
.B(n_2),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_95),
.Y(n_129)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_97),
.Y(n_139)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_20),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_98),
.B(n_5),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_66),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_99),
.B(n_124),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_57),
.A2(n_44),
.B1(n_42),
.B2(n_35),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_100),
.A2(n_138),
.B1(n_149),
.B2(n_158),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_55),
.A2(n_26),
.B1(n_45),
.B2(n_43),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_105),
.A2(n_130),
.B1(n_60),
.B2(n_81),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_56),
.B(n_42),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_108),
.B(n_132),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_68),
.A2(n_37),
.B1(n_29),
.B2(n_18),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_111),
.A2(n_141),
.B1(n_157),
.B2(n_96),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_75),
.A2(n_44),
.B1(n_35),
.B2(n_37),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_114),
.A2(n_116),
.B1(n_127),
.B2(n_134),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_58),
.A2(n_83),
.B1(n_79),
.B2(n_80),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_74),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_85),
.A2(n_29),
.B1(n_41),
.B2(n_45),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_71),
.A2(n_26),
.B1(n_45),
.B2(n_43),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_59),
.B(n_77),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_87),
.A2(n_41),
.B1(n_43),
.B2(n_20),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_67),
.A2(n_20),
.B1(n_28),
.B2(n_46),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_63),
.B(n_5),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_7),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_69),
.A2(n_20),
.B1(n_46),
.B2(n_27),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_151),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_70),
.B(n_7),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_L g157 ( 
.A1(n_91),
.A2(n_78),
.B1(n_76),
.B2(n_89),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_95),
.A2(n_20),
.B1(n_46),
.B2(n_27),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_109),
.B(n_93),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_159),
.B(n_164),
.Y(n_225)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_107),
.Y(n_160)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_160),
.Y(n_245)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_107),
.Y(n_162)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_162),
.Y(n_232)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_165),
.Y(n_220)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_101),
.Y(n_167)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_167),
.Y(n_239)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_101),
.Y(n_168)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_168),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_155),
.A2(n_65),
.B1(n_64),
.B2(n_54),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_169),
.A2(n_192),
.B1(n_203),
.B2(n_154),
.Y(n_235)
);

OAI21xp33_ASAP7_75t_SL g254 ( 
.A1(n_171),
.A2(n_173),
.B(n_201),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_106),
.A2(n_82),
.B1(n_84),
.B2(n_92),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_172),
.A2(n_175),
.B1(n_183),
.B2(n_202),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_147),
.Y(n_174)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_174),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_106),
.A2(n_97),
.B1(n_52),
.B2(n_51),
.Y(n_175)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_102),
.Y(n_176)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_176),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_53),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_178),
.B(n_179),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_132),
.B(n_53),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_128),
.B(n_7),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_180),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_129),
.B(n_8),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_181),
.Y(n_247)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_123),
.Y(n_182)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_182),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_100),
.A2(n_49),
.B1(n_86),
.B2(n_20),
.Y(n_183)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_184),
.Y(n_249)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_102),
.Y(n_185)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_185),
.Y(n_253)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_115),
.Y(n_186)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_186),
.Y(n_260)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_120),
.Y(n_187)
);

BUFx2_ASAP7_75t_SL g233 ( 
.A(n_187),
.Y(n_233)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_188),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_121),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_189),
.B(n_194),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_133),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_190),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_103),
.B(n_8),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_191),
.B(n_193),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_L g192 ( 
.A1(n_157),
.A2(n_88),
.B1(n_47),
.B2(n_50),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_110),
.B(n_9),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_108),
.B(n_9),
.Y(n_194)
);

INVx11_ASAP7_75t_L g195 ( 
.A(n_118),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_195),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_110),
.B(n_10),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_196),
.B(n_198),
.Y(n_252)
);

AND2x4_ASAP7_75t_L g197 ( 
.A(n_113),
.B(n_88),
.Y(n_197)
);

NAND2xp33_ASAP7_75t_SL g250 ( 
.A(n_197),
.B(n_212),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_122),
.B(n_11),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_133),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_199),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_113),
.B(n_11),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_206),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_119),
.A2(n_47),
.B1(n_13),
.B2(n_14),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_131),
.A2(n_47),
.B1(n_13),
.B2(n_14),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_141),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_125),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_204),
.B(n_205),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_139),
.B(n_15),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_140),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_115),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_207),
.B(n_211),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_119),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_208),
.A2(n_140),
.B(n_126),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_119),
.B(n_15),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_209),
.B(n_215),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_131),
.B(n_16),
.C(n_17),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_210),
.B(n_200),
.C(n_197),
.Y(n_255)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_136),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_153),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_156),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_214),
.Y(n_223)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_156),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_104),
.B(n_16),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_142),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_216),
.A2(n_126),
.B1(n_144),
.B2(n_142),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_175),
.A2(n_120),
.B(n_148),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_217),
.A2(n_227),
.B(n_236),
.Y(n_268)
);

A2O1A1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_163),
.A2(n_137),
.B(n_152),
.C(n_144),
.Y(n_218)
);

A2O1A1Ixp33_ASAP7_75t_L g287 ( 
.A1(n_218),
.A2(n_263),
.B(n_188),
.C(n_182),
.Y(n_287)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_224),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_179),
.A2(n_143),
.B(n_148),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_173),
.A2(n_152),
.B1(n_137),
.B2(n_147),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_228),
.A2(n_237),
.B1(n_246),
.B2(n_261),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_231),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_235),
.B(n_259),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_163),
.A2(n_104),
.B(n_117),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_178),
.A2(n_136),
.B1(n_117),
.B2(n_135),
.Y(n_237)
);

MAJx2_ASAP7_75t_L g243 ( 
.A(n_164),
.B(n_135),
.C(n_146),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_243),
.B(n_256),
.C(n_255),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_166),
.A2(n_112),
.B1(n_118),
.B2(n_143),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_244),
.A2(n_235),
.B1(n_217),
.B2(n_227),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_172),
.A2(n_112),
.B1(n_16),
.B2(n_17),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_161),
.A2(n_17),
.B(n_169),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_248),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_213),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_194),
.B(n_165),
.Y(n_256)
);

OAI32xp33_ASAP7_75t_L g259 ( 
.A1(n_177),
.A2(n_170),
.A3(n_205),
.B1(n_197),
.B2(n_209),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_166),
.A2(n_183),
.B1(n_210),
.B2(n_192),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_203),
.A2(n_206),
.B1(n_204),
.B2(n_189),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_262),
.A2(n_216),
.B1(n_207),
.B2(n_186),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_197),
.A2(n_187),
.B(n_162),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_167),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_270),
.B(n_277),
.Y(n_316)
);

NAND2xp33_ASAP7_75t_R g271 ( 
.A(n_219),
.B(n_174),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_271),
.A2(n_233),
.B(n_251),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_174),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_274),
.B(n_278),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_223),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_275),
.B(n_297),
.Y(n_334)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_245),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_276),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_219),
.B(n_168),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_220),
.Y(n_279)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_279),
.Y(n_318)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_220),
.Y(n_280)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_280),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_263),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_281),
.B(n_289),
.Y(n_351)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_229),
.Y(n_282)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_282),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_250),
.B(n_214),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_283),
.B(n_298),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_284),
.B(n_306),
.C(n_260),
.Y(n_315)
);

FAx1_ASAP7_75t_SL g285 ( 
.A(n_243),
.B(n_160),
.CI(n_195),
.CON(n_285),
.SN(n_285)
);

OAI32xp33_ASAP7_75t_L g335 ( 
.A1(n_285),
.A2(n_266),
.A3(n_253),
.B1(n_251),
.B2(n_231),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_261),
.A2(n_230),
.B1(n_254),
.B2(n_228),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_286),
.A2(n_294),
.B1(n_269),
.B2(n_278),
.Y(n_340)
);

A2O1A1Ixp33_ASAP7_75t_SL g322 ( 
.A1(n_287),
.A2(n_303),
.B(n_309),
.C(n_233),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_288),
.A2(n_290),
.B1(n_295),
.B2(n_302),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_223),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_259),
.A2(n_190),
.B1(n_199),
.B2(n_211),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_229),
.Y(n_291)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_291),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_225),
.B(n_176),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_292),
.B(n_293),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_258),
.B(n_236),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_230),
.A2(n_190),
.B1(n_199),
.B2(n_185),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_244),
.A2(n_248),
.B1(n_258),
.B2(n_257),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_247),
.B(n_212),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_296),
.B(n_300),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_240),
.B(n_184),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_264),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_299),
.B(n_304),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_221),
.B(n_264),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_239),
.Y(n_301)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_301),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_257),
.A2(n_243),
.B1(n_262),
.B2(n_240),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_225),
.B(n_234),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_237),
.B(n_218),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_234),
.B(n_252),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_305),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_252),
.B(n_265),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_260),
.Y(n_308)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_308),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_241),
.A2(n_265),
.B1(n_238),
.B2(n_249),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_238),
.B(n_232),
.Y(n_310)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_310),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_246),
.A2(n_226),
.B1(n_241),
.B2(n_266),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_311),
.A2(n_266),
.B1(n_222),
.B2(n_253),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_232),
.B(n_245),
.Y(n_312)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_312),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_284),
.B(n_249),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_313),
.B(n_324),
.C(n_330),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_315),
.B(n_280),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_322),
.A2(n_336),
.B(n_339),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_299),
.B(n_242),
.C(n_239),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_310),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_328),
.B(n_333),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_293),
.B(n_242),
.C(n_222),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_331),
.A2(n_343),
.B1(n_347),
.B2(n_301),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_306),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_332),
.B(n_337),
.C(n_338),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_312),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_335),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_270),
.B(n_273),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_273),
.B(n_298),
.C(n_277),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_340),
.A2(n_304),
.B1(n_311),
.B2(n_275),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_286),
.A2(n_290),
.B1(n_269),
.B2(n_288),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_308),
.Y(n_344)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_344),
.Y(n_358)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_279),
.Y(n_345)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_345),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_295),
.A2(n_273),
.B1(n_268),
.B2(n_304),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_283),
.B(n_268),
.C(n_274),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_348),
.B(n_317),
.C(n_313),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_287),
.A2(n_272),
.B(n_271),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_349),
.A2(n_350),
.B(n_303),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_274),
.A2(n_283),
.B(n_281),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_296),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_353),
.B(n_300),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_355),
.A2(n_357),
.B1(n_371),
.B2(n_372),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_334),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_356),
.B(n_359),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_343),
.A2(n_289),
.B1(n_307),
.B2(n_294),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_341),
.B(n_297),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_317),
.B(n_292),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_360),
.B(n_381),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_329),
.B(n_285),
.Y(n_363)
);

AO21x1_ASAP7_75t_L g396 ( 
.A1(n_363),
.A2(n_369),
.B(n_382),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_364),
.B(n_370),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_365),
.B(n_386),
.C(n_366),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_352),
.B(n_305),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_367),
.B(n_373),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_321),
.A2(n_285),
.B1(n_303),
.B2(n_267),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_368),
.A2(n_377),
.B1(n_384),
.B2(n_360),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_346),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_340),
.A2(n_321),
.B1(n_347),
.B2(n_351),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_338),
.A2(n_267),
.B1(n_282),
.B2(n_291),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_346),
.B(n_276),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_323),
.Y(n_374)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_374),
.Y(n_398)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_325),
.Y(n_376)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_376),
.Y(n_407)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_318),
.Y(n_378)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_378),
.Y(n_411)
);

AOI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_348),
.A2(n_339),
.B1(n_320),
.B2(n_342),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_379),
.A2(n_320),
.B(n_327),
.Y(n_395)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_319),
.Y(n_380)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_380),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_316),
.B(n_314),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_349),
.A2(n_331),
.B1(n_314),
.B2(n_329),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_383),
.A2(n_339),
.B1(n_336),
.B2(n_322),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_350),
.A2(n_316),
.B1(n_314),
.B2(n_335),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_315),
.B(n_332),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_385),
.B(n_386),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_337),
.B(n_324),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_387),
.A2(n_322),
.B(n_369),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_375),
.B(n_330),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_388),
.B(n_405),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_389),
.A2(n_397),
.B1(n_399),
.B2(n_400),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_390),
.A2(n_395),
.B(n_389),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_365),
.B(n_326),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_392),
.B(n_394),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_381),
.B(n_322),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_371),
.A2(n_320),
.B1(n_327),
.B2(n_355),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_354),
.A2(n_383),
.B1(n_357),
.B2(n_382),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_372),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_400),
.B(n_401),
.Y(n_418)
);

OA22x2_ASAP7_75t_L g401 ( 
.A1(n_354),
.A2(n_387),
.B1(n_384),
.B2(n_368),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_402),
.A2(n_406),
.B1(n_393),
.B2(n_399),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_404),
.B(n_410),
.C(n_415),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_359),
.B(n_361),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_366),
.A2(n_358),
.B1(n_380),
.B2(n_362),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_385),
.B(n_361),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_408),
.B(n_412),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_363),
.B(n_358),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_362),
.B(n_378),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_374),
.B(n_376),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_416),
.B(n_391),
.C(n_410),
.Y(n_428)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_415),
.Y(n_417)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_417),
.Y(n_446)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_416),
.Y(n_419)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_419),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_403),
.B(n_409),
.Y(n_421)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_421),
.Y(n_452)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_422),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_423),
.A2(n_441),
.B1(n_422),
.B2(n_438),
.Y(n_443)
);

BUFx24_ASAP7_75t_SL g424 ( 
.A(n_414),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_424),
.B(n_404),
.Y(n_442)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_398),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_425),
.B(n_430),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_428),
.B(n_426),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_429),
.A2(n_436),
.B(n_439),
.Y(n_454)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_407),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_406),
.B(n_408),
.Y(n_431)
);

NAND3xp33_ASAP7_75t_L g460 ( 
.A(n_431),
.B(n_435),
.C(n_437),
.Y(n_460)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_411),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_432),
.B(n_433),
.Y(n_453)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_413),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_392),
.B(n_402),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_390),
.A2(n_396),
.B(n_397),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_401),
.B(n_412),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_401),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_438),
.B(n_439),
.Y(n_457)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_401),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_391),
.B(n_396),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_440),
.B(n_420),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_394),
.A2(n_393),
.B1(n_397),
.B2(n_400),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_442),
.B(n_434),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_443),
.A2(n_456),
.B1(n_433),
.B2(n_434),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_444),
.B(n_445),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g447 ( 
.A(n_421),
.B(n_418),
.Y(n_447)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_447),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_429),
.A2(n_418),
.B(n_436),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_450),
.Y(n_471)
);

BUFx12_ASAP7_75t_L g451 ( 
.A(n_417),
.Y(n_451)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_451),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_454),
.B(n_450),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_426),
.B(n_428),
.C(n_420),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_455),
.B(n_444),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_423),
.A2(n_419),
.B1(n_441),
.B2(n_427),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_425),
.B(n_430),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_458),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_432),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_461),
.B(n_448),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_462),
.B(n_470),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_463),
.A2(n_472),
.B1(n_451),
.B2(n_461),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_457),
.B(n_446),
.Y(n_464)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_464),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_466),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_468),
.A2(n_453),
.B(n_451),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_459),
.A2(n_449),
.B1(n_457),
.B2(n_446),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_469),
.B(n_464),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_443),
.A2(n_459),
.B1(n_456),
.B2(n_447),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_452),
.B(n_460),
.Y(n_474)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_474),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_452),
.B(n_449),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_476),
.B(n_477),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_455),
.B(n_445),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_463),
.B(n_454),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_482),
.B(n_490),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_465),
.B(n_458),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_483),
.B(n_465),
.Y(n_494)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_484),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_469),
.A2(n_451),
.B(n_448),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_485),
.B(n_488),
.Y(n_497)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_486),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_467),
.B(n_453),
.C(n_473),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_471),
.A2(n_475),
.B(n_464),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_489),
.A2(n_466),
.B1(n_479),
.B2(n_478),
.Y(n_498)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_494),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_480),
.B(n_472),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_495),
.B(n_496),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_488),
.B(n_473),
.Y(n_496)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_498),
.Y(n_504)
);

FAx1_ASAP7_75t_SL g499 ( 
.A(n_489),
.B(n_482),
.CI(n_484),
.CON(n_499),
.SN(n_499)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_499),
.B(n_485),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_493),
.B(n_487),
.C(n_490),
.Y(n_501)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_501),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_493),
.B(n_486),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_502),
.Y(n_507)
);

A2O1A1Ixp33_ASAP7_75t_SL g508 ( 
.A1(n_505),
.A2(n_501),
.B(n_504),
.C(n_500),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_508),
.A2(n_497),
.B(n_481),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_506),
.B(n_503),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_509),
.B(n_510),
.Y(n_511)
);

OA21x2_ASAP7_75t_SL g512 ( 
.A1(n_511),
.A2(n_491),
.B(n_492),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_512),
.B(n_491),
.C(n_507),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_513),
.B(n_502),
.Y(n_514)
);


endmodule