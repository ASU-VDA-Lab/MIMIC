module fake_jpeg_18256_n_60 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_60);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_60;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_32;

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_26),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_39),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_10),
.B1(n_23),
.B2(n_20),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_36),
.B1(n_29),
.B2(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_27),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_4),
.Y(n_40)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_44),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_30),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_28),
.B(n_25),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_30),
.B1(n_28),
.B2(n_39),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_47),
.A2(n_50),
.B1(n_51),
.B2(n_43),
.Y(n_53)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_41),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_50),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_48),
.A2(n_38),
.B1(n_35),
.B2(n_7),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_55),
.B(n_52),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_13),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_16),
.B(n_19),
.Y(n_58)
);

AOI322xp5_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_11),
.A3(n_18),
.B1(n_8),
.B2(n_9),
.C1(n_24),
.C2(n_17),
.Y(n_59)
);

OAI211xp5_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_5),
.B(n_6),
.C(n_58),
.Y(n_60)
);


endmodule