module fake_jpeg_31329_n_413 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_413);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_413;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx4f_ASAP7_75t_SL g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_45),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_30),
.B(n_15),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_46),
.B(n_14),
.Y(n_124)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_24),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_48),
.B(n_66),
.Y(n_131)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_50),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_1),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_81),
.Y(n_99)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_53),
.B(n_59),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_43),
.B(n_2),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_56),
.B(n_34),
.C(n_31),
.Y(n_113)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_24),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_62),
.B(n_73),
.Y(n_125)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_63),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_24),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_16),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_71),
.Y(n_127)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_28),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_28),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_74),
.B(n_80),
.Y(n_126)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

BUFx16f_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

CKINVDCx6p67_ASAP7_75t_R g110 ( 
.A(n_76),
.Y(n_110)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_41),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

NAND2xp33_ASAP7_75t_SL g119 ( 
.A(n_83),
.B(n_84),
.Y(n_119)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_47),
.B(n_30),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_121),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_63),
.A2(n_41),
.B1(n_39),
.B2(n_29),
.Y(n_96)
);

AO21x1_ASAP7_75t_L g174 ( 
.A1(n_96),
.A2(n_97),
.B(n_102),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_75),
.A2(n_29),
.B1(n_33),
.B2(n_35),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_52),
.A2(n_40),
.B(n_37),
.C(n_35),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_101),
.B(n_124),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_69),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_65),
.A2(n_33),
.B1(n_18),
.B2(n_22),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_106),
.A2(n_130),
.B1(n_61),
.B2(n_60),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_50),
.A2(n_18),
.B1(n_20),
.B2(n_22),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_109),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_12),
.C(n_11),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g115 ( 
.A1(n_56),
.A2(n_31),
.B(n_27),
.Y(n_115)
);

OR2x4_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_19),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_70),
.A2(n_27),
.B1(n_26),
.B2(n_23),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_117),
.A2(n_122),
.B1(n_128),
.B2(n_45),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_56),
.A2(n_26),
.B1(n_23),
.B2(n_20),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_59),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_76),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_68),
.A2(n_19),
.B1(n_14),
.B2(n_13),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_72),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_L g130 ( 
.A1(n_55),
.A2(n_19),
.B1(n_4),
.B2(n_5),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_132),
.B(n_135),
.Y(n_200)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_85),
.Y(n_134)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

AND2x4_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_76),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_113),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_141),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_84),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_144),
.Y(n_180)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_138),
.Y(n_192)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_139),
.Y(n_206)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_140),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_99),
.B(n_81),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_101),
.A2(n_77),
.B1(n_71),
.B2(n_54),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_142),
.A2(n_123),
.B1(n_116),
.B2(n_112),
.Y(n_193)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_143),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_86),
.B(n_82),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_145),
.A2(n_148),
.B1(n_165),
.B2(n_167),
.Y(n_190)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_146),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_110),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_154),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_93),
.A2(n_79),
.B1(n_57),
.B2(n_51),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_149),
.A2(n_151),
.B(n_152),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_87),
.Y(n_150)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_150),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_114),
.A2(n_67),
.B1(n_64),
.B2(n_58),
.Y(n_152)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_87),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_131),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_155),
.B(n_177),
.C(n_165),
.Y(n_204)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_88),
.Y(n_156)
);

INVx13_ASAP7_75t_L g202 ( 
.A(n_156),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_157),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_95),
.Y(n_158)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_12),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_162),
.Y(n_188)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_89),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_109),
.B(n_12),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_166),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_95),
.Y(n_164)
);

INVx13_ASAP7_75t_L g212 ( 
.A(n_164),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_115),
.A2(n_11),
.B1(n_4),
.B2(n_5),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_88),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_93),
.A2(n_11),
.B1(n_5),
.B2(n_7),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_112),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_169),
.A2(n_103),
.B1(n_107),
.B2(n_94),
.Y(n_201)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_111),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_173),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_127),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_171),
.A2(n_175),
.B1(n_158),
.B2(n_150),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_120),
.B(n_3),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_130),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_110),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_127),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_90),
.Y(n_176)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_176),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_90),
.B(n_9),
.C(n_98),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_98),
.Y(n_178)
);

INVx13_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

AND2x6_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_110),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_184),
.B(n_186),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_141),
.B(n_104),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_191),
.B(n_194),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_193),
.A2(n_203),
.B1(n_208),
.B2(n_186),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_136),
.B(n_104),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_159),
.A2(n_129),
.B1(n_123),
.B2(n_116),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_196),
.A2(n_201),
.B1(n_210),
.B2(n_217),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_168),
.A2(n_129),
.B1(n_103),
.B2(n_107),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_207),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_111),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_174),
.A2(n_149),
.B1(n_135),
.B2(n_132),
.Y(n_208)
);

A2O1A1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_135),
.A2(n_91),
.B(n_133),
.C(n_174),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_209),
.B(n_213),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_135),
.A2(n_91),
.B1(n_177),
.B2(n_175),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_155),
.B(n_156),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_211),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_140),
.B(n_171),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_218),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_134),
.B(n_138),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_191),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_139),
.B(n_178),
.Y(n_218)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_220),
.Y(n_221)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_221),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_183),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_223),
.B(n_235),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_224),
.B(n_226),
.Y(n_258)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_215),
.Y(n_225)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_225),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_218),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_208),
.A2(n_157),
.B(n_143),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_227),
.A2(n_244),
.B(n_219),
.Y(n_278)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_198),
.Y(n_228)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_228),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_230),
.B(n_240),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_210),
.A2(n_153),
.B1(n_164),
.B2(n_170),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_233),
.A2(n_231),
.B1(n_251),
.B2(n_223),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_234),
.B(n_247),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_180),
.B(n_176),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_188),
.B(n_205),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_238),
.Y(n_263)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_182),
.Y(n_239)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_239),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_198),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_185),
.Y(n_241)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_241),
.Y(n_279)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_185),
.Y(n_242)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_242),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_207),
.B(n_194),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_246),
.Y(n_266)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_182),
.Y(n_245)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_245),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_195),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_216),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_203),
.B(n_181),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_249),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_200),
.B(n_181),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_200),
.B(n_214),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_254),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_190),
.A2(n_200),
.B1(n_217),
.B2(n_213),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_251),
.A2(n_192),
.B1(n_216),
.B2(n_206),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_209),
.A2(n_201),
.B(n_193),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_253),
.A2(n_179),
.B(n_199),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_204),
.B(n_190),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_192),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_212),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_184),
.A2(n_199),
.B1(n_183),
.B2(n_220),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_256),
.A2(n_212),
.B1(n_219),
.B2(n_253),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_259),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_179),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_260),
.B(n_271),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_225),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_202),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_262),
.B(n_264),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_237),
.B(n_202),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_236),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_265),
.B(n_276),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_202),
.Y(n_271)
);

FAx1_ASAP7_75t_SL g273 ( 
.A(n_249),
.B(n_219),
.CI(n_189),
.CON(n_273),
.SN(n_273)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_280),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_189),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_227),
.C(n_232),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_206),
.Y(n_276)
);

AO21x1_ASAP7_75t_L g301 ( 
.A1(n_278),
.A2(n_283),
.B(n_242),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_240),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_281),
.A2(n_287),
.B1(n_223),
.B2(n_221),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_222),
.B(n_212),
.Y(n_283)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_286),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_234),
.A2(n_248),
.B1(n_254),
.B2(n_256),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_288),
.A2(n_229),
.B1(n_238),
.B2(n_228),
.Y(n_299)
);

AOI211xp5_ASAP7_75t_SL g289 ( 
.A1(n_259),
.A2(n_244),
.B(n_232),
.C(n_222),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_289),
.A2(n_297),
.B(n_301),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_290),
.B(n_284),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_291),
.B(n_292),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_286),
.Y(n_292)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_272),
.Y(n_296)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_296),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_231),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_243),
.C(n_229),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_298),
.B(n_308),
.C(n_263),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_299),
.A2(n_305),
.B1(n_270),
.B2(n_261),
.Y(n_322)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_272),
.Y(n_300)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_300),
.Y(n_325)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_279),
.Y(n_303)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_303),
.Y(n_326)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_279),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_304),
.B(n_306),
.Y(n_334)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_282),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_266),
.B(n_263),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_307),
.B(n_311),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_275),
.B(n_241),
.C(n_245),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_257),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_310),
.B(n_312),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_266),
.B(n_255),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_285),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_282),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_313),
.Y(n_323)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_257),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_315),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_264),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_317),
.B(n_318),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_262),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_290),
.B(n_288),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_319),
.B(n_320),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_274),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_322),
.B(n_329),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_324),
.B(n_335),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_294),
.A2(n_281),
.B1(n_258),
.B2(n_269),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_327),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_297),
.A2(n_270),
.B1(n_268),
.B2(n_273),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_289),
.A2(n_273),
.B(n_269),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_332),
.A2(n_311),
.B(n_302),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_295),
.A2(n_283),
.B1(n_270),
.B2(n_268),
.Y(n_333)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_333),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_298),
.B(n_284),
.C(n_267),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_336),
.B(n_337),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_307),
.B(n_267),
.Y(n_337)
);

BUFx12f_ASAP7_75t_SL g339 ( 
.A(n_321),
.Y(n_339)
);

INVx11_ASAP7_75t_L g359 ( 
.A(n_339),
.Y(n_359)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_334),
.Y(n_344)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_344),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_338),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_346),
.B(n_351),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_328),
.A2(n_297),
.B1(n_309),
.B2(n_299),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_347),
.A2(n_322),
.B1(n_329),
.B2(n_309),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_350),
.B(n_293),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_330),
.B(n_310),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_331),
.B(n_292),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_352),
.B(n_355),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_336),
.B(n_291),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_353),
.B(n_354),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_316),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_325),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_324),
.B(n_315),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_356),
.B(n_357),
.Y(n_360)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_326),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_358),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_342),
.B(n_319),
.C(n_335),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_361),
.B(n_364),
.C(n_367),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_339),
.A2(n_321),
.B(n_301),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_362),
.A2(n_345),
.B(n_341),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_343),
.A2(n_332),
.B(n_293),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_363),
.B(n_371),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_340),
.B(n_320),
.C(n_337),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_349),
.B(n_348),
.C(n_318),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_341),
.A2(n_343),
.B1(n_347),
.B2(n_351),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_369),
.A2(n_354),
.B1(n_300),
.B2(n_303),
.Y(n_382)
);

XNOR2x1_ASAP7_75t_L g370 ( 
.A(n_348),
.B(n_317),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_370),
.B(n_357),
.C(n_355),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_365),
.B(n_344),
.Y(n_373)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_373),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_360),
.B(n_346),
.Y(n_375)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_375),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_359),
.B(n_350),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_376),
.B(n_378),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_359),
.B(n_352),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_379),
.B(n_362),
.Y(n_391)
);

OA21x2_ASAP7_75t_SL g380 ( 
.A1(n_366),
.A2(n_345),
.B(n_323),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_380),
.B(n_382),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_381),
.B(n_361),
.C(n_372),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_360),
.B(n_296),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_384),
.B(n_368),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_381),
.B(n_366),
.Y(n_387)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_387),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_388),
.B(n_390),
.Y(n_396)
);

MAJx2_ASAP7_75t_L g397 ( 
.A(n_391),
.B(n_363),
.C(n_368),
.Y(n_397)
);

INVx6_ASAP7_75t_L g392 ( 
.A(n_379),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_392),
.A2(n_394),
.B(n_377),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_374),
.B(n_372),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_391),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_395),
.B(n_400),
.Y(n_407)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_397),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_394),
.B(n_374),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_398),
.B(n_399),
.C(n_364),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_385),
.A2(n_383),
.B(n_377),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_387),
.Y(n_401)
);

AOI322xp5_ASAP7_75t_L g405 ( 
.A1(n_401),
.A2(n_371),
.A3(n_367),
.B1(n_358),
.B2(n_370),
.C1(n_304),
.C2(n_277),
.Y(n_405)
);

AOI322xp5_ASAP7_75t_L g403 ( 
.A1(n_402),
.A2(n_393),
.A3(n_389),
.B1(n_369),
.B2(n_386),
.C1(n_306),
.C2(n_313),
.Y(n_403)
);

AOI322xp5_ASAP7_75t_L g410 ( 
.A1(n_403),
.A2(n_405),
.A3(n_397),
.B1(n_277),
.B2(n_247),
.C1(n_239),
.C2(n_221),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_404),
.B(n_396),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_407),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_408),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_411),
.B(n_409),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_412),
.B(n_406),
.C(n_410),
.Y(n_413)
);


endmodule