module fake_netlist_1_9478_n_37 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_10, n_8, n_0, n_37);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_10;
input n_8;
input n_0;
output n_37;
wire n_20;
wire n_36;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_17;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
BUFx6f_ASAP7_75t_L g15 ( .A(n_13), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_6), .Y(n_16) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_0), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_12), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_10), .Y(n_19) );
NOR2xp67_ASAP7_75t_L g20 ( .A(n_1), .B(n_4), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_11), .Y(n_21) );
CKINVDCx11_ASAP7_75t_R g22 ( .A(n_17), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_16), .Y(n_23) );
AOI22xp5_ASAP7_75t_SL g24 ( .A1(n_17), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_24) );
AOI21xp5_ASAP7_75t_L g25 ( .A1(n_23), .A2(n_18), .B(n_21), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_23), .B(n_19), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
OR2x2_ASAP7_75t_L g28 ( .A(n_25), .B(n_24), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
OAI22xp33_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_28), .B1(n_22), .B2(n_24), .Y(n_30) );
AOI22xp33_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_16), .B1(n_20), .B2(n_19), .Y(n_31) );
OAI211xp5_ASAP7_75t_SL g32 ( .A1(n_31), .A2(n_2), .B(n_3), .C(n_5), .Y(n_32) );
NAND2xp5_ASAP7_75t_L g33 ( .A(n_30), .B(n_3), .Y(n_33) );
OAI221xp5_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_15), .B1(n_7), .B2(n_8), .C(n_6), .Y(n_34) );
OAI211xp5_ASAP7_75t_L g35 ( .A1(n_32), .A2(n_15), .B(n_8), .C(n_14), .Y(n_35) );
HB1xp67_ASAP7_75t_L g36 ( .A(n_34), .Y(n_36) );
AOI22xp5_ASAP7_75t_SL g37 ( .A1(n_36), .A2(n_15), .B1(n_35), .B2(n_9), .Y(n_37) );
endmodule