module fake_jpeg_4021_n_61 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_61);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_61;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

INVx8_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

INVx6_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_0),
.B(n_8),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_0),
.B(n_5),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_19),
.A2(n_21),
.B1(n_11),
.B2(n_16),
.Y(n_29)
);

OAI21xp33_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_1),
.B(n_2),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_20),
.B(n_22),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_11),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_15),
.B(n_3),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_14),
.B(n_5),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_29),
.A2(n_33),
.B1(n_21),
.B2(n_9),
.Y(n_40)
);

NAND2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_18),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_30),
.A2(n_22),
.B(n_25),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_12),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_19),
.A2(n_16),
.B1(n_9),
.B2(n_10),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_10),
.C(n_13),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_13),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_38),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_33),
.B1(n_26),
.B2(n_28),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_40),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_41),
.Y(n_47)
);

A2O1A1O1Ixp25_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_12),
.B(n_32),
.C(n_9),
.D(n_27),
.Y(n_43)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_36),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_53),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_39),
.C(n_38),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_51),
.C(n_52),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_40),
.C(n_32),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_35),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_35),
.C(n_27),
.Y(n_53)
);

NOR2x1_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_43),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_5),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_17),
.B(n_18),
.Y(n_57)
);

INVxp33_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_54),
.B1(n_17),
.B2(n_55),
.Y(n_60)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_58),
.B(n_12),
.C(n_56),
.Y(n_61)
);


endmodule