module real_aes_16602_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_756;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_839;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
wire n_869;
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_0), .Y(n_239) );
AND2x4_ASAP7_75t_L g104 ( .A(n_1), .B(n_105), .Y(n_104) );
BUFx3_ASAP7_75t_L g180 ( .A(n_2), .Y(n_180) );
INVx1_ASAP7_75t_L g105 ( .A(n_3), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_4), .B(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g869 ( .A(n_4), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_5), .B(n_152), .Y(n_151) );
BUFx2_ASAP7_75t_L g112 ( .A(n_6), .Y(n_112) );
OR2x2_ASAP7_75t_L g121 ( .A(n_6), .B(n_20), .Y(n_121) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_7), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_8), .B(n_174), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_9), .B(n_174), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_10), .B(n_199), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_11), .A2(n_79), .B1(n_149), .B2(n_174), .Y(n_248) );
OAI21x1_ASAP7_75t_L g144 ( .A1(n_12), .A2(n_33), .B(n_145), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_13), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_14), .B(n_189), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g535 ( .A(n_15), .Y(n_535) );
AO32x2_ASAP7_75t_L g245 ( .A1(n_16), .A2(n_166), .A3(n_167), .B1(n_246), .B2(n_249), .Y(n_245) );
AO32x1_ASAP7_75t_L g283 ( .A1(n_16), .A2(n_166), .A3(n_167), .B1(n_246), .B2(n_249), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_17), .B(n_520), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_18), .B(n_166), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g548 ( .A(n_19), .Y(n_548) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_20), .Y(n_110) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_21), .A2(n_39), .B1(n_177), .B2(n_189), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g247 ( .A1(n_22), .A2(n_87), .B1(n_149), .B2(n_157), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_23), .B(n_156), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g539 ( .A(n_24), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_25), .B(n_212), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_26), .A2(n_58), .B1(n_157), .B2(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_27), .B(n_174), .Y(n_590) );
INVx2_ASAP7_75t_L g855 ( .A(n_28), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_29), .B(n_153), .Y(n_621) );
BUFx3_ASAP7_75t_L g108 ( .A(n_30), .Y(n_108) );
INVx1_ASAP7_75t_L g119 ( .A(n_30), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_31), .B(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_32), .B(n_526), .Y(n_627) );
AND2x2_ASAP7_75t_L g541 ( .A(n_34), .B(n_526), .Y(n_541) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_35), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_36), .B(n_211), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_37), .B(n_520), .Y(n_519) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_38), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_40), .B(n_553), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g210 ( .A1(n_41), .A2(n_73), .B1(n_211), .B2(n_212), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_42), .B(n_254), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_43), .A2(n_190), .B(n_237), .C(n_534), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g173 ( .A1(n_44), .A2(n_75), .B1(n_149), .B2(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g145 ( .A(n_45), .Y(n_145) );
AND2x4_ASAP7_75t_L g163 ( .A(n_46), .B(n_164), .Y(n_163) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_47), .A2(n_48), .B1(n_157), .B2(n_177), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_49), .B(n_166), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_50), .B(n_526), .Y(n_565) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_51), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_52), .B(n_157), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_53), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g164 ( .A(n_54), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_55), .B(n_166), .Y(n_165) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_56), .A2(n_237), .B(n_238), .C(n_240), .Y(n_236) );
NAND3xp33_ASAP7_75t_L g161 ( .A(n_57), .B(n_149), .C(n_159), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g601 ( .A(n_59), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_60), .B(n_166), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_61), .B(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g242 ( .A(n_62), .B(n_243), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_63), .Y(n_258) );
NAND3xp33_ASAP7_75t_L g622 ( .A(n_64), .B(n_153), .C(n_189), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g215 ( .A1(n_65), .A2(n_91), .B1(n_174), .B2(n_211), .Y(n_215) );
INVx2_ASAP7_75t_L g154 ( .A(n_66), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_67), .B(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_68), .B(n_518), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_69), .B(n_174), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_70), .B(n_214), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g858 ( .A1(n_71), .A2(n_859), .B1(n_870), .B2(n_874), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_72), .A2(n_100), .B1(n_113), .B2(n_879), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_74), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_76), .B(n_193), .Y(n_575) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_77), .Y(n_115) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_78), .A2(n_86), .B1(n_520), .B2(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_80), .B(n_174), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_81), .B(n_159), .Y(n_158) );
NAND2xp33_ASAP7_75t_SL g564 ( .A(n_82), .B(n_152), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_83), .B(n_187), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g176 ( .A1(n_84), .A2(n_98), .B1(n_157), .B2(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_85), .B(n_212), .Y(n_269) );
AOI22xp33_ASAP7_75t_SL g123 ( .A1(n_88), .A2(n_124), .B1(n_849), .B2(n_850), .Y(n_123) );
INVx1_ASAP7_75t_SL g850 ( .A(n_88), .Y(n_850) );
INVx1_ASAP7_75t_L g107 ( .A(n_89), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g864 ( .A(n_89), .B(n_865), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_90), .B(n_199), .Y(n_275) );
NAND2xp33_ASAP7_75t_L g573 ( .A(n_92), .B(n_152), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_93), .B(n_526), .Y(n_525) );
NAND3xp33_ASAP7_75t_L g561 ( .A(n_94), .B(n_152), .C(n_214), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_95), .B(n_518), .Y(n_592) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_96), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_97), .B(n_520), .Y(n_523) );
BUFx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
AND2x4_ASAP7_75t_L g101 ( .A(n_102), .B(n_109), .Y(n_101) );
AND2x6_ASAP7_75t_L g880 ( .A(n_102), .B(n_109), .Y(n_880) );
NOR3x1_ASAP7_75t_L g102 ( .A(n_103), .B(n_106), .C(n_108), .Y(n_102) );
INVx2_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
AND3x2_ASAP7_75t_L g117 ( .A(n_106), .B(n_118), .C(n_120), .Y(n_117) );
BUFx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g128 ( .A(n_107), .Y(n_128) );
INVx1_ASAP7_75t_L g857 ( .A(n_108), .Y(n_857) );
NOR2x1_ASAP7_75t_L g878 ( .A(n_108), .B(n_121), .Y(n_878) );
NOR2x1p5_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OR2x6_ASAP7_75t_L g113 ( .A(n_114), .B(n_122), .Y(n_113) );
AOI31xp33_ASAP7_75t_L g868 ( .A1(n_114), .A2(n_130), .A3(n_861), .B(n_869), .Y(n_868) );
NOR2x1_ASAP7_75t_SL g114 ( .A(n_115), .B(n_116), .Y(n_114) );
INVx4_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g865 ( .A(n_119), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_120), .B(n_857), .Y(n_856) );
AND2x6_ASAP7_75t_SL g863 ( .A(n_120), .B(n_864), .Y(n_863) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI21xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_851), .B(n_858), .Y(n_122) );
INVx1_ASAP7_75t_L g849 ( .A(n_124), .Y(n_849) );
OA21x2_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_129), .B(n_505), .Y(n_124) );
INVx8_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
BUFx12f_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_128), .Y(n_127) );
BUFx8_ASAP7_75t_SL g848 ( .A(n_128), .Y(n_848) );
AND2x2_ASAP7_75t_L g877 ( .A(n_128), .B(n_878), .Y(n_877) );
BUFx2_ASAP7_75t_L g867 ( .A(n_129), .Y(n_867) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OR2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_415), .Y(n_130) );
NAND4xp25_ASAP7_75t_L g131 ( .A(n_132), .B(n_320), .C(n_347), .D(n_383), .Y(n_131) );
AOI221x1_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_225), .B1(n_259), .B2(n_295), .C(n_299), .Y(n_132) );
NAND3xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_201), .C(n_223), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_168), .Y(n_136) );
INVx2_ASAP7_75t_L g260 ( .A(n_137), .Y(n_260) );
AND2x2_ASAP7_75t_L g433 ( .A(n_137), .B(n_377), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_137), .B(n_224), .Y(n_442) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g448 ( .A(n_138), .Y(n_448) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g293 ( .A(n_139), .Y(n_293) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OR2x2_ASAP7_75t_L g376 ( .A(n_140), .B(n_222), .Y(n_376) );
OAI21x1_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_146), .B(n_165), .Y(n_140) );
OAI21xp5_ASAP7_75t_L g305 ( .A1(n_141), .A2(n_146), .B(n_165), .Y(n_305) );
OAI21x1_ASAP7_75t_L g514 ( .A1(n_141), .A2(n_515), .B(n_525), .Y(n_514) );
OAI21xp5_ASAP7_75t_L g545 ( .A1(n_141), .A2(n_546), .B(n_554), .Y(n_545) );
OAI21x1_ASAP7_75t_L g644 ( .A1(n_141), .A2(n_546), .B(n_554), .Y(n_644) );
OAI21xp33_ASAP7_75t_SL g735 ( .A1(n_141), .A2(n_515), .B(n_525), .Y(n_735) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g526 ( .A(n_142), .Y(n_526) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g200 ( .A(n_143), .Y(n_200) );
INVx2_ASAP7_75t_L g220 ( .A(n_143), .Y(n_220) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_144), .Y(n_167) );
OAI21x1_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_155), .B(n_162), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_151), .B(n_153), .Y(n_147) );
INVx2_ASAP7_75t_SL g212 ( .A(n_149), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_149), .B(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_150), .Y(n_152) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_150), .Y(n_157) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_150), .Y(n_174) );
INVx1_ASAP7_75t_L g177 ( .A(n_150), .Y(n_177) );
INVx1_ASAP7_75t_L g187 ( .A(n_150), .Y(n_187) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_150), .Y(n_189) );
INVx1_ASAP7_75t_L g211 ( .A(n_150), .Y(n_211) );
INVx1_ASAP7_75t_L g237 ( .A(n_150), .Y(n_237) );
INVx3_ASAP7_75t_L g518 ( .A(n_150), .Y(n_518) );
INVx1_ASAP7_75t_L g521 ( .A(n_150), .Y(n_521) );
INVx2_ASAP7_75t_L g553 ( .A(n_152), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g172 ( .A1(n_153), .A2(n_173), .B1(n_175), .B2(n_176), .Y(n_172) );
INVx6_ASAP7_75t_L g175 ( .A(n_153), .Y(n_175) );
OAI22xp5_ASAP7_75t_L g246 ( .A1(n_153), .A2(n_190), .B1(n_247), .B2(n_248), .Y(n_246) );
O2A1O1Ixp5_ASAP7_75t_L g547 ( .A1(n_153), .A2(n_186), .B(n_548), .C(n_549), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g591 ( .A1(n_153), .A2(n_592), .B(n_593), .Y(n_591) );
BUFx8_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g160 ( .A(n_154), .Y(n_160) );
INVx2_ASAP7_75t_L g195 ( .A(n_154), .Y(n_195) );
INVx1_ASAP7_75t_L g214 ( .A(n_154), .Y(n_214) );
OAI21xp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_158), .B(n_161), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
OAI22xp33_ASAP7_75t_L g538 ( .A1(n_157), .A2(n_518), .B1(n_539), .B2(n_540), .Y(n_538) );
INVx2_ASAP7_75t_L g598 ( .A(n_157), .Y(n_598) );
OAI21xp5_ASAP7_75t_L g620 ( .A1(n_157), .A2(n_621), .B(n_622), .Y(n_620) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
BUFx4f_ASAP7_75t_L g190 ( .A(n_160), .Y(n_190) );
AOI31xp67_ASAP7_75t_L g170 ( .A1(n_162), .A2(n_171), .A3(n_172), .B(n_178), .Y(n_170) );
OAI21x1_ASAP7_75t_L g183 ( .A1(n_162), .A2(n_184), .B(n_191), .Y(n_183) );
OAI21x1_ASAP7_75t_L g515 ( .A1(n_162), .A2(n_516), .B(n_522), .Y(n_515) );
OAI21x1_ASAP7_75t_L g546 ( .A1(n_162), .A2(n_547), .B(n_550), .Y(n_546) );
OAI21x1_ASAP7_75t_L g558 ( .A1(n_162), .A2(n_559), .B(n_562), .Y(n_558) );
AND2x4_ASAP7_75t_SL g578 ( .A(n_162), .B(n_167), .Y(n_578) );
OAI21x1_ASAP7_75t_L g587 ( .A1(n_162), .A2(n_588), .B(n_591), .Y(n_587) );
OAI21x1_ASAP7_75t_L g619 ( .A1(n_162), .A2(n_620), .B(n_623), .Y(n_619) );
BUFx10_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g217 ( .A(n_163), .Y(n_217) );
INVx1_ASAP7_75t_L g241 ( .A(n_163), .Y(n_241) );
AO31x2_ASAP7_75t_L g251 ( .A1(n_163), .A2(n_208), .A3(n_252), .B(n_257), .Y(n_251) );
BUFx10_ASAP7_75t_L g531 ( .A(n_163), .Y(n_531) );
INVx2_ASAP7_75t_L g171 ( .A(n_166), .Y(n_171) );
INVx4_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_167), .B(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g182 ( .A(n_167), .Y(n_182) );
BUFx3_ASAP7_75t_L g208 ( .A(n_167), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_167), .B(n_258), .Y(n_257) );
INVx2_ASAP7_75t_SL g266 ( .A(n_167), .Y(n_266) );
INVx1_ASAP7_75t_SL g557 ( .A(n_167), .Y(n_557) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_168), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_168), .B(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g446 ( .A(n_168), .Y(n_446) );
AND2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_181), .Y(n_168) );
AND2x2_ASAP7_75t_L g224 ( .A(n_169), .B(n_207), .Y(n_224) );
INVx2_ASAP7_75t_L g302 ( .A(n_169), .Y(n_302) );
AND2x2_ASAP7_75t_L g367 ( .A(n_169), .B(n_305), .Y(n_367) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g222 ( .A(n_170), .Y(n_222) );
INVx3_ASAP7_75t_L g274 ( .A(n_174), .Y(n_274) );
OAI21xp5_ASAP7_75t_L g559 ( .A1(n_174), .A2(n_560), .B(n_561), .Y(n_559) );
INVx1_ASAP7_75t_L g626 ( .A(n_174), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g209 ( .A1(n_175), .A2(n_210), .B1(n_213), .B2(n_215), .Y(n_209) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_175), .A2(n_253), .B1(n_255), .B2(n_256), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_175), .A2(n_272), .B(n_273), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_175), .A2(n_537), .B1(n_597), .B2(n_599), .Y(n_596) );
INVx1_ASAP7_75t_L g196 ( .A(n_177), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g232 ( .A1(n_177), .A2(n_189), .B1(n_233), .B2(n_234), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g294 ( .A(n_181), .Y(n_294) );
AND2x2_ASAP7_75t_L g304 ( .A(n_181), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g366 ( .A(n_181), .B(n_207), .Y(n_366) );
OA21x2_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_198), .Y(n_181) );
OA21x2_ASAP7_75t_L g204 ( .A1(n_182), .A2(n_183), .B(n_198), .Y(n_204) );
OAI21x1_ASAP7_75t_L g586 ( .A1(n_182), .A2(n_587), .B(n_594), .Y(n_586) );
OAI21x1_ASAP7_75t_L g618 ( .A1(n_182), .A2(n_619), .B(n_627), .Y(n_618) );
OA21x2_ASAP7_75t_L g630 ( .A1(n_182), .A2(n_619), .B(n_627), .Y(n_630) );
OAI21x1_ASAP7_75t_L g633 ( .A1(n_182), .A2(n_587), .B(n_594), .Y(n_633) );
O2A1O1Ixp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_188), .C(n_190), .Y(n_184) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g254 ( .A(n_189), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_190), .A2(n_517), .B(n_519), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_190), .A2(n_563), .B(n_564), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_190), .A2(n_572), .B(n_573), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_190), .A2(n_589), .B(n_590), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_194), .B1(n_196), .B2(n_197), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_193), .A2(n_551), .B(n_552), .Y(n_550) );
INVx2_ASAP7_75t_SL g193 ( .A(n_194), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_194), .A2(n_575), .B1(n_576), .B2(n_577), .Y(n_574) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
BUFx3_ASAP7_75t_L g240 ( .A(n_195), .Y(n_240) );
INVx2_ASAP7_75t_L g229 ( .A(n_199), .Y(n_229) );
NOR2xp67_ASAP7_75t_SL g529 ( .A(n_199), .B(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AO31x2_ASAP7_75t_L g595 ( .A1(n_200), .A2(n_531), .A3(n_596), .B(n_600), .Y(n_595) );
INVx1_ASAP7_75t_L g331 ( .A(n_201), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_202), .B(n_205), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_203), .B(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_203), .B(n_346), .Y(n_345) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_203), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_203), .B(n_401), .Y(n_408) );
INVx2_ASAP7_75t_SL g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g377 ( .A(n_204), .B(n_352), .Y(n_377) );
OR2x2_ASAP7_75t_L g379 ( .A(n_204), .B(n_305), .Y(n_379) );
INVx1_ASAP7_75t_L g438 ( .A(n_204), .Y(n_438) );
BUFx2_ASAP7_75t_L g452 ( .A(n_204), .Y(n_452) );
OR2x2_ASAP7_75t_L g480 ( .A(n_204), .B(n_207), .Y(n_480) );
INVx1_ASAP7_75t_L g499 ( .A(n_205), .Y(n_499) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g346 ( .A(n_206), .Y(n_346) );
OR2x2_ASAP7_75t_L g359 ( .A(n_206), .B(n_360), .Y(n_359) );
OR2x2_ASAP7_75t_L g378 ( .A(n_206), .B(n_379), .Y(n_378) );
OR2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_221), .Y(n_206) );
INVx2_ASAP7_75t_L g298 ( .A(n_207), .Y(n_298) );
AND2x2_ASAP7_75t_L g314 ( .A(n_207), .B(n_221), .Y(n_314) );
INVx1_ASAP7_75t_L g352 ( .A(n_207), .Y(n_352) );
INVx1_ASAP7_75t_L g395 ( .A(n_207), .Y(n_395) );
AND2x2_ASAP7_75t_L g437 ( .A(n_207), .B(n_438), .Y(n_437) );
AO31x2_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .A3(n_216), .B(n_218), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_211), .B(n_239), .Y(n_238) );
INVx1_ASAP7_75t_SL g213 ( .A(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g235 ( .A(n_214), .Y(n_235) );
INVx2_ASAP7_75t_SL g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_SL g249 ( .A(n_217), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
INVx2_ASAP7_75t_L g243 ( .A(n_220), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_220), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g493 ( .A(n_223), .Y(n_493) );
AND2x4_ASAP7_75t_L g431 ( .A(n_224), .B(n_291), .Y(n_431) );
INVx2_ASAP7_75t_L g460 ( .A(n_224), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_224), .B(n_452), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_225), .B(n_450), .Y(n_449) );
AND2x4_ASAP7_75t_L g225 ( .A(n_226), .B(n_244), .Y(n_225) );
AND2x2_ASAP7_75t_L g371 ( .A(n_226), .B(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g392 ( .A(n_226), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
OR2x2_ASAP7_75t_L g263 ( .A(n_227), .B(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g287 ( .A(n_227), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g318 ( .A(n_227), .Y(n_318) );
AND2x2_ASAP7_75t_L g358 ( .A(n_227), .B(n_250), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_227), .B(n_342), .Y(n_399) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g311 ( .A(n_228), .Y(n_311) );
AOI21x1_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_242), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_236), .B(n_241), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_232), .B(n_235), .Y(n_231) );
AOI21x1_ASAP7_75t_L g623 ( .A1(n_235), .A2(n_624), .B(n_625), .Y(n_623) );
INVx1_ASAP7_75t_L g576 ( .A(n_237), .Y(n_576) );
INVx2_ASAP7_75t_L g256 ( .A(n_240), .Y(n_256) );
INVx2_ASAP7_75t_L g537 ( .A(n_240), .Y(n_537) );
INVx3_ASAP7_75t_L g277 ( .A(n_244), .Y(n_277) );
AND2x2_ASAP7_75t_L g322 ( .A(n_244), .B(n_317), .Y(n_322) );
AND2x2_ASAP7_75t_L g477 ( .A(n_244), .B(n_281), .Y(n_477) );
AND2x4_ASAP7_75t_L g244 ( .A(n_245), .B(n_250), .Y(n_244) );
INVx1_ASAP7_75t_L g328 ( .A(n_245), .Y(n_328) );
AND2x2_ASAP7_75t_L g356 ( .A(n_245), .B(n_264), .Y(n_356) );
OAI21x1_ASAP7_75t_L g267 ( .A1(n_249), .A2(n_268), .B(n_271), .Y(n_267) );
AND2x4_ASAP7_75t_L g309 ( .A(n_250), .B(n_310), .Y(n_309) );
INVx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g282 ( .A(n_251), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g319 ( .A(n_251), .B(n_283), .Y(n_319) );
AND2x2_ASAP7_75t_L g329 ( .A(n_251), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_251), .B(n_264), .Y(n_381) );
AND2x2_ASAP7_75t_L g387 ( .A(n_251), .B(n_311), .Y(n_387) );
AOI21x1_ASAP7_75t_L g268 ( .A1(n_256), .A2(n_269), .B(n_270), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_256), .A2(n_523), .B(n_524), .Y(n_522) );
OAI21xp33_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_261), .B(n_278), .Y(n_259) );
OAI21xp33_ASAP7_75t_L g420 ( .A1(n_260), .A2(n_421), .B(n_425), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_260), .B(n_451), .Y(n_498) );
NAND2x1_ASAP7_75t_SL g261 ( .A(n_262), .B(n_276), .Y(n_261) );
INVx1_ASAP7_75t_L g504 ( .A(n_262), .Y(n_504) );
INVx3_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
BUFx2_ASAP7_75t_L g281 ( .A(n_264), .Y(n_281) );
INVx2_ASAP7_75t_L g286 ( .A(n_264), .Y(n_286) );
INVxp67_ASAP7_75t_L g307 ( .A(n_264), .Y(n_307) );
AND2x2_ASAP7_75t_L g327 ( .A(n_264), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g338 ( .A(n_264), .B(n_339), .Y(n_338) );
INVx3_ASAP7_75t_L g342 ( .A(n_264), .Y(n_342) );
INVx1_ASAP7_75t_L g360 ( .A(n_264), .Y(n_360) );
OR2x2_ASAP7_75t_L g393 ( .A(n_264), .B(n_328), .Y(n_393) );
INVx1_ASAP7_75t_L g464 ( .A(n_264), .Y(n_464) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OAI21x1_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_267), .B(n_275), .Y(n_265) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OAI21xp33_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_284), .B(n_289), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OAI22xp33_ASAP7_75t_L g402 ( .A1(n_280), .A2(n_403), .B1(n_405), .B2(n_408), .Y(n_402) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_281), .B(n_329), .Y(n_363) );
BUFx2_ASAP7_75t_L g422 ( .A(n_281), .Y(n_422) );
INVx2_ASAP7_75t_L g372 ( .A(n_282), .Y(n_372) );
OR2x2_ASAP7_75t_L g456 ( .A(n_282), .B(n_286), .Y(n_456) );
INVx1_ASAP7_75t_L g288 ( .A(n_283), .Y(n_288) );
INVx1_ASAP7_75t_L g337 ( .A(n_283), .Y(n_337) );
NOR2x1p5_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
INVxp67_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_286), .Y(n_407) );
OR2x2_ASAP7_75t_L g491 ( .A(n_286), .B(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g494 ( .A(n_286), .B(n_329), .Y(n_494) );
INVxp67_ASAP7_75t_SL g457 ( .A(n_287), .Y(n_457) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_291), .B(n_351), .Y(n_413) );
AND2x2_ASAP7_75t_L g503 ( .A(n_291), .B(n_301), .Y(n_503) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g412 ( .A(n_292), .B(n_301), .Y(n_412) );
NAND2x1p5_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
AND2x2_ASAP7_75t_L g369 ( .A(n_293), .B(n_302), .Y(n_369) );
AND2x2_ASAP7_75t_L g404 ( .A(n_293), .B(n_298), .Y(n_404) );
INVxp67_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g323 ( .A(n_296), .B(n_304), .Y(n_323) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx2_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g463 ( .A(n_298), .B(n_464), .Y(n_463) );
OAI22xp33_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_306), .B1(n_312), .B2(n_315), .Y(n_299) );
O2A1O1Ixp33_ASAP7_75t_L g500 ( .A1(n_300), .A2(n_501), .B(n_502), .C(n_504), .Y(n_500) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g351 ( .A(n_302), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g419 ( .A(n_302), .Y(n_419) );
OR2x2_ASAP7_75t_L g466 ( .A(n_303), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
AND2x2_ASAP7_75t_L g321 ( .A(n_307), .B(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g424 ( .A(n_310), .Y(n_424) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g330 ( .A(n_311), .Y(n_330) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_311), .Y(n_339) );
INVx1_ASAP7_75t_L g411 ( .A(n_311), .Y(n_411) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g467 ( .A(n_314), .Y(n_467) );
AND2x2_ASAP7_75t_L g489 ( .A(n_314), .B(n_452), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_315), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g341 ( .A(n_319), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g397 ( .A(n_319), .B(n_398), .Y(n_397) );
INVx2_ASAP7_75t_SL g492 ( .A(n_319), .Y(n_492) );
AOI221xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_323), .B1(n_324), .B2(n_331), .C(n_332), .Y(n_320) );
INVxp67_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
INVx2_ASAP7_75t_L g414 ( .A(n_327), .Y(n_414) );
BUFx2_ASAP7_75t_L g434 ( .A(n_329), .Y(n_434) );
AOI21xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_340), .B(n_343), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_335), .B(n_338), .Y(n_334) );
AND2x2_ASAP7_75t_L g476 ( .A(n_335), .B(n_398), .Y(n_476) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g382 ( .A(n_337), .Y(n_382) );
AND2x2_ASAP7_75t_L g472 ( .A(n_337), .B(n_342), .Y(n_472) );
INVx1_ASAP7_75t_L g355 ( .A(n_339), .Y(n_355) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AOI211xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_349), .B(n_361), .C(n_373), .Y(n_347) );
OAI22xp33_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_353), .B1(n_357), .B2(n_359), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
BUFx2_ASAP7_75t_L g389 ( .A(n_356), .Y(n_389) );
AND2x2_ASAP7_75t_L g482 ( .A(n_356), .B(n_424), .Y(n_482) );
OAI21xp33_ASAP7_75t_L g485 ( .A1(n_357), .A2(n_486), .B(n_488), .Y(n_485) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI22xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_364), .B1(n_368), .B2(n_370), .Y(n_361) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_364), .B(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVxp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x4_ASAP7_75t_L g436 ( .A(n_369), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x4_ASAP7_75t_L g423 ( .A(n_372), .B(n_424), .Y(n_423) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_372), .Y(n_439) );
AOI21xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_378), .B(n_380), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_375), .B(n_377), .Y(n_374) );
AND2x2_ASAP7_75t_L g450 ( .A(n_375), .B(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g487 ( .A(n_375), .B(n_452), .Y(n_487) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g401 ( .A(n_376), .Y(n_401) );
OR2x2_ASAP7_75t_L g479 ( .A(n_376), .B(n_480), .Y(n_479) );
OR2x2_ASAP7_75t_L g394 ( .A(n_379), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g426 ( .A(n_379), .Y(n_426) );
OR2x2_ASAP7_75t_L g459 ( .A(n_379), .B(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g430 ( .A(n_380), .Y(n_430) );
OR2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
NOR3xp33_ASAP7_75t_L g383 ( .A(n_384), .B(n_402), .C(n_409), .Y(n_383) );
OAI322xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_388), .A3(n_390), .B1(n_392), .B2(n_394), .C1(n_396), .C2(n_400), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
A2O1A1Ixp33_ASAP7_75t_L g461 ( .A1(n_386), .A2(n_426), .B(n_462), .C(n_465), .Y(n_461) );
BUFx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g406 ( .A(n_387), .B(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g443 ( .A(n_387), .Y(n_443) );
AND2x4_ASAP7_75t_L g471 ( .A(n_387), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI32xp33_ASAP7_75t_L g440 ( .A1(n_389), .A2(n_427), .A3(n_441), .B1(n_443), .B2(n_444), .Y(n_440) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g427 ( .A(n_393), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_395), .B(n_448), .Y(n_447) );
INVxp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
O2A1O1Ixp33_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_412), .B(n_413), .C(n_414), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_416), .B(n_473), .Y(n_415) );
AOI211xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_420), .B(n_428), .C(n_453), .Y(n_416) );
INVxp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
O2A1O1Ixp33_ASAP7_75t_SL g495 ( .A1(n_421), .A2(n_496), .B(n_497), .C(n_499), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
OAI31xp33_ASAP7_75t_L g475 ( .A1(n_423), .A2(n_476), .A3(n_477), .B(n_478), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
INVx2_ASAP7_75t_L g435 ( .A(n_427), .Y(n_435) );
NAND4xp25_ASAP7_75t_SL g428 ( .A(n_429), .B(n_432), .C(n_440), .D(n_449), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
AOI32xp33_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_434), .A3(n_435), .B1(n_436), .B2(n_439), .Y(n_432) );
INVx1_ASAP7_75t_L g484 ( .A(n_436), .Y(n_484) );
INVx1_ASAP7_75t_L g496 ( .A(n_439), .Y(n_496) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NAND3xp33_ASAP7_75t_L g453 ( .A(n_454), .B(n_461), .C(n_468), .Y(n_453) );
OAI21xp5_ASAP7_75t_SL g454 ( .A1(n_455), .A2(n_457), .B(n_458), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_462), .B(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_471), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NOR4xp25_ASAP7_75t_L g473 ( .A(n_474), .B(n_485), .C(n_495), .D(n_500), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_481), .Y(n_474) );
OAI21xp33_ASAP7_75t_L g481 ( .A1(n_476), .A2(n_482), .B(n_483), .Y(n_481) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_490), .B1(n_493), .B2(n_494), .Y(n_488) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_492), .Y(n_501) );
INVxp67_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_848), .Y(n_505) );
NAND2x1p5_ASAP7_75t_L g506 ( .A(n_507), .B(n_743), .Y(n_506) );
NOR2x1_ASAP7_75t_L g507 ( .A(n_508), .B(n_678), .Y(n_507) );
NAND3xp33_ASAP7_75t_L g508 ( .A(n_509), .B(n_602), .C(n_651), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_542), .B(n_566), .C(n_583), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
OR2x2_ASAP7_75t_L g817 ( .A(n_511), .B(n_736), .Y(n_817) );
OR2x2_ASAP7_75t_L g828 ( .A(n_511), .B(n_829), .Y(n_828) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_512), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g719 ( .A(n_512), .B(n_609), .Y(n_719) );
AND2x2_ASAP7_75t_L g840 ( .A(n_512), .B(n_650), .Y(n_840) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_527), .Y(n_512) );
INVx2_ASAP7_75t_L g670 ( .A(n_513), .Y(n_670) );
AND2x2_ASAP7_75t_L g685 ( .A(n_513), .B(n_637), .Y(n_685) );
AND2x2_ASAP7_75t_L g694 ( .A(n_513), .B(n_568), .Y(n_694) );
AND2x2_ASAP7_75t_L g763 ( .A(n_513), .B(n_649), .Y(n_763) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g581 ( .A(n_514), .Y(n_581) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g734 ( .A(n_527), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g582 ( .A(n_528), .B(n_556), .Y(n_582) );
INVx2_ASAP7_75t_L g607 ( .A(n_528), .Y(n_607) );
AOI21x1_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_532), .B(n_541), .Y(n_528) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_536), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
AND2x2_ASAP7_75t_L g771 ( .A(n_542), .B(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_555), .Y(n_543) );
INVx1_ASAP7_75t_L g791 ( .A(n_544), .Y(n_791) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g629 ( .A(n_545), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g712 ( .A(n_545), .B(n_618), .Y(n_712) );
AND2x2_ASAP7_75t_L g638 ( .A(n_555), .B(n_581), .Y(n_638) );
INVxp67_ASAP7_75t_L g787 ( .A(n_555), .Y(n_787) );
OR2x2_ASAP7_75t_L g829 ( .A(n_555), .B(n_568), .Y(n_829) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g611 ( .A(n_556), .Y(n_611) );
OAI21x1_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_558), .B(n_565), .Y(n_556) );
AND2x4_ASAP7_75t_L g566 ( .A(n_567), .B(n_579), .Y(n_566) );
INVx1_ASAP7_75t_L g684 ( .A(n_567), .Y(n_684) );
AND2x2_ASAP7_75t_L g838 ( .A(n_567), .B(n_734), .Y(n_838) );
BUFx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g610 ( .A(n_568), .Y(n_610) );
INVx4_ASAP7_75t_L g649 ( .A(n_568), .Y(n_649) );
AND2x4_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
OAI21x1_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_574), .B(n_578), .Y(n_570) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
AND2x2_ASAP7_75t_L g665 ( .A(n_580), .B(n_648), .Y(n_665) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g702 ( .A(n_581), .B(n_650), .Y(n_702) );
INVx2_ASAP7_75t_L g668 ( .A(n_582), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_582), .B(n_673), .Y(n_836) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_585), .B(n_749), .Y(n_748) );
BUFx2_ASAP7_75t_L g821 ( .A(n_585), .Y(n_821) );
AND2x2_ASAP7_75t_L g835 ( .A(n_585), .B(n_657), .Y(n_835) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_595), .Y(n_585) );
INVx1_ASAP7_75t_L g616 ( .A(n_586), .Y(n_616) );
AND2x2_ASAP7_75t_L g770 ( .A(n_586), .B(n_677), .Y(n_770) );
OR2x2_ASAP7_75t_L g807 ( .A(n_586), .B(n_595), .Y(n_807) );
AND2x2_ASAP7_75t_L g617 ( .A(n_595), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g631 ( .A(n_595), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g677 ( .A(n_595), .Y(n_677) );
OR2x2_ASAP7_75t_L g690 ( .A(n_595), .B(n_630), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_595), .B(n_630), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_612), .B(n_634), .Y(n_602) );
INVxp67_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AOI31xp33_ASAP7_75t_L g680 ( .A1(n_604), .A2(n_681), .A3(n_683), .B(n_686), .Y(n_680) );
OR2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_608), .Y(n_604) );
AND2x2_ASAP7_75t_L g693 ( .A(n_605), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g703 ( .A(n_606), .Y(n_703) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_606), .Y(n_709) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g637 ( .A(n_607), .Y(n_637) );
AND2x2_ASAP7_75t_L g666 ( .A(n_607), .B(n_650), .Y(n_666) );
INVx2_ASAP7_75t_L g716 ( .A(n_607), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_608), .B(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g741 ( .A(n_609), .B(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_L g790 ( .A(n_609), .B(n_791), .Y(n_790) );
AOI33xp33_ASAP7_75t_L g845 ( .A1(n_609), .A2(n_675), .A3(n_685), .B1(n_712), .B2(n_821), .B3(n_846), .Y(n_845) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx2_ASAP7_75t_L g650 ( .A(n_611), .Y(n_650) );
INVx1_ASAP7_75t_L g737 ( .A(n_611), .Y(n_737) );
INVxp67_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_614), .B(n_628), .Y(n_613) );
INVx2_ASAP7_75t_L g645 ( .A(n_614), .Y(n_645) );
AND2x2_ASAP7_75t_L g726 ( .A(n_614), .B(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_617), .Y(n_614) );
INVx1_ASAP7_75t_L g688 ( .A(n_615), .Y(n_688) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g756 ( .A(n_616), .B(n_643), .Y(n_756) );
AND2x2_ASAP7_75t_L g706 ( .A(n_617), .B(n_700), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_617), .B(n_724), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_617), .B(n_756), .Y(n_805) );
AND2x2_ASAP7_75t_L g642 ( .A(n_618), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g661 ( .A(n_618), .B(n_656), .Y(n_661) );
INVx1_ASAP7_75t_L g676 ( .A(n_618), .Y(n_676) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
INVx1_ASAP7_75t_L g731 ( .A(n_629), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_629), .B(n_824), .Y(n_826) );
AND2x2_ASAP7_75t_L g839 ( .A(n_629), .B(n_655), .Y(n_839) );
AND2x2_ASAP7_75t_L g657 ( .A(n_630), .B(n_643), .Y(n_657) );
INVx2_ASAP7_75t_L g639 ( .A(n_631), .Y(n_639) );
AND2x2_ASAP7_75t_L g753 ( .A(n_631), .B(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_L g812 ( .A(n_631), .B(n_724), .Y(n_812) );
BUFx2_ASAP7_75t_L g794 ( .A(n_632), .Y(n_794) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
BUFx3_ASAP7_75t_L g656 ( .A(n_633), .Y(n_656) );
OAI32xp33_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_639), .A3(n_640), .B1(n_645), .B2(n_646), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
INVx2_ASAP7_75t_L g742 ( .A(n_637), .Y(n_742) );
AND2x2_ASAP7_75t_L g772 ( .A(n_637), .B(n_694), .Y(n_772) );
AND2x2_ASAP7_75t_L g714 ( .A(n_638), .B(n_715), .Y(n_714) );
AND3x2_ASAP7_75t_L g721 ( .A(n_638), .B(n_648), .C(n_716), .Y(n_721) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_641), .A2(n_663), .B1(n_672), .B2(n_674), .Y(n_671) );
OAI322xp33_ASAP7_75t_L g819 ( .A1(n_641), .A2(n_740), .A3(n_820), .B1(n_821), .B2(n_822), .C1(n_823), .C2(n_826), .Y(n_819) );
INVx2_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g841 ( .A(n_642), .B(n_824), .Y(n_841) );
INVxp67_ASAP7_75t_SL g660 ( .A(n_643), .Y(n_660) );
INVxp67_ASAP7_75t_SL g700 ( .A(n_643), .Y(n_700) );
BUFx3_ASAP7_75t_L g724 ( .A(n_643), .Y(n_724) );
INVx1_ASAP7_75t_L g750 ( .A(n_643), .Y(n_750) );
INVx1_ASAP7_75t_L g754 ( .A(n_643), .Y(n_754) );
INVx3_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g708 ( .A(n_647), .B(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .Y(n_647) );
INVx1_ASAP7_75t_L g759 ( .A(n_648), .Y(n_759) );
NAND2xp5_ASAP7_75t_SL g810 ( .A(n_648), .B(n_716), .Y(n_810) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2x1_ASAP7_75t_L g669 ( .A(n_649), .B(n_670), .Y(n_669) );
BUFx2_ASAP7_75t_L g673 ( .A(n_649), .Y(n_673) );
AND2x2_ASAP7_75t_L g715 ( .A(n_649), .B(n_716), .Y(n_715) );
OR2x2_ASAP7_75t_L g736 ( .A(n_649), .B(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_650), .B(n_763), .Y(n_820) );
O2A1O1Ixp33_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_658), .B(n_662), .C(n_671), .Y(n_651) );
INVxp67_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AOI31xp33_ASAP7_75t_L g813 ( .A1(n_653), .A2(n_814), .A3(n_816), .B(n_817), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_654), .B(n_657), .Y(n_653) );
AND2x4_ASAP7_75t_L g766 ( .A(n_654), .B(n_675), .Y(n_766) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_655), .Y(n_698) );
INVx3_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NOR2xp67_ASAP7_75t_L g782 ( .A(n_656), .B(n_676), .Y(n_782) );
BUFx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AND2x4_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
NAND2x1_ASAP7_75t_L g662 ( .A(n_663), .B(n_667), .Y(n_662) );
INVx3_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AND2x4_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
INVx1_ASAP7_75t_L g822 ( .A(n_665), .Y(n_822) );
AND2x2_ASAP7_75t_L g682 ( .A(n_666), .B(n_673), .Y(n_682) );
OAI22xp33_ASAP7_75t_L g751 ( .A1(n_667), .A2(n_752), .B1(n_755), .B2(n_757), .Y(n_751) );
OR2x6_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
INVx1_ASAP7_75t_SL g809 ( .A(n_670), .Y(n_809) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g779 ( .A(n_675), .B(n_724), .Y(n_779) );
INVx2_ASAP7_75t_L g825 ( .A(n_675), .Y(n_825) );
AND2x4_ASAP7_75t_L g833 ( .A(n_675), .B(n_754), .Y(n_833) );
AND2x4_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
NAND3xp33_ASAP7_75t_L g678 ( .A(n_679), .B(n_695), .C(n_725), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_680), .B(n_691), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_682), .B(n_812), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
AND2x4_ASAP7_75t_L g746 ( .A(n_684), .B(n_701), .Y(n_746) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_687), .B(n_693), .Y(n_692) );
AND2x4_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
AND2x2_ASAP7_75t_L g777 ( .A(n_689), .B(n_756), .Y(n_777) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_690), .Y(n_697) );
INVx1_ASAP7_75t_L g815 ( .A(n_690), .Y(n_815) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g844 ( .A(n_693), .Y(n_844) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_694), .Y(n_729) );
AOI211xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_701), .B(n_704), .C(n_717), .Y(n_695) );
NOR3x1_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .C(n_699), .Y(n_696) );
NAND2x1_ASAP7_75t_L g765 ( .A(n_699), .B(n_766), .Y(n_765) );
BUFx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NOR2x1p5_ASAP7_75t_SL g701 ( .A(n_702), .B(n_703), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_707), .B1(n_710), .B2(n_713), .Y(n_704) );
INVxp67_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g798 ( .A(n_709), .Y(n_798) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
BUFx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g793 ( .A(n_712), .B(n_794), .Y(n_793) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g847 ( .A(n_715), .Y(n_847) );
AOI21xp33_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_720), .B(n_722), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g801 ( .A(n_722), .Y(n_801) );
OR2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
INVx2_ASAP7_75t_L g728 ( .A(n_724), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_724), .B(n_782), .Y(n_781) );
AOI21xp33_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_729), .B(n_730), .Y(n_725) );
INVxp67_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_728), .B(n_815), .Y(n_814) );
OAI22xp33_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_732), .B1(n_738), .B2(n_740), .Y(n_730) );
OR2x2_ASAP7_75t_L g732 ( .A(n_733), .B(n_736), .Y(n_732) );
INVx1_ASAP7_75t_L g783 ( .A(n_733), .Y(n_783) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g758 ( .A(n_734), .B(n_759), .Y(n_758) );
BUFx2_ASAP7_75t_L g775 ( .A(n_735), .Y(n_775) );
INVx1_ASAP7_75t_L g795 ( .A(n_736), .Y(n_795) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
NOR2x1_ASAP7_75t_L g743 ( .A(n_744), .B(n_799), .Y(n_743) );
NAND3xp33_ASAP7_75t_SL g744 ( .A(n_745), .B(n_760), .C(n_773), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_747), .B(n_751), .Y(n_745) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
OR2x2_ASAP7_75t_L g806 ( .A(n_749), .B(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
NAND2x1p5_ASAP7_75t_L g803 ( .A(n_758), .B(n_786), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_764), .B1(n_767), .B2(n_771), .Y(n_760) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx2_ASAP7_75t_L g816 ( .A(n_766), .Y(n_816) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
OAI21xp33_ASAP7_75t_L g788 ( .A1(n_768), .A2(n_789), .B(n_792), .Y(n_788) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
AOI22xp5_ASAP7_75t_L g773 ( .A1(n_774), .A2(n_784), .B1(n_788), .B2(n_796), .Y(n_773) );
OAI21xp33_ASAP7_75t_L g774 ( .A1(n_775), .A2(n_776), .B(n_778), .Y(n_774) );
INVxp67_ASAP7_75t_SL g776 ( .A(n_777), .Y(n_776) );
OAI21xp5_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_780), .B(n_783), .Y(n_778) );
INVx1_ASAP7_75t_L g843 ( .A(n_779), .Y(n_843) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g832 ( .A(n_782), .Y(n_832) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
BUFx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_793), .B(n_795), .Y(n_792) );
INVx2_ASAP7_75t_L g824 ( .A(n_794), .Y(n_824) );
INVxp67_ASAP7_75t_SL g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_800), .B(n_818), .Y(n_799) );
AOI211xp5_ASAP7_75t_L g800 ( .A1(n_801), .A2(n_802), .B(n_804), .C(n_813), .Y(n_800) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
A2O1A1Ixp33_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_806), .B(n_808), .C(n_811), .Y(n_804) );
OR2x2_ASAP7_75t_L g808 ( .A(n_809), .B(n_810), .Y(n_808) );
NOR3xp33_ASAP7_75t_L g818 ( .A(n_819), .B(n_827), .C(n_842), .Y(n_818) );
OR2x2_ASAP7_75t_L g823 ( .A(n_824), .B(n_825), .Y(n_823) );
OAI221xp5_ASAP7_75t_L g827 ( .A1(n_828), .A2(n_830), .B1(n_834), .B2(n_836), .C(n_837), .Y(n_827) );
NOR2xp67_ASAP7_75t_L g830 ( .A(n_831), .B(n_833), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx2_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_838), .A2(n_839), .B1(n_840), .B2(n_841), .Y(n_837) );
OAI21xp33_ASAP7_75t_SL g842 ( .A1(n_843), .A2(n_844), .B(n_845), .Y(n_842) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
CKINVDCx5p33_ASAP7_75t_R g851 ( .A(n_852), .Y(n_851) );
BUFx12f_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
AND2x6_ASAP7_75t_SL g853 ( .A(n_854), .B(n_856), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx3_ASAP7_75t_L g873 ( .A(n_855), .Y(n_873) );
NOR2xp33_ASAP7_75t_L g875 ( .A(n_855), .B(n_876), .Y(n_875) );
OAI21x1_ASAP7_75t_L g859 ( .A1(n_860), .A2(n_866), .B(n_868), .Y(n_859) );
INVx5_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
BUFx2_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
INVx2_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
BUFx6f_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
CKINVDCx11_ASAP7_75t_R g871 ( .A(n_872), .Y(n_871) );
BUFx6f_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
BUFx10_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
CKINVDCx14_ASAP7_75t_R g879 ( .A(n_880), .Y(n_879) );
endmodule