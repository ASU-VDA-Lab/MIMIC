module fake_jpeg_4521_n_309 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_309);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_309;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_SL g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_38),
.Y(n_59)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_39),
.B(n_44),
.Y(n_85)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_26),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_42),
.B(n_47),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_7),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_22),
.B(n_28),
.Y(n_73)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_0),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_45),
.B(n_32),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_26),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_48),
.A2(n_35),
.B1(n_20),
.B2(n_34),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_52),
.B(n_60),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_21),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_53),
.B(n_66),
.Y(n_112)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_56),
.Y(n_108)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_48),
.A2(n_20),
.B1(n_34),
.B2(n_35),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_58),
.A2(n_17),
.B1(n_16),
.B2(n_18),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_49),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_22),
.C(n_19),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_61),
.A2(n_89),
.B1(n_29),
.B2(n_17),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_20),
.B1(n_35),
.B2(n_34),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_62),
.A2(n_86),
.B1(n_88),
.B2(n_29),
.Y(n_105)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_65),
.Y(n_110)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_21),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_67),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_70),
.Y(n_113)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_73),
.Y(n_114)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_74),
.Y(n_124)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_75),
.B(n_77),
.Y(n_126)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

AND2x4_ASAP7_75t_L g82 ( 
.A(n_36),
.B(n_23),
.Y(n_82)
);

OR2x2_ASAP7_75t_SL g119 ( 
.A(n_82),
.B(n_98),
.Y(n_119)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_39),
.A2(n_24),
.B1(n_32),
.B2(n_30),
.Y(n_89)
);

CKINVDCx12_ASAP7_75t_R g90 ( 
.A(n_41),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_94),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_40),
.B(n_25),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_91),
.B(n_92),
.Y(n_130)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_40),
.B(n_25),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_96),
.Y(n_107)
);

CKINVDCx9p33_ASAP7_75t_R g94 ( 
.A(n_41),
.Y(n_94)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_100),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_41),
.B(n_30),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_36),
.B(n_19),
.Y(n_99)
);

NAND2x1_ASAP7_75t_SL g128 ( 
.A(n_99),
.B(n_33),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_36),
.B(n_24),
.Y(n_100)
);

AO22x1_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_23),
.B1(n_18),
.B2(n_29),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_101),
.A2(n_87),
.B(n_64),
.Y(n_157)
);

OA22x2_ASAP7_75t_L g102 ( 
.A1(n_82),
.A2(n_23),
.B1(n_18),
.B2(n_29),
.Y(n_102)
);

AO22x2_ASAP7_75t_L g133 ( 
.A1(n_102),
.A2(n_81),
.B1(n_83),
.B2(n_94),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_123),
.B1(n_127),
.B2(n_86),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_106),
.A2(n_72),
.B1(n_60),
.B2(n_17),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_61),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_95),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_89),
.A2(n_17),
.B1(n_16),
.B2(n_18),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g125 ( 
.A(n_82),
.B(n_23),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_SL g134 ( 
.A(n_125),
.B(n_83),
.C(n_98),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_58),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_131),
.A2(n_149),
.B1(n_154),
.B2(n_102),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_99),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_135),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_133),
.A2(n_147),
.B1(n_152),
.B2(n_163),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_134),
.A2(n_157),
.B(n_125),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_85),
.Y(n_136)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_136),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_70),
.Y(n_137)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_59),
.Y(n_138)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_138),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_62),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_140),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_68),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_145),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_142),
.A2(n_144),
.B(n_146),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_117),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_143),
.B(n_153),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_18),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_18),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_54),
.B1(n_80),
.B2(n_77),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_156),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_54),
.B1(n_88),
.B2(n_69),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_76),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_150),
.B(n_151),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_68),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_127),
.A2(n_52),
.B1(n_16),
.B2(n_78),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_106),
.A2(n_64),
.B1(n_76),
.B2(n_84),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_155),
.A2(n_166),
.B1(n_120),
.B2(n_118),
.Y(n_189)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_104),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_107),
.B(n_33),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_159),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_107),
.B(n_130),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_160),
.B(n_165),
.Y(n_198)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_104),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_161),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_110),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_164),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_128),
.A2(n_33),
.B1(n_84),
.B2(n_8),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_110),
.B(n_125),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_102),
.A2(n_33),
.B1(n_87),
.B2(n_2),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_167),
.A2(n_146),
.B1(n_133),
.B2(n_157),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_125),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_170),
.A2(n_180),
.B(n_184),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_172),
.A2(n_155),
.B1(n_133),
.B2(n_151),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_102),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_187),
.C(n_188),
.Y(n_205)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_175),
.B(n_185),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_162),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_177),
.B(n_183),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_101),
.B(n_121),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_140),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_101),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_139),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_135),
.B(n_129),
.C(n_124),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_121),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_189),
.A2(n_6),
.B1(n_12),
.B2(n_11),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_129),
.C(n_124),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_200),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_142),
.A2(n_120),
.B1(n_118),
.B2(n_122),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_194),
.A2(n_199),
.B1(n_166),
.B2(n_152),
.Y(n_206)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_195),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_154),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_197),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_142),
.A2(n_122),
.B1(n_111),
.B2(n_103),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_144),
.B(n_121),
.Y(n_200)
);

A2O1A1O1Ixp25_ASAP7_75t_L g201 ( 
.A1(n_167),
.A2(n_144),
.B(n_146),
.C(n_134),
.D(n_133),
.Y(n_201)
);

NOR3xp33_ASAP7_75t_SL g237 ( 
.A(n_201),
.B(n_209),
.C(n_180),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_202),
.A2(n_225),
.B(n_179),
.Y(n_231)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_212),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_210),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_172),
.A2(n_191),
.B1(n_194),
.B2(n_199),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_103),
.C(n_10),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_173),
.A2(n_111),
.B1(n_104),
.B2(n_87),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_215),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_176),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_173),
.B(n_0),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_217),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_0),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_171),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_224),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_191),
.A2(n_116),
.B1(n_1),
.B2(n_2),
.Y(n_219)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_219),
.Y(n_229)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_220),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_190),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_222)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_222),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_169),
.B(n_2),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_196),
.B(n_3),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_213),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_235),
.C(n_240),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_231),
.B(n_232),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_215),
.B(n_168),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_211),
.A2(n_201),
.B1(n_219),
.B2(n_206),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_233),
.A2(n_238),
.B(n_245),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_188),
.C(n_174),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_237),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_223),
.A2(n_170),
.B(n_184),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_169),
.C(n_200),
.Y(n_240)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_246),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_218),
.A2(n_184),
.B1(n_170),
.B2(n_169),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_226),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_189),
.C(n_186),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_208),
.C(n_223),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_229),
.A2(n_227),
.B1(n_242),
.B2(n_239),
.Y(n_250)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_250),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_228),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_254),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_240),
.C(n_233),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_224),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_258),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_203),
.Y(n_256)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_256),
.Y(n_274)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_234),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_230),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_261),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_230),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_210),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_262),
.B(n_242),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_229),
.A2(n_214),
.B(n_216),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_263),
.A2(n_243),
.B(n_231),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_175),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_268),
.C(n_275),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_266),
.A2(n_259),
.B1(n_254),
.B2(n_220),
.Y(n_280)
);

AOI321xp33_ASAP7_75t_L g267 ( 
.A1(n_260),
.A2(n_245),
.A3(n_243),
.B1(n_237),
.B2(n_207),
.C(n_227),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_271),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_247),
.C(n_241),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_241),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_249),
.B(n_181),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_195),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_217),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_272),
.A2(n_261),
.B1(n_255),
.B2(n_258),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_277),
.A2(n_279),
.B(n_280),
.Y(n_296)
);

AOI211xp5_ASAP7_75t_L g278 ( 
.A1(n_267),
.A2(n_248),
.B(n_260),
.C(n_239),
.Y(n_278)
);

AOI322xp5_ASAP7_75t_L g290 ( 
.A1(n_278),
.A2(n_275),
.A3(n_269),
.B1(n_182),
.B2(n_7),
.C1(n_9),
.C2(n_10),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_276),
.A2(n_253),
.B1(n_263),
.B2(n_257),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_204),
.C(n_222),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_14),
.Y(n_294)
);

OAI31xp67_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_225),
.A3(n_198),
.B(n_11),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_283),
.B(n_274),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_285),
.Y(n_292)
);

NAND2xp67_ASAP7_75t_SL g287 ( 
.A(n_270),
.B(n_3),
.Y(n_287)
);

AO21x1_ASAP7_75t_L g293 ( 
.A1(n_287),
.A2(n_182),
.B(n_9),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_288),
.B(n_295),
.Y(n_302)
);

NAND3xp33_ASAP7_75t_L g289 ( 
.A(n_287),
.B(n_265),
.C(n_271),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_289),
.A2(n_290),
.B(n_291),
.Y(n_299)
);

MAJx2_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_269),
.C(n_286),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_293),
.Y(n_298)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_294),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g295 ( 
.A(n_285),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_279),
.B1(n_280),
.B2(n_282),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_300),
.C(n_3),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_281),
.C(n_286),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_300),
.A2(n_288),
.B(n_278),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_304),
.C(n_305),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_299),
.A2(n_14),
.B(n_4),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_305),
.A2(n_301),
.B1(n_298),
.B2(n_297),
.Y(n_306)
);

AOI31xp67_ASAP7_75t_L g308 ( 
.A1(n_306),
.A2(n_302),
.A3(n_14),
.B(n_5),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_307),
.Y(n_309)
);


endmodule