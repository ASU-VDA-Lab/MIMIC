module fake_jpeg_10940_n_19 (n_3, n_2, n_1, n_0, n_4, n_5, n_19);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_19;

wire n_13;
wire n_10;
wire n_6;
wire n_14;
wire n_18;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

BUFx4f_ASAP7_75t_SL g6 ( 
.A(n_0),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_4),
.Y(n_7)
);

INVx5_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_8),
.Y(n_9)
);

XNOR2x1_ASAP7_75t_L g11 ( 
.A(n_9),
.B(n_10),
.Y(n_11)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_9),
.B(n_6),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_12),
.B(n_6),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_11),
.B(n_7),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_L g16 ( 
.A1(n_13),
.A2(n_14),
.B(n_0),
.Y(n_16)
);

INVxp33_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

NOR2xp67_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_16),
.Y(n_17)
);

O2A1O1Ixp33_ASAP7_75t_SL g18 ( 
.A1(n_17),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_18),
.A2(n_1),
.B(n_2),
.Y(n_19)
);


endmodule