module fake_ariane_1747_n_2027 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2027);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2027;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1860;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_330;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_236;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g204 ( 
.A(n_123),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_69),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_159),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_71),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_183),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_117),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_82),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_130),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_28),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_2),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_120),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_129),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_201),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_108),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_48),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_62),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_127),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_74),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_11),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_134),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_65),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_104),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_188),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_142),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_124),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_190),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_55),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_193),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_26),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_40),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_157),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_28),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_122),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_41),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_8),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_137),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_26),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_1),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_148),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_4),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_16),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_113),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_75),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_60),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_9),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_191),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_34),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_30),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_111),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_54),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_69),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_78),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_95),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_165),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_86),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_149),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_170),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_1),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_20),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_187),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_119),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_68),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_109),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_160),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_179),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_63),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_38),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_147),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_24),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_21),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_184),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_155),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_161),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_107),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_162),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_33),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_41),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_143),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_178),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_25),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_48),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_38),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_23),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_169),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_24),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_97),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_0),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_85),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_198),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_136),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_46),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_9),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_15),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_118),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_150),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_37),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_180),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_84),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_98),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_10),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_88),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_7),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_105),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_168),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_2),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_135),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_64),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_23),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_37),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_110),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_42),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_30),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_156),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_5),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_186),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_141),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_83),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_60),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_61),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_93),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_151),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_0),
.Y(n_326)
);

BUFx10_ASAP7_75t_L g327 ( 
.A(n_196),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_43),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_57),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_185),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_52),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_194),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_94),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_154),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_32),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_173),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_56),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_77),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_21),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_39),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_19),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_203),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_4),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_132),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_58),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_56),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_114),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_138),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_13),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_45),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_89),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_43),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_125),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_53),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_46),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_17),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_54),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_200),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_174),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_32),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_199),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_34),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_133),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_139),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_45),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_36),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_126),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_106),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_144),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_19),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_61),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_175),
.Y(n_372)
);

BUFx10_ASAP7_75t_L g373 ( 
.A(n_140),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_42),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_167),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_80),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_18),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_18),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_181),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_112),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_14),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_116),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_177),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_59),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_72),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_121),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_68),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_17),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_202),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_63),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_16),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_11),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_158),
.Y(n_393)
);

BUFx10_ASAP7_75t_L g394 ( 
.A(n_53),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_99),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_90),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_192),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_145),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_131),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_103),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_171),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_81),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_44),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_40),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_39),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_29),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_25),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_49),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_7),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_100),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_6),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_240),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_402),
.B(n_3),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_242),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_242),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_247),
.Y(n_416)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_255),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_317),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_242),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_242),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_242),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_300),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_306),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_322),
.Y(n_424)
);

INVxp67_ASAP7_75t_SL g425 ( 
.A(n_255),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_334),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_251),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_263),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_306),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_331),
.Y(n_430)
);

INVxp67_ASAP7_75t_SL g431 ( 
.A(n_263),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_306),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_306),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_306),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_262),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_284),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_390),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_340),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_390),
.Y(n_439)
);

INVxp67_ASAP7_75t_SL g440 ( 
.A(n_271),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_390),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_327),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_390),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_346),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_266),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_390),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_391),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_391),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_327),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_391),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_270),
.Y(n_451)
);

INVxp33_ASAP7_75t_L g452 ( 
.A(n_212),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_273),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_205),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_285),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_286),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_287),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_391),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_327),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_373),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_391),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_214),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_289),
.Y(n_463)
);

BUFx3_ASAP7_75t_L g464 ( 
.A(n_214),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_315),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_291),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_295),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_315),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_373),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_296),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_377),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_377),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_407),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_407),
.Y(n_474)
);

NOR2xp67_ASAP7_75t_L g475 ( 
.A(n_339),
.B(n_3),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_257),
.Y(n_476)
);

NOR2xp67_ASAP7_75t_L g477 ( 
.A(n_339),
.B(n_5),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_257),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_282),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_373),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_282),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_297),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_304),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_394),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_290),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_204),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_271),
.B(n_6),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_316),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_290),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_318),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_394),
.Y(n_491)
);

INVxp33_ASAP7_75t_SL g492 ( 
.A(n_411),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_321),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_335),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_394),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_321),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_336),
.Y(n_497)
);

INVxp33_ASAP7_75t_L g498 ( 
.A(n_225),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_205),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_213),
.Y(n_500)
);

NOR2xp67_ASAP7_75t_L g501 ( 
.A(n_223),
.B(n_8),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_213),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_231),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_336),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_352),
.B(n_10),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_337),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_219),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_215),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_352),
.Y(n_509)
);

NAND2xp33_ASAP7_75t_R g510 ( 
.A(n_206),
.B(n_73),
.Y(n_510)
);

NOR2xp67_ASAP7_75t_L g511 ( 
.A(n_280),
.B(n_12),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_343),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_349),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_219),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_363),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_220),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_363),
.Y(n_517)
);

INVxp67_ASAP7_75t_SL g518 ( 
.A(n_370),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_410),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_370),
.Y(n_520)
);

BUFx8_ASAP7_75t_L g521 ( 
.A(n_509),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_462),
.B(n_218),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_437),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_437),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_437),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_437),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_486),
.B(n_234),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_462),
.B(n_232),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_414),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_414),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_423),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_415),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_423),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_415),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_508),
.B(n_237),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_419),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_505),
.B(n_217),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_433),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_433),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_419),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_461),
.Y(n_541)
);

AND2x6_ASAP7_75t_L g542 ( 
.A(n_505),
.B(n_230),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_430),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_413),
.B(n_410),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_461),
.Y(n_545)
);

AND3x2_ASAP7_75t_L g546 ( 
.A(n_422),
.B(n_241),
.C(n_238),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_508),
.B(n_256),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_420),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_420),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_421),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_421),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_475),
.B(n_217),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_429),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_486),
.B(n_245),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_429),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_432),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_464),
.B(n_226),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_509),
.B(n_248),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_520),
.B(n_274),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_432),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_434),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_434),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_439),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_439),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_508),
.B(n_259),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_441),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_464),
.B(n_260),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_499),
.A2(n_411),
.B1(n_409),
.B2(n_254),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_441),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_443),
.Y(n_570)
);

BUFx8_ASAP7_75t_L g571 ( 
.A(n_520),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_SL g572 ( 
.A1(n_427),
.A2(n_409),
.B1(n_220),
.B2(n_406),
.Y(n_572)
);

NAND2xp33_ASAP7_75t_SL g573 ( 
.A(n_452),
.B(n_233),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_464),
.B(n_261),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_443),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_446),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_498),
.B(n_281),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_446),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_447),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_447),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_448),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_448),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_450),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_450),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_458),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_458),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_417),
.B(n_226),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_476),
.B(n_275),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_476),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_478),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_478),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_479),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_479),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_475),
.B(n_229),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_481),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_481),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_485),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_485),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_489),
.Y(n_599)
);

OA21x2_ASAP7_75t_L g600 ( 
.A1(n_489),
.A2(n_292),
.B(n_288),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_425),
.B(n_309),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_477),
.B(n_229),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_493),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_428),
.B(n_431),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_519),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_519),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_493),
.B(n_293),
.Y(n_607)
);

INVx4_ASAP7_75t_L g608 ( 
.A(n_542),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_557),
.B(n_435),
.Y(n_609)
);

INVxp67_ASAP7_75t_SL g610 ( 
.A(n_522),
.Y(n_610)
);

INVx5_ASAP7_75t_L g611 ( 
.A(n_542),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_604),
.B(n_440),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_604),
.B(n_445),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_529),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_557),
.B(n_451),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_542),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_529),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_530),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_604),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_577),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_524),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_544),
.B(n_492),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_521),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_524),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_577),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_596),
.Y(n_626)
);

AND2x6_ASAP7_75t_L g627 ( 
.A(n_537),
.B(n_230),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_524),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_525),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_530),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_521),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_527),
.B(n_518),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_544),
.B(n_453),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_526),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_537),
.A2(n_573),
.B1(n_577),
.B2(n_542),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_526),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_573),
.A2(n_510),
.B1(n_455),
.B2(n_457),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_532),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_526),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_532),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_587),
.B(n_456),
.Y(n_641)
);

BUFx4f_ASAP7_75t_L g642 ( 
.A(n_542),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_525),
.Y(n_643)
);

CKINVDCx16_ASAP7_75t_R g644 ( 
.A(n_543),
.Y(n_644)
);

XNOR2xp5_ASAP7_75t_L g645 ( 
.A(n_572),
.B(n_436),
.Y(n_645)
);

OR2x6_ASAP7_75t_L g646 ( 
.A(n_572),
.B(n_477),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_596),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_525),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_587),
.B(n_463),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_603),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_601),
.A2(n_466),
.B1(n_470),
.B2(n_467),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_603),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_523),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_537),
.B(n_482),
.Y(n_654)
);

INVx8_ASAP7_75t_L g655 ( 
.A(n_542),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_603),
.Y(n_656)
);

OAI21xp33_ASAP7_75t_SL g657 ( 
.A1(n_552),
.A2(n_511),
.B(n_501),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_537),
.A2(n_422),
.B1(n_444),
.B2(n_487),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_537),
.B(n_483),
.Y(n_659)
);

CKINVDCx6p67_ASAP7_75t_R g660 ( 
.A(n_543),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_592),
.Y(n_661)
);

AND2x6_ASAP7_75t_L g662 ( 
.A(n_601),
.B(n_230),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_601),
.B(n_488),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_592),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_552),
.B(n_490),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_594),
.B(n_494),
.Y(n_666)
);

BUFx2_ASAP7_75t_L g667 ( 
.A(n_521),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_523),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_523),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_542),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_523),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_590),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_527),
.B(n_454),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_594),
.B(n_506),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_558),
.B(n_512),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_523),
.Y(n_676)
);

XOR2xp5_ASAP7_75t_SL g677 ( 
.A(n_521),
.B(n_500),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_590),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_527),
.B(n_503),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_602),
.B(n_513),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_602),
.B(n_424),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_521),
.Y(n_682)
);

INVx5_ASAP7_75t_L g683 ( 
.A(n_542),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_549),
.Y(n_684)
);

BUFx3_ASAP7_75t_L g685 ( 
.A(n_542),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_526),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_593),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_549),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_567),
.B(n_496),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_567),
.B(n_496),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_549),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_549),
.Y(n_692)
);

INVx5_ASAP7_75t_L g693 ( 
.A(n_542),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_574),
.B(n_589),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_549),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_554),
.B(n_502),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_558),
.B(n_507),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_534),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_534),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_558),
.B(n_426),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_589),
.Y(n_701)
);

BUFx10_ASAP7_75t_L g702 ( 
.A(n_546),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_600),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_555),
.Y(n_704)
);

NAND2xp33_ASAP7_75t_L g705 ( 
.A(n_526),
.B(n_230),
.Y(n_705)
);

BUFx4f_ASAP7_75t_L g706 ( 
.A(n_600),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_559),
.B(n_206),
.Y(n_707)
);

BUFx10_ASAP7_75t_L g708 ( 
.A(n_546),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_589),
.B(n_591),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_555),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_559),
.B(n_207),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_536),
.Y(n_712)
);

OR2x6_ASAP7_75t_L g713 ( 
.A(n_554),
.B(n_501),
.Y(n_713)
);

INVx5_ASAP7_75t_L g714 ( 
.A(n_526),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_555),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_555),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_536),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_555),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_SL g719 ( 
.A(n_571),
.B(n_442),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_581),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_526),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_535),
.B(n_449),
.Y(n_722)
);

INVxp67_ASAP7_75t_L g723 ( 
.A(n_568),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_593),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_540),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_589),
.B(n_497),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_559),
.B(n_207),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_581),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_581),
.Y(n_729)
);

NAND2xp33_ASAP7_75t_SL g730 ( 
.A(n_535),
.B(n_459),
.Y(n_730)
);

NAND3xp33_ASAP7_75t_L g731 ( 
.A(n_547),
.B(n_236),
.C(n_233),
.Y(n_731)
);

INVx4_ASAP7_75t_L g732 ( 
.A(n_600),
.Y(n_732)
);

BUFx2_ASAP7_75t_L g733 ( 
.A(n_571),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_547),
.B(n_460),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_571),
.B(n_208),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_590),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_565),
.B(n_469),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_568),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_581),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_540),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_565),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_571),
.B(n_208),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_581),
.Y(n_743)
);

INVx4_ASAP7_75t_L g744 ( 
.A(n_600),
.Y(n_744)
);

BUFx10_ASAP7_75t_L g745 ( 
.A(n_595),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_548),
.Y(n_746)
);

NAND2xp33_ASAP7_75t_R g747 ( 
.A(n_600),
.B(n_480),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_589),
.B(n_591),
.Y(n_748)
);

AND2x6_ASAP7_75t_L g749 ( 
.A(n_554),
.B(n_230),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_591),
.B(n_465),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_591),
.B(n_504),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_526),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_591),
.Y(n_753)
);

BUFx6f_ASAP7_75t_SL g754 ( 
.A(n_571),
.Y(n_754)
);

INVx8_ASAP7_75t_L g755 ( 
.A(n_590),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_588),
.B(n_209),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_642),
.B(n_590),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_641),
.B(n_522),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_621),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_614),
.Y(n_760)
);

OAI22xp33_ASAP7_75t_L g761 ( 
.A1(n_723),
.A2(n_511),
.B1(n_516),
.B2(n_514),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_621),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_637),
.B(n_209),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_651),
.B(n_210),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_622),
.A2(n_599),
.B1(n_595),
.B2(n_600),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_624),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_619),
.A2(n_599),
.B1(n_211),
.B2(n_216),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_738),
.A2(n_597),
.B1(n_605),
.B2(n_598),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_619),
.A2(n_597),
.B1(n_605),
.B2(n_598),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_610),
.B(n_528),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_624),
.Y(n_771)
);

INVxp33_ASAP7_75t_L g772 ( 
.A(n_645),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_670),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_741),
.B(n_528),
.Y(n_774)
);

OAI22xp33_ASAP7_75t_L g775 ( 
.A1(n_646),
.A2(n_328),
.B1(n_312),
.B2(n_239),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_614),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_694),
.A2(n_748),
.B(n_709),
.Y(n_777)
);

CKINVDCx20_ASAP7_75t_R g778 ( 
.A(n_644),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_609),
.B(n_597),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_615),
.B(n_598),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_628),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_649),
.B(n_605),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_629),
.Y(n_783)
);

INVxp67_ASAP7_75t_SL g784 ( 
.A(n_670),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_617),
.Y(n_785)
);

INVxp67_ASAP7_75t_SL g786 ( 
.A(n_685),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_629),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_612),
.B(n_722),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_612),
.B(n_606),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_612),
.B(n_606),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_617),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_613),
.B(n_588),
.Y(n_792)
);

INVxp67_ASAP7_75t_L g793 ( 
.A(n_734),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_737),
.B(n_620),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_642),
.B(n_590),
.Y(n_795)
);

INVxp67_ASAP7_75t_L g796 ( 
.A(n_700),
.Y(n_796)
);

AOI22xp5_ASAP7_75t_L g797 ( 
.A1(n_633),
.A2(n_211),
.B1(n_216),
.B2(n_210),
.Y(n_797)
);

OR2x2_ASAP7_75t_L g798 ( 
.A(n_660),
.B(n_412),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_620),
.B(n_606),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_642),
.B(n_590),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_625),
.B(n_607),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_643),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_625),
.B(n_607),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_643),
.Y(n_804)
);

NAND2xp33_ASAP7_75t_L g805 ( 
.A(n_655),
.B(n_221),
.Y(n_805)
);

INVx6_ASAP7_75t_L g806 ( 
.A(n_745),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_667),
.B(n_416),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_685),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_660),
.B(n_484),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_618),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_654),
.B(n_659),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_663),
.B(n_350),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_702),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_648),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_745),
.Y(n_815)
);

BUFx6f_ASAP7_75t_SL g816 ( 
.A(n_702),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_648),
.Y(n_817)
);

BUFx6f_ASAP7_75t_SL g818 ( 
.A(n_702),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_666),
.B(n_680),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_635),
.B(n_590),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_SL g821 ( 
.A(n_754),
.B(n_418),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_608),
.B(n_222),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_632),
.B(n_504),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_679),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_618),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_675),
.B(n_665),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_674),
.B(n_354),
.Y(n_827)
);

INVxp67_ASAP7_75t_SL g828 ( 
.A(n_703),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_679),
.Y(n_829)
);

INVxp67_ASAP7_75t_L g830 ( 
.A(n_681),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_608),
.B(n_222),
.Y(n_831)
);

NAND3xp33_ASAP7_75t_L g832 ( 
.A(n_658),
.B(n_239),
.C(n_236),
.Y(n_832)
);

HB1xp67_ASAP7_75t_L g833 ( 
.A(n_679),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_632),
.B(n_515),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_707),
.B(n_355),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_689),
.B(n_515),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_690),
.B(n_517),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_645),
.Y(n_838)
);

NOR2xp67_ASAP7_75t_L g839 ( 
.A(n_623),
.B(n_517),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_630),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_638),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_750),
.B(n_550),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_638),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_750),
.B(n_553),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_661),
.B(n_553),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_640),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_746),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_746),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_664),
.B(n_556),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_655),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_608),
.B(n_224),
.Y(n_851)
);

NAND3xp33_ASAP7_75t_L g852 ( 
.A(n_731),
.B(n_249),
.C(n_244),
.Y(n_852)
);

INVx2_ASAP7_75t_SL g853 ( 
.A(n_708),
.Y(n_853)
);

NAND2xp33_ASAP7_75t_L g854 ( 
.A(n_655),
.B(n_224),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_698),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_687),
.B(n_556),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_711),
.B(n_356),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_719),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_708),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_673),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_727),
.B(n_756),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_713),
.A2(n_228),
.B1(n_235),
.B2(n_227),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_755),
.A2(n_563),
.B(n_560),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_684),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_698),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_701),
.B(n_753),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_655),
.Y(n_867)
);

NOR3xp33_ASAP7_75t_L g868 ( 
.A(n_697),
.B(n_313),
.C(n_311),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_616),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_684),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_708),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_724),
.B(n_560),
.Y(n_872)
);

INVxp67_ASAP7_75t_L g873 ( 
.A(n_673),
.Y(n_873)
);

NOR2xp67_ASAP7_75t_SL g874 ( 
.A(n_611),
.B(n_244),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_616),
.B(n_227),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_701),
.B(n_357),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_616),
.B(n_228),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_672),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_696),
.B(n_491),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_699),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_688),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_753),
.B(n_362),
.Y(n_882)
);

INVxp33_ASAP7_75t_L g883 ( 
.A(n_696),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_699),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_662),
.B(n_563),
.Y(n_885)
);

OAI221xp5_ASAP7_75t_L g886 ( 
.A1(n_646),
.A2(n_392),
.B1(n_323),
.B2(n_326),
.C(n_329),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_706),
.B(n_235),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_688),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_623),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_713),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_713),
.Y(n_891)
);

AND2x6_ASAP7_75t_SL g892 ( 
.A(n_646),
.B(n_341),
.Y(n_892)
);

NOR3xp33_ASAP7_75t_L g893 ( 
.A(n_657),
.B(n_360),
.C(n_345),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_667),
.B(n_495),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_713),
.A2(n_253),
.B1(n_246),
.B2(n_243),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_706),
.A2(n_586),
.B(n_585),
.C(n_566),
.Y(n_896)
);

NAND3x1_ASAP7_75t_L g897 ( 
.A(n_677),
.B(n_438),
.C(n_371),
.Y(n_897)
);

NOR2x1p5_ASAP7_75t_L g898 ( 
.A(n_631),
.B(n_249),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_662),
.B(n_566),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_691),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_652),
.B(n_366),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_652),
.B(n_243),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_662),
.B(n_569),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_631),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_656),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_656),
.B(n_246),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_662),
.B(n_569),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_735),
.B(n_252),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_742),
.B(n_252),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_712),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_691),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_626),
.B(n_254),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_733),
.B(n_253),
.Y(n_913)
);

OAI22xp5_ASAP7_75t_L g914 ( 
.A1(n_647),
.A2(n_374),
.B1(n_381),
.B2(n_406),
.Y(n_914)
);

INVxp33_ASAP7_75t_L g915 ( 
.A(n_733),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_662),
.B(n_570),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_692),
.Y(n_917)
);

NAND2x1_ASAP7_75t_L g918 ( 
.A(n_634),
.B(n_586),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_611),
.B(n_683),
.Y(n_919)
);

INVx4_ASAP7_75t_L g920 ( 
.A(n_611),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_662),
.B(n_570),
.Y(n_921)
);

INVx4_ASAP7_75t_L g922 ( 
.A(n_611),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_819),
.B(n_682),
.Y(n_923)
);

O2A1O1Ixp5_ASAP7_75t_L g924 ( 
.A1(n_819),
.A2(n_717),
.B(n_725),
.C(n_712),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_850),
.Y(n_925)
);

OAI321xp33_ASAP7_75t_L g926 ( 
.A1(n_886),
.A2(n_646),
.A3(n_365),
.B1(n_408),
.B2(n_387),
.C(n_468),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_779),
.A2(n_703),
.B(n_755),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_780),
.A2(n_755),
.B(n_650),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_777),
.A2(n_755),
.B(n_636),
.Y(n_929)
);

OR2x2_ASAP7_75t_L g930 ( 
.A(n_860),
.B(n_879),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_758),
.B(n_811),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_758),
.B(n_682),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_883),
.B(n_465),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_811),
.A2(n_725),
.B1(n_740),
.B2(n_717),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_850),
.Y(n_935)
);

OAI22xp5_ASAP7_75t_L g936 ( 
.A1(n_760),
.A2(n_785),
.B1(n_791),
.B2(n_776),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_850),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_782),
.A2(n_636),
.B(n_634),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_828),
.A2(n_887),
.B(n_795),
.Y(n_939)
);

NAND2x1p5_ASAP7_75t_L g940 ( 
.A(n_773),
.B(n_611),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_887),
.A2(n_795),
.B(n_757),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_869),
.B(n_672),
.Y(n_942)
);

INVx1_ASAP7_75t_SL g943 ( 
.A(n_778),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_896),
.A2(n_744),
.B(n_732),
.Y(n_944)
);

NOR2xp67_ASAP7_75t_L g945 ( 
.A(n_830),
.B(n_726),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_788),
.B(n_754),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_800),
.A2(n_686),
.B(n_639),
.Y(n_947)
);

O2A1O1Ixp5_ASAP7_75t_L g948 ( 
.A1(n_822),
.A2(n_740),
.B(n_744),
.C(n_732),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_864),
.A2(n_686),
.B(n_639),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_864),
.A2(n_752),
.B(n_721),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_794),
.B(n_627),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_870),
.A2(n_752),
.B(n_721),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_850),
.Y(n_953)
);

AOI21xp33_ASAP7_75t_L g954 ( 
.A1(n_908),
.A2(n_747),
.B(n_909),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_810),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_870),
.A2(n_752),
.B(n_721),
.Y(n_956)
);

OAI21xp5_ASAP7_75t_L g957 ( 
.A1(n_765),
.A2(n_744),
.B(n_732),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_792),
.B(n_627),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_881),
.A2(n_695),
.B(n_692),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_869),
.B(n_672),
.Y(n_960)
);

NAND2xp33_ASAP7_75t_SL g961 ( 
.A(n_815),
.B(n_754),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_792),
.B(n_627),
.Y(n_962)
);

A2O1A1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_826),
.A2(n_715),
.B(n_743),
.C(n_739),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_L g964 ( 
.A1(n_825),
.A2(n_653),
.B1(n_676),
.B2(n_669),
.Y(n_964)
);

BUFx8_ASAP7_75t_L g965 ( 
.A(n_816),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_869),
.B(n_672),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_888),
.A2(n_710),
.B(n_704),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_873),
.A2(n_751),
.B(n_671),
.C(n_676),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_824),
.B(n_468),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_829),
.B(n_471),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_815),
.B(n_826),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_840),
.A2(n_653),
.B1(n_671),
.B2(n_669),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_847),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_869),
.B(n_889),
.Y(n_974)
);

AOI21xp33_ASAP7_75t_L g975 ( 
.A1(n_908),
.A2(n_668),
.B(n_710),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_L g976 ( 
.A1(n_841),
.A2(n_668),
.B1(n_743),
.B2(n_739),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_796),
.B(n_730),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_867),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_867),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_774),
.B(n_627),
.Y(n_980)
);

O2A1O1Ixp5_ASAP7_75t_L g981 ( 
.A1(n_822),
.A2(n_718),
.B(n_715),
.C(n_716),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_833),
.B(n_730),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_888),
.A2(n_718),
.B(n_716),
.Y(n_983)
);

AND2x2_ASAP7_75t_SL g984 ( 
.A(n_805),
.B(n_677),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_801),
.B(n_720),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_L g986 ( 
.A1(n_832),
.A2(n_627),
.B1(n_749),
.B2(n_585),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_803),
.B(n_627),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_867),
.B(n_672),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_842),
.A2(n_728),
.B(n_729),
.C(n_575),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_770),
.B(n_729),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_900),
.A2(n_736),
.B(n_678),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_823),
.B(n_749),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_911),
.A2(n_917),
.B(n_875),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_843),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_834),
.B(n_749),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_L g996 ( 
.A1(n_911),
.A2(n_714),
.B(n_693),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_917),
.A2(n_736),
.B(n_678),
.Y(n_997)
);

O2A1O1Ixp5_ASAP7_75t_L g998 ( 
.A1(n_831),
.A2(n_583),
.B(n_576),
.C(n_580),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_863),
.A2(n_714),
.B(n_693),
.Y(n_999)
);

CKINVDCx8_ASAP7_75t_R g1000 ( 
.A(n_807),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_789),
.B(n_749),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_894),
.B(n_471),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_831),
.A2(n_736),
.B(n_678),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_844),
.A2(n_576),
.B(n_580),
.C(n_583),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_861),
.B(n_678),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_875),
.A2(n_736),
.B(n_714),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_773),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_827),
.A2(n_736),
.B(n_298),
.C(n_364),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_827),
.A2(n_302),
.B(n_395),
.C(n_398),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_790),
.B(n_749),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_861),
.B(n_374),
.Y(n_1011)
);

BUFx2_ASAP7_75t_L g1012 ( 
.A(n_904),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_876),
.B(n_683),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_891),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_882),
.B(n_683),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_909),
.A2(n_332),
.B(n_342),
.C(n_347),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_847),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_878),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_915),
.B(n_378),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_848),
.A2(n_855),
.B(n_846),
.Y(n_1020)
);

BUFx8_ASAP7_75t_SL g1021 ( 
.A(n_816),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_848),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_865),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_882),
.B(n_683),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_877),
.A2(n_714),
.B(n_693),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_877),
.A2(n_714),
.B(n_693),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_808),
.B(n_683),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_901),
.B(n_378),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_878),
.B(n_368),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_880),
.B(n_381),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_884),
.B(n_384),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_759),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_808),
.B(n_368),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_910),
.A2(n_705),
.B(n_582),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_806),
.A2(n_388),
.B1(n_384),
.B2(n_403),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_851),
.A2(n_375),
.B(n_372),
.Y(n_1036)
);

BUFx4f_ASAP7_75t_L g1037 ( 
.A(n_806),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_866),
.A2(n_382),
.B(n_375),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_806),
.B(n_388),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_878),
.B(n_382),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_878),
.B(n_383),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_799),
.B(n_403),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_768),
.B(n_404),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_761),
.B(n_404),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_807),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_866),
.A2(n_385),
.B(n_383),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_768),
.B(n_405),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_918),
.A2(n_385),
.B(n_386),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_845),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_797),
.A2(n_405),
.B1(n_301),
.B2(n_307),
.Y(n_1050)
);

AOI21x1_ASAP7_75t_L g1051 ( 
.A1(n_820),
.A2(n_548),
.B(n_579),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_798),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_849),
.A2(n_389),
.B(n_393),
.Y(n_1053)
);

INVxp67_ASAP7_75t_SL g1054 ( 
.A(n_784),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_835),
.A2(n_401),
.B(n_380),
.C(n_310),
.Y(n_1055)
);

CKINVDCx8_ASAP7_75t_R g1056 ( 
.A(n_892),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_905),
.B(n_393),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_813),
.B(n_396),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_905),
.B(n_396),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_856),
.A2(n_397),
.B(n_399),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_872),
.A2(n_854),
.B(n_762),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_839),
.B(n_397),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_862),
.B(n_399),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_853),
.B(n_400),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_859),
.B(n_541),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_809),
.Y(n_1066)
);

AO21x1_ASAP7_75t_L g1067 ( 
.A1(n_836),
.A2(n_379),
.B(n_369),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_766),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_871),
.B(n_541),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_912),
.B(n_541),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_786),
.A2(n_376),
.B1(n_278),
.B2(n_308),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_766),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_890),
.B(n_250),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_771),
.A2(n_344),
.B(n_264),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_771),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_812),
.B(n_283),
.Y(n_1076)
);

AOI21x1_ASAP7_75t_L g1077 ( 
.A1(n_885),
.A2(n_548),
.B(n_579),
.Y(n_1077)
);

O2A1O1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_764),
.A2(n_584),
.B(n_562),
.C(n_561),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_781),
.A2(n_348),
.B(n_265),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_898),
.B(n_472),
.Y(n_1080)
);

AOI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_835),
.A2(n_353),
.B1(n_267),
.B2(n_268),
.Y(n_1081)
);

OAI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_781),
.A2(n_584),
.B(n_562),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_783),
.A2(n_802),
.B(n_787),
.Y(n_1083)
);

INVx4_ASAP7_75t_L g1084 ( 
.A(n_818),
.Y(n_1084)
);

AOI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_857),
.A2(n_258),
.B1(n_269),
.B2(n_272),
.Y(n_1085)
);

AO21x1_ASAP7_75t_L g1086 ( 
.A1(n_837),
.A2(n_584),
.B(n_561),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_787),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_912),
.B(n_541),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_802),
.A2(n_814),
.B(n_817),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_812),
.B(n_12),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_804),
.A2(n_358),
.B(n_277),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_804),
.A2(n_359),
.B(n_279),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_814),
.A2(n_817),
.B(n_902),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_769),
.B(n_541),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_899),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_821),
.B(n_472),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_895),
.B(n_551),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_965),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_1037),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_1002),
.B(n_772),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_931),
.B(n_893),
.Y(n_1101)
);

NAND3xp33_ASAP7_75t_SL g1102 ( 
.A(n_1090),
.B(n_857),
.C(n_767),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_925),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_934),
.A2(n_906),
.B(n_913),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_955),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_1084),
.B(n_858),
.Y(n_1106)
);

NOR2x1_ASAP7_75t_R g1107 ( 
.A(n_1012),
.B(n_838),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_932),
.B(n_775),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_925),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_973),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_1090),
.A2(n_852),
.B1(n_763),
.B2(n_897),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_930),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1049),
.B(n_868),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_923),
.B(n_818),
.Y(n_1114)
);

INVx2_ASAP7_75t_SL g1115 ( 
.A(n_1037),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1011),
.A2(n_907),
.B1(n_921),
.B2(n_903),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_927),
.A2(n_929),
.B(n_990),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_994),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1011),
.A2(n_916),
.B1(n_914),
.B2(n_561),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1017),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_1028),
.A2(n_474),
.B(n_473),
.C(n_562),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_965),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_985),
.B(n_920),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1022),
.Y(n_1124)
);

AOI22xp33_ASAP7_75t_L g1125 ( 
.A1(n_954),
.A2(n_922),
.B1(n_920),
.B2(n_473),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_936),
.A2(n_474),
.B1(n_545),
.B2(n_539),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_1076),
.B(n_874),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_1076),
.B(n_276),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_1014),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1023),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_985),
.B(n_922),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_925),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_1021),
.Y(n_1133)
);

INVx2_ASAP7_75t_SL g1134 ( 
.A(n_1084),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_943),
.Y(n_1135)
);

AND2x6_ASAP7_75t_L g1136 ( 
.A(n_925),
.B(n_338),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_1050),
.A2(n_545),
.B(n_539),
.C(n_919),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_1009),
.A2(n_545),
.B1(n_564),
.B2(n_551),
.Y(n_1138)
);

NAND3xp33_ASAP7_75t_L g1139 ( 
.A(n_1044),
.B(n_578),
.C(n_564),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_941),
.A2(n_333),
.B(n_299),
.Y(n_1140)
);

AOI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1044),
.A2(n_294),
.B1(n_303),
.B2(n_305),
.Y(n_1141)
);

OR2x6_ASAP7_75t_L g1142 ( 
.A(n_1045),
.B(n_545),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_977),
.B(n_314),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_1000),
.Y(n_1144)
);

AND2x2_ASAP7_75t_SL g1145 ( 
.A(n_984),
.B(n_338),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_926),
.B(n_319),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_977),
.B(n_971),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_939),
.A2(n_361),
.B(n_324),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1032),
.Y(n_1149)
);

AND2x4_ASAP7_75t_SL g1150 ( 
.A(n_1014),
.B(n_531),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1068),
.Y(n_1151)
);

OA21x2_ASAP7_75t_L g1152 ( 
.A1(n_1086),
.A2(n_367),
.B(n_325),
.Y(n_1152)
);

INVx1_ASAP7_75t_SL g1153 ( 
.A(n_1066),
.Y(n_1153)
);

INVx4_ASAP7_75t_L g1154 ( 
.A(n_935),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1061),
.A2(n_320),
.B(n_330),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_969),
.B(n_531),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_938),
.A2(n_338),
.B(n_351),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1016),
.A2(n_578),
.B1(n_564),
.B2(n_551),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_SL g1159 ( 
.A(n_1056),
.B(n_531),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1005),
.B(n_551),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1072),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_957),
.A2(n_338),
.B(n_351),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_945),
.B(n_578),
.Y(n_1163)
);

AOI33xp33_ASAP7_75t_L g1164 ( 
.A1(n_1080),
.A2(n_13),
.A3(n_14),
.B1(n_15),
.B2(n_20),
.B3(n_22),
.Y(n_1164)
);

NOR3xp33_ASAP7_75t_L g1165 ( 
.A(n_1063),
.B(n_22),
.C(n_27),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1054),
.B(n_578),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_SL g1167 ( 
.A(n_984),
.B(n_533),
.Y(n_1167)
);

OAI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_944),
.A2(n_578),
.B(n_564),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1013),
.A2(n_338),
.B(n_351),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_970),
.B(n_538),
.Y(n_1170)
);

NOR2xp67_ASAP7_75t_L g1171 ( 
.A(n_1039),
.B(n_101),
.Y(n_1171)
);

CKINVDCx20_ASAP7_75t_R g1172 ( 
.A(n_1052),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_933),
.B(n_531),
.Y(n_1173)
);

OR2x2_ASAP7_75t_L g1174 ( 
.A(n_1030),
.B(n_538),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1015),
.A2(n_351),
.B(n_564),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1054),
.B(n_578),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_982),
.B(n_27),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1024),
.A2(n_351),
.B(n_564),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_928),
.A2(n_578),
.B(n_564),
.Y(n_1179)
);

OAI21xp33_ASAP7_75t_L g1180 ( 
.A1(n_1081),
.A2(n_578),
.B(n_551),
.Y(n_1180)
);

NAND3xp33_ASAP7_75t_L g1181 ( 
.A(n_1055),
.B(n_551),
.C(n_538),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_SL g1182 ( 
.A1(n_989),
.A2(n_29),
.B(n_31),
.C(n_33),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1020),
.A2(n_538),
.B1(n_533),
.B2(n_531),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1042),
.A2(n_31),
.B(n_35),
.C(n_36),
.Y(n_1184)
);

OAI22x1_ASAP7_75t_L g1185 ( 
.A1(n_982),
.A2(n_35),
.B1(n_44),
.B2(n_47),
.Y(n_1185)
);

AOI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1019),
.A2(n_538),
.B1(n_533),
.B2(n_531),
.Y(n_1186)
);

INVx1_ASAP7_75t_SL g1187 ( 
.A(n_1096),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1035),
.B(n_47),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_946),
.B(n_538),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1051),
.A2(n_538),
.B(n_533),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1075),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1073),
.B(n_531),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1007),
.B(n_49),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1058),
.B(n_50),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1007),
.B(n_50),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_974),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1043),
.A2(n_51),
.B1(n_52),
.B2(n_55),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1064),
.B(n_51),
.Y(n_1198)
);

AOI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1077),
.A2(n_115),
.B(n_189),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1073),
.B(n_57),
.Y(n_1200)
);

O2A1O1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1031),
.A2(n_58),
.B(n_59),
.C(n_62),
.Y(n_1201)
);

OAI21xp33_ASAP7_75t_SL g1202 ( 
.A1(n_1057),
.A2(n_1059),
.B(n_958),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_935),
.B(n_64),
.Y(n_1203)
);

AOI221xp5_ASAP7_75t_L g1204 ( 
.A1(n_1047),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.C(n_70),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_1018),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_937),
.B(n_66),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_947),
.A2(n_950),
.B(n_949),
.Y(n_1207)
);

INVx2_ASAP7_75t_SL g1208 ( 
.A(n_1018),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1071),
.B(n_67),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_1018),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_952),
.A2(n_146),
.B(n_76),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1087),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_956),
.A2(n_152),
.B(n_79),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_962),
.B(n_70),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_924),
.A2(n_87),
.B(n_91),
.C(n_92),
.Y(n_1215)
);

O2A1O1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_1008),
.A2(n_96),
.B(n_102),
.C(n_128),
.Y(n_1216)
);

O2A1O1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1057),
.A2(n_153),
.B(n_163),
.C(n_164),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1095),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1085),
.B(n_197),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1094),
.Y(n_1220)
);

AOI21x1_ASAP7_75t_L g1221 ( 
.A1(n_993),
.A2(n_166),
.B(n_172),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_980),
.B(n_176),
.Y(n_1222)
);

OAI21xp33_ASAP7_75t_L g1223 ( 
.A1(n_1038),
.A2(n_182),
.B(n_1046),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1065),
.Y(n_1224)
);

BUFx4f_ASAP7_75t_L g1225 ( 
.A(n_935),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_963),
.B(n_987),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1070),
.A2(n_1088),
.B1(n_951),
.B2(n_976),
.Y(n_1227)
);

INVx4_ASAP7_75t_L g1228 ( 
.A(n_935),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_SL g1229 ( 
.A1(n_986),
.A2(n_1069),
.B1(n_1018),
.B2(n_992),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1059),
.B(n_1062),
.Y(n_1230)
);

AO22x1_ASAP7_75t_L g1231 ( 
.A1(n_937),
.A2(n_978),
.B1(n_979),
.B2(n_953),
.Y(n_1231)
);

A2O1A1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_975),
.A2(n_968),
.B(n_995),
.C(n_1093),
.Y(n_1232)
);

A2O1A1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_998),
.A2(n_948),
.B(n_1060),
.C(n_1053),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1083),
.B(n_1089),
.Y(n_1234)
);

HB1xp67_ASAP7_75t_L g1235 ( 
.A(n_1029),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1003),
.A2(n_997),
.B(n_991),
.Y(n_1236)
);

BUFx12f_ASAP7_75t_L g1237 ( 
.A(n_940),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_953),
.B(n_979),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_978),
.B(n_967),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1078),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_R g1241 ( 
.A(n_961),
.B(n_1001),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_959),
.B(n_983),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1082),
.Y(n_1243)
);

AOI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1029),
.A2(n_1041),
.B1(n_1040),
.B2(n_1033),
.Y(n_1244)
);

AND2x2_ASAP7_75t_SL g1245 ( 
.A(n_986),
.B(n_1010),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_942),
.A2(n_960),
.B(n_966),
.Y(n_1246)
);

OAI22x1_ASAP7_75t_L g1247 ( 
.A1(n_1209),
.A2(n_1041),
.B1(n_1040),
.B2(n_1097),
.Y(n_1247)
);

AO31x2_ASAP7_75t_L g1248 ( 
.A1(n_1232),
.A2(n_1067),
.A3(n_1006),
.B(n_972),
.Y(n_1248)
);

AO32x2_ASAP7_75t_L g1249 ( 
.A1(n_1111),
.A2(n_964),
.A3(n_981),
.B1(n_1004),
.B2(n_1097),
.Y(n_1249)
);

AND2x4_ASAP7_75t_L g1250 ( 
.A(n_1099),
.B(n_988),
.Y(n_1250)
);

O2A1O1Ixp33_ASAP7_75t_SL g1251 ( 
.A1(n_1101),
.A2(n_988),
.B(n_942),
.C(n_960),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1145),
.A2(n_1036),
.B1(n_1048),
.B2(n_1079),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1101),
.B(n_1091),
.Y(n_1253)
);

O2A1O1Ixp33_ASAP7_75t_SL g1254 ( 
.A1(n_1193),
.A2(n_966),
.B(n_999),
.C(n_1027),
.Y(n_1254)
);

AO31x2_ASAP7_75t_L g1255 ( 
.A1(n_1162),
.A2(n_1025),
.A3(n_1026),
.B(n_1074),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1168),
.A2(n_996),
.B(n_1034),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1108),
.B(n_1092),
.Y(n_1257)
);

BUFx2_ASAP7_75t_L g1258 ( 
.A(n_1135),
.Y(n_1258)
);

INVx5_ASAP7_75t_L g1259 ( 
.A(n_1099),
.Y(n_1259)
);

AOI221xp5_ASAP7_75t_L g1260 ( 
.A1(n_1111),
.A2(n_940),
.B1(n_1177),
.B2(n_1188),
.C(n_1143),
.Y(n_1260)
);

HB1xp67_ASAP7_75t_L g1261 ( 
.A(n_1112),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1168),
.A2(n_1117),
.B(n_1227),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1172),
.Y(n_1263)
);

O2A1O1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1194),
.A2(n_1198),
.B(n_1127),
.C(n_1147),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1105),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1227),
.A2(n_1207),
.B(n_1131),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1118),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1123),
.A2(n_1131),
.B(n_1242),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1187),
.B(n_1100),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1114),
.A2(n_1244),
.B1(n_1113),
.B2(n_1104),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1129),
.B(n_1113),
.Y(n_1271)
);

AOI21xp33_ASAP7_75t_L g1272 ( 
.A1(n_1202),
.A2(n_1230),
.B(n_1121),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1123),
.A2(n_1242),
.B(n_1180),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1160),
.A2(n_1178),
.B(n_1175),
.Y(n_1274)
);

NOR2xp67_ASAP7_75t_L g1275 ( 
.A(n_1115),
.B(n_1099),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1190),
.A2(n_1236),
.B(n_1234),
.Y(n_1276)
);

O2A1O1Ixp33_ASAP7_75t_SL g1277 ( 
.A1(n_1193),
.A2(n_1195),
.B(n_1215),
.C(n_1182),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1153),
.B(n_1200),
.Y(n_1278)
);

AOI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1219),
.A2(n_1141),
.B1(n_1165),
.B2(n_1196),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1160),
.A2(n_1176),
.B(n_1166),
.Y(n_1280)
);

O2A1O1Ixp33_ASAP7_75t_L g1281 ( 
.A1(n_1184),
.A2(n_1201),
.B(n_1235),
.C(n_1204),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1218),
.B(n_1130),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1214),
.A2(n_1139),
.B(n_1246),
.Y(n_1283)
);

AO31x2_ASAP7_75t_L g1284 ( 
.A1(n_1234),
.A2(n_1169),
.A3(n_1233),
.B(n_1226),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1144),
.B(n_1106),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1106),
.B(n_1224),
.Y(n_1286)
);

AOI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1167),
.A2(n_1185),
.B1(n_1142),
.B2(n_1206),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1166),
.A2(n_1176),
.B(n_1223),
.Y(n_1288)
);

NAND2x1p5_ASAP7_75t_L g1289 ( 
.A(n_1098),
.B(n_1122),
.Y(n_1289)
);

AO31x2_ASAP7_75t_L g1290 ( 
.A1(n_1226),
.A2(n_1222),
.A3(n_1157),
.B(n_1243),
.Y(n_1290)
);

CKINVDCx20_ASAP7_75t_R g1291 ( 
.A(n_1133),
.Y(n_1291)
);

AOI221xp5_ASAP7_75t_SL g1292 ( 
.A1(n_1197),
.A2(n_1203),
.B1(n_1195),
.B2(n_1119),
.C(n_1214),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1222),
.A2(n_1239),
.B(n_1189),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1221),
.A2(n_1179),
.B(n_1199),
.Y(n_1294)
);

OAI22x1_ASAP7_75t_L g1295 ( 
.A1(n_1206),
.A2(n_1212),
.B1(n_1134),
.B2(n_1146),
.Y(n_1295)
);

OAI22x1_ASAP7_75t_L g1296 ( 
.A1(n_1164),
.A2(n_1152),
.B1(n_1156),
.B2(n_1170),
.Y(n_1296)
);

NAND3xp33_ASAP7_75t_SL g1297 ( 
.A(n_1217),
.B(n_1216),
.C(n_1159),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1110),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1119),
.A2(n_1116),
.B(n_1240),
.Y(n_1299)
);

OAI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1116),
.A2(n_1140),
.B(n_1126),
.Y(n_1300)
);

AO31x2_ASAP7_75t_L g1301 ( 
.A1(n_1183),
.A2(n_1158),
.A3(n_1138),
.B(n_1151),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1142),
.B(n_1173),
.Y(n_1302)
);

NAND2x1_ASAP7_75t_L g1303 ( 
.A(n_1154),
.B(n_1228),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1107),
.B(n_1142),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_L g1305 ( 
.A(n_1237),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1120),
.B(n_1149),
.Y(n_1306)
);

O2A1O1Ixp33_ASAP7_75t_SL g1307 ( 
.A1(n_1238),
.A2(n_1163),
.B(n_1208),
.C(n_1174),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1124),
.A2(n_1161),
.B1(n_1170),
.B2(n_1156),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1126),
.Y(n_1309)
);

AO22x2_ASAP7_75t_L g1310 ( 
.A1(n_1158),
.A2(n_1181),
.B1(n_1138),
.B2(n_1192),
.Y(n_1310)
);

AND2x4_ASAP7_75t_L g1311 ( 
.A(n_1205),
.B(n_1150),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1103),
.B(n_1109),
.Y(n_1312)
);

BUFx2_ASAP7_75t_SL g1313 ( 
.A(n_1136),
.Y(n_1313)
);

AOI221x1_ASAP7_75t_L g1314 ( 
.A1(n_1229),
.A2(n_1211),
.B1(n_1213),
.B2(n_1183),
.C(n_1148),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1231),
.B(n_1103),
.Y(n_1315)
);

NAND3xp33_ASAP7_75t_L g1316 ( 
.A(n_1155),
.B(n_1152),
.C(n_1171),
.Y(n_1316)
);

OA21x2_ASAP7_75t_L g1317 ( 
.A1(n_1186),
.A2(n_1125),
.B(n_1245),
.Y(n_1317)
);

O2A1O1Ixp33_ASAP7_75t_L g1318 ( 
.A1(n_1137),
.A2(n_1109),
.B(n_1132),
.C(n_1241),
.Y(n_1318)
);

O2A1O1Ixp33_ASAP7_75t_SL g1319 ( 
.A1(n_1154),
.A2(n_1228),
.B(n_1210),
.C(n_1136),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1210),
.B(n_1136),
.Y(n_1320)
);

BUFx2_ASAP7_75t_L g1321 ( 
.A(n_1136),
.Y(n_1321)
);

INVx2_ASAP7_75t_SL g1322 ( 
.A(n_1136),
.Y(n_1322)
);

AO32x2_ASAP7_75t_L g1323 ( 
.A1(n_1111),
.A2(n_1229),
.A3(n_1227),
.B1(n_1126),
.B2(n_1158),
.Y(n_1323)
);

AO31x2_ASAP7_75t_L g1324 ( 
.A1(n_1232),
.A2(n_1086),
.A3(n_1162),
.B(n_1117),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1101),
.B(n_931),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1190),
.A2(n_1236),
.B(n_1117),
.Y(n_1326)
);

OA21x2_ASAP7_75t_L g1327 ( 
.A1(n_1117),
.A2(n_1168),
.B(n_1236),
.Y(n_1327)
);

BUFx10_ASAP7_75t_L g1328 ( 
.A(n_1133),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1133),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_SL g1330 ( 
.A(n_1127),
.B(n_923),
.Y(n_1330)
);

INVx3_ASAP7_75t_L g1331 ( 
.A(n_1225),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1099),
.B(n_1115),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1105),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1168),
.A2(n_931),
.B(n_1162),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1168),
.A2(n_931),
.B(n_1162),
.Y(n_1335)
);

NOR2xp67_ASAP7_75t_L g1336 ( 
.A(n_1115),
.B(n_1084),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1168),
.A2(n_931),
.B(n_1162),
.Y(n_1337)
);

AO31x2_ASAP7_75t_L g1338 ( 
.A1(n_1232),
.A2(n_1086),
.A3(n_1162),
.B(n_1117),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1190),
.A2(n_1236),
.B(n_1117),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_SL g1340 ( 
.A(n_1127),
.B(n_923),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_SL g1341 ( 
.A(n_1127),
.B(n_923),
.Y(n_1341)
);

O2A1O1Ixp33_ASAP7_75t_SL g1342 ( 
.A1(n_1102),
.A2(n_931),
.B(n_1101),
.C(n_923),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1101),
.B(n_931),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1190),
.A2(n_1236),
.B(n_1117),
.Y(n_1344)
);

O2A1O1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1102),
.A2(n_819),
.B(n_793),
.C(n_931),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1101),
.B(n_931),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1168),
.A2(n_931),
.B(n_1162),
.Y(n_1347)
);

AOI221x1_ASAP7_75t_L g1348 ( 
.A1(n_1102),
.A2(n_954),
.B1(n_1111),
.B2(n_1090),
.C(n_1185),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1099),
.Y(n_1349)
);

AOI221xp5_ASAP7_75t_L g1350 ( 
.A1(n_1108),
.A2(n_723),
.B1(n_738),
.B2(n_761),
.C(n_568),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1220),
.Y(n_1351)
);

AOI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1128),
.A2(n_819),
.B1(n_1108),
.B2(n_1076),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1101),
.B(n_931),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1101),
.B(n_931),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1168),
.A2(n_931),
.B(n_1162),
.Y(n_1355)
);

NOR4xp25_ASAP7_75t_L g1356 ( 
.A(n_1102),
.B(n_1111),
.C(n_1164),
.D(n_1209),
.Y(n_1356)
);

AOI221xp5_ASAP7_75t_SL g1357 ( 
.A1(n_1188),
.A2(n_1090),
.B1(n_1050),
.B2(n_1177),
.C(n_1209),
.Y(n_1357)
);

INVx1_ASAP7_75t_SL g1358 ( 
.A(n_1172),
.Y(n_1358)
);

OAI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1128),
.A2(n_819),
.B(n_931),
.Y(n_1359)
);

AO31x2_ASAP7_75t_L g1360 ( 
.A1(n_1232),
.A2(n_1086),
.A3(n_1162),
.B(n_1117),
.Y(n_1360)
);

OR2x2_ASAP7_75t_L g1361 ( 
.A(n_1112),
.B(n_1153),
.Y(n_1361)
);

AO31x2_ASAP7_75t_L g1362 ( 
.A1(n_1232),
.A2(n_1086),
.A3(n_1162),
.B(n_1117),
.Y(n_1362)
);

NAND3xp33_ASAP7_75t_L g1363 ( 
.A(n_1128),
.B(n_819),
.C(n_1090),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1191),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_SL g1365 ( 
.A1(n_1104),
.A2(n_1214),
.B(n_1195),
.Y(n_1365)
);

BUFx4f_ASAP7_75t_SL g1366 ( 
.A(n_1098),
.Y(n_1366)
);

AOI211x1_ASAP7_75t_L g1367 ( 
.A1(n_1102),
.A2(n_1101),
.B(n_1050),
.C(n_886),
.Y(n_1367)
);

A2O1A1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1102),
.A2(n_819),
.B(n_931),
.C(n_1090),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1168),
.A2(n_931),
.B(n_1162),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1168),
.A2(n_931),
.B(n_1162),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_1225),
.Y(n_1371)
);

INVxp67_ASAP7_75t_L g1372 ( 
.A(n_1129),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1172),
.Y(n_1373)
);

AO32x2_ASAP7_75t_L g1374 ( 
.A1(n_1111),
.A2(n_1229),
.A3(n_1227),
.B1(n_1126),
.B2(n_1158),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_1112),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1168),
.A2(n_931),
.B(n_1162),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1112),
.B(n_1153),
.Y(n_1377)
);

AOI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1162),
.A2(n_1117),
.B(n_1207),
.Y(n_1378)
);

BUFx2_ASAP7_75t_SL g1379 ( 
.A(n_1172),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1168),
.A2(n_931),
.B(n_1162),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1101),
.B(n_931),
.Y(n_1381)
);

NOR2xp33_ASAP7_75t_L g1382 ( 
.A(n_1128),
.B(n_819),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1128),
.B(n_819),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1101),
.B(n_931),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1168),
.A2(n_931),
.B(n_1162),
.Y(n_1385)
);

INVxp67_ASAP7_75t_L g1386 ( 
.A(n_1129),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1190),
.A2(n_1236),
.B(n_1117),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1101),
.B(n_931),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1128),
.A2(n_819),
.B(n_931),
.Y(n_1389)
);

AO31x2_ASAP7_75t_L g1390 ( 
.A1(n_1232),
.A2(n_1086),
.A3(n_1162),
.B(n_1117),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_SL g1391 ( 
.A(n_1127),
.B(n_923),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1100),
.B(n_738),
.Y(n_1392)
);

AO221x2_ASAP7_75t_L g1393 ( 
.A1(n_1185),
.A2(n_1111),
.B1(n_568),
.B2(n_572),
.C(n_775),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1108),
.A2(n_931),
.B1(n_819),
.B2(n_932),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1168),
.A2(n_931),
.B(n_1162),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1168),
.A2(n_931),
.B(n_1162),
.Y(n_1396)
);

BUFx4f_ASAP7_75t_SL g1397 ( 
.A(n_1098),
.Y(n_1397)
);

INVx6_ASAP7_75t_SL g1398 ( 
.A(n_1106),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1191),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1190),
.A2(n_1236),
.B(n_1117),
.Y(n_1400)
);

OAI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1352),
.A2(n_1383),
.B(n_1382),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1393),
.A2(n_1363),
.B1(n_1260),
.B2(n_1350),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_L g1403 ( 
.A(n_1305),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1265),
.Y(n_1404)
);

OAI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1368),
.A2(n_1389),
.B(n_1359),
.Y(n_1405)
);

CKINVDCx20_ASAP7_75t_R g1406 ( 
.A(n_1291),
.Y(n_1406)
);

BUFx3_ASAP7_75t_L g1407 ( 
.A(n_1373),
.Y(n_1407)
);

BUFx4f_ASAP7_75t_SL g1408 ( 
.A(n_1398),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_1366),
.Y(n_1409)
);

INVx1_ASAP7_75t_SL g1410 ( 
.A(n_1312),
.Y(n_1410)
);

AOI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1393),
.A2(n_1357),
.B1(n_1394),
.B2(n_1356),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_SL g1412 ( 
.A1(n_1270),
.A2(n_1346),
.B1(n_1343),
.B2(n_1353),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1392),
.A2(n_1279),
.B1(n_1278),
.B2(n_1269),
.Y(n_1413)
);

INVx2_ASAP7_75t_SL g1414 ( 
.A(n_1305),
.Y(n_1414)
);

INVx6_ASAP7_75t_L g1415 ( 
.A(n_1305),
.Y(n_1415)
);

CKINVDCx20_ASAP7_75t_R g1416 ( 
.A(n_1397),
.Y(n_1416)
);

INVx6_ASAP7_75t_L g1417 ( 
.A(n_1259),
.Y(n_1417)
);

AOI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1325),
.A2(n_1384),
.B1(n_1381),
.B2(n_1354),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1388),
.A2(n_1351),
.B1(n_1341),
.B2(n_1391),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1267),
.Y(n_1420)
);

BUFx2_ASAP7_75t_L g1421 ( 
.A(n_1398),
.Y(n_1421)
);

INVx6_ASAP7_75t_L g1422 ( 
.A(n_1259),
.Y(n_1422)
);

BUFx10_ASAP7_75t_L g1423 ( 
.A(n_1329),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_SL g1424 ( 
.A1(n_1317),
.A2(n_1300),
.B1(n_1299),
.B2(n_1348),
.Y(n_1424)
);

AOI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1330),
.A2(n_1340),
.B1(n_1287),
.B2(n_1271),
.Y(n_1425)
);

CKINVDCx20_ASAP7_75t_R g1426 ( 
.A(n_1258),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1333),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1351),
.A2(n_1298),
.B1(n_1399),
.B2(n_1364),
.Y(n_1428)
);

INVx1_ASAP7_75t_SL g1429 ( 
.A(n_1315),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1296),
.A2(n_1247),
.B1(n_1308),
.B2(n_1317),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1264),
.A2(n_1367),
.B1(n_1309),
.B2(n_1345),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1257),
.A2(n_1385),
.B1(n_1376),
.B2(n_1370),
.Y(n_1432)
);

INVxp67_ASAP7_75t_SL g1433 ( 
.A(n_1273),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1334),
.A2(n_1369),
.B1(n_1355),
.B2(n_1347),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1282),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1306),
.Y(n_1436)
);

CKINVDCx14_ASAP7_75t_R g1437 ( 
.A(n_1328),
.Y(n_1437)
);

INVx1_ASAP7_75t_SL g1438 ( 
.A(n_1261),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1375),
.B(n_1361),
.Y(n_1439)
);

INVx6_ASAP7_75t_L g1440 ( 
.A(n_1328),
.Y(n_1440)
);

INVx6_ASAP7_75t_L g1441 ( 
.A(n_1349),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1377),
.Y(n_1442)
);

CKINVDCx20_ASAP7_75t_R g1443 ( 
.A(n_1379),
.Y(n_1443)
);

BUFx8_ASAP7_75t_L g1444 ( 
.A(n_1349),
.Y(n_1444)
);

AND2x4_ASAP7_75t_L g1445 ( 
.A(n_1320),
.B(n_1311),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1286),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_1289),
.Y(n_1447)
);

OAI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1253),
.A2(n_1302),
.B1(n_1372),
.B2(n_1386),
.Y(n_1448)
);

CKINVDCx20_ASAP7_75t_R g1449 ( 
.A(n_1358),
.Y(n_1449)
);

CKINVDCx11_ASAP7_75t_R g1450 ( 
.A(n_1332),
.Y(n_1450)
);

BUFx3_ASAP7_75t_L g1451 ( 
.A(n_1285),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1311),
.Y(n_1452)
);

INVx1_ASAP7_75t_SL g1453 ( 
.A(n_1321),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1250),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1295),
.Y(n_1455)
);

INVx4_ASAP7_75t_SL g1456 ( 
.A(n_1322),
.Y(n_1456)
);

BUFx10_ASAP7_75t_L g1457 ( 
.A(n_1304),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_1332),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1342),
.B(n_1268),
.Y(n_1459)
);

OAI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1314),
.A2(n_1272),
.B1(n_1374),
.B2(n_1323),
.Y(n_1460)
);

INVx6_ASAP7_75t_L g1461 ( 
.A(n_1275),
.Y(n_1461)
);

INVx6_ASAP7_75t_L g1462 ( 
.A(n_1336),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1331),
.Y(n_1463)
);

OAI22x1_ASAP7_75t_SL g1464 ( 
.A1(n_1331),
.A2(n_1371),
.B1(n_1323),
.B2(n_1374),
.Y(n_1464)
);

CKINVDCx20_ASAP7_75t_R g1465 ( 
.A(n_1371),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1303),
.Y(n_1466)
);

INVx3_ASAP7_75t_SL g1467 ( 
.A(n_1310),
.Y(n_1467)
);

INVx1_ASAP7_75t_SL g1468 ( 
.A(n_1313),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1297),
.A2(n_1310),
.B1(n_1365),
.B2(n_1252),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1316),
.A2(n_1380),
.B1(n_1337),
.B2(n_1396),
.Y(n_1470)
);

NAND2x1p5_ASAP7_75t_L g1471 ( 
.A(n_1280),
.B(n_1294),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1335),
.A2(n_1395),
.B1(n_1288),
.B2(n_1256),
.Y(n_1472)
);

INVx6_ASAP7_75t_L g1473 ( 
.A(n_1319),
.Y(n_1473)
);

INVx4_ASAP7_75t_L g1474 ( 
.A(n_1327),
.Y(n_1474)
);

BUFx2_ASAP7_75t_L g1475 ( 
.A(n_1249),
.Y(n_1475)
);

OAI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1262),
.A2(n_1281),
.B1(n_1266),
.B2(n_1283),
.Y(n_1476)
);

CKINVDCx14_ASAP7_75t_R g1477 ( 
.A(n_1292),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1290),
.B(n_1293),
.Y(n_1478)
);

BUFx10_ASAP7_75t_L g1479 ( 
.A(n_1318),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1301),
.B(n_1290),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1274),
.A2(n_1327),
.B1(n_1249),
.B2(n_1277),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1307),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1276),
.A2(n_1400),
.B1(n_1387),
.B2(n_1344),
.Y(n_1483)
);

NAND2x1p5_ASAP7_75t_L g1484 ( 
.A(n_1378),
.B(n_1339),
.Y(n_1484)
);

INVx2_ASAP7_75t_SL g1485 ( 
.A(n_1248),
.Y(n_1485)
);

OAI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1301),
.A2(n_1254),
.B1(n_1251),
.B2(n_1248),
.Y(n_1486)
);

BUFx8_ASAP7_75t_L g1487 ( 
.A(n_1301),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1326),
.A2(n_1284),
.B1(n_1324),
.B2(n_1338),
.Y(n_1488)
);

INVx3_ASAP7_75t_L g1489 ( 
.A(n_1324),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1338),
.A2(n_1360),
.B1(n_1362),
.B2(n_1390),
.Y(n_1490)
);

INVx8_ASAP7_75t_L g1491 ( 
.A(n_1360),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1362),
.Y(n_1492)
);

CKINVDCx8_ASAP7_75t_R g1493 ( 
.A(n_1255),
.Y(n_1493)
);

CKINVDCx20_ASAP7_75t_R g1494 ( 
.A(n_1291),
.Y(n_1494)
);

BUFx2_ASAP7_75t_SL g1495 ( 
.A(n_1291),
.Y(n_1495)
);

OAI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1352),
.A2(n_1383),
.B1(n_1382),
.B2(n_1363),
.Y(n_1496)
);

CKINVDCx11_ASAP7_75t_R g1497 ( 
.A(n_1291),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1284),
.Y(n_1498)
);

BUFx6f_ASAP7_75t_L g1499 ( 
.A(n_1305),
.Y(n_1499)
);

CKINVDCx11_ASAP7_75t_R g1500 ( 
.A(n_1291),
.Y(n_1500)
);

INVx8_ASAP7_75t_L g1501 ( 
.A(n_1259),
.Y(n_1501)
);

NAND2x1p5_ASAP7_75t_L g1502 ( 
.A(n_1259),
.B(n_1225),
.Y(n_1502)
);

INVxp67_ASAP7_75t_L g1503 ( 
.A(n_1271),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1265),
.Y(n_1504)
);

CKINVDCx11_ASAP7_75t_R g1505 ( 
.A(n_1291),
.Y(n_1505)
);

BUFx8_ASAP7_75t_L g1506 ( 
.A(n_1263),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1265),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1393),
.A2(n_954),
.B1(n_1383),
.B2(n_1382),
.Y(n_1508)
);

INVx6_ASAP7_75t_L g1509 ( 
.A(n_1305),
.Y(n_1509)
);

CKINVDCx14_ASAP7_75t_R g1510 ( 
.A(n_1291),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_SL g1511 ( 
.A1(n_1382),
.A2(n_1383),
.B1(n_1352),
.B2(n_1363),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_1373),
.Y(n_1512)
);

CKINVDCx20_ASAP7_75t_R g1513 ( 
.A(n_1291),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1382),
.B(n_1383),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1352),
.A2(n_1382),
.B1(n_1383),
.B2(n_931),
.Y(n_1515)
);

BUFx2_ASAP7_75t_L g1516 ( 
.A(n_1398),
.Y(n_1516)
);

CKINVDCx11_ASAP7_75t_R g1517 ( 
.A(n_1291),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_SL g1518 ( 
.A1(n_1393),
.A2(n_1145),
.B1(n_1383),
.B2(n_1382),
.Y(n_1518)
);

AOI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1382),
.A2(n_1383),
.B1(n_1352),
.B2(n_1363),
.Y(n_1519)
);

OAI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1352),
.A2(n_1383),
.B1(n_1382),
.B2(n_1363),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1265),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_1329),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1265),
.Y(n_1523)
);

CKINVDCx6p67_ASAP7_75t_R g1524 ( 
.A(n_1291),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1393),
.A2(n_954),
.B1(n_1383),
.B2(n_1382),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1265),
.Y(n_1526)
);

AOI21xp5_ASAP7_75t_L g1527 ( 
.A1(n_1262),
.A2(n_1266),
.B(n_1334),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1265),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1393),
.A2(n_954),
.B1(n_1383),
.B2(n_1382),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_SL g1530 ( 
.A1(n_1393),
.A2(n_1145),
.B1(n_1383),
.B2(n_1382),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1265),
.Y(n_1531)
);

BUFx6f_ASAP7_75t_L g1532 ( 
.A(n_1305),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_L g1533 ( 
.A(n_1438),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1480),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1404),
.Y(n_1535)
);

OA21x2_ASAP7_75t_L g1536 ( 
.A1(n_1527),
.A2(n_1481),
.B(n_1470),
.Y(n_1536)
);

OAI21x1_ASAP7_75t_L g1537 ( 
.A1(n_1527),
.A2(n_1484),
.B(n_1471),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1420),
.Y(n_1538)
);

BUFx3_ASAP7_75t_L g1539 ( 
.A(n_1473),
.Y(n_1539)
);

BUFx4f_ASAP7_75t_SL g1540 ( 
.A(n_1409),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1503),
.B(n_1418),
.Y(n_1541)
);

INVx2_ASAP7_75t_SL g1542 ( 
.A(n_1473),
.Y(n_1542)
);

INVx3_ASAP7_75t_L g1543 ( 
.A(n_1474),
.Y(n_1543)
);

OAI21x1_ASAP7_75t_L g1544 ( 
.A1(n_1484),
.A2(n_1471),
.B(n_1434),
.Y(n_1544)
);

CKINVDCx6p67_ASAP7_75t_R g1545 ( 
.A(n_1416),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1514),
.B(n_1401),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_1497),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1410),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1427),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1475),
.B(n_1503),
.Y(n_1550)
);

OAI21x1_ASAP7_75t_L g1551 ( 
.A1(n_1434),
.A2(n_1432),
.B(n_1483),
.Y(n_1551)
);

OA21x2_ASAP7_75t_L g1552 ( 
.A1(n_1472),
.A2(n_1478),
.B(n_1459),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1504),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1439),
.Y(n_1554)
);

INVx4_ASAP7_75t_SL g1555 ( 
.A(n_1467),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1507),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1521),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1523),
.Y(n_1558)
);

INVx4_ASAP7_75t_L g1559 ( 
.A(n_1479),
.Y(n_1559)
);

BUFx3_ASAP7_75t_L g1560 ( 
.A(n_1442),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1526),
.Y(n_1561)
);

AO21x2_ASAP7_75t_L g1562 ( 
.A1(n_1460),
.A2(n_1486),
.B(n_1478),
.Y(n_1562)
);

OR2x6_ASAP7_75t_L g1563 ( 
.A(n_1491),
.B(n_1485),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1518),
.A2(n_1530),
.B1(n_1477),
.B2(n_1508),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1528),
.Y(n_1565)
);

BUFx10_ASAP7_75t_L g1566 ( 
.A(n_1440),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1531),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1498),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_L g1569 ( 
.A(n_1401),
.B(n_1511),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1424),
.B(n_1498),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1492),
.Y(n_1571)
);

NAND3xp33_ASAP7_75t_SL g1572 ( 
.A(n_1519),
.B(n_1518),
.C(n_1530),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1492),
.Y(n_1573)
);

OAI21x1_ASAP7_75t_L g1574 ( 
.A1(n_1432),
.A2(n_1476),
.B(n_1459),
.Y(n_1574)
);

BUFx2_ASAP7_75t_SL g1575 ( 
.A(n_1479),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1433),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1418),
.B(n_1412),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1433),
.Y(n_1578)
);

BUFx3_ASAP7_75t_L g1579 ( 
.A(n_1444),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1456),
.B(n_1453),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1487),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1487),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1429),
.B(n_1448),
.Y(n_1583)
);

OAI21x1_ASAP7_75t_L g1584 ( 
.A1(n_1476),
.A2(n_1489),
.B(n_1488),
.Y(n_1584)
);

OAI21x1_ASAP7_75t_L g1585 ( 
.A1(n_1490),
.A2(n_1469),
.B(n_1482),
.Y(n_1585)
);

BUFx2_ASAP7_75t_L g1586 ( 
.A(n_1474),
.Y(n_1586)
);

OA21x2_ASAP7_75t_L g1587 ( 
.A1(n_1430),
.A2(n_1405),
.B(n_1455),
.Y(n_1587)
);

OAI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1515),
.A2(n_1519),
.B(n_1520),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1412),
.B(n_1515),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1491),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1448),
.B(n_1491),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1493),
.Y(n_1592)
);

INVx4_ASAP7_75t_L g1593 ( 
.A(n_1501),
.Y(n_1593)
);

OAI221xp5_ASAP7_75t_L g1594 ( 
.A1(n_1525),
.A2(n_1529),
.B1(n_1402),
.B2(n_1511),
.C(n_1411),
.Y(n_1594)
);

AOI21x1_ASAP7_75t_L g1595 ( 
.A1(n_1431),
.A2(n_1405),
.B(n_1452),
.Y(n_1595)
);

OAI21xp5_ASAP7_75t_L g1596 ( 
.A1(n_1496),
.A2(n_1411),
.B(n_1431),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1486),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1464),
.Y(n_1598)
);

INVx3_ASAP7_75t_L g1599 ( 
.A(n_1466),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1456),
.B(n_1453),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1436),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1413),
.A2(n_1454),
.B1(n_1446),
.B2(n_1425),
.Y(n_1602)
);

INVx3_ASAP7_75t_L g1603 ( 
.A(n_1468),
.Y(n_1603)
);

BUFx2_ASAP7_75t_L g1604 ( 
.A(n_1468),
.Y(n_1604)
);

OA21x2_ASAP7_75t_L g1605 ( 
.A1(n_1425),
.A2(n_1435),
.B(n_1428),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1419),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1451),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_SL g1608 ( 
.A1(n_1461),
.A2(n_1462),
.B1(n_1408),
.B2(n_1458),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1445),
.Y(n_1609)
);

INVx2_ASAP7_75t_SL g1610 ( 
.A(n_1444),
.Y(n_1610)
);

OR2x6_ASAP7_75t_L g1611 ( 
.A(n_1501),
.B(n_1417),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_1465),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1407),
.B(n_1512),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1463),
.B(n_1457),
.Y(n_1614)
);

INVx2_ASAP7_75t_SL g1615 ( 
.A(n_1422),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1441),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1462),
.Y(n_1617)
);

BUFx2_ASAP7_75t_L g1618 ( 
.A(n_1506),
.Y(n_1618)
);

INVx4_ASAP7_75t_L g1619 ( 
.A(n_1502),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1461),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1457),
.B(n_1403),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1532),
.Y(n_1622)
);

OAI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1502),
.A2(n_1449),
.B(n_1426),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1421),
.B(n_1516),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1499),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1499),
.Y(n_1626)
);

OA21x2_ASAP7_75t_L g1627 ( 
.A1(n_1574),
.A2(n_1414),
.B(n_1522),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1554),
.B(n_1548),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1546),
.B(n_1510),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1560),
.B(n_1495),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1560),
.B(n_1532),
.Y(n_1631)
);

A2O1A1Ixp33_ASAP7_75t_L g1632 ( 
.A1(n_1569),
.A2(n_1564),
.B(n_1572),
.C(n_1594),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1533),
.Y(n_1633)
);

INVx3_ASAP7_75t_L g1634 ( 
.A(n_1580),
.Y(n_1634)
);

O2A1O1Ixp33_ASAP7_75t_L g1635 ( 
.A1(n_1588),
.A2(n_1437),
.B(n_1447),
.C(n_1443),
.Y(n_1635)
);

OR2x6_ASAP7_75t_L g1636 ( 
.A(n_1591),
.B(n_1563),
.Y(n_1636)
);

INVx4_ASAP7_75t_L g1637 ( 
.A(n_1559),
.Y(n_1637)
);

AOI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1577),
.A2(n_1450),
.B1(n_1415),
.B2(n_1509),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1598),
.A2(n_1506),
.B1(n_1415),
.B2(n_1509),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1541),
.B(n_1440),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1604),
.B(n_1524),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1607),
.B(n_1423),
.Y(n_1642)
);

AO21x1_ASAP7_75t_L g1643 ( 
.A1(n_1589),
.A2(n_1500),
.B(n_1505),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1550),
.B(n_1423),
.Y(n_1644)
);

OR2x6_ASAP7_75t_L g1645 ( 
.A(n_1591),
.B(n_1517),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1550),
.B(n_1406),
.Y(n_1646)
);

AOI21xp33_ASAP7_75t_L g1647 ( 
.A1(n_1596),
.A2(n_1494),
.B(n_1513),
.Y(n_1647)
);

OR2x6_ASAP7_75t_L g1648 ( 
.A(n_1563),
.B(n_1580),
.Y(n_1648)
);

AO32x2_ASAP7_75t_L g1649 ( 
.A1(n_1559),
.A2(n_1542),
.A3(n_1615),
.B1(n_1610),
.B2(n_1619),
.Y(n_1649)
);

AO32x2_ASAP7_75t_L g1650 ( 
.A1(n_1559),
.A2(n_1542),
.A3(n_1615),
.B1(n_1610),
.B2(n_1619),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_1545),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1576),
.B(n_1578),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1535),
.Y(n_1653)
);

OA21x2_ASAP7_75t_L g1654 ( 
.A1(n_1574),
.A2(n_1551),
.B(n_1537),
.Y(n_1654)
);

BUFx6f_ASAP7_75t_L g1655 ( 
.A(n_1539),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1535),
.Y(n_1656)
);

NOR2x1_ASAP7_75t_SL g1657 ( 
.A(n_1611),
.B(n_1575),
.Y(n_1657)
);

BUFx3_ASAP7_75t_L g1658 ( 
.A(n_1540),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1603),
.B(n_1612),
.Y(n_1659)
);

OAI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1595),
.A2(n_1583),
.B(n_1597),
.Y(n_1660)
);

A2O1A1Ixp33_ASAP7_75t_L g1661 ( 
.A1(n_1570),
.A2(n_1606),
.B(n_1585),
.C(n_1539),
.Y(n_1661)
);

NOR2x1_ASAP7_75t_L g1662 ( 
.A(n_1559),
.B(n_1575),
.Y(n_1662)
);

O2A1O1Ixp33_ASAP7_75t_L g1663 ( 
.A1(n_1562),
.A2(n_1536),
.B(n_1587),
.C(n_1624),
.Y(n_1663)
);

INVx3_ASAP7_75t_L g1664 ( 
.A(n_1600),
.Y(n_1664)
);

AND2x4_ASAP7_75t_L g1665 ( 
.A(n_1600),
.B(n_1581),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1602),
.A2(n_1595),
.B1(n_1618),
.B2(n_1613),
.Y(n_1666)
);

CKINVDCx20_ASAP7_75t_R g1667 ( 
.A(n_1547),
.Y(n_1667)
);

A2O1A1Ixp33_ASAP7_75t_L g1668 ( 
.A1(n_1585),
.A2(n_1623),
.B(n_1584),
.C(n_1592),
.Y(n_1668)
);

BUFx4f_ASAP7_75t_SL g1669 ( 
.A(n_1579),
.Y(n_1669)
);

OAI211xp5_ASAP7_75t_L g1670 ( 
.A1(n_1536),
.A2(n_1587),
.B(n_1552),
.C(n_1551),
.Y(n_1670)
);

NOR2x1_ASAP7_75t_L g1671 ( 
.A(n_1579),
.B(n_1599),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_1547),
.Y(n_1672)
);

INVxp67_ASAP7_75t_L g1673 ( 
.A(n_1617),
.Y(n_1673)
);

AO32x2_ASAP7_75t_L g1674 ( 
.A1(n_1619),
.A2(n_1587),
.A3(n_1593),
.B1(n_1605),
.B2(n_1562),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1618),
.B(n_1566),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1621),
.B(n_1614),
.Y(n_1676)
);

HB1xp67_ASAP7_75t_L g1677 ( 
.A(n_1538),
.Y(n_1677)
);

OAI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1584),
.A2(n_1536),
.B(n_1587),
.Y(n_1678)
);

INVxp67_ASAP7_75t_L g1679 ( 
.A(n_1617),
.Y(n_1679)
);

AO32x2_ASAP7_75t_L g1680 ( 
.A1(n_1619),
.A2(n_1593),
.A3(n_1605),
.B1(n_1534),
.B2(n_1601),
.Y(n_1680)
);

NOR2x1_ASAP7_75t_SL g1681 ( 
.A(n_1611),
.B(n_1593),
.Y(n_1681)
);

A2O1A1Ixp33_ASAP7_75t_L g1682 ( 
.A1(n_1620),
.A2(n_1608),
.B(n_1582),
.C(n_1590),
.Y(n_1682)
);

INVx1_ASAP7_75t_SL g1683 ( 
.A(n_1622),
.Y(n_1683)
);

AOI221xp5_ASAP7_75t_L g1684 ( 
.A1(n_1549),
.A2(n_1553),
.B1(n_1558),
.B2(n_1557),
.C(n_1556),
.Y(n_1684)
);

OAI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1536),
.A2(n_1552),
.B(n_1605),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1625),
.B(n_1626),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1537),
.A2(n_1544),
.B(n_1586),
.Y(n_1687)
);

INVx3_ASAP7_75t_L g1688 ( 
.A(n_1654),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1653),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1656),
.Y(n_1690)
);

BUFx3_ASAP7_75t_L g1691 ( 
.A(n_1645),
.Y(n_1691)
);

AOI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1632),
.A2(n_1609),
.B1(n_1555),
.B2(n_1558),
.Y(n_1692)
);

HB1xp67_ASAP7_75t_L g1693 ( 
.A(n_1633),
.Y(n_1693)
);

INVx1_ASAP7_75t_SL g1694 ( 
.A(n_1683),
.Y(n_1694)
);

BUFx2_ASAP7_75t_L g1695 ( 
.A(n_1649),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1648),
.B(n_1543),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1652),
.Y(n_1697)
);

NOR2x1_ASAP7_75t_SL g1698 ( 
.A(n_1645),
.B(n_1611),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1677),
.Y(n_1699)
);

INVxp33_ASAP7_75t_L g1700 ( 
.A(n_1657),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1678),
.B(n_1565),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1680),
.Y(n_1702)
);

BUFx6f_ASAP7_75t_L g1703 ( 
.A(n_1627),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1685),
.B(n_1556),
.Y(n_1704)
);

BUFx2_ASAP7_75t_L g1705 ( 
.A(n_1649),
.Y(n_1705)
);

BUFx2_ASAP7_75t_L g1706 ( 
.A(n_1649),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1680),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1685),
.B(n_1557),
.Y(n_1708)
);

BUFx2_ASAP7_75t_L g1709 ( 
.A(n_1650),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1680),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1645),
.A2(n_1567),
.B1(n_1561),
.B2(n_1553),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1634),
.B(n_1664),
.Y(n_1712)
);

INVxp67_ASAP7_75t_SL g1713 ( 
.A(n_1663),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1684),
.B(n_1568),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1684),
.B(n_1568),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1634),
.B(n_1664),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1674),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1659),
.B(n_1676),
.Y(n_1718)
);

HB1xp67_ASAP7_75t_L g1719 ( 
.A(n_1628),
.Y(n_1719)
);

INVxp67_ASAP7_75t_SL g1720 ( 
.A(n_1663),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1674),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1644),
.B(n_1683),
.Y(n_1722)
);

INVx4_ASAP7_75t_L g1723 ( 
.A(n_1691),
.Y(n_1723)
);

NAND4xp25_ASAP7_75t_L g1724 ( 
.A(n_1695),
.B(n_1647),
.C(n_1629),
.D(n_1644),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1688),
.Y(n_1725)
);

INVxp67_ASAP7_75t_L g1726 ( 
.A(n_1699),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1688),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1695),
.B(n_1674),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1697),
.B(n_1704),
.Y(n_1729)
);

NOR2x1_ASAP7_75t_L g1730 ( 
.A(n_1691),
.B(n_1671),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1695),
.B(n_1630),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1689),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1699),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1688),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1689),
.Y(n_1735)
);

OAI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1713),
.A2(n_1666),
.B(n_1660),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1688),
.Y(n_1737)
);

BUFx6f_ASAP7_75t_L g1738 ( 
.A(n_1703),
.Y(n_1738)
);

AOI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1713),
.A2(n_1670),
.B(n_1687),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1698),
.B(n_1665),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1719),
.B(n_1646),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1688),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1719),
.B(n_1660),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1689),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1690),
.Y(n_1745)
);

BUFx2_ASAP7_75t_L g1746 ( 
.A(n_1705),
.Y(n_1746)
);

AOI21xp33_ASAP7_75t_L g1747 ( 
.A1(n_1720),
.A2(n_1666),
.B(n_1670),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1705),
.B(n_1686),
.Y(n_1748)
);

INVxp67_ASAP7_75t_L g1749 ( 
.A(n_1693),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1690),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1706),
.B(n_1650),
.Y(n_1751)
);

INVx5_ASAP7_75t_SL g1752 ( 
.A(n_1703),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1704),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1693),
.B(n_1640),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1697),
.B(n_1640),
.Y(n_1755)
);

AND2x4_ASAP7_75t_L g1756 ( 
.A(n_1698),
.B(n_1665),
.Y(n_1756)
);

NOR2x1_ASAP7_75t_L g1757 ( 
.A(n_1691),
.B(n_1662),
.Y(n_1757)
);

BUFx3_ASAP7_75t_L g1758 ( 
.A(n_1691),
.Y(n_1758)
);

OAI31xp33_ASAP7_75t_SL g1759 ( 
.A1(n_1711),
.A2(n_1647),
.A3(n_1675),
.B(n_1641),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1706),
.B(n_1631),
.Y(n_1760)
);

OR2x2_ASAP7_75t_L g1761 ( 
.A(n_1722),
.B(n_1668),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1709),
.B(n_1642),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1690),
.Y(n_1763)
);

OAI33xp33_ASAP7_75t_L g1764 ( 
.A1(n_1714),
.A2(n_1635),
.A3(n_1673),
.B1(n_1679),
.B2(n_1571),
.B3(n_1573),
.Y(n_1764)
);

NOR2x1_ASAP7_75t_L g1765 ( 
.A(n_1709),
.B(n_1637),
.Y(n_1765)
);

OAI33xp33_ASAP7_75t_L g1766 ( 
.A1(n_1714),
.A2(n_1635),
.A3(n_1573),
.B1(n_1651),
.B2(n_1616),
.B3(n_1672),
.Y(n_1766)
);

HB1xp67_ASAP7_75t_L g1767 ( 
.A(n_1704),
.Y(n_1767)
);

INVx3_ASAP7_75t_L g1768 ( 
.A(n_1703),
.Y(n_1768)
);

NAND3xp33_ASAP7_75t_L g1769 ( 
.A(n_1720),
.B(n_1661),
.C(n_1638),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1718),
.B(n_1650),
.Y(n_1770)
);

AOI22xp33_ASAP7_75t_SL g1771 ( 
.A1(n_1702),
.A2(n_1681),
.B1(n_1655),
.B2(n_1636),
.Y(n_1771)
);

INVx1_ASAP7_75t_SL g1772 ( 
.A(n_1694),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1724),
.B(n_1643),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1751),
.B(n_1712),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1732),
.Y(n_1775)
);

AND2x4_ASAP7_75t_SL g1776 ( 
.A(n_1740),
.B(n_1696),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1751),
.B(n_1712),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1732),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1738),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1729),
.B(n_1708),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1733),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1735),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1753),
.B(n_1716),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1738),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1735),
.Y(n_1785)
);

AND2x4_ASAP7_75t_L g1786 ( 
.A(n_1740),
.B(n_1756),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1753),
.B(n_1716),
.Y(n_1787)
);

NOR2x1_ASAP7_75t_L g1788 ( 
.A(n_1723),
.B(n_1694),
.Y(n_1788)
);

INVx1_ASAP7_75t_SL g1789 ( 
.A(n_1772),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1729),
.B(n_1708),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1738),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1738),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1744),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1738),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1744),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1738),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1725),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1726),
.B(n_1708),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1767),
.B(n_1702),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1726),
.B(n_1701),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1767),
.B(n_1702),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1740),
.B(n_1756),
.Y(n_1802)
);

AND2x4_ASAP7_75t_SL g1803 ( 
.A(n_1740),
.B(n_1756),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1725),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1755),
.B(n_1701),
.Y(n_1805)
);

INVx1_ASAP7_75t_SL g1806 ( 
.A(n_1772),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1770),
.B(n_1702),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1725),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1724),
.B(n_1669),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1746),
.B(n_1743),
.Y(n_1810)
);

INVx3_ASAP7_75t_L g1811 ( 
.A(n_1752),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1746),
.B(n_1717),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1745),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1770),
.B(n_1707),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1755),
.B(n_1749),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1728),
.B(n_1707),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1803),
.B(n_1762),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1775),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1803),
.B(n_1762),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1803),
.B(n_1731),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1803),
.B(n_1731),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1775),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1815),
.B(n_1743),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1778),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1797),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1797),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1797),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1815),
.B(n_1728),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1778),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1797),
.Y(n_1830)
);

INVx2_ASAP7_75t_SL g1831 ( 
.A(n_1776),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1810),
.B(n_1749),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1776),
.B(n_1760),
.Y(n_1833)
);

OR2x2_ASAP7_75t_L g1834 ( 
.A(n_1810),
.B(n_1805),
.Y(n_1834)
);

OAI31xp33_ASAP7_75t_L g1835 ( 
.A1(n_1773),
.A2(n_1769),
.A3(n_1747),
.B(n_1761),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1776),
.B(n_1760),
.Y(n_1836)
);

NOR2xp33_ASAP7_75t_L g1837 ( 
.A(n_1809),
.B(n_1667),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1782),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1782),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1785),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1776),
.B(n_1723),
.Y(n_1841)
);

NAND3xp33_ASAP7_75t_L g1842 ( 
.A(n_1773),
.B(n_1759),
.C(n_1739),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1804),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1785),
.Y(n_1844)
);

OR2x2_ASAP7_75t_L g1845 ( 
.A(n_1810),
.B(n_1805),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1786),
.B(n_1723),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1789),
.B(n_1728),
.Y(n_1847)
);

OAI21xp33_ASAP7_75t_SL g1848 ( 
.A1(n_1788),
.A2(n_1759),
.B(n_1765),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1789),
.B(n_1733),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1793),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1786),
.B(n_1723),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1804),
.Y(n_1852)
);

CKINVDCx16_ASAP7_75t_R g1853 ( 
.A(n_1809),
.Y(n_1853)
);

OR2x2_ASAP7_75t_L g1854 ( 
.A(n_1798),
.B(n_1754),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1786),
.B(n_1748),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1806),
.B(n_1781),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1786),
.B(n_1748),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1793),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1806),
.B(n_1750),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1781),
.B(n_1763),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1795),
.Y(n_1861)
);

BUFx2_ASAP7_75t_L g1862 ( 
.A(n_1788),
.Y(n_1862)
);

HB1xp67_ASAP7_75t_L g1863 ( 
.A(n_1812),
.Y(n_1863)
);

OR2x6_ASAP7_75t_L g1864 ( 
.A(n_1842),
.B(n_1739),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1834),
.B(n_1800),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1834),
.B(n_1800),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1820),
.B(n_1786),
.Y(n_1867)
);

NAND2x1p5_ASAP7_75t_L g1868 ( 
.A(n_1862),
.B(n_1730),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1820),
.B(n_1802),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1821),
.B(n_1802),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1818),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1825),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_L g1873 ( 
.A(n_1842),
.B(n_1766),
.Y(n_1873)
);

HB1xp67_ASAP7_75t_L g1874 ( 
.A(n_1863),
.Y(n_1874)
);

AOI22xp33_ASAP7_75t_L g1875 ( 
.A1(n_1835),
.A2(n_1747),
.B1(n_1736),
.B2(n_1769),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1818),
.Y(n_1876)
);

AND2x4_ASAP7_75t_L g1877 ( 
.A(n_1831),
.B(n_1802),
.Y(n_1877)
);

AND2x4_ASAP7_75t_L g1878 ( 
.A(n_1831),
.B(n_1802),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1822),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1835),
.B(n_1761),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1845),
.B(n_1798),
.Y(n_1881)
);

OAI22xp33_ASAP7_75t_L g1882 ( 
.A1(n_1847),
.A2(n_1736),
.B1(n_1692),
.B2(n_1715),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1856),
.B(n_1783),
.Y(n_1883)
);

NAND4xp25_ASAP7_75t_L g1884 ( 
.A(n_1856),
.B(n_1765),
.C(n_1794),
.D(n_1792),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1832),
.B(n_1783),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1845),
.B(n_1780),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1832),
.B(n_1783),
.Y(n_1887)
);

AOI21xp33_ASAP7_75t_L g1888 ( 
.A1(n_1848),
.A2(n_1812),
.B(n_1791),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1821),
.B(n_1817),
.Y(n_1889)
);

NOR2xp33_ASAP7_75t_SL g1890 ( 
.A(n_1837),
.B(n_1766),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1849),
.B(n_1787),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1849),
.B(n_1787),
.Y(n_1892)
);

A2O1A1Ixp33_ASAP7_75t_L g1893 ( 
.A1(n_1848),
.A2(n_1816),
.B(n_1707),
.C(n_1710),
.Y(n_1893)
);

INVxp67_ASAP7_75t_L g1894 ( 
.A(n_1859),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1817),
.B(n_1802),
.Y(n_1895)
);

NOR2xp67_ASAP7_75t_L g1896 ( 
.A(n_1831),
.B(n_1811),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1819),
.B(n_1807),
.Y(n_1897)
);

INVx1_ASAP7_75t_SL g1898 ( 
.A(n_1853),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1819),
.B(n_1807),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1823),
.B(n_1787),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1853),
.B(n_1658),
.Y(n_1901)
);

INVx1_ASAP7_75t_SL g1902 ( 
.A(n_1841),
.Y(n_1902)
);

AOI31xp33_ASAP7_75t_L g1903 ( 
.A1(n_1898),
.A2(n_1851),
.A3(n_1846),
.B(n_1841),
.Y(n_1903)
);

AOI221xp5_ASAP7_75t_L g1904 ( 
.A1(n_1873),
.A2(n_1828),
.B1(n_1847),
.B2(n_1764),
.C(n_1816),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1873),
.B(n_1863),
.Y(n_1905)
);

OAI21xp5_ASAP7_75t_SL g1906 ( 
.A1(n_1875),
.A2(n_1862),
.B(n_1851),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1874),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1875),
.B(n_1823),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1901),
.B(n_1846),
.Y(n_1909)
);

NAND4xp25_ASAP7_75t_SL g1910 ( 
.A(n_1893),
.B(n_1828),
.C(n_1857),
.D(n_1855),
.Y(n_1910)
);

O2A1O1Ixp33_ASAP7_75t_L g1911 ( 
.A1(n_1864),
.A2(n_1812),
.B(n_1859),
.C(n_1860),
.Y(n_1911)
);

AOI21xp33_ASAP7_75t_L g1912 ( 
.A1(n_1864),
.A2(n_1824),
.B(n_1822),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1901),
.B(n_1855),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_SL g1914 ( 
.A(n_1882),
.B(n_1833),
.Y(n_1914)
);

OR2x2_ASAP7_75t_L g1915 ( 
.A(n_1864),
.B(n_1854),
.Y(n_1915)
);

AOI221x1_ASAP7_75t_L g1916 ( 
.A1(n_1880),
.A2(n_1860),
.B1(n_1861),
.B2(n_1858),
.C(n_1824),
.Y(n_1916)
);

OAI21xp33_ASAP7_75t_L g1917 ( 
.A1(n_1864),
.A2(n_1854),
.B(n_1857),
.Y(n_1917)
);

AOI21xp5_ASAP7_75t_L g1918 ( 
.A1(n_1893),
.A2(n_1764),
.B(n_1715),
.Y(n_1918)
);

OAI211xp5_ASAP7_75t_SL g1919 ( 
.A1(n_1888),
.A2(n_1861),
.B(n_1858),
.C(n_1829),
.Y(n_1919)
);

AOI22xp33_ASAP7_75t_L g1920 ( 
.A1(n_1890),
.A2(n_1882),
.B1(n_1721),
.B2(n_1717),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1874),
.Y(n_1921)
);

INVxp67_ASAP7_75t_L g1922 ( 
.A(n_1871),
.Y(n_1922)
);

INVxp67_ASAP7_75t_L g1923 ( 
.A(n_1876),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1879),
.Y(n_1924)
);

OAI221xp5_ASAP7_75t_L g1925 ( 
.A1(n_1884),
.A2(n_1721),
.B1(n_1717),
.B2(n_1707),
.C(n_1710),
.Y(n_1925)
);

O2A1O1Ixp33_ASAP7_75t_L g1926 ( 
.A1(n_1894),
.A2(n_1829),
.B(n_1850),
.C(n_1844),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1872),
.Y(n_1927)
);

INVx1_ASAP7_75t_SL g1928 ( 
.A(n_1902),
.Y(n_1928)
);

NAND4xp25_ASAP7_75t_SL g1929 ( 
.A(n_1867),
.B(n_1833),
.C(n_1836),
.D(n_1799),
.Y(n_1929)
);

AOI221xp5_ASAP7_75t_L g1930 ( 
.A1(n_1872),
.A2(n_1816),
.B1(n_1717),
.B2(n_1721),
.C(n_1710),
.Y(n_1930)
);

AOI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1885),
.A2(n_1839),
.B(n_1838),
.Y(n_1931)
);

A2O1A1Ixp33_ASAP7_75t_L g1932 ( 
.A1(n_1918),
.A2(n_1721),
.B(n_1710),
.C(n_1807),
.Y(n_1932)
);

OAI21xp5_ASAP7_75t_SL g1933 ( 
.A1(n_1906),
.A2(n_1868),
.B(n_1889),
.Y(n_1933)
);

O2A1O1Ixp5_ASAP7_75t_L g1934 ( 
.A1(n_1914),
.A2(n_1877),
.B(n_1878),
.C(n_1887),
.Y(n_1934)
);

INVx3_ASAP7_75t_L g1935 ( 
.A(n_1913),
.Y(n_1935)
);

OAI21xp5_ASAP7_75t_L g1936 ( 
.A1(n_1920),
.A2(n_1896),
.B(n_1868),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1909),
.Y(n_1937)
);

OAI21xp33_ASAP7_75t_L g1938 ( 
.A1(n_1910),
.A2(n_1883),
.B(n_1900),
.Y(n_1938)
);

OR2x2_ASAP7_75t_L g1939 ( 
.A(n_1928),
.B(n_1865),
.Y(n_1939)
);

OAI211xp5_ASAP7_75t_L g1940 ( 
.A1(n_1916),
.A2(n_1870),
.B(n_1867),
.C(n_1895),
.Y(n_1940)
);

AOI322xp5_ASAP7_75t_L g1941 ( 
.A1(n_1908),
.A2(n_1814),
.A3(n_1801),
.B1(n_1799),
.B2(n_1899),
.C1(n_1897),
.C2(n_1891),
.Y(n_1941)
);

OR2x2_ASAP7_75t_L g1942 ( 
.A(n_1905),
.B(n_1915),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1917),
.B(n_1870),
.Y(n_1943)
);

OAI21xp33_ASAP7_75t_L g1944 ( 
.A1(n_1904),
.A2(n_1929),
.B(n_1919),
.Y(n_1944)
);

OAI21xp5_ASAP7_75t_SL g1945 ( 
.A1(n_1919),
.A2(n_1878),
.B(n_1877),
.Y(n_1945)
);

OAI21xp5_ASAP7_75t_SL g1946 ( 
.A1(n_1903),
.A2(n_1878),
.B(n_1877),
.Y(n_1946)
);

NAND2xp33_ASAP7_75t_R g1947 ( 
.A(n_1907),
.B(n_1869),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1921),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1924),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1931),
.B(n_1866),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1927),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1922),
.Y(n_1952)
);

AOI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1930),
.A2(n_1703),
.B1(n_1814),
.B2(n_1692),
.Y(n_1953)
);

NAND2xp33_ASAP7_75t_L g1954 ( 
.A(n_1912),
.B(n_1881),
.Y(n_1954)
);

NOR2xp33_ASAP7_75t_L g1955 ( 
.A(n_1935),
.B(n_1922),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1932),
.B(n_1923),
.Y(n_1956)
);

HB1xp67_ASAP7_75t_L g1957 ( 
.A(n_1935),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1937),
.B(n_1836),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1950),
.B(n_1923),
.Y(n_1959)
);

XNOR2x1_ASAP7_75t_L g1960 ( 
.A(n_1942),
.B(n_1814),
.Y(n_1960)
);

OAI22xp33_ASAP7_75t_SL g1961 ( 
.A1(n_1939),
.A2(n_1925),
.B1(n_1936),
.B2(n_1953),
.Y(n_1961)
);

AOI22xp5_ASAP7_75t_L g1962 ( 
.A1(n_1944),
.A2(n_1947),
.B1(n_1933),
.B2(n_1954),
.Y(n_1962)
);

O2A1O1Ixp33_ASAP7_75t_L g1963 ( 
.A1(n_1933),
.A2(n_1911),
.B(n_1926),
.C(n_1892),
.Y(n_1963)
);

AOI221xp5_ASAP7_75t_L g1964 ( 
.A1(n_1934),
.A2(n_1825),
.B1(n_1852),
.B2(n_1826),
.C(n_1827),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1948),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1952),
.B(n_1886),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1951),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1949),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1938),
.B(n_1774),
.Y(n_1969)
);

NOR3xp33_ASAP7_75t_L g1970 ( 
.A(n_1945),
.B(n_1826),
.C(n_1825),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1960),
.B(n_1943),
.Y(n_1971)
);

INVxp67_ASAP7_75t_L g1972 ( 
.A(n_1957),
.Y(n_1972)
);

AOI21xp5_ASAP7_75t_L g1973 ( 
.A1(n_1956),
.A2(n_1945),
.B(n_1946),
.Y(n_1973)
);

O2A1O1Ixp5_ASAP7_75t_L g1974 ( 
.A1(n_1956),
.A2(n_1940),
.B(n_1830),
.C(n_1827),
.Y(n_1974)
);

AOI221xp5_ASAP7_75t_SL g1975 ( 
.A1(n_1963),
.A2(n_1941),
.B1(n_1838),
.B2(n_1850),
.C(n_1844),
.Y(n_1975)
);

NAND5xp2_ASAP7_75t_L g1976 ( 
.A(n_1962),
.B(n_1700),
.C(n_1639),
.D(n_1771),
.E(n_1799),
.Y(n_1976)
);

NAND3xp33_ASAP7_75t_L g1977 ( 
.A(n_1955),
.B(n_1852),
.C(n_1827),
.Y(n_1977)
);

NOR2x1_ASAP7_75t_L g1978 ( 
.A(n_1959),
.B(n_1839),
.Y(n_1978)
);

INVx1_ASAP7_75t_SL g1979 ( 
.A(n_1966),
.Y(n_1979)
);

OAI21x1_ASAP7_75t_SL g1980 ( 
.A1(n_1969),
.A2(n_1840),
.B(n_1830),
.Y(n_1980)
);

BUFx6f_ASAP7_75t_L g1981 ( 
.A(n_1968),
.Y(n_1981)
);

NAND3xp33_ASAP7_75t_L g1982 ( 
.A(n_1970),
.B(n_1852),
.C(n_1830),
.Y(n_1982)
);

NOR3x1_ASAP7_75t_L g1983 ( 
.A(n_1965),
.B(n_1967),
.C(n_1958),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1964),
.B(n_1774),
.Y(n_1984)
);

NOR2xp33_ASAP7_75t_L g1985 ( 
.A(n_1961),
.B(n_1840),
.Y(n_1985)
);

OAI22xp5_ASAP7_75t_L g1986 ( 
.A1(n_1979),
.A2(n_1811),
.B1(n_1801),
.B2(n_1752),
.Y(n_1986)
);

OAI211xp5_ASAP7_75t_L g1987 ( 
.A1(n_1973),
.A2(n_1811),
.B(n_1801),
.C(n_1779),
.Y(n_1987)
);

NAND3xp33_ASAP7_75t_SL g1988 ( 
.A(n_1974),
.B(n_1771),
.C(n_1682),
.Y(n_1988)
);

OAI211xp5_ASAP7_75t_SL g1989 ( 
.A1(n_1972),
.A2(n_1811),
.B(n_1779),
.C(n_1792),
.Y(n_1989)
);

OAI211xp5_ASAP7_75t_SL g1990 ( 
.A1(n_1971),
.A2(n_1811),
.B(n_1779),
.C(n_1792),
.Y(n_1990)
);

NAND3xp33_ASAP7_75t_L g1991 ( 
.A(n_1981),
.B(n_1843),
.C(n_1826),
.Y(n_1991)
);

NAND3xp33_ASAP7_75t_SL g1992 ( 
.A(n_1985),
.B(n_1843),
.C(n_1784),
.Y(n_1992)
);

AOI21xp5_ASAP7_75t_L g1993 ( 
.A1(n_1978),
.A2(n_1843),
.B(n_1784),
.Y(n_1993)
);

AOI211xp5_ASAP7_75t_L g1994 ( 
.A1(n_1975),
.A2(n_1711),
.B(n_1784),
.C(n_1779),
.Y(n_1994)
);

NAND4xp25_ASAP7_75t_SL g1995 ( 
.A(n_1984),
.B(n_1977),
.C(n_1982),
.D(n_1983),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_SL g1996 ( 
.A(n_1987),
.B(n_1981),
.Y(n_1996)
);

OAI211xp5_ASAP7_75t_L g1997 ( 
.A1(n_1992),
.A2(n_1981),
.B(n_1980),
.C(n_1976),
.Y(n_1997)
);

AOI221xp5_ASAP7_75t_L g1998 ( 
.A1(n_1995),
.A2(n_1703),
.B1(n_1768),
.B2(n_1804),
.C(n_1808),
.Y(n_1998)
);

AOI221xp5_ASAP7_75t_L g1999 ( 
.A1(n_1988),
.A2(n_1703),
.B1(n_1768),
.B2(n_1804),
.C(n_1808),
.Y(n_1999)
);

OAI22xp33_ASAP7_75t_L g2000 ( 
.A1(n_1991),
.A2(n_1703),
.B1(n_1796),
.B2(n_1784),
.Y(n_2000)
);

AOI221xp5_ASAP7_75t_L g2001 ( 
.A1(n_1990),
.A2(n_1989),
.B1(n_1993),
.B2(n_1994),
.C(n_1986),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_SL g2002 ( 
.A(n_1987),
.B(n_1792),
.Y(n_2002)
);

INVxp67_ASAP7_75t_L g2003 ( 
.A(n_1995),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1996),
.Y(n_2004)
);

NOR2x1_ASAP7_75t_L g2005 ( 
.A(n_1997),
.B(n_1794),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_2003),
.Y(n_2006)
);

NOR2x1_ASAP7_75t_L g2007 ( 
.A(n_2002),
.B(n_1794),
.Y(n_2007)
);

NOR2x1p5_ASAP7_75t_L g2008 ( 
.A(n_2001),
.B(n_1794),
.Y(n_2008)
);

NOR2xp33_ASAP7_75t_R g2009 ( 
.A(n_1998),
.B(n_1566),
.Y(n_2009)
);

AOI21xp5_ASAP7_75t_L g2010 ( 
.A1(n_2006),
.A2(n_1999),
.B(n_2000),
.Y(n_2010)
);

NOR3xp33_ASAP7_75t_L g2011 ( 
.A(n_2004),
.B(n_1796),
.C(n_1791),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_2005),
.B(n_1796),
.Y(n_2012)
);

AOI221xp5_ASAP7_75t_L g2013 ( 
.A1(n_2009),
.A2(n_1796),
.B1(n_1791),
.B2(n_1703),
.C(n_1808),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_2012),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_2011),
.Y(n_2015)
);

OAI22x1_ASAP7_75t_L g2016 ( 
.A1(n_2015),
.A2(n_2008),
.B1(n_2007),
.B2(n_2010),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_SL g2017 ( 
.A(n_2016),
.B(n_2014),
.Y(n_2017)
);

XNOR2x1_ASAP7_75t_L g2018 ( 
.A(n_2016),
.B(n_2013),
.Y(n_2018)
);

AOI221xp5_ASAP7_75t_L g2019 ( 
.A1(n_2017),
.A2(n_1808),
.B1(n_1727),
.B2(n_1734),
.C(n_1737),
.Y(n_2019)
);

OAI22xp5_ASAP7_75t_L g2020 ( 
.A1(n_2018),
.A2(n_1790),
.B1(n_1780),
.B2(n_1777),
.Y(n_2020)
);

AOI21xp5_ASAP7_75t_L g2021 ( 
.A1(n_2020),
.A2(n_2019),
.B(n_1790),
.Y(n_2021)
);

AO221x1_ASAP7_75t_L g2022 ( 
.A1(n_2020),
.A2(n_1768),
.B1(n_1703),
.B2(n_1813),
.C(n_1795),
.Y(n_2022)
);

OAI22x1_ASAP7_75t_L g2023 ( 
.A1(n_2022),
.A2(n_1730),
.B1(n_1757),
.B2(n_1741),
.Y(n_2023)
);

OAI21xp5_ASAP7_75t_L g2024 ( 
.A1(n_2023),
.A2(n_2021),
.B(n_1777),
.Y(n_2024)
);

OAI22xp33_ASAP7_75t_L g2025 ( 
.A1(n_2024),
.A2(n_1768),
.B1(n_1734),
.B2(n_1737),
.Y(n_2025)
);

AOI221xp5_ASAP7_75t_L g2026 ( 
.A1(n_2025),
.A2(n_1742),
.B1(n_1734),
.B2(n_1737),
.C(n_1727),
.Y(n_2026)
);

AOI211xp5_ASAP7_75t_L g2027 ( 
.A1(n_2026),
.A2(n_1758),
.B(n_1566),
.C(n_1727),
.Y(n_2027)
);


endmodule