module fake_jpeg_14061_n_91 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_91);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_91;

wire n_10;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_4),
.B(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_1),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_30),
.Y(n_33)
);

AOI21xp33_ASAP7_75t_L g26 ( 
.A1(n_12),
.A2(n_1),
.B(n_2),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_28),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_19),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_3),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_10),
.B(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_23),
.A2(n_20),
.B1(n_18),
.B2(n_16),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_32),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_16),
.B1(n_11),
.B2(n_21),
.Y(n_38)
);

NOR2x1_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_41),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_25),
.A2(n_11),
.B1(n_13),
.B2(n_20),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_22),
.A2(n_13),
.B1(n_6),
.B2(n_8),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_46),
.B(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_5),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_48),
.A2(n_34),
.B1(n_23),
.B2(n_24),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_5),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_49),
.B(n_51),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_22),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_6),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

OR2x4_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_27),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_24),
.B1(n_37),
.B2(n_44),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_52),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_63),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_43),
.B(n_37),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_64),
.A2(n_45),
.B(n_54),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_69),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_68),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_48),
.C(n_45),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_72),
.Y(n_73)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_55),
.B(n_51),
.Y(n_71)
);

NOR4xp25_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_57),
.C(n_61),
.D(n_63),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_43),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_74),
.A2(n_69),
.B(n_27),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_57),
.B1(n_60),
.B2(n_29),
.Y(n_76)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_69),
.B1(n_72),
.B2(n_66),
.Y(n_78)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_77),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_27),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_73),
.C(n_77),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_83),
.B(n_84),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_75),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_80),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_84),
.B(n_82),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_86),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_89),
.A2(n_9),
.B(n_29),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_90),
.B(n_29),
.Y(n_91)
);


endmodule