module fake_jpeg_7078_n_80 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_80);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_80;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_8;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_1),
.B(n_6),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_7),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_7),
.B(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_15),
.B1(n_8),
.B2(n_11),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_21),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_14),
.B(n_2),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_21),
.B(n_14),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_13),
.C(n_11),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_18),
.B(n_13),
.Y(n_29)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_17),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g28 ( 
.A(n_24),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_30),
.B(n_6),
.Y(n_45)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_12),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_23),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_34),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_23),
.A2(n_8),
.B1(n_15),
.B2(n_26),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_35),
.A2(n_20),
.B1(n_26),
.B2(n_9),
.Y(n_44)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_44),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_41),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_30),
.B(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_31),
.B1(n_33),
.B2(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_52),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_49),
.B(n_53),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_24),
.C(n_17),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_55),
.B(n_3),
.Y(n_63)
);

NOR3xp33_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_43),
.C(n_39),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_57),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_50),
.C(n_48),
.Y(n_64)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

AOI221xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_24),
.B1(n_19),
.B2(n_4),
.C(n_3),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_61),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_49),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_58),
.B(n_62),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_60),
.B1(n_56),
.B2(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_65),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_70),
.A2(n_64),
.B(n_68),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_66),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_72),
.A2(n_73),
.B1(n_54),
.B2(n_38),
.Y(n_75)
);

OAI21x1_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_24),
.B(n_4),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_76),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_78),
.B(n_4),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_19),
.Y(n_80)
);


endmodule