module fake_aes_7297_n_26 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_26);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_26;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
INVx1_ASAP7_75t_L g13 ( .A(n_9), .Y(n_13) );
NOR2x1_ASAP7_75t_L g14 ( .A(n_1), .B(n_3), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_12), .Y(n_15) );
OAI21x1_ASAP7_75t_L g16 ( .A1(n_0), .A2(n_4), .B(n_8), .Y(n_16) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_0), .Y(n_17) );
AOI21xp5_ASAP7_75t_L g18 ( .A1(n_13), .A2(n_5), .B(n_6), .Y(n_18) );
AOI21x1_ASAP7_75t_L g19 ( .A1(n_15), .A2(n_7), .B(n_10), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_20), .B(n_18), .Y(n_21) );
BUFx6f_ASAP7_75t_SL g22 ( .A(n_21), .Y(n_22) );
NOR4xp75_ASAP7_75t_SL g23 ( .A(n_22), .B(n_16), .C(n_2), .D(n_1), .Y(n_23) );
CKINVDCx5p33_ASAP7_75t_R g24 ( .A(n_23), .Y(n_24) );
OAI22x1_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_17), .B1(n_23), .B2(n_14), .Y(n_25) );
AOI22xp5_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_17), .B1(n_2), .B2(n_11), .Y(n_26) );
endmodule