module fake_jpeg_7646_n_208 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_208);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_13),
.B(n_6),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_32),
.Y(n_39)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_34),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_36),
.B(n_21),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_12),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_16),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_15),
.B1(n_17),
.B2(n_24),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_38),
.A2(n_42),
.B1(n_26),
.B2(n_18),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_29),
.A2(n_15),
.B1(n_16),
.B2(n_24),
.Y(n_42)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_50),
.B(n_10),
.Y(n_63)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_52),
.B(n_19),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_54),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_27),
.B(n_0),
.Y(n_54)
);

OAI32xp33_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_30),
.A3(n_20),
.B1(n_25),
.B2(n_28),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_55),
.A2(n_62),
.B1(n_70),
.B2(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_57),
.Y(n_72)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVxp67_ASAP7_75t_SL g85 ( 
.A(n_58),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_43),
.B(n_19),
.Y(n_60)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_63),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_20),
.B1(n_26),
.B2(n_18),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_41),
.A2(n_25),
.B1(n_20),
.B2(n_7),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_64),
.A2(n_47),
.B1(n_46),
.B2(n_49),
.Y(n_86)
);

NAND3xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_54),
.C(n_53),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_7),
.C(n_12),
.Y(n_79)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_44),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_41),
.A2(n_20),
.B1(n_28),
.B2(n_2),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_65),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_73),
.B(n_77),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_43),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_82),
.Y(n_90)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_85),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_68),
.Y(n_77)
);

OR2x6_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_66),
.Y(n_101)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_69),
.B1(n_55),
.B2(n_42),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_45),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_62),
.A2(n_45),
.B(n_39),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_86),
.B(n_56),
.C(n_57),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_48),
.Y(n_87)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_91),
.A2(n_92),
.B1(n_104),
.B2(n_57),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_67),
.B1(n_61),
.B2(n_71),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_94),
.B(n_95),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_87),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_72),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_74),
.Y(n_111)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_75),
.B(n_59),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_99),
.A2(n_101),
.B(n_102),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_71),
.B(n_39),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_60),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_82),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_73),
.A2(n_71),
.B1(n_70),
.B2(n_68),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_84),
.B1(n_83),
.B2(n_75),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_81),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_107),
.C(n_119),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_90),
.C(n_95),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_77),
.Y(n_109)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_113),
.Y(n_131)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_89),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_93),
.B(n_78),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_114),
.B(n_117),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_85),
.Y(n_116)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_118),
.A2(n_120),
.B(n_105),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_72),
.C(n_78),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_91),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_101),
.C(n_104),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_122),
.B(n_82),
.Y(n_134)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_117),
.A2(n_105),
.B1(n_96),
.B2(n_100),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_126),
.A2(n_49),
.B1(n_76),
.B2(n_28),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_101),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_137),
.C(n_138),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_94),
.Y(n_128)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_129),
.A2(n_132),
.B1(n_135),
.B2(n_123),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_121),
.Y(n_130)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_118),
.A2(n_101),
.B1(n_105),
.B2(n_104),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_139),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_105),
.B1(n_104),
.B2(n_101),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_101),
.C(n_88),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_108),
.B(n_88),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_110),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_147),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_144),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_136),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_152),
.C(n_153),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_127),
.B(n_115),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_132),
.A2(n_120),
.B1(n_115),
.B2(n_79),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_145),
.A2(n_151),
.B1(n_128),
.B2(n_34),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_124),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_133),
.A2(n_122),
.B1(n_97),
.B2(n_76),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_154),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_114),
.C(n_88),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_49),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_8),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_164),
.Y(n_173)
);

AOI321xp33_ASAP7_75t_L g158 ( 
.A1(n_150),
.A2(n_128),
.A3(n_34),
.B1(n_32),
.B2(n_31),
.C(n_4),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_11),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_154),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_162),
.A2(n_3),
.B(n_5),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_9),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_34),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_31),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_10),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_167),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_7),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_163),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_155),
.B(n_149),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_169),
.A2(n_3),
.B(n_6),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_179),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_144),
.C(n_145),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_176),
.C(n_177),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_178),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_34),
.C(n_32),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_156),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_158),
.C(n_31),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_160),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_180),
.A2(n_182),
.B(n_1),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_162),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_185),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_161),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_177),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_170),
.A2(n_3),
.B1(n_6),
.B2(n_11),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_187),
.B(n_1),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_172),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_176),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_191),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_193),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_192),
.B(n_32),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_1),
.C(n_32),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_195),
.A2(n_183),
.B(n_31),
.Y(n_196)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_196),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_199),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_194),
.B(n_195),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_200),
.B(n_190),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_202),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_203),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_201),
.C(n_197),
.Y(n_206)
);

BUFx24_ASAP7_75t_SL g207 ( 
.A(n_206),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_204),
.Y(n_208)
);


endmodule