module fake_jpeg_2053_n_51 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_51);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_51;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_5),
.B(n_2),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_2),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_21),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_9),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_18),
.A2(n_19),
.B1(n_26),
.B2(n_20),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_8),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_23),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_11),
.A2(n_1),
.B(n_7),
.C(n_13),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

NOR2x1p5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_25),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_15),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_10),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_19),
.A2(n_10),
.B1(n_14),
.B2(n_23),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_29),
.B1(n_33),
.B2(n_20),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_17),
.A2(n_14),
.B1(n_24),
.B2(n_21),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_34),
.B(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_30),
.B(n_28),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

AO22x1_ASAP7_75t_SL g37 ( 
.A1(n_33),
.A2(n_27),
.B1(n_32),
.B2(n_22),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_37),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_27),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_32),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_38),
.A2(n_34),
.B1(n_37),
.B2(n_36),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_44),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_41),
.B(n_32),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_44),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_48),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_42),
.Y(n_48)
);

AOI321xp33_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_29),
.A3(n_31),
.B1(n_37),
.B2(n_38),
.C(n_30),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_37),
.Y(n_51)
);


endmodule