module fake_jpeg_8186_n_52 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_52);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_52;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_24;
wire n_26;
wire n_36;
wire n_17;
wire n_31;
wire n_25;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_12),
.B(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_3),
.B(n_11),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_13),
.Y(n_26)
);

INVx3_ASAP7_75t_SL g27 ( 
.A(n_0),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_5),
.B(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx4_ASAP7_75t_SL g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_20),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_35),
.C(n_36),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_10),
.B1(n_21),
.B2(n_19),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_33),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_31),
.Y(n_39)
);

OR2x4_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_16),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_25),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_40),
.C(n_29),
.Y(n_45)
);

NOR3xp33_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_46),
.C(n_38),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_36),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_40),
.B1(n_41),
.B2(n_24),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_48),
.B1(n_22),
.B2(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_49),
.B(n_23),
.Y(n_50)
);

AOI322xp5_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_21),
.A3(n_26),
.B1(n_32),
.B2(n_18),
.C1(n_42),
.C2(n_37),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_32),
.C(n_26),
.Y(n_52)
);


endmodule