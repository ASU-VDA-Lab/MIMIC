module fake_ariane_393_n_2019 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2019);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2019;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_967;
wire n_274;
wire n_337;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_928;
wire n_253;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_136),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_104),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_2),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_54),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_75),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_35),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_105),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_91),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_51),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_48),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_192),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_112),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_132),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_89),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_27),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_150),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_65),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g213 ( 
.A(n_118),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g214 ( 
.A(n_2),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_115),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_45),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_160),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_191),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_31),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_177),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_155),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_8),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_61),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_123),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_23),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_83),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_21),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_106),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_12),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_48),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_121),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_181),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_142),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_31),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_159),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_76),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_37),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_64),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_43),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_3),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_100),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_39),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_145),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_87),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_124),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_97),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_81),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_164),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_90),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_92),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_73),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_157),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_175),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_133),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_190),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_163),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_152),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_82),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_126),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_149),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_36),
.Y(n_261)
);

BUFx10_ASAP7_75t_L g262 ( 
.A(n_169),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_30),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_67),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_10),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_18),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_32),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_60),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_38),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_36),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_189),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_114),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_1),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_173),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_171),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_53),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_96),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_21),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_6),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_166),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_70),
.Y(n_281)
);

BUFx10_ASAP7_75t_L g282 ( 
.A(n_45),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_11),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_130),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_40),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_78),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_1),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_16),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_59),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_139),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_7),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_49),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_188),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_128),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_101),
.Y(n_295)
);

BUFx10_ASAP7_75t_L g296 ( 
.A(n_46),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_156),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_27),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_24),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_15),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_18),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_16),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_24),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_174),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_193),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_111),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_144),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_143),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_108),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_183),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_88),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_46),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_32),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_44),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_56),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_60),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_116),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_176),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_69),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_57),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_70),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_19),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_110),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_13),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_85),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_25),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_68),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_137),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_147),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_134),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_84),
.Y(n_331)
);

BUFx5_ASAP7_75t_L g332 ( 
.A(n_57),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_99),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_138),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_64),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_3),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_135),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_65),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_117),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_12),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_41),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_113),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_58),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_161),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_13),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_153),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_151),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_0),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_148),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_98),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_80),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_68),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_11),
.Y(n_353)
);

INVx4_ASAP7_75t_R g354 ( 
.A(n_102),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_75),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_178),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_131),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_37),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_67),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_42),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_120),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_17),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_51),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_47),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_47),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_154),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_26),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_179),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_52),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_17),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_180),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_29),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_58),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_14),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_15),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_52),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_93),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_71),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_6),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_69),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_44),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_28),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_158),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_127),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_74),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_22),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_19),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_172),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_332),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_332),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_207),
.B(n_0),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_276),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_332),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_332),
.B(n_4),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_332),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_332),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_195),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_332),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_208),
.Y(n_399)
);

INVxp33_ASAP7_75t_SL g400 ( 
.A(n_263),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_332),
.Y(n_401)
);

INVxp33_ASAP7_75t_SL g402 ( 
.A(n_199),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_217),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_218),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_226),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_332),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_255),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_310),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_344),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_385),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_385),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_207),
.Y(n_412)
);

INVxp67_ASAP7_75t_SL g413 ( 
.A(n_267),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_268),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_350),
.Y(n_415)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_267),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_209),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_209),
.B(n_4),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_377),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_205),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_273),
.Y(n_421)
);

BUFx10_ASAP7_75t_L g422 ( 
.A(n_274),
.Y(n_422)
);

INVxp67_ASAP7_75t_SL g423 ( 
.A(n_273),
.Y(n_423)
);

CKINVDCx14_ASAP7_75t_R g424 ( 
.A(n_262),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_215),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_210),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_215),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_221),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_204),
.Y(n_429)
);

BUFx6f_ASAP7_75t_SL g430 ( 
.A(n_262),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_270),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_307),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_221),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_228),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_287),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_228),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_235),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_212),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_291),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_R g440 ( 
.A(n_388),
.B(n_196),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g441 ( 
.A(n_262),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_216),
.Y(n_442)
);

NOR2xp67_ASAP7_75t_L g443 ( 
.A(n_198),
.B(n_5),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_325),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_235),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_245),
.Y(n_446)
);

NOR2xp67_ASAP7_75t_L g447 ( 
.A(n_198),
.B(n_5),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_320),
.Y(n_448)
);

INVxp67_ASAP7_75t_SL g449 ( 
.A(n_336),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_222),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_245),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_225),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_246),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_227),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_272),
.B(n_7),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_369),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_246),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_247),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_230),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_247),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_336),
.Y(n_461)
);

INVxp67_ASAP7_75t_SL g462 ( 
.A(n_268),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_248),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_268),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_248),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_268),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_258),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_258),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_259),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_238),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_197),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_259),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g473 ( 
.A(n_268),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_271),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_301),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_271),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_277),
.B(n_284),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_239),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_240),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_277),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_284),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_242),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_290),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_381),
.Y(n_484)
);

OA21x2_ASAP7_75t_L g485 ( 
.A1(n_394),
.A2(n_329),
.B(n_290),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_389),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_432),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_389),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_432),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_444),
.B(n_422),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_432),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_390),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_390),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_411),
.Y(n_494)
);

CKINVDCx11_ASAP7_75t_R g495 ( 
.A(n_429),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_475),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_475),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_462),
.B(n_329),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_393),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_475),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g501 ( 
.A(n_441),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_475),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_400),
.A2(n_410),
.B1(n_441),
.B2(n_455),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_396),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_432),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_432),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_393),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_432),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_479),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_395),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_392),
.B(n_219),
.Y(n_511)
);

NAND2xp33_ASAP7_75t_L g512 ( 
.A(n_412),
.B(n_301),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_410),
.B(n_229),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_396),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_412),
.B(n_301),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_395),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_398),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_399),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_471),
.A2(n_223),
.B1(n_313),
.B2(n_229),
.Y(n_519)
);

NAND2xp33_ASAP7_75t_R g520 ( 
.A(n_420),
.B(n_387),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_398),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_401),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_401),
.Y(n_523)
);

NAND2xp33_ASAP7_75t_L g524 ( 
.A(n_417),
.B(n_301),
.Y(n_524)
);

OA21x2_ASAP7_75t_L g525 ( 
.A1(n_417),
.A2(n_339),
.B(n_331),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_461),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_473),
.B(n_331),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_406),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_477),
.B(n_339),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_406),
.Y(n_530)
);

BUFx8_ASAP7_75t_L g531 ( 
.A(n_430),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_392),
.B(n_219),
.Y(n_532)
);

BUFx8_ASAP7_75t_L g533 ( 
.A(n_430),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_444),
.B(n_301),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_414),
.Y(n_535)
);

OA21x2_ASAP7_75t_L g536 ( 
.A1(n_425),
.A2(n_366),
.B(n_361),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_425),
.B(n_361),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_414),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_427),
.B(n_366),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_464),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_427),
.B(n_300),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_464),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_466),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_466),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_428),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_428),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_433),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_422),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_433),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_434),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_434),
.B(n_368),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_422),
.B(n_201),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_436),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_436),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_SL g555 ( 
.A(n_430),
.B(n_214),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_437),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_437),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_445),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_445),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_446),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_446),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_451),
.B(n_453),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_451),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_453),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_530),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_554),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_554),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_517),
.Y(n_568)
);

INVx5_ASAP7_75t_L g569 ( 
.A(n_487),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_530),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_554),
.Y(n_571)
);

NAND2xp33_ASAP7_75t_L g572 ( 
.A(n_548),
.B(n_426),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_485),
.A2(n_418),
.B1(n_391),
.B2(n_443),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_530),
.Y(n_574)
);

INVxp67_ASAP7_75t_SL g575 ( 
.A(n_537),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_517),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_490),
.B(n_438),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_519),
.A2(n_447),
.B1(n_313),
.B2(n_251),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_554),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_530),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_554),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_485),
.A2(n_519),
.B1(n_534),
.B2(n_525),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_517),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_562),
.B(n_413),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g585 ( 
.A(n_494),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_554),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_517),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_526),
.B(n_407),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_554),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_521),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_548),
.B(n_402),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_485),
.A2(n_458),
.B1(n_460),
.B2(n_457),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_548),
.B(n_490),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_554),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_485),
.A2(n_458),
.B1(n_460),
.B2(n_457),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_555),
.A2(n_265),
.B1(n_269),
.B2(n_266),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_564),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_564),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_521),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_521),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_564),
.Y(n_601)
);

NAND2xp33_ASAP7_75t_L g602 ( 
.A(n_529),
.B(n_564),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_564),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_564),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_521),
.Y(n_605)
);

BUFx8_ASAP7_75t_SL g606 ( 
.A(n_518),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_504),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_494),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_504),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_504),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_534),
.B(n_424),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_504),
.Y(n_612)
);

BUFx6f_ASAP7_75t_SL g613 ( 
.A(n_531),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_555),
.B(n_442),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_504),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_514),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_562),
.B(n_416),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_485),
.A2(n_465),
.B1(n_467),
.B2(n_463),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_495),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_552),
.B(n_450),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_564),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_485),
.A2(n_465),
.B1(n_467),
.B2(n_463),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_516),
.Y(n_623)
);

CKINVDCx16_ASAP7_75t_R g624 ( 
.A(n_501),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_564),
.Y(n_625)
);

BUFx8_ASAP7_75t_SL g626 ( 
.A(n_518),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_509),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_560),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_513),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_530),
.Y(n_630)
);

BUFx2_ASAP7_75t_L g631 ( 
.A(n_509),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_514),
.Y(n_632)
);

BUFx2_ASAP7_75t_L g633 ( 
.A(n_526),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_495),
.Y(n_634)
);

AND2x6_ASAP7_75t_L g635 ( 
.A(n_562),
.B(n_368),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_513),
.B(n_452),
.Y(n_636)
);

BUFx4f_ASAP7_75t_L g637 ( 
.A(n_525),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_516),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_560),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_525),
.A2(n_469),
.B1(n_472),
.B2(n_468),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_560),
.Y(n_641)
);

INVx4_ASAP7_75t_L g642 ( 
.A(n_525),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_561),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_561),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_516),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_513),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_516),
.Y(n_647)
);

INVx4_ASAP7_75t_L g648 ( 
.A(n_525),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_561),
.Y(n_649)
);

OAI22x1_ASAP7_75t_L g650 ( 
.A1(n_503),
.A2(n_415),
.B1(n_419),
.B2(n_409),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_516),
.Y(n_651)
);

INVx1_ASAP7_75t_SL g652 ( 
.A(n_501),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_503),
.A2(n_278),
.B1(n_288),
.B2(n_279),
.Y(n_653)
);

AO22x2_ASAP7_75t_L g654 ( 
.A1(n_529),
.A2(n_468),
.B1(n_472),
.B2(n_469),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_516),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_516),
.Y(n_656)
);

BUFx8_ASAP7_75t_SL g657 ( 
.A(n_511),
.Y(n_657)
);

BUFx6f_ASAP7_75t_SL g658 ( 
.A(n_531),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_563),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_552),
.B(n_454),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_516),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_486),
.B(n_474),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_486),
.Y(n_663)
);

AND2x6_ASAP7_75t_L g664 ( 
.A(n_515),
.B(n_371),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_563),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_486),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_541),
.B(n_421),
.Y(n_667)
);

INVx5_ASAP7_75t_L g668 ( 
.A(n_487),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_488),
.Y(n_669)
);

INVxp67_ASAP7_75t_SL g670 ( 
.A(n_514),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_488),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_563),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_488),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_492),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_514),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_492),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_531),
.B(n_459),
.Y(n_677)
);

NAND3xp33_ASAP7_75t_SL g678 ( 
.A(n_537),
.B(n_478),
.C(n_470),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_498),
.B(n_482),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_545),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_531),
.B(n_440),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_492),
.Y(n_682)
);

NAND2xp33_ASAP7_75t_L g683 ( 
.A(n_549),
.B(n_474),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_531),
.B(n_422),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_541),
.B(n_423),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_545),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_493),
.B(n_476),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_493),
.B(n_476),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_531),
.B(n_480),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_493),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_499),
.B(n_480),
.Y(n_691)
);

XOR2xp5_ASAP7_75t_L g692 ( 
.A(n_511),
.B(n_397),
.Y(n_692)
);

HB1xp67_ASAP7_75t_L g693 ( 
.A(n_520),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_499),
.B(n_481),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_499),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_533),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_507),
.B(n_481),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_545),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_498),
.B(n_449),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_514),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_514),
.Y(n_701)
);

INVxp67_ASAP7_75t_SL g702 ( 
.A(n_514),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_545),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_507),
.B(n_483),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_546),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_507),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_510),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_546),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_511),
.B(n_483),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_514),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_546),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_541),
.B(n_214),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_533),
.B(n_289),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_510),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_546),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_547),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_547),
.Y(n_717)
);

BUFx6f_ASAP7_75t_SL g718 ( 
.A(n_629),
.Y(n_718)
);

BUFx5_ASAP7_75t_L g719 ( 
.A(n_565),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_593),
.B(n_533),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_663),
.Y(n_721)
);

A2O1A1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_575),
.A2(n_550),
.B(n_549),
.C(n_522),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_628),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_575),
.B(n_533),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_679),
.B(n_533),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_637),
.B(n_510),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_699),
.B(n_533),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_628),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_591),
.B(n_550),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_584),
.B(n_532),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_637),
.B(n_522),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_584),
.B(n_532),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_629),
.B(n_527),
.Y(n_733)
);

OAI221xp5_ASAP7_75t_L g734 ( 
.A1(n_578),
.A2(n_520),
.B1(n_237),
.B2(n_319),
.C(n_261),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_639),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_584),
.B(n_611),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_637),
.B(n_522),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_627),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_646),
.A2(n_551),
.B1(n_539),
.B2(n_547),
.Y(n_739)
);

AND2x4_ASAP7_75t_L g740 ( 
.A(n_584),
.B(n_532),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_639),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_637),
.B(n_523),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_565),
.B(n_523),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_641),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_616),
.Y(n_745)
);

OR2x2_ASAP7_75t_L g746 ( 
.A(n_627),
.B(n_527),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_620),
.B(n_528),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_660),
.B(n_528),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_565),
.B(n_523),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_616),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_669),
.Y(n_751)
);

OAI22xp33_ASAP7_75t_L g752 ( 
.A1(n_596),
.A2(n_551),
.B1(n_539),
.B2(n_321),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_635),
.A2(n_525),
.B1(n_536),
.B2(n_547),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_712),
.B(n_553),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_663),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_666),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_646),
.B(n_553),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_712),
.B(n_553),
.Y(n_758)
);

A2O1A1Ixp33_ASAP7_75t_L g759 ( 
.A1(n_573),
.A2(n_553),
.B(n_557),
.C(n_556),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_617),
.B(n_556),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_617),
.B(n_556),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_667),
.B(n_556),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_667),
.B(n_685),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_570),
.B(n_557),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_570),
.B(n_557),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_685),
.B(n_557),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_SL g767 ( 
.A1(n_653),
.A2(n_435),
.B1(n_439),
.B2(n_431),
.Y(n_767)
);

OR2x2_ASAP7_75t_L g768 ( 
.A(n_631),
.B(n_633),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_635),
.B(n_558),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_635),
.B(n_558),
.Y(n_770)
);

HB1xp67_ASAP7_75t_L g771 ( 
.A(n_633),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_570),
.B(n_558),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_693),
.B(n_403),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_574),
.B(n_558),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_635),
.B(n_559),
.Y(n_775)
);

NAND2xp33_ASAP7_75t_SL g776 ( 
.A(n_613),
.B(n_559),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_641),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_635),
.B(n_559),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_635),
.B(n_559),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_635),
.B(n_515),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_670),
.A2(n_536),
.B(n_497),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_635),
.B(n_515),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_572),
.B(n_515),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_643),
.Y(n_784)
);

A2O1A1Ixp33_ASAP7_75t_L g785 ( 
.A1(n_643),
.A2(n_515),
.B(n_496),
.C(n_500),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_577),
.B(n_515),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_644),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_631),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_574),
.B(n_371),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_616),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_644),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_649),
.Y(n_792)
);

NOR3xp33_ASAP7_75t_L g793 ( 
.A(n_636),
.B(n_200),
.C(n_197),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_574),
.B(n_496),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_709),
.B(n_536),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_580),
.B(n_497),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_649),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_673),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_616),
.Y(n_799)
);

NOR2xp67_ASAP7_75t_L g800 ( 
.A(n_596),
.B(n_535),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_659),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_659),
.Y(n_802)
);

NAND3xp33_ASAP7_75t_L g803 ( 
.A(n_653),
.B(n_298),
.C(n_292),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_585),
.B(n_404),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_665),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_709),
.B(n_536),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_673),
.Y(n_807)
);

AOI22xp5_ASAP7_75t_L g808 ( 
.A1(n_678),
.A2(n_536),
.B1(n_274),
.B2(n_328),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_580),
.B(n_500),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_669),
.B(n_536),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_669),
.B(n_502),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_614),
.B(n_299),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_671),
.B(n_502),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_671),
.B(n_323),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_678),
.B(n_303),
.Y(n_815)
);

INVxp67_ASAP7_75t_L g816 ( 
.A(n_692),
.Y(n_816)
);

OAI22xp33_ASAP7_75t_L g817 ( 
.A1(n_578),
.A2(n_358),
.B1(n_321),
.B2(n_335),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_671),
.B(n_662),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_662),
.B(n_357),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_665),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_608),
.B(n_405),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_673),
.Y(n_822)
);

INVx4_ASAP7_75t_L g823 ( 
.A(n_613),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_580),
.B(n_201),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_588),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_630),
.B(n_280),
.Y(n_826)
);

BUFx5_ASAP7_75t_L g827 ( 
.A(n_630),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_624),
.B(n_312),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_606),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_672),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_687),
.B(n_535),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_642),
.A2(n_491),
.B(n_489),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_672),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_687),
.B(n_535),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_624),
.B(n_314),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_680),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_674),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_688),
.B(n_691),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_688),
.B(n_691),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_683),
.A2(n_524),
.B1(n_512),
.B2(n_408),
.Y(n_840)
);

INVxp67_ASAP7_75t_L g841 ( 
.A(n_692),
.Y(n_841)
);

INVx4_ASAP7_75t_L g842 ( 
.A(n_613),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_696),
.B(n_315),
.Y(n_843)
);

OR2x6_ASAP7_75t_L g844 ( 
.A(n_650),
.B(n_300),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_694),
.B(n_535),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_694),
.B(n_697),
.Y(n_846)
);

NAND2xp33_ASAP7_75t_SL g847 ( 
.A(n_613),
.B(n_316),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_630),
.B(n_280),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_697),
.B(n_535),
.Y(n_849)
);

NAND2xp33_ASAP7_75t_L g850 ( 
.A(n_674),
.B(n_324),
.Y(n_850)
);

OR2x2_ASAP7_75t_L g851 ( 
.A(n_588),
.B(n_448),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_674),
.Y(n_852)
);

NAND2xp33_ASAP7_75t_L g853 ( 
.A(n_676),
.B(n_326),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_704),
.B(n_544),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_704),
.B(n_544),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_654),
.A2(n_358),
.B1(n_335),
.B2(n_348),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_642),
.B(n_295),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_642),
.B(n_295),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_680),
.Y(n_859)
);

BUFx2_ASAP7_75t_L g860 ( 
.A(n_657),
.Y(n_860)
);

OR2x6_ASAP7_75t_SL g861 ( 
.A(n_626),
.B(n_338),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_676),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_686),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_686),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_582),
.B(n_544),
.Y(n_865)
);

OAI22xp33_ASAP7_75t_L g866 ( 
.A1(n_652),
.A2(n_355),
.B1(n_234),
.B2(n_237),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_676),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_592),
.B(n_544),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_677),
.B(n_340),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_664),
.A2(n_512),
.B1(n_524),
.B2(n_254),
.Y(n_870)
);

INVxp67_ASAP7_75t_L g871 ( 
.A(n_652),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_616),
.Y(n_872)
);

NOR2xp67_ASAP7_75t_L g873 ( 
.A(n_696),
.B(n_544),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_698),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_698),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_642),
.B(n_304),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_682),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_654),
.A2(n_648),
.B1(n_664),
.B2(n_618),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_682),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_648),
.B(n_304),
.Y(n_880)
);

AOI22xp5_ASAP7_75t_L g881 ( 
.A1(n_664),
.A2(n_252),
.B1(n_257),
.B2(n_256),
.Y(n_881)
);

INVxp67_ASAP7_75t_L g882 ( 
.A(n_650),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_654),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_713),
.B(n_341),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_682),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_595),
.B(n_540),
.Y(n_886)
);

INVxp33_ASAP7_75t_L g887 ( 
.A(n_619),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_838),
.A2(n_702),
.B(n_602),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_747),
.A2(n_690),
.B1(n_706),
.B2(n_695),
.Y(n_889)
);

OAI21xp33_ASAP7_75t_L g890 ( 
.A1(n_729),
.A2(n_733),
.B(n_815),
.Y(n_890)
);

AOI21x1_ASAP7_75t_L g891 ( 
.A1(n_857),
.A2(n_705),
.B(n_703),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_723),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_719),
.B(n_648),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_733),
.B(n_622),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_763),
.A2(n_664),
.B1(n_684),
.B2(n_681),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_757),
.B(n_654),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_829),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_757),
.B(n_654),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_736),
.B(n_640),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_738),
.B(n_456),
.Y(n_900)
);

AO21x2_ASAP7_75t_L g901 ( 
.A1(n_865),
.A2(n_689),
.B(n_703),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_839),
.A2(n_710),
.B(n_700),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_748),
.A2(n_690),
.B1(n_706),
.B2(n_695),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_771),
.Y(n_904)
);

NOR2x1_ASAP7_75t_L g905 ( 
.A(n_746),
.B(n_648),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_721),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_L g907 ( 
.A1(n_856),
.A2(n_664),
.B1(n_695),
.B2(n_690),
.Y(n_907)
);

O2A1O1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_752),
.A2(n_706),
.B(n_714),
.C(n_707),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_788),
.B(n_707),
.Y(n_909)
);

A2O1A1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_815),
.A2(n_707),
.B(n_714),
.C(n_708),
.Y(n_910)
);

INVx1_ASAP7_75t_SL g911 ( 
.A(n_768),
.Y(n_911)
);

INVxp67_ASAP7_75t_L g912 ( 
.A(n_771),
.Y(n_912)
);

NOR3xp33_ASAP7_75t_L g913 ( 
.A(n_825),
.B(n_234),
.C(n_200),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_719),
.B(n_714),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_730),
.B(n_716),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_L g916 ( 
.A1(n_832),
.A2(n_576),
.B(n_568),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_732),
.B(n_716),
.Y(n_917)
);

OAI21x1_ASAP7_75t_L g918 ( 
.A1(n_781),
.A2(n_638),
.B(n_623),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_846),
.A2(n_710),
.B(n_700),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_719),
.B(n_616),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_728),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_735),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_726),
.A2(n_710),
.B(n_700),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_754),
.B(n_664),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_726),
.A2(n_710),
.B(n_700),
.Y(n_925)
);

OAI21xp5_ASAP7_75t_L g926 ( 
.A1(n_810),
.A2(n_576),
.B(n_568),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_741),
.Y(n_927)
);

NAND3xp33_ASAP7_75t_SL g928 ( 
.A(n_734),
.B(n_634),
.C(n_484),
.Y(n_928)
);

A2O1A1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_786),
.A2(n_716),
.B(n_708),
.C(n_711),
.Y(n_929)
);

BUFx2_ASAP7_75t_L g930 ( 
.A(n_804),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_758),
.B(n_664),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_740),
.B(n_871),
.Y(n_932)
);

OAI321xp33_ASAP7_75t_L g933 ( 
.A1(n_817),
.A2(n_319),
.A3(n_360),
.B1(n_363),
.B2(n_372),
.C(n_302),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_744),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_740),
.A2(n_664),
.B1(n_716),
.B2(n_711),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_731),
.A2(n_638),
.B(n_623),
.Y(n_936)
);

A2O1A1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_777),
.A2(n_715),
.B(n_717),
.C(n_705),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_819),
.B(n_715),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_755),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_756),
.Y(n_940)
);

O2A1O1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_752),
.A2(n_717),
.B(n_609),
.C(n_610),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_745),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_786),
.A2(n_609),
.B(n_610),
.C(n_607),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_760),
.B(n_607),
.Y(n_944)
);

AO21x1_ASAP7_75t_L g945 ( 
.A1(n_725),
.A2(n_567),
.B(n_566),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_784),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_761),
.B(n_607),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_808),
.A2(n_609),
.B(n_610),
.C(n_612),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_787),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_818),
.A2(n_751),
.B1(n_792),
.B2(n_791),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_821),
.B(n_773),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_773),
.B(n_214),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_737),
.A2(n_647),
.B(n_645),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_851),
.B(n_282),
.Y(n_954)
);

NOR2x1p5_ASAP7_75t_L g955 ( 
.A(n_803),
.B(n_261),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_762),
.B(n_612),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_751),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_766),
.B(n_612),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_742),
.A2(n_647),
.B(n_645),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_739),
.B(n_615),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_742),
.A2(n_655),
.B(n_651),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_767),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_823),
.B(n_615),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_831),
.A2(n_655),
.B(n_651),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_797),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_719),
.B(n_632),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_801),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_802),
.Y(n_968)
);

INVxp67_ASAP7_75t_SL g969 ( 
.A(n_795),
.Y(n_969)
);

O2A1O1Ixp5_ASAP7_75t_L g970 ( 
.A1(n_720),
.A2(n_599),
.B(n_583),
.C(n_587),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_745),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_798),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_745),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_834),
.A2(n_655),
.B(n_651),
.Y(n_974)
);

AOI21x1_ASAP7_75t_L g975 ( 
.A1(n_857),
.A2(n_567),
.B(n_566),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_719),
.B(n_632),
.Y(n_976)
);

AO21x1_ASAP7_75t_L g977 ( 
.A1(n_858),
.A2(n_579),
.B(n_571),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_845),
.A2(n_656),
.B(n_661),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_849),
.A2(n_656),
.B(n_661),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_805),
.Y(n_980)
);

NOR2xp67_ASAP7_75t_L g981 ( 
.A(n_869),
.B(n_615),
.Y(n_981)
);

INVx4_ASAP7_75t_L g982 ( 
.A(n_718),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_854),
.A2(n_656),
.B(n_661),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_814),
.B(n_568),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_855),
.A2(n_661),
.B(n_583),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_858),
.A2(n_583),
.B(n_576),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_743),
.A2(n_590),
.B(n_587),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_727),
.B(n_587),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_743),
.A2(n_599),
.B(n_590),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_745),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_869),
.B(n_590),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_749),
.A2(n_600),
.B(n_599),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_820),
.B(n_600),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_750),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_830),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_750),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_749),
.A2(n_605),
.B(n_600),
.Y(n_997)
);

INVx2_ASAP7_75t_SL g998 ( 
.A(n_860),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_816),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_833),
.B(n_605),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_806),
.A2(n_605),
.B(n_579),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_876),
.A2(n_880),
.B(n_813),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_718),
.B(n_581),
.Y(n_1003)
);

OAI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_876),
.A2(n_586),
.B(n_571),
.Y(n_1004)
);

INVx3_ASAP7_75t_L g1005 ( 
.A(n_750),
.Y(n_1005)
);

AOI33xp33_ASAP7_75t_L g1006 ( 
.A1(n_817),
.A2(n_283),
.A3(n_281),
.B1(n_285),
.B2(n_302),
.B3(n_322),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_750),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_724),
.B(n_581),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_841),
.B(n_282),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_880),
.A2(n_589),
.B(n_586),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_SL g1011 ( 
.A(n_887),
.B(n_658),
.Y(n_1011)
);

OR2x6_ASAP7_75t_L g1012 ( 
.A(n_883),
.B(n_844),
.Y(n_1012)
);

INVx4_ASAP7_75t_L g1013 ( 
.A(n_790),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_884),
.B(n_812),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_823),
.B(n_581),
.Y(n_1015)
);

NOR2xp67_ASAP7_75t_L g1016 ( 
.A(n_884),
.B(n_581),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_836),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_811),
.A2(n_594),
.B(n_589),
.Y(n_1018)
);

NOR2x1_ASAP7_75t_L g1019 ( 
.A(n_800),
.B(n_597),
.Y(n_1019)
);

OAI21xp33_ASAP7_75t_L g1020 ( 
.A1(n_812),
.A2(n_353),
.B(n_345),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_859),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_764),
.A2(n_598),
.B(n_594),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_764),
.A2(n_603),
.B(n_598),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_828),
.B(n_597),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_863),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_856),
.B(n_597),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_765),
.A2(n_604),
.B(n_603),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_765),
.A2(n_621),
.B(n_604),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_722),
.B(n_597),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_864),
.B(n_874),
.Y(n_1030)
);

O2A1O1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_772),
.A2(n_281),
.B(n_264),
.C(n_283),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_719),
.B(n_632),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_L g1033 ( 
.A1(n_878),
.A2(n_322),
.B1(n_264),
.B2(n_360),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_772),
.A2(n_625),
.B(n_621),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_878),
.A2(n_601),
.B1(n_625),
.B2(n_658),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_R g1036 ( 
.A(n_847),
.B(n_658),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_774),
.A2(n_796),
.B(n_794),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_774),
.A2(n_601),
.B(n_632),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_875),
.B(n_601),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_827),
.B(n_632),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_807),
.B(n_601),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_822),
.B(n_837),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_852),
.B(n_862),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_759),
.A2(n_374),
.B(n_327),
.C(n_343),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_753),
.A2(n_491),
.B(n_489),
.Y(n_1045)
);

INVx2_ASAP7_75t_SL g1046 ( 
.A(n_835),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_867),
.B(n_632),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_882),
.B(n_675),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_794),
.A2(n_701),
.B(n_675),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_789),
.A2(n_372),
.B(n_285),
.C(n_363),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_780),
.B(n_675),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_769),
.A2(n_355),
.B(n_327),
.C(n_374),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_782),
.B(n_675),
.Y(n_1053)
);

HB1xp67_ASAP7_75t_L g1054 ( 
.A(n_770),
.Y(n_1054)
);

INVxp33_ASAP7_75t_SL g1055 ( 
.A(n_840),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_877),
.B(n_675),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_879),
.B(n_675),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_885),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_827),
.B(n_701),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_796),
.B(n_701),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_809),
.A2(n_701),
.B(n_668),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_827),
.B(n_783),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_868),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_809),
.A2(n_701),
.B(n_668),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_789),
.A2(n_386),
.B(n_352),
.C(n_343),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_827),
.B(n_701),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_785),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_775),
.A2(n_668),
.B(n_569),
.Y(n_1068)
);

OAI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_753),
.A2(n_779),
.B(n_778),
.Y(n_1069)
);

A2O1A1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_850),
.A2(n_348),
.B(n_352),
.C(n_386),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_827),
.B(n_359),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_827),
.B(n_362),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_886),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_853),
.A2(n_311),
.B(n_342),
.C(n_380),
.Y(n_1074)
);

INVx4_ASAP7_75t_L g1075 ( 
.A(n_790),
.Y(n_1075)
);

O2A1O1Ixp5_ASAP7_75t_L g1076 ( 
.A1(n_824),
.A2(n_508),
.B(n_489),
.C(n_491),
.Y(n_1076)
);

INVx5_ASAP7_75t_L g1077 ( 
.A(n_942),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_1014),
.B(n_866),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_911),
.B(n_866),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_890),
.A2(n_881),
.B1(n_790),
.B2(n_872),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_909),
.B(n_793),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_918),
.A2(n_826),
.B(n_824),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_1055),
.B(n_843),
.Y(n_1083)
);

O2A1O1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_912),
.A2(n_848),
.B(n_826),
.C(n_844),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_1062),
.A2(n_799),
.B(n_790),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_969),
.B(n_799),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_1070),
.A2(n_848),
.B(n_844),
.C(n_342),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_969),
.B(n_799),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_894),
.B(n_799),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_904),
.B(n_861),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_904),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_909),
.A2(n_873),
.B(n_776),
.C(n_870),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_932),
.B(n_872),
.Y(n_1093)
);

INVx8_ASAP7_75t_L g1094 ( 
.A(n_897),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_900),
.B(n_872),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_888),
.A2(n_872),
.B(n_668),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_942),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_L g1098 ( 
.A1(n_928),
.A2(n_296),
.B1(n_282),
.B2(n_658),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_SL g1099 ( 
.A1(n_1003),
.A2(n_489),
.B(n_491),
.C(n_505),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1033),
.B(n_842),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_920),
.A2(n_668),
.B(n_569),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_SL g1102 ( 
.A1(n_1003),
.A2(n_505),
.B(n_506),
.C(n_508),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_906),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_1033),
.A2(n_378),
.B1(n_364),
.B2(n_365),
.Y(n_1104)
);

O2A1O1Ixp5_ASAP7_75t_L g1105 ( 
.A1(n_945),
.A2(n_842),
.B(n_505),
.C(n_506),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_920),
.A2(n_668),
.B(n_569),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_966),
.A2(n_668),
.B(n_569),
.Y(n_1107)
);

HB1xp67_ASAP7_75t_L g1108 ( 
.A(n_930),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_954),
.B(n_367),
.Y(n_1109)
);

INVx3_ASAP7_75t_L g1110 ( 
.A(n_1015),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_966),
.A2(n_569),
.B(n_505),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_1020),
.A2(n_311),
.B(n_325),
.C(n_538),
.Y(n_1112)
);

NAND3xp33_ASAP7_75t_L g1113 ( 
.A(n_1074),
.B(n_370),
.C(n_379),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_976),
.A2(n_569),
.B(n_506),
.Y(n_1114)
);

O2A1O1Ixp5_ASAP7_75t_SL g1115 ( 
.A1(n_976),
.A2(n_543),
.B(n_540),
.C(n_538),
.Y(n_1115)
);

AOI21xp33_ASAP7_75t_L g1116 ( 
.A1(n_896),
.A2(n_543),
.B(n_538),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_908),
.A2(n_373),
.B(n_375),
.C(n_376),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_942),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_915),
.A2(n_917),
.B(n_1053),
.C(n_1051),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_999),
.B(n_382),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_1070),
.A2(n_506),
.B(n_508),
.C(n_542),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1032),
.A2(n_569),
.B(n_508),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_892),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_951),
.B(n_296),
.Y(n_1124)
);

INVx4_ASAP7_75t_L g1125 ( 
.A(n_982),
.Y(n_1125)
);

O2A1O1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_910),
.A2(n_542),
.B(n_296),
.C(n_10),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1032),
.A2(n_297),
.B(n_203),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1040),
.A2(n_1066),
.B(n_1059),
.Y(n_1128)
);

BUFx8_ASAP7_75t_L g1129 ( 
.A(n_998),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_962),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_921),
.Y(n_1131)
);

OAI22x1_ASAP7_75t_L g1132 ( 
.A1(n_955),
.A2(n_294),
.B1(n_384),
.B2(n_383),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1040),
.A2(n_293),
.B(n_206),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_922),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_927),
.Y(n_1135)
);

NOR2xp67_ASAP7_75t_L g1136 ( 
.A(n_982),
.B(n_542),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_1009),
.B(n_202),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1059),
.A2(n_306),
.B(n_220),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_910),
.A2(n_542),
.B(n_286),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_934),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_946),
.B(n_8),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_949),
.B(n_9),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_1012),
.Y(n_1143)
);

OR2x6_ASAP7_75t_L g1144 ( 
.A(n_1012),
.B(n_307),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1073),
.B(n_213),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_939),
.Y(n_1146)
);

AOI221xp5_ASAP7_75t_L g1147 ( 
.A1(n_913),
.A2(n_231),
.B1(n_224),
.B2(n_232),
.C(n_211),
.Y(n_1147)
);

HB1xp67_ASAP7_75t_L g1148 ( 
.A(n_1012),
.Y(n_1148)
);

INVx4_ASAP7_75t_L g1149 ( 
.A(n_942),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_952),
.B(n_233),
.Y(n_1150)
);

NAND2xp33_ASAP7_75t_SL g1151 ( 
.A(n_1036),
.B(n_236),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1066),
.A2(n_317),
.B(n_356),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_965),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_907),
.A2(n_241),
.B1(n_243),
.B2(n_244),
.Y(n_1154)
);

CKINVDCx11_ASAP7_75t_R g1155 ( 
.A(n_971),
.Y(n_1155)
);

BUFx4f_ASAP7_75t_L g1156 ( 
.A(n_1046),
.Y(n_1156)
);

O2A1O1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_950),
.A2(n_9),
.B(n_14),
.C(n_20),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_913),
.A2(n_318),
.B1(n_249),
.B2(n_351),
.Y(n_1158)
);

A2O1A1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_915),
.A2(n_309),
.B(n_250),
.C(n_349),
.Y(n_1159)
);

BUFx12f_ASAP7_75t_L g1160 ( 
.A(n_971),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_967),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_968),
.B(n_20),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_971),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1006),
.B(n_22),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_902),
.A2(n_330),
.B(n_260),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_919),
.A2(n_916),
.B(n_1008),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_907),
.A2(n_333),
.B1(n_253),
.B2(n_347),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_980),
.B(n_23),
.Y(n_1168)
);

INVx8_ASAP7_75t_L g1169 ( 
.A(n_1015),
.Y(n_1169)
);

HB1xp67_ASAP7_75t_L g1170 ( 
.A(n_1048),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_R g1171 ( 
.A(n_1011),
.B(n_275),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_995),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_1013),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1017),
.B(n_25),
.Y(n_1174)
);

INVx2_ASAP7_75t_SL g1175 ( 
.A(n_1021),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1044),
.A2(n_26),
.B(n_28),
.C(n_29),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_R g1177 ( 
.A(n_990),
.B(n_305),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_971),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1025),
.B(n_917),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_938),
.B(n_1048),
.Y(n_1180)
);

AOI21x1_ASAP7_75t_L g1181 ( 
.A1(n_975),
.A2(n_487),
.B(n_213),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_973),
.Y(n_1182)
);

INVx2_ASAP7_75t_SL g1183 ( 
.A(n_973),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1030),
.A2(n_308),
.B1(n_334),
.B2(n_337),
.Y(n_1184)
);

A2O1A1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1051),
.A2(n_346),
.B(n_307),
.C(n_487),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_898),
.B(n_30),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_957),
.B(n_33),
.Y(n_1187)
);

INVx3_ASAP7_75t_L g1188 ( 
.A(n_1013),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1054),
.A2(n_307),
.B1(n_213),
.B2(n_354),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1024),
.B(n_33),
.Y(n_1190)
);

O2A1O1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1044),
.A2(n_34),
.B(n_35),
.C(n_38),
.Y(n_1191)
);

O2A1O1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_929),
.A2(n_34),
.B(n_39),
.C(n_40),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_988),
.A2(n_487),
.B(n_307),
.Y(n_1193)
);

INVx4_ASAP7_75t_L g1194 ( 
.A(n_973),
.Y(n_1194)
);

XOR2x2_ASAP7_75t_L g1195 ( 
.A(n_1024),
.B(n_41),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_893),
.A2(n_487),
.B(n_103),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_1036),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_1054),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_893),
.A2(n_487),
.B(n_95),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_899),
.B(n_42),
.Y(n_1200)
);

INVx4_ASAP7_75t_L g1201 ( 
.A(n_973),
.Y(n_1201)
);

OR2x6_ASAP7_75t_L g1202 ( 
.A(n_963),
.B(n_1069),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_994),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_914),
.A2(n_487),
.B(n_107),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_935),
.A2(n_43),
.B1(n_49),
.B2(n_50),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_940),
.A2(n_213),
.B1(n_53),
.B2(n_54),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1063),
.B(n_213),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1045),
.A2(n_213),
.B(n_119),
.Y(n_1208)
);

AOI21x1_ASAP7_75t_L g1209 ( 
.A1(n_891),
.A2(n_213),
.B(n_122),
.Y(n_1209)
);

NOR3x1_ASAP7_75t_L g1210 ( 
.A(n_1071),
.B(n_50),
.C(n_55),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_895),
.B(n_213),
.Y(n_1211)
);

AOI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1053),
.A2(n_213),
.B1(n_56),
.B2(n_59),
.Y(n_1212)
);

INVx1_ASAP7_75t_SL g1213 ( 
.A(n_994),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1075),
.B(n_55),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_957),
.B(n_61),
.Y(n_1215)
);

BUFx8_ASAP7_75t_L g1216 ( 
.A(n_994),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_933),
.B(n_62),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_936),
.A2(n_129),
.B(n_187),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1072),
.B(n_62),
.Y(n_1219)
);

INVxp67_ASAP7_75t_SL g1220 ( 
.A(n_994),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_972),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_1007),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_944),
.B(n_63),
.Y(n_1223)
);

O2A1O1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_889),
.A2(n_63),
.B(n_66),
.C(n_71),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_905),
.A2(n_981),
.B1(n_1067),
.B2(n_924),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_914),
.A2(n_141),
.B(n_186),
.Y(n_1226)
);

INVxp67_ASAP7_75t_L g1227 ( 
.A(n_1058),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1042),
.Y(n_1228)
);

O2A1O1Ixp33_ASAP7_75t_SL g1229 ( 
.A1(n_937),
.A2(n_960),
.B(n_943),
.C(n_993),
.Y(n_1229)
);

O2A1O1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_903),
.A2(n_66),
.B(n_72),
.C(n_73),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1000),
.A2(n_72),
.B1(n_74),
.B2(n_77),
.Y(n_1231)
);

INVx2_ASAP7_75t_SL g1232 ( 
.A(n_1007),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_964),
.A2(n_79),
.B(n_86),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1043),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_947),
.B(n_94),
.Y(n_1235)
);

AND2x4_ASAP7_75t_L g1236 ( 
.A(n_1075),
.B(n_963),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_990),
.B(n_109),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1041),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1052),
.B(n_194),
.Y(n_1239)
);

CKINVDCx6p67_ASAP7_75t_R g1240 ( 
.A(n_1094),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1119),
.A2(n_1229),
.B(n_1166),
.Y(n_1241)
);

CKINVDCx11_ASAP7_75t_R g1242 ( 
.A(n_1094),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1208),
.A2(n_970),
.B(n_961),
.Y(n_1243)
);

AO21x1_ASAP7_75t_L g1244 ( 
.A1(n_1078),
.A2(n_991),
.B(n_1035),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1079),
.B(n_1052),
.Y(n_1245)
);

A2O1A1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1219),
.A2(n_1126),
.B(n_1087),
.C(n_1190),
.Y(n_1246)
);

O2A1O1Ixp33_ASAP7_75t_SL g1247 ( 
.A1(n_1179),
.A2(n_937),
.B(n_931),
.C(n_1029),
.Y(n_1247)
);

INVx1_ASAP7_75t_SL g1248 ( 
.A(n_1155),
.Y(n_1248)
);

CKINVDCx20_ASAP7_75t_R g1249 ( 
.A(n_1129),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1123),
.Y(n_1250)
);

INVx1_ASAP7_75t_SL g1251 ( 
.A(n_1091),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1086),
.A2(n_1002),
.B(n_1001),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1081),
.A2(n_956),
.B1(n_958),
.B2(n_1026),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1180),
.B(n_1170),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1228),
.B(n_996),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1195),
.B(n_1065),
.Y(n_1256)
);

A2O1A1Ixp33_ASAP7_75t_L g1257 ( 
.A1(n_1212),
.A2(n_1016),
.B(n_1050),
.C(n_1031),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1082),
.A2(n_959),
.B(n_953),
.Y(n_1258)
);

NAND3xp33_ASAP7_75t_SL g1259 ( 
.A(n_1158),
.B(n_941),
.C(n_977),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1131),
.Y(n_1260)
);

O2A1O1Ixp33_ASAP7_75t_SL g1261 ( 
.A1(n_1159),
.A2(n_1039),
.B(n_1037),
.C(n_1060),
.Y(n_1261)
);

INVx3_ASAP7_75t_L g1262 ( 
.A(n_1160),
.Y(n_1262)
);

OR2x2_ASAP7_75t_L g1263 ( 
.A(n_1108),
.B(n_996),
.Y(n_1263)
);

OAI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1200),
.A2(n_948),
.B(n_985),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1086),
.A2(n_1088),
.B(n_1085),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1146),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1128),
.A2(n_974),
.B(n_1010),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1088),
.A2(n_926),
.B(n_983),
.Y(n_1268)
);

AOI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1209),
.A2(n_984),
.B(n_1049),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1235),
.A2(n_978),
.B(n_979),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1234),
.B(n_1005),
.Y(n_1271)
);

AO31x2_ASAP7_75t_L g1272 ( 
.A1(n_1193),
.A2(n_1185),
.A3(n_1089),
.B(n_1080),
.Y(n_1272)
);

AOI32xp33_ASAP7_75t_L g1273 ( 
.A1(n_1104),
.A2(n_1019),
.A3(n_1060),
.B1(n_1005),
.B2(n_1056),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1096),
.A2(n_1047),
.B(n_1057),
.Y(n_1274)
);

A2O1A1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1157),
.A2(n_1004),
.B(n_997),
.C(n_987),
.Y(n_1275)
);

OAI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1205),
.A2(n_1007),
.B1(n_989),
.B2(n_992),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1198),
.B(n_1007),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1218),
.A2(n_1115),
.B(n_1105),
.Y(n_1278)
);

AO21x2_ASAP7_75t_L g1279 ( 
.A1(n_1139),
.A2(n_986),
.B(n_901),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1134),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1130),
.B(n_901),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1135),
.Y(n_1282)
);

AO31x2_ASAP7_75t_L g1283 ( 
.A1(n_1089),
.A2(n_1018),
.A3(n_925),
.B(n_923),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1140),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1124),
.A2(n_1022),
.B1(n_1027),
.B2(n_1028),
.Y(n_1285)
);

BUFx10_ASAP7_75t_L g1286 ( 
.A(n_1090),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1080),
.A2(n_1038),
.B(n_1068),
.Y(n_1287)
);

INVx1_ASAP7_75t_SL g1288 ( 
.A(n_1143),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1205),
.A2(n_1034),
.B1(n_1023),
.B2(n_1061),
.Y(n_1289)
);

AOI221x1_ASAP7_75t_L g1290 ( 
.A1(n_1231),
.A2(n_1064),
.B1(n_1076),
.B2(n_146),
.C(n_162),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1196),
.A2(n_125),
.B(n_140),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_1083),
.B(n_165),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1092),
.A2(n_168),
.B(n_170),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1101),
.A2(n_182),
.B(n_184),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1199),
.A2(n_185),
.B(n_1111),
.Y(n_1295)
);

BUFx10_ASAP7_75t_L g1296 ( 
.A(n_1120),
.Y(n_1296)
);

INVx4_ASAP7_75t_L g1297 ( 
.A(n_1094),
.Y(n_1297)
);

AO21x2_ASAP7_75t_L g1298 ( 
.A1(n_1139),
.A2(n_1116),
.B(n_1225),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1106),
.A2(n_1107),
.B(n_1223),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1153),
.Y(n_1300)
);

O2A1O1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1109),
.A2(n_1230),
.B(n_1224),
.C(n_1231),
.Y(n_1301)
);

O2A1O1Ixp33_ASAP7_75t_SL g1302 ( 
.A1(n_1117),
.A2(n_1223),
.B(n_1215),
.C(n_1099),
.Y(n_1302)
);

BUFx2_ASAP7_75t_L g1303 ( 
.A(n_1129),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1114),
.A2(n_1122),
.B(n_1204),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1233),
.A2(n_1102),
.B(n_1226),
.Y(n_1305)
);

OAI22x1_ASAP7_75t_L g1306 ( 
.A1(n_1095),
.A2(n_1175),
.B1(n_1150),
.B2(n_1148),
.Y(n_1306)
);

OA21x2_ASAP7_75t_L g1307 ( 
.A1(n_1211),
.A2(n_1116),
.B(n_1145),
.Y(n_1307)
);

AO21x2_ASAP7_75t_L g1308 ( 
.A1(n_1145),
.A2(n_1207),
.B(n_1186),
.Y(n_1308)
);

AO31x2_ASAP7_75t_L g1309 ( 
.A1(n_1207),
.A2(n_1112),
.A3(n_1238),
.B(n_1221),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1161),
.B(n_1172),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1141),
.A2(n_1174),
.B1(n_1162),
.B2(n_1142),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1121),
.A2(n_1173),
.B(n_1188),
.Y(n_1312)
);

OAI22x1_ASAP7_75t_L g1313 ( 
.A1(n_1137),
.A2(n_1239),
.B1(n_1214),
.B2(n_1164),
.Y(n_1313)
);

BUFx12f_ASAP7_75t_L g1314 ( 
.A(n_1197),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1173),
.A2(n_1188),
.B(n_1084),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1202),
.A2(n_1220),
.B(n_1213),
.Y(n_1316)
);

INVx1_ASAP7_75t_SL g1317 ( 
.A(n_1093),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1192),
.A2(n_1168),
.B(n_1136),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1202),
.A2(n_1213),
.B(n_1077),
.Y(n_1319)
);

OA21x2_ASAP7_75t_L g1320 ( 
.A1(n_1100),
.A2(n_1165),
.B(n_1189),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1176),
.A2(n_1191),
.B(n_1110),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_1156),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1127),
.A2(n_1152),
.B(n_1133),
.Y(n_1323)
);

A2O1A1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1113),
.A2(n_1217),
.B(n_1187),
.C(n_1167),
.Y(n_1324)
);

A2O1A1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1147),
.A2(n_1098),
.B(n_1206),
.C(n_1184),
.Y(n_1325)
);

OAI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1202),
.A2(n_1138),
.B(n_1184),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1077),
.A2(n_1154),
.B(n_1194),
.Y(n_1327)
);

AO21x1_ASAP7_75t_L g1328 ( 
.A1(n_1154),
.A2(n_1237),
.B(n_1214),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1156),
.B(n_1227),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1077),
.A2(n_1169),
.B(n_1232),
.Y(n_1330)
);

A2O1A1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1104),
.A2(n_1237),
.B(n_1236),
.C(n_1151),
.Y(n_1331)
);

CKINVDCx20_ASAP7_75t_R g1332 ( 
.A(n_1216),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1077),
.A2(n_1201),
.B(n_1194),
.Y(n_1333)
);

INVxp67_ASAP7_75t_L g1334 ( 
.A(n_1132),
.Y(n_1334)
);

NAND3xp33_ASAP7_75t_L g1335 ( 
.A(n_1097),
.B(n_1118),
.C(n_1182),
.Y(n_1335)
);

BUFx8_ASAP7_75t_L g1336 ( 
.A(n_1097),
.Y(n_1336)
);

AO31x2_ASAP7_75t_L g1337 ( 
.A1(n_1149),
.A2(n_1201),
.A3(n_1210),
.B(n_1144),
.Y(n_1337)
);

INVxp67_ASAP7_75t_L g1338 ( 
.A(n_1144),
.Y(n_1338)
);

BUFx2_ASAP7_75t_L g1339 ( 
.A(n_1177),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1149),
.A2(n_1097),
.B(n_1118),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_1125),
.B(n_1144),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1169),
.B(n_1171),
.Y(n_1342)
);

AO31x2_ASAP7_75t_L g1343 ( 
.A1(n_1125),
.A2(n_1118),
.A3(n_1163),
.B(n_1222),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1169),
.A2(n_1183),
.B(n_1178),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1203),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1163),
.A2(n_1178),
.B(n_1182),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1163),
.A2(n_1178),
.B(n_1182),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1222),
.A2(n_1119),
.B(n_1229),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_SL g1349 ( 
.A1(n_1222),
.A2(n_596),
.B(n_591),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1119),
.A2(n_1229),
.B(n_890),
.Y(n_1350)
);

A2O1A1Ixp33_ASAP7_75t_L g1351 ( 
.A1(n_1219),
.A2(n_1014),
.B(n_890),
.C(n_1078),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1180),
.B(n_890),
.Y(n_1352)
);

INVxp67_ASAP7_75t_L g1353 ( 
.A(n_1108),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1179),
.A2(n_1033),
.B1(n_890),
.B2(n_1014),
.Y(n_1354)
);

NOR2xp67_ASAP7_75t_SL g1355 ( 
.A(n_1160),
.B(n_829),
.Y(n_1355)
);

OA21x2_ASAP7_75t_L g1356 ( 
.A1(n_1105),
.A2(n_1166),
.B(n_945),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1119),
.A2(n_910),
.B(n_890),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_1129),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1123),
.Y(n_1359)
);

AND2x4_ASAP7_75t_L g1360 ( 
.A(n_1110),
.B(n_1143),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1208),
.A2(n_1181),
.B(n_918),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1079),
.B(n_738),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1119),
.A2(n_1229),
.B(n_890),
.Y(n_1363)
);

INVx3_ASAP7_75t_L g1364 ( 
.A(n_1160),
.Y(n_1364)
);

BUFx8_ASAP7_75t_L g1365 ( 
.A(n_1160),
.Y(n_1365)
);

AO21x1_ASAP7_75t_L g1366 ( 
.A1(n_1078),
.A2(n_1014),
.B(n_1219),
.Y(n_1366)
);

BUFx10_ASAP7_75t_L g1367 ( 
.A(n_1090),
.Y(n_1367)
);

AOI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1078),
.A2(n_518),
.B1(n_1014),
.B2(n_1055),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1123),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_L g1370 ( 
.A(n_1083),
.B(n_518),
.Y(n_1370)
);

AO31x2_ASAP7_75t_L g1371 ( 
.A1(n_1166),
.A2(n_945),
.A3(n_977),
.B(n_910),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1180),
.B(n_890),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1119),
.A2(n_1229),
.B(n_890),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1103),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1079),
.B(n_771),
.Y(n_1375)
);

AND2x4_ASAP7_75t_L g1376 ( 
.A(n_1110),
.B(n_1143),
.Y(n_1376)
);

OAI22x1_ASAP7_75t_L g1377 ( 
.A1(n_1079),
.A2(n_596),
.B1(n_653),
.B2(n_503),
.Y(n_1377)
);

INVxp67_ASAP7_75t_L g1378 ( 
.A(n_1108),
.Y(n_1378)
);

INVxp67_ASAP7_75t_SL g1379 ( 
.A(n_1086),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1179),
.A2(n_1033),
.B1(n_890),
.B2(n_1014),
.Y(n_1380)
);

AOI221xp5_ASAP7_75t_L g1381 ( 
.A1(n_1078),
.A2(n_734),
.B1(n_400),
.B2(n_1079),
.C(n_752),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1119),
.A2(n_1229),
.B(n_890),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1119),
.A2(n_1229),
.B(n_890),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1123),
.Y(n_1384)
);

INVx1_ASAP7_75t_SL g1385 ( 
.A(n_1155),
.Y(n_1385)
);

CKINVDCx6p67_ASAP7_75t_R g1386 ( 
.A(n_1094),
.Y(n_1386)
);

AO31x2_ASAP7_75t_L g1387 ( 
.A1(n_1166),
.A2(n_945),
.A3(n_977),
.B(n_910),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1119),
.A2(n_1229),
.B(n_890),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1119),
.A2(n_910),
.B(n_890),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_SL g1390 ( 
.A(n_1083),
.B(n_1014),
.Y(n_1390)
);

NOR2xp33_ASAP7_75t_L g1391 ( 
.A(n_1083),
.B(n_518),
.Y(n_1391)
);

OA21x2_ASAP7_75t_L g1392 ( 
.A1(n_1105),
.A2(n_1166),
.B(n_945),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1108),
.Y(n_1393)
);

OAI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1119),
.A2(n_910),
.B(n_890),
.Y(n_1394)
);

INVx5_ASAP7_75t_L g1395 ( 
.A(n_1094),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1119),
.A2(n_1229),
.B(n_890),
.Y(n_1396)
);

AOI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1078),
.A2(n_518),
.B1(n_1014),
.B2(n_1055),
.Y(n_1397)
);

OAI221xp5_ASAP7_75t_L g1398 ( 
.A1(n_1078),
.A2(n_1014),
.B1(n_890),
.B2(n_596),
.C(n_825),
.Y(n_1398)
);

AOI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1078),
.A2(n_518),
.B1(n_1014),
.B2(n_1055),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1103),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1119),
.A2(n_1229),
.B(n_890),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_1155),
.Y(n_1402)
);

O2A1O1Ixp33_ASAP7_75t_SL g1403 ( 
.A1(n_1119),
.A2(n_1014),
.B(n_1179),
.C(n_890),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1110),
.B(n_1143),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1377),
.A2(n_1256),
.B1(n_1381),
.B2(n_1245),
.Y(n_1405)
);

INVx6_ASAP7_75t_L g1406 ( 
.A(n_1336),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1313),
.A2(n_1366),
.B1(n_1354),
.B2(n_1380),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1368),
.A2(n_1397),
.B1(n_1399),
.B2(n_1370),
.Y(n_1408)
);

CKINVDCx11_ASAP7_75t_R g1409 ( 
.A(n_1249),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1354),
.A2(n_1380),
.B1(n_1398),
.B2(n_1311),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_1242),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1250),
.Y(n_1412)
);

CKINVDCx11_ASAP7_75t_R g1413 ( 
.A(n_1332),
.Y(n_1413)
);

OAI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1362),
.A2(n_1349),
.B1(n_1254),
.B2(n_1372),
.Y(n_1414)
);

BUFx10_ASAP7_75t_L g1415 ( 
.A(n_1402),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1260),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1311),
.A2(n_1375),
.B1(n_1244),
.B2(n_1328),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_1395),
.Y(n_1418)
);

CKINVDCx6p67_ASAP7_75t_R g1419 ( 
.A(n_1395),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1298),
.A2(n_1390),
.B1(n_1281),
.B2(n_1391),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_1314),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1298),
.A2(n_1334),
.B1(n_1357),
.B2(n_1389),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1280),
.Y(n_1423)
);

INVx6_ASAP7_75t_L g1424 ( 
.A(n_1336),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_SL g1425 ( 
.A1(n_1326),
.A2(n_1357),
.B1(n_1389),
.B2(n_1394),
.Y(n_1425)
);

INVx1_ASAP7_75t_SL g1426 ( 
.A(n_1339),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1282),
.Y(n_1427)
);

NAND2xp33_ASAP7_75t_SL g1428 ( 
.A(n_1402),
.B(n_1297),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1394),
.A2(n_1259),
.B1(n_1306),
.B2(n_1254),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1284),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1253),
.A2(n_1373),
.B1(n_1382),
.B2(n_1401),
.Y(n_1431)
);

INVx1_ASAP7_75t_SL g1432 ( 
.A(n_1322),
.Y(n_1432)
);

BUFx4f_ASAP7_75t_SL g1433 ( 
.A(n_1365),
.Y(n_1433)
);

INVx2_ASAP7_75t_SL g1434 ( 
.A(n_1365),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_SL g1435 ( 
.A1(n_1326),
.A2(n_1296),
.B1(n_1253),
.B2(n_1388),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_SL g1436 ( 
.A1(n_1351),
.A2(n_1331),
.B(n_1246),
.Y(n_1436)
);

INVx1_ASAP7_75t_SL g1437 ( 
.A(n_1296),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1300),
.Y(n_1438)
);

BUFx10_ASAP7_75t_L g1439 ( 
.A(n_1402),
.Y(n_1439)
);

BUFx4f_ASAP7_75t_SL g1440 ( 
.A(n_1240),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1350),
.A2(n_1383),
.B1(n_1363),
.B2(n_1396),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1359),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1386),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1352),
.A2(n_1372),
.B1(n_1308),
.B2(n_1369),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1303),
.Y(n_1445)
);

CKINVDCx8_ASAP7_75t_R g1446 ( 
.A(n_1358),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1251),
.B(n_1393),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1353),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1384),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_SL g1450 ( 
.A1(n_1352),
.A2(n_1320),
.B1(n_1286),
.B2(n_1367),
.Y(n_1450)
);

CKINVDCx20_ASAP7_75t_R g1451 ( 
.A(n_1248),
.Y(n_1451)
);

OAI22x1_ASAP7_75t_L g1452 ( 
.A1(n_1288),
.A2(n_1251),
.B1(n_1338),
.B2(n_1341),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1308),
.A2(n_1317),
.B1(n_1400),
.B2(n_1266),
.Y(n_1453)
);

CKINVDCx6p67_ASAP7_75t_R g1454 ( 
.A(n_1248),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1349),
.A2(n_1325),
.B1(n_1324),
.B2(n_1301),
.Y(n_1455)
);

CKINVDCx11_ASAP7_75t_R g1456 ( 
.A(n_1385),
.Y(n_1456)
);

INVx6_ASAP7_75t_L g1457 ( 
.A(n_1297),
.Y(n_1457)
);

CKINVDCx20_ASAP7_75t_R g1458 ( 
.A(n_1385),
.Y(n_1458)
);

BUFx6f_ASAP7_75t_SL g1459 ( 
.A(n_1286),
.Y(n_1459)
);

BUFx3_ASAP7_75t_L g1460 ( 
.A(n_1262),
.Y(n_1460)
);

CKINVDCx11_ASAP7_75t_R g1461 ( 
.A(n_1367),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1317),
.A2(n_1374),
.B1(n_1379),
.B2(n_1292),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1307),
.A2(n_1279),
.B1(n_1320),
.B2(n_1271),
.Y(n_1463)
);

CKINVDCx11_ASAP7_75t_R g1464 ( 
.A(n_1288),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1255),
.Y(n_1465)
);

BUFx4f_ASAP7_75t_L g1466 ( 
.A(n_1341),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1360),
.B(n_1376),
.Y(n_1467)
);

BUFx12f_ASAP7_75t_L g1468 ( 
.A(n_1263),
.Y(n_1468)
);

INVx4_ASAP7_75t_L g1469 ( 
.A(n_1262),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1255),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1378),
.B(n_1277),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1307),
.A2(n_1279),
.B1(n_1271),
.B2(n_1321),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1345),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1404),
.B(n_1403),
.Y(n_1474)
);

OAI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1257),
.A2(n_1241),
.B1(n_1348),
.B2(n_1285),
.Y(n_1475)
);

BUFx3_ASAP7_75t_L g1476 ( 
.A(n_1364),
.Y(n_1476)
);

CKINVDCx20_ASAP7_75t_R g1477 ( 
.A(n_1342),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1404),
.B(n_1329),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1264),
.A2(n_1318),
.B1(n_1289),
.B2(n_1293),
.Y(n_1479)
);

OAI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1290),
.A2(n_1364),
.B1(n_1289),
.B2(n_1264),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1316),
.A2(n_1319),
.B1(n_1276),
.B2(n_1265),
.Y(n_1481)
);

INVx3_ASAP7_75t_L g1482 ( 
.A(n_1343),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1275),
.A2(n_1273),
.B1(n_1276),
.B2(n_1335),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1268),
.A2(n_1355),
.B1(n_1335),
.B2(n_1315),
.Y(n_1484)
);

AOI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1247),
.A2(n_1302),
.B1(n_1330),
.B2(n_1344),
.Y(n_1485)
);

BUFx4f_ASAP7_75t_L g1486 ( 
.A(n_1356),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1305),
.A2(n_1299),
.B1(n_1287),
.B2(n_1392),
.Y(n_1487)
);

BUFx12f_ASAP7_75t_L g1488 ( 
.A(n_1343),
.Y(n_1488)
);

AOI22xp5_ASAP7_75t_SL g1489 ( 
.A1(n_1337),
.A2(n_1346),
.B1(n_1347),
.B2(n_1294),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1309),
.Y(n_1490)
);

BUFx12f_ASAP7_75t_L g1491 ( 
.A(n_1337),
.Y(n_1491)
);

INVx6_ASAP7_75t_L g1492 ( 
.A(n_1333),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1337),
.B(n_1340),
.Y(n_1493)
);

INVx6_ASAP7_75t_L g1494 ( 
.A(n_1327),
.Y(n_1494)
);

INVx4_ASAP7_75t_L g1495 ( 
.A(n_1356),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1312),
.Y(n_1496)
);

AOI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1261),
.A2(n_1392),
.B1(n_1291),
.B2(n_1252),
.Y(n_1497)
);

CKINVDCx11_ASAP7_75t_R g1498 ( 
.A(n_1272),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1274),
.A2(n_1323),
.B1(n_1270),
.B2(n_1295),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1269),
.A2(n_1387),
.B1(n_1371),
.B2(n_1272),
.Y(n_1500)
);

INVx3_ASAP7_75t_L g1501 ( 
.A(n_1283),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1387),
.A2(n_1272),
.B1(n_1283),
.B2(n_1278),
.Y(n_1502)
);

INVx1_ASAP7_75t_SL g1503 ( 
.A(n_1267),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1283),
.Y(n_1504)
);

NAND2xp33_ASAP7_75t_SL g1505 ( 
.A(n_1387),
.B(n_1304),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1258),
.B(n_1243),
.Y(n_1506)
);

CKINVDCx20_ASAP7_75t_R g1507 ( 
.A(n_1361),
.Y(n_1507)
);

BUFx10_ASAP7_75t_L g1508 ( 
.A(n_1402),
.Y(n_1508)
);

INVx2_ASAP7_75t_SL g1509 ( 
.A(n_1395),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1375),
.B(n_1256),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1375),
.B(n_1256),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1377),
.A2(n_1256),
.B1(n_1078),
.B2(n_1381),
.Y(n_1512)
);

INVx6_ASAP7_75t_L g1513 ( 
.A(n_1336),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1310),
.Y(n_1514)
);

BUFx2_ASAP7_75t_SL g1515 ( 
.A(n_1332),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_SL g1516 ( 
.A1(n_1256),
.A2(n_767),
.B1(n_1055),
.B2(n_403),
.Y(n_1516)
);

OAI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1368),
.A2(n_1397),
.B1(n_1399),
.B2(n_1245),
.Y(n_1517)
);

BUFx12f_ASAP7_75t_L g1518 ( 
.A(n_1242),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1368),
.A2(n_1397),
.B1(n_1399),
.B2(n_1014),
.Y(n_1519)
);

CKINVDCx11_ASAP7_75t_R g1520 ( 
.A(n_1249),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1310),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1310),
.Y(n_1522)
);

CKINVDCx11_ASAP7_75t_R g1523 ( 
.A(n_1249),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_SL g1524 ( 
.A1(n_1256),
.A2(n_767),
.B1(n_1055),
.B2(n_403),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1377),
.A2(n_1256),
.B1(n_1078),
.B2(n_1381),
.Y(n_1525)
);

BUFx3_ASAP7_75t_L g1526 ( 
.A(n_1336),
.Y(n_1526)
);

CKINVDCx11_ASAP7_75t_R g1527 ( 
.A(n_1249),
.Y(n_1527)
);

BUFx12f_ASAP7_75t_L g1528 ( 
.A(n_1242),
.Y(n_1528)
);

OAI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1368),
.A2(n_1397),
.B1(n_1399),
.B2(n_1245),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_SL g1530 ( 
.A1(n_1256),
.A2(n_767),
.B1(n_1055),
.B2(n_403),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1368),
.A2(n_1397),
.B1(n_1399),
.B2(n_1014),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1377),
.A2(n_1256),
.B1(n_1078),
.B2(n_1381),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1368),
.A2(n_1397),
.B1(n_1399),
.B2(n_1014),
.Y(n_1533)
);

INVx4_ASAP7_75t_L g1534 ( 
.A(n_1242),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1310),
.Y(n_1535)
);

OAI22xp33_ASAP7_75t_R g1536 ( 
.A1(n_1370),
.A2(n_1391),
.B1(n_851),
.B2(n_200),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1377),
.A2(n_1256),
.B1(n_1078),
.B2(n_1381),
.Y(n_1537)
);

INVx3_ASAP7_75t_L g1538 ( 
.A(n_1336),
.Y(n_1538)
);

BUFx8_ASAP7_75t_SL g1539 ( 
.A(n_1332),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1368),
.A2(n_1397),
.B1(n_1399),
.B2(n_1014),
.Y(n_1540)
);

CKINVDCx14_ASAP7_75t_R g1541 ( 
.A(n_1242),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1375),
.B(n_1256),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_SL g1543 ( 
.A1(n_1256),
.A2(n_767),
.B1(n_1055),
.B2(n_403),
.Y(n_1543)
);

CKINVDCx6p67_ASAP7_75t_R g1544 ( 
.A(n_1395),
.Y(n_1544)
);

CKINVDCx11_ASAP7_75t_R g1545 ( 
.A(n_1249),
.Y(n_1545)
);

BUFx2_ASAP7_75t_SL g1546 ( 
.A(n_1332),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1377),
.A2(n_1256),
.B1(n_1078),
.B2(n_1381),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1310),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1465),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1504),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1420),
.B(n_1422),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1470),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1493),
.B(n_1482),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1447),
.Y(n_1554)
);

INVx3_ASAP7_75t_L g1555 ( 
.A(n_1495),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1420),
.B(n_1422),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1425),
.B(n_1412),
.Y(n_1557)
);

CKINVDCx14_ASAP7_75t_R g1558 ( 
.A(n_1541),
.Y(n_1558)
);

CKINVDCx20_ASAP7_75t_R g1559 ( 
.A(n_1539),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1487),
.A2(n_1499),
.B(n_1479),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1416),
.B(n_1423),
.Y(n_1561)
);

CKINVDCx6p67_ASAP7_75t_R g1562 ( 
.A(n_1518),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1444),
.B(n_1514),
.Y(n_1563)
);

BUFx3_ASAP7_75t_L g1564 ( 
.A(n_1491),
.Y(n_1564)
);

INVx2_ASAP7_75t_SL g1565 ( 
.A(n_1492),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1471),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1427),
.Y(n_1567)
);

AOI21xp33_ASAP7_75t_SL g1568 ( 
.A1(n_1455),
.A2(n_1408),
.B(n_1519),
.Y(n_1568)
);

BUFx2_ASAP7_75t_L g1569 ( 
.A(n_1486),
.Y(n_1569)
);

INVx3_ASAP7_75t_L g1570 ( 
.A(n_1495),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1430),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1448),
.Y(n_1572)
);

INVx2_ASAP7_75t_SL g1573 ( 
.A(n_1492),
.Y(n_1573)
);

AO21x2_ASAP7_75t_L g1574 ( 
.A1(n_1490),
.A2(n_1500),
.B(n_1497),
.Y(n_1574)
);

AOI21x1_ASAP7_75t_L g1575 ( 
.A1(n_1502),
.A2(n_1506),
.B(n_1475),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1521),
.B(n_1522),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1438),
.Y(n_1577)
);

AND2x4_ASAP7_75t_SL g1578 ( 
.A(n_1419),
.B(n_1544),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1501),
.Y(n_1579)
);

OAI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1531),
.A2(n_1533),
.B1(n_1540),
.B2(n_1536),
.Y(n_1580)
);

BUFx12f_ASAP7_75t_L g1581 ( 
.A(n_1413),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1442),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1449),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1548),
.B(n_1535),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1486),
.B(n_1410),
.Y(n_1585)
);

OR2x6_ASAP7_75t_L g1586 ( 
.A(n_1488),
.B(n_1436),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1473),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1496),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1512),
.A2(n_1537),
.B1(n_1532),
.B2(n_1525),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1414),
.B(n_1510),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1410),
.B(n_1444),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1452),
.Y(n_1592)
);

INVx3_ASAP7_75t_L g1593 ( 
.A(n_1492),
.Y(n_1593)
);

INVx3_ASAP7_75t_L g1594 ( 
.A(n_1494),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1483),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1512),
.A2(n_1537),
.B1(n_1532),
.B2(n_1525),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1472),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1472),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1463),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1463),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1503),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1498),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1481),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1547),
.A2(n_1405),
.B1(n_1516),
.B2(n_1524),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1481),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1511),
.B(n_1542),
.Y(n_1606)
);

NOR2x1_ASAP7_75t_SL g1607 ( 
.A(n_1474),
.B(n_1418),
.Y(n_1607)
);

AND2x4_ASAP7_75t_L g1608 ( 
.A(n_1507),
.B(n_1467),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1453),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1453),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1414),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1505),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1407),
.B(n_1429),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1429),
.B(n_1435),
.Y(n_1614)
);

NAND2x1p5_ASAP7_75t_L g1615 ( 
.A(n_1466),
.B(n_1489),
.Y(n_1615)
);

OAI31xp33_ASAP7_75t_L g1616 ( 
.A1(n_1517),
.A2(n_1529),
.A3(n_1547),
.B(n_1405),
.Y(n_1616)
);

AO21x2_ASAP7_75t_L g1617 ( 
.A1(n_1480),
.A2(n_1485),
.B(n_1529),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1480),
.Y(n_1618)
);

INVx1_ASAP7_75t_SL g1619 ( 
.A(n_1464),
.Y(n_1619)
);

AO21x2_ASAP7_75t_L g1620 ( 
.A1(n_1517),
.A2(n_1478),
.B(n_1407),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1431),
.Y(n_1621)
);

NAND2x1_ASAP7_75t_L g1622 ( 
.A(n_1484),
.B(n_1431),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1468),
.Y(n_1623)
);

INVx2_ASAP7_75t_SL g1624 ( 
.A(n_1406),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1467),
.B(n_1417),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1530),
.A2(n_1543),
.B1(n_1417),
.B2(n_1462),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1437),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_1409),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1450),
.Y(n_1629)
);

OR2x6_ASAP7_75t_L g1630 ( 
.A(n_1406),
.B(n_1513),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1441),
.B(n_1479),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1441),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1484),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1499),
.Y(n_1634)
);

OAI21x1_ASAP7_75t_L g1635 ( 
.A1(n_1462),
.A2(n_1538),
.B(n_1509),
.Y(n_1635)
);

INVx4_ASAP7_75t_L g1636 ( 
.A(n_1466),
.Y(n_1636)
);

OAI21x1_ASAP7_75t_L g1637 ( 
.A1(n_1538),
.A2(n_1457),
.B(n_1459),
.Y(n_1637)
);

AOI21x1_ASAP7_75t_L g1638 ( 
.A1(n_1459),
.A2(n_1434),
.B(n_1457),
.Y(n_1638)
);

OAI21x1_ASAP7_75t_L g1639 ( 
.A1(n_1428),
.A2(n_1469),
.B(n_1460),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1426),
.B(n_1476),
.Y(n_1640)
);

AO21x2_ASAP7_75t_L g1641 ( 
.A1(n_1469),
.A2(n_1461),
.B(n_1477),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1446),
.Y(n_1642)
);

OA21x2_ASAP7_75t_L g1643 ( 
.A1(n_1445),
.A2(n_1432),
.B(n_1443),
.Y(n_1643)
);

INVx1_ASAP7_75t_SL g1644 ( 
.A(n_1546),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1424),
.Y(n_1645)
);

INVx3_ASAP7_75t_L g1646 ( 
.A(n_1513),
.Y(n_1646)
);

INVx3_ASAP7_75t_L g1647 ( 
.A(n_1513),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1526),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_L g1649 ( 
.A(n_1568),
.B(n_1454),
.Y(n_1649)
);

NOR2x1_ASAP7_75t_SL g1650 ( 
.A(n_1586),
.B(n_1528),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1566),
.B(n_1526),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1553),
.B(n_1534),
.Y(n_1652)
);

INVxp67_ASAP7_75t_L g1653 ( 
.A(n_1627),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1557),
.B(n_1534),
.Y(n_1654)
);

INVxp67_ASAP7_75t_L g1655 ( 
.A(n_1640),
.Y(n_1655)
);

A2O1A1Ixp33_ASAP7_75t_L g1656 ( 
.A1(n_1616),
.A2(n_1541),
.B(n_1515),
.C(n_1458),
.Y(n_1656)
);

OAI21xp33_ASAP7_75t_L g1657 ( 
.A1(n_1568),
.A2(n_1451),
.B(n_1411),
.Y(n_1657)
);

INVx5_ASAP7_75t_SL g1658 ( 
.A(n_1562),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1554),
.B(n_1421),
.Y(n_1659)
);

OAI211xp5_ASAP7_75t_L g1660 ( 
.A1(n_1616),
.A2(n_1456),
.B(n_1527),
.C(n_1545),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1587),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1553),
.B(n_1415),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1580),
.B(n_1439),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1608),
.B(n_1508),
.Y(n_1664)
);

AOI221xp5_ASAP7_75t_L g1665 ( 
.A1(n_1589),
.A2(n_1508),
.B1(n_1523),
.B2(n_1520),
.C(n_1433),
.Y(n_1665)
);

AO21x2_ASAP7_75t_L g1666 ( 
.A1(n_1633),
.A2(n_1433),
.B(n_1440),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1557),
.B(n_1440),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1567),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1606),
.B(n_1572),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1585),
.B(n_1561),
.Y(n_1670)
);

NAND3xp33_ASAP7_75t_L g1671 ( 
.A(n_1595),
.B(n_1614),
.C(n_1618),
.Y(n_1671)
);

A2O1A1Ixp33_ASAP7_75t_L g1672 ( 
.A1(n_1596),
.A2(n_1613),
.B(n_1591),
.C(n_1622),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1553),
.B(n_1593),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1571),
.B(n_1577),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1595),
.B(n_1584),
.Y(n_1675)
);

CKINVDCx6p67_ASAP7_75t_R g1676 ( 
.A(n_1581),
.Y(n_1676)
);

A2O1A1Ixp33_ASAP7_75t_L g1677 ( 
.A1(n_1613),
.A2(n_1591),
.B(n_1622),
.C(n_1626),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1571),
.Y(n_1678)
);

NAND3xp33_ASAP7_75t_L g1679 ( 
.A(n_1618),
.B(n_1611),
.C(n_1603),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_1581),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1643),
.B(n_1602),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1577),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1588),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1590),
.B(n_1643),
.Y(n_1684)
);

AND2x4_ASAP7_75t_L g1685 ( 
.A(n_1553),
.B(n_1593),
.Y(n_1685)
);

OA21x2_ASAP7_75t_L g1686 ( 
.A1(n_1560),
.A2(n_1634),
.B(n_1575),
.Y(n_1686)
);

OA21x2_ASAP7_75t_L g1687 ( 
.A1(n_1560),
.A2(n_1634),
.B(n_1575),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_1562),
.Y(n_1688)
);

AOI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1617),
.A2(n_1631),
.B(n_1603),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1569),
.B(n_1641),
.Y(n_1690)
);

OAI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1611),
.A2(n_1631),
.B(n_1605),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1569),
.B(n_1641),
.Y(n_1692)
);

A2O1A1Ixp33_ASAP7_75t_L g1693 ( 
.A1(n_1604),
.A2(n_1629),
.B(n_1556),
.C(n_1551),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_SL g1694 ( 
.A1(n_1558),
.A2(n_1619),
.B1(n_1559),
.B2(n_1628),
.Y(n_1694)
);

OAI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1621),
.A2(n_1632),
.B(n_1633),
.Y(n_1695)
);

AOI211xp5_ASAP7_75t_L g1696 ( 
.A1(n_1629),
.A2(n_1556),
.B(n_1551),
.C(n_1621),
.Y(n_1696)
);

AOI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1597),
.A2(n_1598),
.B1(n_1617),
.B2(n_1592),
.C(n_1620),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1641),
.B(n_1648),
.Y(n_1698)
);

AOI221x1_ASAP7_75t_SL g1699 ( 
.A1(n_1632),
.A2(n_1648),
.B1(n_1583),
.B2(n_1582),
.C(n_1549),
.Y(n_1699)
);

INVxp67_ASAP7_75t_L g1700 ( 
.A(n_1642),
.Y(n_1700)
);

OAI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1635),
.A2(n_1639),
.B(n_1637),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_SL g1702 ( 
.A1(n_1630),
.A2(n_1644),
.B1(n_1624),
.B2(n_1586),
.Y(n_1702)
);

OA21x2_ASAP7_75t_L g1703 ( 
.A1(n_1612),
.A2(n_1597),
.B(n_1598),
.Y(n_1703)
);

NOR2x1_ASAP7_75t_R g1704 ( 
.A(n_1624),
.B(n_1646),
.Y(n_1704)
);

OAI211xp5_ASAP7_75t_L g1705 ( 
.A1(n_1612),
.A2(n_1625),
.B(n_1583),
.C(n_1588),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1549),
.B(n_1574),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1620),
.A2(n_1617),
.B1(n_1586),
.B2(n_1599),
.Y(n_1707)
);

AOI221xp5_ASAP7_75t_L g1708 ( 
.A1(n_1620),
.A2(n_1600),
.B1(n_1599),
.B2(n_1576),
.C(n_1609),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1574),
.B(n_1601),
.Y(n_1709)
);

AOI221xp5_ASAP7_75t_L g1710 ( 
.A1(n_1600),
.A2(n_1610),
.B1(n_1609),
.B2(n_1550),
.C(n_1563),
.Y(n_1710)
);

BUFx2_ASAP7_75t_R g1711 ( 
.A(n_1564),
.Y(n_1711)
);

AOI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1586),
.A2(n_1636),
.B1(n_1645),
.B2(n_1615),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1683),
.Y(n_1713)
);

HB1xp67_ASAP7_75t_L g1714 ( 
.A(n_1655),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1668),
.Y(n_1715)
);

INVxp67_ASAP7_75t_SL g1716 ( 
.A(n_1706),
.Y(n_1716)
);

BUFx3_ASAP7_75t_L g1717 ( 
.A(n_1652),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1684),
.B(n_1574),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1684),
.B(n_1550),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1699),
.B(n_1573),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1689),
.B(n_1573),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1670),
.B(n_1570),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1678),
.Y(n_1723)
);

INVx3_ASAP7_75t_SL g1724 ( 
.A(n_1676),
.Y(n_1724)
);

INVxp67_ASAP7_75t_SL g1725 ( 
.A(n_1709),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1703),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1682),
.Y(n_1727)
);

OAI221xp5_ASAP7_75t_L g1728 ( 
.A1(n_1677),
.A2(n_1615),
.B1(n_1630),
.B2(n_1638),
.C(n_1623),
.Y(n_1728)
);

INVx2_ASAP7_75t_SL g1729 ( 
.A(n_1652),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1674),
.Y(n_1730)
);

HB1xp67_ASAP7_75t_L g1731 ( 
.A(n_1661),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1674),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1703),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1675),
.B(n_1565),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1703),
.Y(n_1735)
);

AOI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1697),
.A2(n_1708),
.B1(n_1671),
.B2(n_1707),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1686),
.B(n_1555),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1705),
.B(n_1552),
.Y(n_1738)
);

INVxp67_ASAP7_75t_L g1739 ( 
.A(n_1681),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1673),
.B(n_1594),
.Y(n_1740)
);

INVxp67_ASAP7_75t_L g1741 ( 
.A(n_1698),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1653),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1686),
.B(n_1555),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1669),
.B(n_1607),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1679),
.Y(n_1745)
);

INVx3_ASAP7_75t_L g1746 ( 
.A(n_1673),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1687),
.B(n_1579),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1687),
.B(n_1673),
.Y(n_1748)
);

BUFx2_ASAP7_75t_L g1749 ( 
.A(n_1737),
.Y(n_1749)
);

OAI221xp5_ASAP7_75t_L g1750 ( 
.A1(n_1736),
.A2(n_1672),
.B1(n_1677),
.B2(n_1656),
.C(n_1693),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1719),
.B(n_1687),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1716),
.B(n_1654),
.Y(n_1752)
);

AOI221xp5_ASAP7_75t_L g1753 ( 
.A1(n_1745),
.A2(n_1672),
.B1(n_1656),
.B2(n_1693),
.C(n_1660),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1726),
.Y(n_1754)
);

OAI21x1_ASAP7_75t_L g1755 ( 
.A1(n_1726),
.A2(n_1701),
.B(n_1707),
.Y(n_1755)
);

OA21x2_ASAP7_75t_L g1756 ( 
.A1(n_1726),
.A2(n_1695),
.B(n_1710),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1733),
.Y(n_1757)
);

INVxp67_ASAP7_75t_L g1758 ( 
.A(n_1720),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1748),
.B(n_1690),
.Y(n_1759)
);

OAI221xp5_ASAP7_75t_L g1760 ( 
.A1(n_1745),
.A2(n_1696),
.B1(n_1691),
.B2(n_1665),
.C(n_1663),
.Y(n_1760)
);

INVx1_ASAP7_75t_SL g1761 ( 
.A(n_1720),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1748),
.B(n_1692),
.Y(n_1762)
);

INVxp33_ASAP7_75t_L g1763 ( 
.A(n_1728),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1719),
.B(n_1713),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1716),
.B(n_1651),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1733),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1715),
.Y(n_1767)
);

AND2x4_ASAP7_75t_L g1768 ( 
.A(n_1748),
.B(n_1685),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1718),
.B(n_1685),
.Y(n_1769)
);

INVxp67_ASAP7_75t_L g1770 ( 
.A(n_1742),
.Y(n_1770)
);

AOI211xp5_ASAP7_75t_SL g1771 ( 
.A1(n_1728),
.A2(n_1649),
.B(n_1663),
.C(n_1694),
.Y(n_1771)
);

BUFx6f_ASAP7_75t_L g1772 ( 
.A(n_1737),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1733),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1744),
.B(n_1657),
.Y(n_1774)
);

OAI221xp5_ASAP7_75t_L g1775 ( 
.A1(n_1718),
.A2(n_1721),
.B1(n_1649),
.B2(n_1738),
.C(n_1725),
.Y(n_1775)
);

INVxp67_ASAP7_75t_SL g1776 ( 
.A(n_1747),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1715),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1723),
.Y(n_1778)
);

INVx4_ASAP7_75t_L g1779 ( 
.A(n_1724),
.Y(n_1779)
);

BUFx3_ASAP7_75t_L g1780 ( 
.A(n_1724),
.Y(n_1780)
);

INVxp67_ASAP7_75t_SL g1781 ( 
.A(n_1747),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1723),
.Y(n_1782)
);

INVx5_ASAP7_75t_SL g1783 ( 
.A(n_1740),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1735),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1727),
.Y(n_1785)
);

AOI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1738),
.A2(n_1667),
.B1(n_1702),
.B2(n_1666),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1735),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1739),
.B(n_1722),
.Y(n_1788)
);

HB1xp67_ASAP7_75t_L g1789 ( 
.A(n_1714),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1767),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1768),
.B(n_1776),
.Y(n_1791)
);

NOR2xp67_ASAP7_75t_L g1792 ( 
.A(n_1779),
.B(n_1741),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1789),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1768),
.B(n_1746),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1768),
.B(n_1746),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1767),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1761),
.B(n_1758),
.Y(n_1797)
);

INVxp67_ASAP7_75t_L g1798 ( 
.A(n_1774),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1754),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1768),
.B(n_1746),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1777),
.Y(n_1801)
);

OAI21xp5_ASAP7_75t_L g1802 ( 
.A1(n_1771),
.A2(n_1741),
.B(n_1721),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1754),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1761),
.B(n_1730),
.Y(n_1804)
);

NOR2xp67_ASAP7_75t_L g1805 ( 
.A(n_1779),
.B(n_1746),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1754),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1758),
.B(n_1731),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1777),
.Y(n_1808)
);

INVx2_ASAP7_75t_SL g1809 ( 
.A(n_1780),
.Y(n_1809)
);

NAND2x1_ASAP7_75t_L g1810 ( 
.A(n_1768),
.B(n_1749),
.Y(n_1810)
);

NOR2x1p5_ASAP7_75t_L g1811 ( 
.A(n_1780),
.B(n_1676),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1778),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1788),
.B(n_1729),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1757),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1764),
.B(n_1730),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1788),
.B(n_1729),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1764),
.B(n_1732),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1788),
.B(n_1729),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1783),
.B(n_1717),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1789),
.B(n_1770),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1778),
.Y(n_1821)
);

AND2x4_ASAP7_75t_L g1822 ( 
.A(n_1776),
.B(n_1781),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1782),
.Y(n_1823)
);

INVxp67_ASAP7_75t_L g1824 ( 
.A(n_1774),
.Y(n_1824)
);

BUFx2_ASAP7_75t_L g1825 ( 
.A(n_1779),
.Y(n_1825)
);

INVx4_ASAP7_75t_L g1826 ( 
.A(n_1779),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1782),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1785),
.Y(n_1828)
);

NAND3xp33_ASAP7_75t_L g1829 ( 
.A(n_1771),
.B(n_1700),
.C(n_1743),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1783),
.B(n_1717),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1770),
.B(n_1734),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1751),
.B(n_1732),
.Y(n_1832)
);

AOI22xp33_ASAP7_75t_L g1833 ( 
.A1(n_1829),
.A2(n_1763),
.B1(n_1750),
.B2(n_1753),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1819),
.B(n_1783),
.Y(n_1834)
);

INVxp67_ASAP7_75t_SL g1835 ( 
.A(n_1798),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1819),
.B(n_1783),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1824),
.B(n_1781),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1822),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1830),
.B(n_1783),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1809),
.B(n_1724),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1804),
.B(n_1751),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1804),
.B(n_1797),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1797),
.B(n_1765),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1815),
.B(n_1817),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1790),
.Y(n_1845)
);

AOI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1829),
.A2(n_1750),
.B1(n_1753),
.B2(n_1763),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1830),
.B(n_1783),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1790),
.Y(n_1848)
);

AOI32xp33_ASAP7_75t_L g1849 ( 
.A1(n_1822),
.A2(n_1760),
.A3(n_1775),
.B1(n_1749),
.B2(n_1759),
.Y(n_1849)
);

OR2x6_ASAP7_75t_L g1850 ( 
.A(n_1809),
.B(n_1779),
.Y(n_1850)
);

INVx2_ASAP7_75t_SL g1851 ( 
.A(n_1811),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1796),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1796),
.Y(n_1853)
);

HB1xp67_ASAP7_75t_L g1854 ( 
.A(n_1793),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1807),
.B(n_1765),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1801),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1831),
.B(n_1820),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1801),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1808),
.Y(n_1859)
);

HB1xp67_ASAP7_75t_L g1860 ( 
.A(n_1808),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1791),
.B(n_1780),
.Y(n_1861)
);

NOR2xp33_ASAP7_75t_L g1862 ( 
.A(n_1826),
.B(n_1680),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1791),
.B(n_1813),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1812),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1802),
.B(n_1765),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1815),
.B(n_1769),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1817),
.B(n_1752),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1822),
.Y(n_1868)
);

AOI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1822),
.A2(n_1760),
.B1(n_1786),
.B2(n_1756),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1799),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1812),
.Y(n_1871)
);

INVx1_ASAP7_75t_SL g1872 ( 
.A(n_1825),
.Y(n_1872)
);

OR2x6_ASAP7_75t_L g1873 ( 
.A(n_1811),
.B(n_1637),
.Y(n_1873)
);

CKINVDCx16_ASAP7_75t_R g1874 ( 
.A(n_1826),
.Y(n_1874)
);

CKINVDCx16_ASAP7_75t_R g1875 ( 
.A(n_1826),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1821),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1799),
.Y(n_1877)
);

AND2x4_ASAP7_75t_SL g1878 ( 
.A(n_1791),
.B(n_1662),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1834),
.B(n_1825),
.Y(n_1879)
);

NAND2x1_ASAP7_75t_L g1880 ( 
.A(n_1850),
.B(n_1791),
.Y(n_1880)
);

INVxp67_ASAP7_75t_SL g1881 ( 
.A(n_1835),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1844),
.B(n_1842),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1860),
.Y(n_1883)
);

HB1xp67_ASAP7_75t_L g1884 ( 
.A(n_1854),
.Y(n_1884)
);

NOR2xp33_ASAP7_75t_L g1885 ( 
.A(n_1862),
.B(n_1680),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1845),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1834),
.B(n_1826),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1870),
.Y(n_1888)
);

O2A1O1Ixp33_ASAP7_75t_L g1889 ( 
.A1(n_1833),
.A2(n_1775),
.B(n_1749),
.C(n_1810),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1846),
.B(n_1813),
.Y(n_1890)
);

NOR2x1p5_ASAP7_75t_L g1891 ( 
.A(n_1865),
.B(n_1810),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1870),
.Y(n_1892)
);

INVx3_ASAP7_75t_L g1893 ( 
.A(n_1878),
.Y(n_1893)
);

AOI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1849),
.A2(n_1869),
.B(n_1837),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1877),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1845),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1836),
.B(n_1794),
.Y(n_1897)
);

NAND3xp33_ASAP7_75t_SL g1898 ( 
.A(n_1842),
.B(n_1786),
.C(n_1688),
.Y(n_1898)
);

O2A1O1Ixp33_ASAP7_75t_L g1899 ( 
.A1(n_1857),
.A2(n_1792),
.B(n_1799),
.C(n_1803),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1836),
.B(n_1794),
.Y(n_1900)
);

OR2x2_ASAP7_75t_L g1901 ( 
.A(n_1844),
.B(n_1832),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1848),
.Y(n_1902)
);

INVxp67_ASAP7_75t_L g1903 ( 
.A(n_1840),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1872),
.B(n_1816),
.Y(n_1904)
);

HB1xp67_ASAP7_75t_L g1905 ( 
.A(n_1843),
.Y(n_1905)
);

AND2x4_ASAP7_75t_L g1906 ( 
.A(n_1863),
.B(n_1805),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1855),
.B(n_1867),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1866),
.B(n_1816),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1866),
.B(n_1818),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1839),
.B(n_1795),
.Y(n_1910)
);

INVx1_ASAP7_75t_SL g1911 ( 
.A(n_1874),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1875),
.B(n_1818),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1848),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1853),
.B(n_1821),
.Y(n_1914)
);

OR2x2_ASAP7_75t_L g1915 ( 
.A(n_1841),
.B(n_1832),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1882),
.Y(n_1916)
);

NOR3xp33_ASAP7_75t_SL g1917 ( 
.A(n_1881),
.B(n_1688),
.C(n_1852),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_SL g1918 ( 
.A(n_1889),
.B(n_1894),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1882),
.Y(n_1919)
);

AOI21xp33_ASAP7_75t_L g1920 ( 
.A1(n_1899),
.A2(n_1868),
.B(n_1838),
.Y(n_1920)
);

OR2x2_ASAP7_75t_L g1921 ( 
.A(n_1901),
.B(n_1856),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1879),
.B(n_1861),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1886),
.Y(n_1923)
);

AOI21xp33_ASAP7_75t_L g1924 ( 
.A1(n_1890),
.A2(n_1868),
.B(n_1838),
.Y(n_1924)
);

OAI22xp5_ASAP7_75t_L g1925 ( 
.A1(n_1891),
.A2(n_1878),
.B1(n_1850),
.B2(n_1792),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1886),
.Y(n_1926)
);

AOI22xp33_ASAP7_75t_L g1927 ( 
.A1(n_1905),
.A2(n_1756),
.B1(n_1877),
.B2(n_1755),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1896),
.Y(n_1928)
);

INVxp67_ASAP7_75t_L g1929 ( 
.A(n_1884),
.Y(n_1929)
);

OAI21xp5_ASAP7_75t_L g1930 ( 
.A1(n_1898),
.A2(n_1861),
.B(n_1851),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1879),
.B(n_1839),
.Y(n_1931)
);

OAI31xp33_ASAP7_75t_SL g1932 ( 
.A1(n_1911),
.A2(n_1847),
.A3(n_1863),
.B(n_1800),
.Y(n_1932)
);

OAI221xp5_ASAP7_75t_L g1933 ( 
.A1(n_1911),
.A2(n_1873),
.B1(n_1841),
.B2(n_1851),
.C(n_1756),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1897),
.B(n_1847),
.Y(n_1934)
);

OAI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1891),
.A2(n_1850),
.B1(n_1805),
.B2(n_1873),
.Y(n_1935)
);

INVx1_ASAP7_75t_SL g1936 ( 
.A(n_1887),
.Y(n_1936)
);

AOI22xp5_ASAP7_75t_L g1937 ( 
.A1(n_1888),
.A2(n_1756),
.B1(n_1873),
.B2(n_1755),
.Y(n_1937)
);

OAI221xp5_ASAP7_75t_L g1938 ( 
.A1(n_1915),
.A2(n_1873),
.B1(n_1756),
.B2(n_1871),
.C(n_1852),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1907),
.B(n_1858),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1896),
.Y(n_1940)
);

XNOR2xp5_ASAP7_75t_L g1941 ( 
.A(n_1887),
.B(n_1638),
.Y(n_1941)
);

OAI211xp5_ASAP7_75t_SL g1942 ( 
.A1(n_1903),
.A2(n_1871),
.B(n_1876),
.C(n_1864),
.Y(n_1942)
);

OAI22xp5_ASAP7_75t_L g1943 ( 
.A1(n_1918),
.A2(n_1893),
.B1(n_1912),
.B2(n_1909),
.Y(n_1943)
);

OAI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1918),
.A2(n_1893),
.B1(n_1908),
.B2(n_1904),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1916),
.Y(n_1945)
);

INVx1_ASAP7_75t_SL g1946 ( 
.A(n_1936),
.Y(n_1946)
);

NOR2xp33_ASAP7_75t_SL g1947 ( 
.A(n_1931),
.B(n_1885),
.Y(n_1947)
);

AOI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1938),
.A2(n_1895),
.B1(n_1888),
.B2(n_1892),
.Y(n_1948)
);

OR2x2_ASAP7_75t_L g1949 ( 
.A(n_1919),
.B(n_1901),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1921),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1934),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1921),
.Y(n_1952)
);

OR2x2_ASAP7_75t_L g1953 ( 
.A(n_1939),
.B(n_1915),
.Y(n_1953)
);

OAI22xp5_ASAP7_75t_L g1954 ( 
.A1(n_1933),
.A2(n_1893),
.B1(n_1880),
.B2(n_1906),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1923),
.Y(n_1955)
);

AOI22xp5_ASAP7_75t_L g1956 ( 
.A1(n_1937),
.A2(n_1888),
.B1(n_1892),
.B2(n_1895),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1931),
.B(n_1883),
.Y(n_1957)
);

OR2x2_ASAP7_75t_L g1958 ( 
.A(n_1929),
.B(n_1883),
.Y(n_1958)
);

AOI22xp5_ASAP7_75t_L g1959 ( 
.A1(n_1924),
.A2(n_1895),
.B1(n_1892),
.B2(n_1902),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1934),
.B(n_1897),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1926),
.Y(n_1961)
);

AOI31xp33_ASAP7_75t_SL g1962 ( 
.A1(n_1920),
.A2(n_1914),
.A3(n_1893),
.B(n_1659),
.Y(n_1962)
);

OAI22xp5_ASAP7_75t_L g1963 ( 
.A1(n_1917),
.A2(n_1880),
.B1(n_1906),
.B2(n_1910),
.Y(n_1963)
);

OAI22xp5_ASAP7_75t_L g1964 ( 
.A1(n_1930),
.A2(n_1906),
.B1(n_1910),
.B2(n_1900),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1951),
.B(n_1922),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1960),
.B(n_1922),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1949),
.Y(n_1967)
);

INVxp67_ASAP7_75t_L g1968 ( 
.A(n_1947),
.Y(n_1968)
);

INVxp67_ASAP7_75t_SL g1969 ( 
.A(n_1957),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1946),
.B(n_1932),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1950),
.B(n_1900),
.Y(n_1971)
);

AOI22xp5_ASAP7_75t_L g1972 ( 
.A1(n_1948),
.A2(n_1927),
.B1(n_1941),
.B2(n_1942),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_SL g1973 ( 
.A(n_1959),
.B(n_1944),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1958),
.Y(n_1974)
);

INVx2_ASAP7_75t_SL g1975 ( 
.A(n_1952),
.Y(n_1975)
);

OAI31xp33_ASAP7_75t_L g1976 ( 
.A1(n_1954),
.A2(n_1927),
.A3(n_1935),
.B(n_1925),
.Y(n_1976)
);

O2A1O1Ixp33_ASAP7_75t_L g1977 ( 
.A1(n_1973),
.A2(n_1962),
.B(n_1943),
.C(n_1945),
.Y(n_1977)
);

NOR2xp33_ASAP7_75t_L g1978 ( 
.A(n_1968),
.B(n_1953),
.Y(n_1978)
);

AOI22xp33_ASAP7_75t_SL g1979 ( 
.A1(n_1970),
.A2(n_1964),
.B1(n_1963),
.B2(n_1961),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_SL g1980 ( 
.A(n_1967),
.B(n_1955),
.Y(n_1980)
);

NOR4xp25_ASAP7_75t_L g1981 ( 
.A(n_1973),
.B(n_1940),
.C(n_1928),
.D(n_1902),
.Y(n_1981)
);

NOR3xp33_ASAP7_75t_L g1982 ( 
.A(n_1969),
.B(n_1974),
.C(n_1975),
.Y(n_1982)
);

OR2x2_ASAP7_75t_L g1983 ( 
.A(n_1965),
.B(n_1959),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1971),
.B(n_1956),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1971),
.B(n_1966),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_L g1986 ( 
.A(n_1975),
.B(n_1850),
.Y(n_1986)
);

AOI222xp33_ASAP7_75t_L g1987 ( 
.A1(n_1984),
.A2(n_1972),
.B1(n_1913),
.B2(n_1976),
.C1(n_1803),
.C2(n_1806),
.Y(n_1987)
);

NOR3xp33_ASAP7_75t_SL g1988 ( 
.A(n_1978),
.B(n_1913),
.C(n_1658),
.Y(n_1988)
);

A2O1A1Ixp33_ASAP7_75t_L g1989 ( 
.A1(n_1977),
.A2(n_1906),
.B(n_1859),
.C(n_1755),
.Y(n_1989)
);

AOI221xp5_ASAP7_75t_L g1990 ( 
.A1(n_1981),
.A2(n_1803),
.B1(n_1806),
.B2(n_1814),
.C(n_1766),
.Y(n_1990)
);

AOI21xp33_ASAP7_75t_L g1991 ( 
.A1(n_1983),
.A2(n_1814),
.B(n_1806),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1985),
.B(n_1823),
.Y(n_1992)
);

AOI221xp5_ASAP7_75t_L g1993 ( 
.A1(n_1989),
.A2(n_1982),
.B1(n_1980),
.B2(n_1979),
.C(n_1986),
.Y(n_1993)
);

AOI22xp5_ASAP7_75t_L g1994 ( 
.A1(n_1987),
.A2(n_1666),
.B1(n_1814),
.B2(n_1658),
.Y(n_1994)
);

OAI211xp5_ASAP7_75t_L g1995 ( 
.A1(n_1988),
.A2(n_1658),
.B(n_1800),
.C(n_1795),
.Y(n_1995)
);

AOI211xp5_ASAP7_75t_L g1996 ( 
.A1(n_1992),
.A2(n_1759),
.B(n_1762),
.C(n_1772),
.Y(n_1996)
);

AOI221xp5_ASAP7_75t_L g1997 ( 
.A1(n_1991),
.A2(n_1784),
.B1(n_1773),
.B2(n_1787),
.C(n_1757),
.Y(n_1997)
);

NOR3xp33_ASAP7_75t_L g1998 ( 
.A(n_1990),
.B(n_1646),
.C(n_1647),
.Y(n_1998)
);

NAND4xp75_ASAP7_75t_L g1999 ( 
.A(n_1993),
.B(n_1650),
.C(n_1759),
.D(n_1762),
.Y(n_1999)
);

AND5x1_ASAP7_75t_L g2000 ( 
.A(n_1994),
.B(n_1712),
.C(n_1711),
.D(n_1578),
.E(n_1647),
.Y(n_2000)
);

NOR2xp33_ASAP7_75t_L g2001 ( 
.A(n_1995),
.B(n_1578),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1996),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1998),
.Y(n_2003)
);

INVxp33_ASAP7_75t_L g2004 ( 
.A(n_2001),
.Y(n_2004)
);

NOR4xp75_ASAP7_75t_L g2005 ( 
.A(n_1999),
.B(n_1646),
.C(n_1647),
.D(n_1769),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_2001),
.B(n_2002),
.Y(n_2006)
);

NAND4xp25_ASAP7_75t_L g2007 ( 
.A(n_2006),
.B(n_2003),
.C(n_2000),
.D(n_1997),
.Y(n_2007)
);

INVx2_ASAP7_75t_L g2008 ( 
.A(n_2007),
.Y(n_2008)
);

AND2x4_ASAP7_75t_L g2009 ( 
.A(n_2008),
.B(n_2005),
.Y(n_2009)
);

INVx3_ASAP7_75t_SL g2010 ( 
.A(n_2008),
.Y(n_2010)
);

CKINVDCx20_ASAP7_75t_R g2011 ( 
.A(n_2010),
.Y(n_2011)
);

AO22x2_ASAP7_75t_L g2012 ( 
.A1(n_2009),
.A2(n_2004),
.B1(n_1828),
.B2(n_1827),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_2011),
.Y(n_2013)
);

NOR2x1p5_ASAP7_75t_L g2014 ( 
.A(n_2012),
.B(n_2004),
.Y(n_2014)
);

AOI21xp5_ASAP7_75t_L g2015 ( 
.A1(n_2013),
.A2(n_1578),
.B(n_1828),
.Y(n_2015)
);

AOI21xp33_ASAP7_75t_L g2016 ( 
.A1(n_2015),
.A2(n_2014),
.B(n_1766),
.Y(n_2016)
);

OAI22xp33_ASAP7_75t_SL g2017 ( 
.A1(n_2016),
.A2(n_1827),
.B1(n_1823),
.B2(n_1646),
.Y(n_2017)
);

AOI221xp5_ASAP7_75t_L g2018 ( 
.A1(n_2017),
.A2(n_1647),
.B1(n_1762),
.B2(n_1772),
.C(n_1787),
.Y(n_2018)
);

AOI211xp5_ASAP7_75t_L g2019 ( 
.A1(n_2018),
.A2(n_1639),
.B(n_1704),
.C(n_1664),
.Y(n_2019)
);


endmodule