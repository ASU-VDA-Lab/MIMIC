module real_jpeg_24822_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_57;
wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_38;
wire n_35;
wire n_33;
wire n_50;
wire n_29;
wire n_55;
wire n_49;
wire n_52;
wire n_10;
wire n_9;
wire n_31;
wire n_58;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_60;
wire n_44;
wire n_46;
wire n_59;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_51;
wire n_45;
wire n_25;
wire n_61;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_39;
wire n_36;
wire n_40;
wire n_41;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_26;
wire n_48;
wire n_30;
wire n_56;
wire n_16;
wire n_15;
wire n_13;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_1),
.A2(n_13),
.B1(n_14),
.B2(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_3),
.A2(n_20),
.B1(n_22),
.B2(n_32),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_3),
.B(n_14),
.C(n_15),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_3),
.A2(n_18),
.B1(n_52),
.B2(n_55),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_4),
.A2(n_13),
.B1(n_14),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_5),
.A2(n_13),
.B1(n_14),
.B2(n_21),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_5),
.A2(n_21),
.B1(n_52),
.B2(n_55),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_39),
.Y(n_8)
);

OAI21xp5_ASAP7_75t_SL g9 ( 
.A1(n_10),
.A2(n_30),
.B(n_38),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_19),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_11),
.B(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_18),
.Y(n_11)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_12),
.B(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g12 ( 
.A1(n_13),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_13),
.B(n_34),
.Y(n_33)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_15),
.A2(n_17),
.B1(n_52),
.B2(n_55),
.Y(n_57)
);

BUFx24_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_22),
.B1(n_26),
.B2(n_28),
.Y(n_19)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_23),
.A2(n_42),
.B1(n_43),
.B2(n_46),
.Y(n_41)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_26),
.Y(n_42)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_60),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_49),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_49),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_52),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);


endmodule