module fake_jpeg_10018_n_18 (n_3, n_2, n_1, n_0, n_4, n_18);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_18;

wire n_13;
wire n_11;
wire n_14;
wire n_17;
wire n_16;
wire n_10;
wire n_12;
wire n_8;
wire n_9;
wire n_15;
wire n_6;
wire n_5;
wire n_7;

BUFx6f_ASAP7_75t_L g5 ( 
.A(n_0),
.Y(n_5)
);

NOR2xp33_ASAP7_75t_SL g6 ( 
.A(n_1),
.B(n_2),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_8),
.Y(n_9)
);

NAND2xp33_ASAP7_75t_SL g12 ( 
.A(n_9),
.B(n_11),
.Y(n_12)
);

AND2x6_ASAP7_75t_L g10 ( 
.A(n_7),
.B(n_0),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_10),
.B(n_11),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_6),
.B(n_0),
.Y(n_11)
);

AO22x1_ASAP7_75t_L g14 ( 
.A1(n_13),
.A2(n_7),
.B1(n_3),
.B2(n_4),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g16 ( 
.A1(n_14),
.A2(n_15),
.B(n_13),
.Y(n_16)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

AOI22xp33_ASAP7_75t_L g17 ( 
.A1(n_16),
.A2(n_8),
.B1(n_5),
.B2(n_3),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_17),
.A2(n_5),
.B(n_1),
.Y(n_18)
);


endmodule