module fake_jpeg_1697_n_319 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_10),
.B(n_11),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_29),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g137 ( 
.A(n_46),
.Y(n_137)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_47),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_49),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_20),
.Y(n_50)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_34),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_53),
.B(n_61),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_54),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_55),
.A2(n_45),
.B1(n_50),
.B2(n_38),
.Y(n_93)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_29),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g134 ( 
.A(n_57),
.Y(n_134)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_1),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_37),
.B(n_1),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_82),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_4),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_64),
.B(n_77),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_33),
.A2(n_4),
.B(n_5),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_67),
.B(n_36),
.C(n_41),
.Y(n_119)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_75),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_76),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_17),
.B(n_26),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g94 ( 
.A(n_79),
.B(n_83),
.Y(n_94)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_80),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_81),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_21),
.B(n_6),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_22),
.B(n_6),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_86),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_85),
.B(n_87),
.Y(n_136)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_SL g117 ( 
.A1(n_88),
.A2(n_19),
.B(n_35),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_26),
.B(n_6),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_7),
.Y(n_102)
);

OA22x2_ASAP7_75t_L g165 ( 
.A1(n_93),
.A2(n_83),
.B1(n_81),
.B2(n_76),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_56),
.B(n_27),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_95),
.B(n_102),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_27),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_110),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_30),
.C(n_36),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_55),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_31),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_47),
.B(n_31),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_122),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_48),
.A2(n_30),
.B1(n_45),
.B2(n_35),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_115),
.A2(n_120),
.B1(n_72),
.B2(n_74),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_117),
.A2(n_94),
.B(n_93),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_119),
.B(n_15),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_54),
.A2(n_41),
.B1(n_19),
.B2(n_40),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_7),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_73),
.B(n_8),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_131),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_51),
.B(n_9),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_59),
.B(n_11),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_11),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_78),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_133),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_60),
.A2(n_19),
.B1(n_40),
.B2(n_39),
.Y(n_135)
);

OA22x2_ASAP7_75t_SL g177 ( 
.A1(n_135),
.A2(n_19),
.B1(n_25),
.B2(n_39),
.Y(n_177)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_142),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_143),
.B(n_44),
.Y(n_210)
);

FAx1_ASAP7_75t_SL g144 ( 
.A(n_106),
.B(n_52),
.CI(n_88),
.CON(n_144),
.SN(n_144)
);

MAJIxp5_ASAP7_75t_SL g206 ( 
.A(n_144),
.B(n_171),
.C(n_25),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_135),
.A2(n_58),
.B1(n_87),
.B2(n_65),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_145),
.Y(n_195)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_146),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_91),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_147),
.Y(n_197)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_148),
.Y(n_200)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_97),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_154),
.Y(n_183)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_151),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_152),
.Y(n_193)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_91),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_157),
.Y(n_187)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_158),
.B(n_159),
.Y(n_207)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_160),
.B(n_166),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_137),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_161),
.B(n_162),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_138),
.Y(n_162)
);

INVx13_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_163),
.B(n_164),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_165),
.A2(n_139),
.B1(n_125),
.B2(n_101),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_136),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_168),
.A2(n_140),
.B(n_108),
.Y(n_194)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_104),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_172),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_90),
.B(n_13),
.Y(n_170)
);

NOR2xp67_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_173),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_107),
.B(n_15),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_109),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_175),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_121),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_178),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_177),
.A2(n_182),
.B1(n_127),
.B2(n_99),
.Y(n_184)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_109),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_100),
.B(n_16),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_180),
.Y(n_192)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_128),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_136),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_113),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_184),
.A2(n_202),
.B1(n_172),
.B2(n_165),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_168),
.A2(n_115),
.B1(n_126),
.B2(n_139),
.Y(n_185)
);

AO22x1_ASAP7_75t_L g227 ( 
.A1(n_185),
.A2(n_204),
.B1(n_209),
.B2(n_138),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_189),
.A2(n_177),
.B1(n_165),
.B2(n_175),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_194),
.A2(n_155),
.B(n_156),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_210),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_143),
.B(n_112),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_208),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_177),
.A2(n_121),
.B1(n_108),
.B2(n_112),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_145),
.A2(n_101),
.B1(n_134),
.B2(n_123),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_153),
.Y(n_231)
);

OAI32xp33_ASAP7_75t_L g208 ( 
.A1(n_144),
.A2(n_96),
.A3(n_19),
.B1(n_98),
.B2(n_123),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_144),
.A2(n_105),
.B1(n_96),
.B2(n_98),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_141),
.B(n_118),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_190),
.Y(n_214)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_214),
.Y(n_244)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_190),
.Y(n_216)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_188),
.Y(n_217)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_217),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_218),
.A2(n_233),
.B1(n_236),
.B2(n_237),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_219),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_203),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_220),
.B(n_221),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_196),
.B(n_149),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_188),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_222),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_155),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_210),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_191),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_224),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_225),
.A2(n_227),
.B1(n_185),
.B2(n_189),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_167),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_226),
.B(n_192),
.Y(n_252)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_186),
.Y(n_228)
);

OAI21xp33_ASAP7_75t_SL g243 ( 
.A1(n_228),
.A2(n_232),
.B(n_235),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_231),
.A2(n_212),
.B(n_206),
.Y(n_239)
);

INVxp67_ASAP7_75t_SL g232 ( 
.A(n_197),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_195),
.A2(n_176),
.B1(n_180),
.B2(n_151),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_187),
.Y(n_234)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_234),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_207),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_186),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_235),
.A2(n_194),
.B(n_195),
.Y(n_238)
);

INVxp67_ASAP7_75t_SL g265 ( 
.A(n_238),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_239),
.B(n_227),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_245),
.B(n_249),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_230),
.A2(n_208),
.B(n_209),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_211),
.C(n_171),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_251),
.C(n_224),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_213),
.C(n_198),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_252),
.A2(n_256),
.B1(n_225),
.B2(n_236),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_215),
.A2(n_202),
.B(n_184),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_255),
.A2(n_227),
.B1(n_228),
.B2(n_237),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_271),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_258),
.A2(n_264),
.B1(n_270),
.B2(n_244),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_215),
.C(n_223),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_266),
.C(n_268),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_242),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_261),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_254),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_256),
.A2(n_218),
.B1(n_217),
.B2(n_222),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_262),
.A2(n_272),
.B1(n_248),
.B2(n_219),
.Y(n_284)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_240),
.Y(n_263)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_263),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_231),
.C(n_216),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_254),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_267),
.A2(n_242),
.B(n_248),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_231),
.C(n_214),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_240),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_255),
.A2(n_220),
.B1(n_204),
.B2(n_221),
.Y(n_272)
);

AOI321xp33_ASAP7_75t_L g275 ( 
.A1(n_266),
.A2(n_239),
.A3(n_249),
.B1(n_246),
.B2(n_244),
.C(n_247),
.Y(n_275)
);

NOR3xp33_ASAP7_75t_SL g288 ( 
.A(n_275),
.B(n_278),
.C(n_259),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_276),
.A2(n_262),
.B1(n_261),
.B2(n_267),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_265),
.A2(n_238),
.B(n_241),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_277),
.A2(n_281),
.B(n_272),
.Y(n_285)
);

NOR4xp25_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_246),
.C(n_253),
.D(n_247),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_243),
.C(n_198),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_283),
.C(n_270),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_183),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_284),
.A2(n_277),
.B1(n_282),
.B2(n_274),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_285),
.A2(n_279),
.B(n_275),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_286),
.A2(n_193),
.B1(n_273),
.B2(n_152),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_284),
.A2(n_258),
.B1(n_271),
.B2(n_263),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_287),
.A2(n_290),
.B1(n_147),
.B2(n_163),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_291),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_294),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_219),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_205),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_293),
.Y(n_302)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_283),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_201),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_296),
.A2(n_298),
.B(n_292),
.Y(n_305)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_297),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_288),
.A2(n_200),
.B(n_197),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_200),
.C(n_105),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_289),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_287),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_306),
.Y(n_308)
);

OAI21x1_ASAP7_75t_L g309 ( 
.A1(n_305),
.A2(n_307),
.B(n_296),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_292),
.Y(n_307)
);

OA21x2_ASAP7_75t_L g312 ( 
.A1(n_309),
.A2(n_307),
.B(n_169),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_304),
.A2(n_286),
.B1(n_301),
.B2(n_299),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_311),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_306),
.A2(n_302),
.B1(n_295),
.B2(n_300),
.Y(n_311)
);

OAI21x1_ASAP7_75t_L g316 ( 
.A1(n_312),
.A2(n_313),
.B(n_308),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_308),
.A2(n_16),
.B(n_44),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_314),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_316),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_315),
.B(n_311),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_44),
.B(n_317),
.Y(n_319)
);


endmodule