module fake_jpeg_117_n_187 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_187);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_21),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_28),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_6),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_34),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_17),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_14),
.B(n_43),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_74),
.Y(n_81)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_60),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_66),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_51),
.B(n_61),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_56),
.B(n_75),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_51),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_83),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_61),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_67),
.C(n_53),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_86),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_76),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_59),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_56),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_64),
.B1(n_66),
.B2(n_62),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_89),
.A2(n_54),
.B1(n_55),
.B2(n_63),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_94),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_78),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_85),
.B(n_48),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_93),
.B(n_0),
.Y(n_111)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_88),
.A2(n_64),
.B1(n_58),
.B2(n_73),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_96),
.A2(n_97),
.B1(n_78),
.B2(n_91),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_88),
.A2(n_67),
.B1(n_53),
.B2(n_48),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_104),
.Y(n_116)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_80),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_101),
.B(n_105),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_80),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_77),
.Y(n_103)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_103),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_79),
.A2(n_55),
.B1(n_54),
.B2(n_57),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_65),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_108),
.B(n_123),
.Y(n_126)
);

AOI32xp33_ASAP7_75t_L g109 ( 
.A1(n_105),
.A2(n_68),
.A3(n_52),
.B1(n_3),
.B2(n_4),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_111),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_98),
.A2(n_0),
.B(n_1),
.C(n_3),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_121),
.Y(n_133)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_47),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_104),
.B(n_1),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_143)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_107),
.A2(n_92),
.B1(n_5),
.B2(n_7),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_136),
.B1(n_145),
.B2(n_132),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_120),
.A2(n_24),
.B1(n_46),
.B2(n_45),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_129),
.A2(n_143),
.B1(n_145),
.B2(n_11),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_132),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_39),
.C(n_38),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_119),
.B(n_116),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_134),
.B(n_146),
.Y(n_154)
);

AO22x1_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_37),
.B1(n_36),
.B2(n_35),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_129),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_33),
.C(n_32),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_23),
.Y(n_155)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_140),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_4),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_8),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_142),
.Y(n_161)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_144),
.Y(n_148)
);

AO21x2_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_30),
.B(n_29),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_133),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_150),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_131),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_151),
.A2(n_156),
.B1(n_159),
.B2(n_145),
.Y(n_165)
);

NOR3xp33_ASAP7_75t_SL g152 ( 
.A(n_135),
.B(n_112),
.C(n_31),
.Y(n_152)
);

AOI221xp5_ASAP7_75t_L g163 ( 
.A1(n_152),
.A2(n_158),
.B1(n_160),
.B2(n_137),
.C(n_14),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_25),
.Y(n_153)
);

OAI32xp33_ASAP7_75t_L g164 ( 
.A1(n_153),
.A2(n_128),
.A3(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_157),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_9),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_138),
.B(n_10),
.Y(n_158)
);

NOR3xp33_ASAP7_75t_SL g160 ( 
.A(n_127),
.B(n_11),
.C(n_12),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_163),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_165),
.Y(n_172)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_168),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_145),
.B(n_15),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_13),
.B(n_18),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_169),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_170),
.A2(n_156),
.B1(n_161),
.B2(n_147),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_173),
.B(n_170),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_162),
.C(n_166),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_176),
.B(n_177),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_162),
.C(n_153),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_175),
.C(n_174),
.Y(n_179)
);

AOI31xp67_ASAP7_75t_SL g181 ( 
.A1(n_179),
.A2(n_152),
.A3(n_172),
.B(n_160),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_181),
.A2(n_172),
.B(n_174),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_182),
.B(n_180),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_183),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_13),
.C(n_18),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_19),
.B(n_20),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_19),
.Y(n_187)
);


endmodule