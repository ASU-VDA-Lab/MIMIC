module fake_jpeg_22905_n_42 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_42);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_42;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx5_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_1),
.B(n_2),
.Y(n_8)
);

CKINVDCx9p33_ASAP7_75t_R g9 ( 
.A(n_4),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_0),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_19),
.Y(n_26)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_3),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_8),
.A2(n_6),
.B(n_3),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_20),
.A2(n_15),
.B(n_23),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_4),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_22),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_6),
.Y(n_22)
);

AND2x6_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_14),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_17),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_12),
.A2(n_13),
.B1(n_7),
.B2(n_14),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_25),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_10),
.A2(n_15),
.B1(n_12),
.B2(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_16),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_10),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_30),
.B(n_29),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_33),
.B(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_36),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

AOI322xp5_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_37),
.A3(n_40),
.B1(n_33),
.B2(n_35),
.C1(n_32),
.C2(n_38),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_39),
.Y(n_42)
);


endmodule