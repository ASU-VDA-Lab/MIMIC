module real_jpeg_10225_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_215;
wire n_166;
wire n_221;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_1),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_1),
.A2(n_55),
.B1(n_56),
.B2(n_65),
.Y(n_67)
);

AOI21xp33_ASAP7_75t_L g136 ( 
.A1(n_1),
.A2(n_8),
.B(n_55),
.Y(n_136)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_4),
.A2(n_36),
.B(n_38),
.C(n_39),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_4),
.B(n_36),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_4),
.A2(n_21),
.B1(n_25),
.B2(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_4),
.A2(n_8),
.B(n_21),
.Y(n_183)
);

BUFx6f_ASAP7_75t_SL g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_7),
.A2(n_36),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_7),
.A2(n_43),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_7),
.A2(n_43),
.B1(n_64),
.B2(n_70),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_7),
.A2(n_21),
.B1(n_25),
.B2(n_43),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_8),
.A2(n_36),
.B1(n_42),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_8),
.A2(n_45),
.B1(n_55),
.B2(n_56),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_8),
.A2(n_45),
.B1(n_64),
.B2(n_70),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_8),
.A2(n_21),
.B1(n_25),
.B2(n_45),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_8),
.B(n_94),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_8),
.B(n_50),
.Y(n_199)
);

O2A1O1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_8),
.A2(n_52),
.B(n_56),
.C(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_9),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_9),
.A2(n_24),
.B1(n_36),
.B2(n_42),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_11),
.A2(n_21),
.B1(n_25),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_11),
.A2(n_32),
.B1(n_36),
.B2(n_42),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_123),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_121),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_100),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_15),
.B(n_100),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_73),
.C(n_82),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_16),
.A2(n_17),
.B1(n_73),
.B2(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_46),
.B1(n_47),
.B2(n_72),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_18),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_33),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_19),
.A2(n_33),
.B1(n_34),
.B2(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_19),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_20),
.Y(n_85)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_28),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_25),
.B(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_26),
.B(n_29),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_27),
.B(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_27),
.A2(n_28),
.B1(n_88),
.B2(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_28),
.A2(n_85),
.B(n_86),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_28),
.B(n_45),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_29),
.A2(n_87),
.B(n_171),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_31),
.B(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_33),
.A2(n_34),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_33),
.A2(n_34),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_34),
.B(n_137),
.C(n_198),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_34),
.B(n_215),
.C(n_221),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_39),
.B1(n_41),
.B2(n_44),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_35),
.B(n_44),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_35),
.A2(n_39),
.B1(n_78),
.B2(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_35),
.B(n_39),
.Y(n_152)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_42),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

OAI21xp33_ASAP7_75t_SL g208 ( 
.A1(n_36),
.A2(n_45),
.B(n_53),
.Y(n_208)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_39),
.A2(n_78),
.B(n_79),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_39),
.B(n_45),
.Y(n_190)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_40),
.A2(n_42),
.B(n_45),
.C(n_183),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_44),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_45),
.A2(n_64),
.B(n_65),
.C(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_61),
.B2(n_62),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_48),
.A2(n_49),
.B1(n_150),
.B2(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_48),
.A2(n_49),
.B1(n_89),
.B2(n_90),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_49),
.B(n_61),
.C(n_72),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_49),
.B(n_93),
.C(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_49),
.B(n_90),
.C(n_210),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_54),
.B(n_57),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_50),
.B(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_50),
.A2(n_54),
.B1(n_99),
.B2(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_51),
.A2(n_52),
.B(n_56),
.C(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_52),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_56),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_55),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_58),
.B(n_98),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_61),
.B(n_105),
.C(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_61),
.A2(n_62),
.B1(n_104),
.B2(n_105),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_71),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_63),
.B(n_67),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B(n_66),
.C(n_67),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_65),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_64),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_67),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_69),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_71),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_73),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_77),
.B2(n_81),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_74),
.A2(n_75),
.B1(n_113),
.B2(n_116),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_77),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_76),
.B(n_88),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_77),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_91),
.B(n_92),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_82),
.B(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_93),
.C(n_96),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_89),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_84),
.A2(n_89),
.B1(n_90),
.B2(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_84),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_89),
.A2(n_90),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_90),
.B(n_182),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_93),
.A2(n_96),
.B1(n_97),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_93),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_93),
.A2(n_128),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_119),
.B2(n_120),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_110),
.B1(n_117),
.B2(n_118),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_103),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_107),
.B(n_109),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_107),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_104),
.A2(n_105),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_105),
.B(n_169),
.C(n_170),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_110),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_113),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_119),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_142),
.B(n_231),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_139),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_125),
.B(n_139),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.C(n_131),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_129),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_131),
.A2(n_132),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_133),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_134),
.A2(n_135),
.B1(n_137),
.B2(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_137),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_137),
.B(n_190),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_137),
.A2(n_166),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_138),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_173),
.Y(n_142)
);

INVxp33_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_158),
.B(n_172),
.Y(n_144)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_145),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_155),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_146),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_146),
.B(n_155),
.Y(n_172)
);

FAx1_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_149),
.CI(n_153),
.CON(n_146),
.SN(n_146)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_150),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_159),
.B(n_160),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.C(n_167),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_161),
.B(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_165),
.A2(n_167),
.B1(n_168),
.B2(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_165),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_169),
.A2(n_170),
.B1(n_186),
.B2(n_218),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_169),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_170),
.B(n_180),
.Y(n_192)
);

NOR3xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_229),
.C(n_230),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_223),
.B(n_228),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_212),
.B(n_222),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_201),
.B(n_211),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_193),
.B(n_200),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_184),
.B(n_192),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_189),
.B(n_191),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_194),
.B(n_195),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_202),
.B(n_203),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_210),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_206),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_209),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_213),
.B(n_214),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_220),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_224),
.B(n_225),
.Y(n_228)
);


endmodule