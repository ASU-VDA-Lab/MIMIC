module fake_jpeg_12485_n_65 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_65);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_65;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_51;
wire n_47;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_32;

INVx2_ASAP7_75t_SL g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_8),
.B(n_4),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_11),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_1),
.B(n_16),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_35),
.Y(n_39)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

OAI21xp33_ASAP7_75t_SL g37 ( 
.A1(n_33),
.A2(n_23),
.B(n_29),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_5),
.B(n_6),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_41),
.Y(n_47)
);

AND2x6_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_14),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_23),
.C(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_2),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_48),
.C(n_50),
.Y(n_57)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_26),
.B1(n_2),
.B2(n_0),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_49),
.A2(n_7),
.B1(n_10),
.B2(n_12),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_51),
.A2(n_52),
.B(n_13),
.Y(n_56)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_38),
.C(n_9),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_55),
.C(n_58),
.Y(n_60)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_57),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_61),
.Y(n_62)
);

AOI322xp5_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_59),
.A3(n_60),
.B1(n_54),
.B2(n_53),
.C1(n_22),
.C2(n_19),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

OA21x2_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_59),
.B(n_20),
.Y(n_65)
);


endmodule