module fake_jpeg_14050_n_557 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_557);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_557;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_4),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_11),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_9),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_61),
.Y(n_178)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_18),
.Y(n_62)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_62),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_63),
.Y(n_133)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_65),
.Y(n_143)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_66),
.Y(n_157)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_68),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_21),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_69),
.B(n_73),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_70),
.Y(n_154)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_71),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_72),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_17),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_74),
.Y(n_160)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_75),
.Y(n_131)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_76),
.Y(n_136)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_77),
.B(n_78),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_21),
.Y(n_78)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_18),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_79),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_80),
.Y(n_147)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_81),
.B(n_84),
.Y(n_151)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_18),
.Y(n_83)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_83),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_23),
.B(n_0),
.Y(n_84)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_85),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_86),
.Y(n_190)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_27),
.B(n_2),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_88),
.B(n_91),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_89),
.Y(n_192)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_90),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_46),
.B(n_2),
.C(n_5),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_92),
.B(n_93),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_46),
.B(n_30),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_43),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_94),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_95),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_26),
.Y(n_97)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

BUFx16f_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_99),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_26),
.Y(n_100)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_32),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_101),
.B(n_102),
.Y(n_183)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_41),
.B(n_2),
.Y(n_102)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_26),
.Y(n_103)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_104),
.Y(n_159)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_105),
.Y(n_172)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_33),
.Y(n_106)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_107),
.Y(n_187)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_36),
.Y(n_108)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_108),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_18),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_109),
.B(n_112),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_40),
.Y(n_110)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_36),
.Y(n_111)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_111),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_21),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_40),
.Y(n_114)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_114),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_115),
.Y(n_189)
);

BUFx10_ASAP7_75t_L g116 ( 
.A(n_40),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_116),
.Y(n_153)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_40),
.Y(n_117)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_37),
.Y(n_118)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_118),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_119),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_21),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_120),
.B(n_31),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_39),
.Y(n_121)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_121),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_23),
.B(n_16),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_2),
.Y(n_164)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_27),
.Y(n_123)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_123),
.Y(n_198)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_39),
.Y(n_124)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_124),
.Y(n_191)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_40),
.Y(n_125)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_125),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_72),
.A2(n_59),
.B1(n_54),
.B2(n_40),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_128),
.A2(n_134),
.B1(n_145),
.B2(n_173),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_63),
.A2(n_95),
.B1(n_70),
.B2(n_121),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_129),
.A2(n_158),
.B1(n_28),
.B2(n_48),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_73),
.B(n_54),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_132),
.B(n_142),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_72),
.A2(n_54),
.B1(n_25),
.B2(n_53),
.Y(n_134)
);

AND2x4_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_38),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_103),
.A2(n_25),
.B1(n_49),
.B2(n_45),
.Y(n_145)
);

AND2x2_ASAP7_75t_SL g146 ( 
.A(n_94),
.B(n_25),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_146),
.B(n_96),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_74),
.A2(n_100),
.B1(n_86),
.B2(n_97),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_162),
.B(n_181),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_164),
.B(n_175),
.Y(n_220)
);

NAND2xp33_ASAP7_75t_SL g168 ( 
.A(n_75),
.B(n_57),
.Y(n_168)
);

OR2x2_ASAP7_75t_SL g235 ( 
.A(n_168),
.B(n_116),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_80),
.A2(n_45),
.B1(n_53),
.B2(n_39),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_105),
.B(n_31),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_174),
.B(n_177),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_109),
.B(n_30),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_85),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_124),
.A2(n_45),
.B1(n_53),
.B2(n_49),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_179),
.A2(n_195),
.B1(n_49),
.B2(n_38),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_61),
.B(n_35),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_180),
.B(n_199),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_113),
.B(n_57),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_107),
.A2(n_45),
.B1(n_53),
.B2(n_49),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_83),
.Y(n_196)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_196),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_90),
.B(n_24),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_117),
.B(n_24),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_200),
.B(n_62),
.Y(n_254)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_115),
.Y(n_203)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_203),
.Y(n_215)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_205),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_140),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_206),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_129),
.A2(n_29),
.B1(n_58),
.B2(n_56),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_207),
.A2(n_245),
.B1(n_195),
.B2(n_138),
.Y(n_292)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_137),
.Y(n_208)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_208),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_135),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_211),
.B(n_223),
.Y(n_278)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_133),
.Y(n_212)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_212),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_159),
.A2(n_80),
.B1(n_89),
.B2(n_96),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_213),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_184),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_216),
.Y(n_310)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_152),
.Y(n_218)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_218),
.Y(n_275)
);

AO22x2_ASAP7_75t_L g219 ( 
.A1(n_158),
.A2(n_116),
.B1(n_125),
.B2(n_119),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_219),
.B(n_235),
.Y(n_277)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_184),
.Y(n_221)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_221),
.Y(n_276)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_161),
.Y(n_222)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_222),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_135),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_171),
.B(n_27),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_224),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_193),
.Y(n_225)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_225),
.Y(n_281)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_191),
.Y(n_226)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_226),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_188),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_227),
.B(n_231),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_228),
.A2(n_263),
.B1(n_230),
.B2(n_272),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_188),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_232),
.B(n_240),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_144),
.Y(n_233)
);

BUFx8_ASAP7_75t_L g282 ( 
.A(n_233),
.Y(n_282)
);

BUFx12f_ASAP7_75t_L g234 ( 
.A(n_156),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_234),
.B(n_237),
.Y(n_295)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_126),
.Y(n_236)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_236),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_181),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_133),
.Y(n_238)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_238),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_165),
.A2(n_89),
.B1(n_51),
.B2(n_37),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_239),
.A2(n_246),
.B1(n_259),
.B2(n_260),
.Y(n_296)
);

INVx13_ASAP7_75t_L g240 ( 
.A(n_127),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_171),
.B(n_98),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_241),
.B(n_242),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_143),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_163),
.Y(n_243)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_243),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_167),
.B(n_51),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_262),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_170),
.A2(n_48),
.B1(n_42),
.B2(n_56),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_131),
.Y(n_247)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_247),
.Y(n_302)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_154),
.Y(n_248)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_248),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_157),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_249),
.B(n_251),
.Y(n_326)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_147),
.Y(n_250)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_250),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_151),
.B(n_42),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_141),
.Y(n_252)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_252),
.Y(n_309)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_201),
.Y(n_253)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_253),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_254),
.B(n_255),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_151),
.B(n_167),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_132),
.B(n_5),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_256),
.B(n_272),
.C(n_153),
.Y(n_299)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_154),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_257),
.B(n_258),
.Y(n_328)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_192),
.Y(n_258)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_149),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_148),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_146),
.A2(n_28),
.B1(n_55),
.B2(n_35),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_261),
.A2(n_269),
.B(n_50),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_166),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_183),
.A2(n_58),
.B1(n_55),
.B2(n_29),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_155),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_264),
.A2(n_265),
.B1(n_267),
.B2(n_268),
.Y(n_303)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_187),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_198),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_270),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_160),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_160),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_189),
.A2(n_50),
.B1(n_47),
.B2(n_21),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_197),
.Y(n_270)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_194),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_271),
.A2(n_185),
.B1(n_176),
.B2(n_138),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_142),
.B(n_6),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_130),
.B(n_6),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_6),
.Y(n_291)
);

AOI32xp33_ASAP7_75t_L g283 ( 
.A1(n_244),
.A2(n_183),
.A3(n_142),
.B1(n_130),
.B2(n_153),
.Y(n_283)
);

FAx1_ASAP7_75t_SL g358 ( 
.A(n_283),
.B(n_240),
.CI(n_259),
.CON(n_358),
.SN(n_358)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_210),
.A2(n_178),
.B1(n_128),
.B2(n_150),
.Y(n_285)
);

OA21x2_ASAP7_75t_L g337 ( 
.A1(n_285),
.A2(n_290),
.B(n_256),
.Y(n_337)
);

O2A1O1Ixp33_ASAP7_75t_L g290 ( 
.A1(n_235),
.A2(n_134),
.B(n_173),
.C(n_179),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_291),
.B(n_7),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_292),
.A2(n_300),
.B1(n_313),
.B2(n_316),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_297),
.A2(n_311),
.B1(n_315),
.B2(n_324),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_231),
.B(n_139),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_298),
.B(n_312),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_299),
.B(n_243),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_245),
.A2(n_261),
.B1(n_219),
.B2(n_209),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_305),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_229),
.B(n_172),
.C(n_136),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_307),
.B(n_317),
.C(n_232),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_219),
.A2(n_186),
.B1(n_190),
.B2(n_169),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_220),
.B(n_272),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_219),
.A2(n_186),
.B1(n_190),
.B2(n_204),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_229),
.A2(n_202),
.B1(n_50),
.B2(n_47),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_217),
.A2(n_50),
.B1(n_47),
.B2(n_9),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_229),
.B(n_50),
.C(n_47),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_318),
.A2(n_271),
.B1(n_250),
.B2(n_248),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_269),
.A2(n_47),
.B1(n_7),
.B2(n_11),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_322),
.A2(n_325),
.B1(n_256),
.B2(n_243),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_232),
.A2(n_6),
.B1(n_7),
.B2(n_12),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_208),
.A2(n_7),
.B1(n_13),
.B2(n_14),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g330 ( 
.A1(n_300),
.A2(n_253),
.B1(n_225),
.B2(n_270),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g375 ( 
.A1(n_330),
.A2(n_314),
.B1(n_274),
.B2(n_309),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_331),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_277),
.A2(n_222),
.B1(n_225),
.B2(n_252),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_332),
.A2(n_354),
.B1(n_366),
.B2(n_325),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_295),
.B(n_234),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_333),
.B(n_336),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_334),
.B(n_335),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_288),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_323),
.B(n_234),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_337),
.A2(n_353),
.B(n_285),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_308),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_338),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_288),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_339),
.B(n_342),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_341),
.B(n_346),
.C(n_351),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_292),
.A2(n_260),
.B1(n_236),
.B2(n_265),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_343),
.B(n_348),
.Y(n_373)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_301),
.Y(n_344)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_344),
.Y(n_371)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_301),
.Y(n_345)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_345),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_307),
.B(n_317),
.C(n_280),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_319),
.Y(n_347)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_347),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_294),
.B(n_226),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_313),
.A2(n_205),
.B1(n_218),
.B2(n_214),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_349),
.B(n_350),
.Y(n_392)
);

OA22x2_ASAP7_75t_L g350 ( 
.A1(n_277),
.A2(n_221),
.B1(n_215),
.B2(n_264),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_280),
.B(n_258),
.C(n_206),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_326),
.B(n_233),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_352),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_277),
.A2(n_212),
.B1(n_257),
.B2(n_268),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_319),
.Y(n_355)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_355),
.Y(n_382)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_281),
.Y(n_356)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_356),
.Y(n_387)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_308),
.Y(n_357)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_357),
.Y(n_390)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_358),
.B(n_299),
.Y(n_388)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_279),
.Y(n_359)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_359),
.Y(n_393)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_279),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_360),
.B(n_363),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_290),
.A2(n_238),
.B1(n_267),
.B2(n_16),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_362),
.B(n_367),
.Y(n_397)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_276),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_278),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_364),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_297),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_281),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_276),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_368),
.B(n_370),
.Y(n_401)
);

INVx6_ASAP7_75t_L g369 ( 
.A(n_328),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_369),
.B(n_302),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_327),
.B(n_14),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_374),
.Y(n_410)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_375),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_376),
.B(n_398),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_337),
.A2(n_287),
.B1(n_298),
.B2(n_322),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_378),
.A2(n_396),
.B1(n_329),
.B2(n_331),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_337),
.A2(n_287),
.B1(n_316),
.B2(n_314),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_383),
.A2(n_362),
.B1(n_334),
.B2(n_343),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_332),
.A2(n_296),
.B(n_318),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_384),
.A2(n_389),
.B(n_394),
.Y(n_425)
);

CKINVDCx14_ASAP7_75t_R g386 ( 
.A(n_348),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_386),
.B(n_350),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_388),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_358),
.A2(n_314),
.B(n_320),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_353),
.A2(n_274),
.B(n_306),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_361),
.A2(n_320),
.B1(n_312),
.B2(n_283),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_335),
.A2(n_306),
.B(n_303),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_350),
.A2(n_293),
.B(n_302),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_399),
.B(n_402),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_341),
.B(n_315),
.C(n_309),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_404),
.B(n_360),
.C(n_359),
.Y(n_428)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_406),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_385),
.B(n_346),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_407),
.B(n_418),
.C(n_428),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_395),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_408),
.B(n_411),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_392),
.A2(n_365),
.B1(n_354),
.B2(n_358),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_409),
.A2(n_413),
.B1(n_415),
.B2(n_417),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_377),
.B(n_369),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_391),
.B(n_340),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_412),
.B(n_429),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_397),
.A2(n_329),
.B1(n_340),
.B2(n_351),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_414),
.A2(n_431),
.B1(n_393),
.B2(n_382),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_397),
.A2(n_392),
.B1(n_384),
.B2(n_399),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_379),
.B(n_368),
.Y(n_416)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_416),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_384),
.A2(n_399),
.B1(n_394),
.B2(n_386),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_385),
.B(n_355),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_381),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_419),
.B(n_427),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_420),
.A2(n_398),
.B1(n_373),
.B2(n_404),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_394),
.A2(n_398),
.B1(n_373),
.B2(n_379),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_424),
.A2(n_378),
.B1(n_383),
.B2(n_400),
.Y(n_453)
);

O2A1O1Ixp33_ASAP7_75t_L g426 ( 
.A1(n_374),
.A2(n_350),
.B(n_347),
.C(n_363),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_426),
.B(n_375),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_395),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_391),
.B(n_344),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_402),
.B(n_367),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_430),
.B(n_371),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_396),
.A2(n_349),
.B1(n_345),
.B2(n_356),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_380),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_432),
.Y(n_458)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_380),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_434),
.B(n_382),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_403),
.B(n_310),
.C(n_286),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_435),
.B(n_385),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_436),
.A2(n_443),
.B1(n_451),
.B2(n_409),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_433),
.A2(n_388),
.B(n_377),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_439),
.B(n_446),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_440),
.B(n_425),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_431),
.A2(n_404),
.B1(n_405),
.B2(n_389),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_407),
.B(n_388),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_445),
.B(n_447),
.Y(n_470)
);

INVxp33_ASAP7_75t_L g446 ( 
.A(n_411),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_418),
.B(n_428),
.Y(n_447)
);

A2O1A1Ixp33_ASAP7_75t_SL g479 ( 
.A1(n_448),
.A2(n_456),
.B(n_426),
.C(n_406),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_449),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_450),
.A2(n_415),
.B1(n_424),
.B2(n_423),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_420),
.A2(n_400),
.B1(n_376),
.B2(n_393),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_453),
.A2(n_423),
.B1(n_422),
.B2(n_408),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_414),
.B(n_383),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_455),
.B(n_457),
.Y(n_476)
);

OAI22x1_ASAP7_75t_L g456 ( 
.A1(n_417),
.A2(n_372),
.B1(n_387),
.B2(n_371),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_435),
.B(n_401),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_433),
.A2(n_401),
.B(n_291),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_412),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_413),
.B(n_372),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_460),
.B(n_462),
.C(n_416),
.Y(n_481)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_461),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_425),
.B(n_387),
.Y(n_462)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_449),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_464),
.B(n_466),
.Y(n_489)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_442),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_467),
.A2(n_473),
.B1(n_381),
.B2(n_357),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_468),
.B(n_482),
.C(n_454),
.Y(n_486)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_458),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_469),
.B(n_474),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_446),
.A2(n_410),
.B(n_421),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_472),
.A2(n_484),
.B(n_293),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_437),
.A2(n_422),
.B(n_421),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_475),
.A2(n_477),
.B1(n_480),
.B2(n_485),
.Y(n_487)
);

CKINVDCx14_ASAP7_75t_R g478 ( 
.A(n_438),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_478),
.B(n_463),
.Y(n_497)
);

O2A1O1Ixp33_ASAP7_75t_L g490 ( 
.A1(n_479),
.A2(n_448),
.B(n_456),
.C(n_462),
.Y(n_490)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_458),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_481),
.B(n_324),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_454),
.B(n_427),
.C(n_430),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_457),
.B(n_429),
.Y(n_483)
);

AO221x1_ASAP7_75t_L g503 ( 
.A1(n_483),
.A2(n_474),
.B1(n_464),
.B2(n_463),
.C(n_484),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_436),
.A2(n_426),
.B(n_432),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_452),
.A2(n_434),
.B1(n_419),
.B2(n_390),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_486),
.B(n_488),
.C(n_491),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_470),
.B(n_447),
.C(n_440),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_490),
.A2(n_502),
.B(n_479),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_470),
.B(n_445),
.C(n_460),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_482),
.B(n_443),
.C(n_455),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_492),
.B(n_495),
.C(n_496),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_471),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_494),
.B(n_481),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_476),
.B(n_451),
.C(n_441),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_476),
.B(n_448),
.C(n_444),
.Y(n_496)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_497),
.Y(n_507)
);

AOI321xp33_ASAP7_75t_L g498 ( 
.A1(n_466),
.A2(n_448),
.A3(n_390),
.B1(n_304),
.B2(n_289),
.C(n_286),
.Y(n_498)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_498),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_499),
.B(n_501),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_500),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_468),
.B(n_304),
.Y(n_501)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_503),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_465),
.B(n_475),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_504),
.B(n_469),
.Y(n_508)
);

NAND4xp25_ASAP7_75t_SL g506 ( 
.A(n_489),
.B(n_282),
.C(n_472),
.D(n_479),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_506),
.B(n_515),
.Y(n_523)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_508),
.Y(n_520)
);

AND2x4_ASAP7_75t_SL g510 ( 
.A(n_493),
.B(n_479),
.Y(n_510)
);

XNOR2x1_ASAP7_75t_L g527 ( 
.A(n_510),
.B(n_501),
.Y(n_527)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_512),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_487),
.B(n_480),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_517),
.A2(n_519),
.B(n_321),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_486),
.B(n_473),
.C(n_485),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_518),
.B(n_492),
.C(n_491),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_502),
.A2(n_479),
.B(n_289),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_514),
.B(n_495),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_521),
.B(n_524),
.Y(n_538)
);

BUFx24_ASAP7_75t_SL g522 ( 
.A(n_507),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g539 ( 
.A(n_522),
.B(n_509),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_SL g525 ( 
.A1(n_516),
.A2(n_490),
.B1(n_500),
.B2(n_498),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_525),
.A2(n_517),
.B(n_508),
.Y(n_536)
);

FAx1_ASAP7_75t_SL g526 ( 
.A(n_512),
.B(n_496),
.CI(n_488),
.CON(n_526),
.SN(n_526)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_526),
.B(n_531),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_527),
.B(n_510),
.C(n_518),
.Y(n_533)
);

INVx11_ASAP7_75t_L g528 ( 
.A(n_506),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_528),
.A2(n_530),
.B1(n_505),
.B2(n_511),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_519),
.A2(n_499),
.B1(n_381),
.B2(n_338),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_533),
.B(n_521),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_534),
.B(n_537),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_523),
.A2(n_520),
.B(n_529),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_535),
.A2(n_536),
.B1(n_526),
.B2(n_510),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_528),
.B(n_514),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_539),
.B(n_540),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_524),
.B(n_509),
.C(n_513),
.Y(n_540)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_542),
.Y(n_551)
);

A2O1A1Ixp33_ASAP7_75t_SL g543 ( 
.A1(n_532),
.A2(n_527),
.B(n_526),
.C(n_530),
.Y(n_543)
);

AO221x1_ASAP7_75t_L g550 ( 
.A1(n_543),
.A2(n_545),
.B1(n_282),
.B2(n_275),
.C(n_284),
.Y(n_550)
);

NOR3xp33_ASAP7_75t_SL g544 ( 
.A(n_538),
.B(n_537),
.C(n_532),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_544),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_538),
.B(n_513),
.C(n_321),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_L g549 ( 
.A1(n_546),
.A2(n_541),
.B(n_547),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_549),
.A2(n_550),
.B(n_547),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_552),
.A2(n_553),
.B(n_548),
.Y(n_554)
);

MAJx2_ASAP7_75t_L g553 ( 
.A(n_551),
.B(n_543),
.C(n_275),
.Y(n_553)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_554),
.Y(n_555)
);

O2A1O1Ixp33_ASAP7_75t_SL g556 ( 
.A1(n_555),
.A2(n_543),
.B(n_282),
.C(n_284),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_556),
.B(n_282),
.Y(n_557)
);


endmodule