module real_aes_5983_n_3 (n_0, n_2, n_1, n_3);
input n_0;
input n_2;
input n_1;
output n_3;
wire n_4;
wire n_5;
wire n_7;
wire n_9;
wire n_6;
wire n_8;
wire n_10;
wire n_11;
BUFx6f_ASAP7_75t_L g8 ( .A(n_0), .Y(n_8) );
HB1xp67_ASAP7_75t_L g9 ( .A(n_1), .Y(n_9) );
AOI22xp33_ASAP7_75t_L g3 ( .A1(n_2), .A2(n_4), .B1(n_9), .B2(n_10), .Y(n_3) );
HB1xp67_ASAP7_75t_L g4 ( .A(n_5), .Y(n_4) );
INVx2_ASAP7_75t_SL g5 ( .A(n_6), .Y(n_5) );
CKINVDCx14_ASAP7_75t_R g11 ( .A(n_6), .Y(n_11) );
BUFx2_ASAP7_75t_L g6 ( .A(n_7), .Y(n_6) );
HB1xp67_ASAP7_75t_L g7 ( .A(n_8), .Y(n_7) );
CKINVDCx20_ASAP7_75t_R g10 ( .A(n_11), .Y(n_10) );
endmodule