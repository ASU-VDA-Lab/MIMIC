module fake_jpeg_8523_n_303 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_303);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_303;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_299;
wire n_300;
wire n_211;
wire n_294;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_SL g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx8_ASAP7_75t_SL g26 ( 
.A(n_5),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_38),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_24),
.B1(n_27),
.B2(n_20),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_17),
.B1(n_29),
.B2(n_34),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_27),
.B1(n_17),
.B2(n_23),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_45),
.A2(n_59),
.B1(n_21),
.B2(n_22),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_46),
.B(n_47),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_30),
.Y(n_47)
);

INVx2_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_48),
.A2(n_22),
.B(n_31),
.Y(n_82)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_65),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_23),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_62),
.C(n_34),
.Y(n_74)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_66),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_28),
.Y(n_58)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_27),
.B1(n_24),
.B2(n_25),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_23),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_24),
.B1(n_21),
.B2(n_20),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_64),
.A2(n_50),
.B1(n_63),
.B2(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_38),
.B(n_28),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_29),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_67),
.A2(n_79),
.B1(n_81),
.B2(n_83),
.Y(n_108)
);

CKINVDCx6p67_ASAP7_75t_R g69 ( 
.A(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_69),
.Y(n_114)
);

NOR2x1_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_17),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_70),
.A2(n_71),
.B(n_82),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_53),
.A2(n_17),
.B1(n_33),
.B2(n_19),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_77),
.Y(n_99)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_20),
.B1(n_21),
.B2(n_25),
.Y(n_73)
);

OAI32xp33_ASAP7_75t_L g119 ( 
.A1(n_73),
.A2(n_49),
.A3(n_60),
.B1(n_57),
.B2(n_56),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_92),
.Y(n_106)
);

BUFx16f_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_76),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_66),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_65),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_86),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_45),
.A2(n_25),
.B1(n_31),
.B2(n_33),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_44),
.A2(n_19),
.B1(n_32),
.B2(n_18),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_85),
.Y(n_107)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_87),
.A2(n_92),
.B1(n_70),
.B2(n_69),
.Y(n_113)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_63),
.B1(n_61),
.B2(n_56),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_55),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_58),
.Y(n_109)
);

AND2x4_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_32),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_64),
.A2(n_50),
.B1(n_47),
.B2(n_53),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_94),
.A2(n_62),
.B1(n_63),
.B2(n_45),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_46),
.C(n_52),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_104),
.C(n_117),
.Y(n_123)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_111),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_103),
.A2(n_119),
.B1(n_69),
.B2(n_83),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_62),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_109),
.B(n_110),
.Y(n_132)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_85),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_118),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_113),
.A2(n_71),
.B1(n_79),
.B2(n_81),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_62),
.B(n_54),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_115),
.A2(n_91),
.B(n_68),
.Y(n_139)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_116),
.B(n_120),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_60),
.C(n_57),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_76),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_78),
.Y(n_140)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_122),
.B(n_130),
.Y(n_180)
);

OR2x2_ASAP7_75t_SL g124 ( 
.A(n_120),
.B(n_68),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_124),
.B(n_140),
.Y(n_171)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_125),
.B(n_129),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_102),
.A2(n_69),
.B(n_70),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_126),
.A2(n_150),
.B(n_116),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_89),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_137),
.Y(n_160)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_133),
.A2(n_146),
.B1(n_149),
.B2(n_114),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_74),
.C(n_69),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_139),
.Y(n_166)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_139),
.A2(n_143),
.B(n_148),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_80),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_141),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_101),
.Y(n_142)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_84),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_106),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_108),
.A2(n_73),
.B1(n_88),
.B2(n_80),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_145),
.A2(n_114),
.B1(n_72),
.B2(n_106),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_67),
.B1(n_88),
.B2(n_73),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_77),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_147),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_95),
.B(n_73),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_108),
.A2(n_86),
.B1(n_60),
.B2(n_57),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_115),
.A2(n_82),
.B(n_49),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_152),
.B(n_153),
.Y(n_198)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_102),
.B(n_109),
.C(n_113),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_162),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_156),
.A2(n_161),
.B1(n_165),
.B2(n_76),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_127),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_168),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_159),
.B(n_0),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_133),
.A2(n_114),
.B1(n_119),
.B2(n_100),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_149),
.A2(n_146),
.B1(n_134),
.B2(n_123),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_123),
.C(n_136),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_167),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_202)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_122),
.Y(n_168)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_144),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_173),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_124),
.B(n_106),
.Y(n_173)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_174),
.Y(n_194)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_145),
.A2(n_134),
.B1(n_143),
.B2(n_148),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_176),
.A2(n_178),
.B1(n_179),
.B2(n_125),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_106),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_142),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_130),
.A2(n_98),
.B1(n_118),
.B2(n_111),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_148),
.A2(n_112),
.B1(n_96),
.B2(n_97),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_197),
.C(n_200),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_183),
.A2(n_156),
.B1(n_161),
.B2(n_158),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_180),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_187),
.Y(n_220)
);

A2O1A1O1Ixp25_ASAP7_75t_L g186 ( 
.A1(n_164),
.A2(n_150),
.B(n_137),
.C(n_138),
.D(n_129),
.Y(n_186)
);

XNOR2x1_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_189),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_170),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_164),
.A2(n_0),
.B(n_1),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_171),
.B(n_160),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_170),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_195),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_193),
.B(n_204),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_157),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_206),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_142),
.C(n_135),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_199),
.A2(n_167),
.B1(n_155),
.B2(n_162),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_177),
.C(n_159),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_111),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_203),
.C(n_175),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_202),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_165),
.B(n_8),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_176),
.A2(n_8),
.B1(n_15),
.B2(n_13),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_160),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_205),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_223),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_212),
.A2(n_214),
.B(n_216),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_193),
.A2(n_206),
.B(n_181),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_198),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_172),
.Y(n_217)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_217),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_218),
.A2(n_228),
.B1(n_229),
.B2(n_207),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_221),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_226),
.C(n_200),
.Y(n_238)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_224),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_194),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_225),
.B(n_230),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_182),
.B(n_152),
.C(n_163),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_163),
.Y(n_227)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_199),
.A2(n_151),
.B1(n_153),
.B2(n_154),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_183),
.A2(n_171),
.B1(n_151),
.B2(n_154),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_197),
.Y(n_230)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_233),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_231),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_234),
.A2(n_220),
.B(n_210),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_224),
.A2(n_188),
.B(n_191),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_237),
.A2(n_215),
.B1(n_211),
.B2(n_227),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_249),
.C(n_213),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_239),
.B(n_231),
.Y(n_251)
);

AOI21xp33_ASAP7_75t_L g240 ( 
.A1(n_208),
.A2(n_186),
.B(n_203),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_240),
.A2(n_243),
.B1(n_246),
.B2(n_229),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_208),
.A2(n_191),
.B1(n_189),
.B2(n_201),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_168),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_245),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_194),
.Y(n_245)
);

OAI31xp33_ASAP7_75t_L g246 ( 
.A1(n_214),
.A2(n_213),
.A3(n_217),
.B(n_221),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_174),
.C(n_2),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_251),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_253),
.C(n_260),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_226),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_254),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_255),
.A2(n_247),
.B1(n_242),
.B2(n_243),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_256),
.A2(n_262),
.B(n_236),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_235),
.A2(n_211),
.B1(n_223),
.B2(n_215),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_257),
.A2(n_259),
.B1(n_242),
.B2(n_174),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_241),
.A2(n_209),
.B1(n_216),
.B2(n_218),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_222),
.C(n_228),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_232),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_263),
.C(n_8),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_234),
.B(n_220),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_236),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_264),
.A2(n_271),
.B1(n_275),
.B2(n_274),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_246),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_266),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_248),
.Y(n_266)
);

OAI21x1_ASAP7_75t_SL g267 ( 
.A1(n_263),
.A2(n_237),
.B(n_247),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_275),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_268),
.B(n_269),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_249),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_212),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_252),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_273),
.A2(n_258),
.B1(n_259),
.B2(n_257),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_279),
.Y(n_289)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_278),
.Y(n_287)
);

MAJx2_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_253),
.C(n_9),
.Y(n_279)
);

AOI322xp5_ASAP7_75t_L g288 ( 
.A1(n_280),
.A2(n_6),
.A3(n_13),
.B1(n_12),
.B2(n_11),
.C1(n_10),
.C2(n_16),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_7),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_283),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_270),
.A2(n_266),
.B(n_272),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_270),
.A2(n_7),
.B(n_13),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_285),
.B(n_276),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_292),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_281),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_291),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_6),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_286),
.A2(n_276),
.B(n_279),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_296),
.C(n_297),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_286),
.A2(n_284),
.B(n_10),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_1),
.Y(n_297)
);

OAI311xp33_ASAP7_75t_L g299 ( 
.A1(n_293),
.A2(n_289),
.A3(n_2),
.B1(n_3),
.C1(n_4),
.Y(n_299)
);

NAND2xp33_ASAP7_75t_SL g300 ( 
.A(n_299),
.B(n_1),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_300),
.A2(n_294),
.B1(n_298),
.B2(n_4),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_301),
.A2(n_289),
.B(n_3),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_302),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_303)
);


endmodule