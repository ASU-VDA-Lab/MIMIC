module real_aes_12561_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_905;
wire n_503;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_792;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_453;
wire n_374;
wire n_647;
wire n_235;
wire n_932;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_298;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_363;
wire n_182;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_898;
wire n_115;
wire n_604;
wire n_110;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_914;
wire n_203;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_899;
wire n_637;
wire n_526;
wire n_155;
wire n_653;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_922;
wire n_520;
wire n_482;
wire n_633;
wire n_679;
wire n_926;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_516;
wire n_177;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_888;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_911;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
wire n_862;
INVx2_ASAP7_75t_SL g197 ( .A(n_0), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_1), .Y(n_331) );
OA21x2_ASAP7_75t_L g144 ( .A1(n_2), .A2(n_48), .B(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g205 ( .A(n_2), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g304 ( .A(n_3), .B(n_194), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_4), .B(n_236), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g910 ( .A1(n_5), .A2(n_65), .B1(n_911), .B2(n_912), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_5), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_6), .B(n_214), .Y(n_641) );
NAND2xp33_ASAP7_75t_L g658 ( .A(n_7), .B(n_659), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_8), .A2(n_104), .B1(n_924), .B2(n_934), .Y(n_103) );
AND2x2_ASAP7_75t_L g265 ( .A(n_9), .B(n_142), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_10), .B(n_154), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_11), .B(n_120), .Y(n_119) );
NAND3xp33_ASAP7_75t_L g923 ( .A(n_11), .B(n_121), .C(n_129), .Y(n_923) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_12), .B(n_234), .Y(n_601) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_13), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_14), .B(n_276), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g625 ( .A(n_15), .Y(n_625) );
BUFx3_ASAP7_75t_L g152 ( .A(n_16), .Y(n_152) );
INVx1_ASAP7_75t_L g157 ( .A(n_16), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_17), .B(n_141), .Y(n_307) );
A2O1A1Ixp33_ASAP7_75t_L g612 ( .A1(n_18), .A2(n_158), .B(n_216), .C(n_613), .Y(n_612) );
BUFx10_ASAP7_75t_L g127 ( .A(n_19), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_20), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_21), .B(n_154), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_22), .B(n_150), .Y(n_652) );
A2O1A1Ixp33_ASAP7_75t_L g617 ( .A1(n_23), .A2(n_287), .B(n_618), .C(n_620), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_24), .B(n_259), .Y(n_684) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_25), .Y(n_289) );
NAND3xp33_ASAP7_75t_L g241 ( .A(n_26), .B(n_239), .C(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g589 ( .A(n_27), .B(n_170), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_28), .B(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_29), .B(n_141), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_30), .A2(n_75), .B1(n_302), .B2(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g175 ( .A(n_31), .Y(n_175) );
INVx1_ASAP7_75t_L g644 ( .A(n_32), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_33), .B(n_186), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_34), .B(n_302), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_35), .B(n_141), .Y(n_660) );
INVx1_ASAP7_75t_L g116 ( .A(n_36), .Y(n_116) );
AND3x2_ASAP7_75t_L g922 ( .A(n_36), .B(n_124), .C(n_125), .Y(n_922) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_37), .B(n_222), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_38), .B(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g334 ( .A(n_39), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_40), .B(n_141), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_41), .B(n_194), .Y(n_595) );
CKINVDCx5p33_ASAP7_75t_R g614 ( .A(n_42), .Y(n_614) );
AND2x4_ASAP7_75t_L g174 ( .A(n_43), .B(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_44), .B(n_141), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_45), .B(n_170), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_46), .B(n_141), .Y(n_140) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_47), .A2(n_87), .B1(n_234), .B2(n_302), .Y(n_629) );
INVx1_ASAP7_75t_L g204 ( .A(n_48), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_49), .Y(n_260) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_50), .A2(n_193), .B(n_195), .C(n_198), .Y(n_192) );
INVx1_ASAP7_75t_L g145 ( .A(n_51), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_52), .B(n_141), .Y(n_337) );
AND2x4_ASAP7_75t_L g932 ( .A(n_53), .B(n_933), .Y(n_932) );
INVx3_ASAP7_75t_L g286 ( .A(n_54), .Y(n_286) );
OAI21xp5_ASAP7_75t_L g904 ( .A1(n_55), .A2(n_905), .B(n_913), .Y(n_904) );
INVx1_ASAP7_75t_L g915 ( .A(n_55), .Y(n_915) );
NOR2xp67_ASAP7_75t_L g117 ( .A(n_56), .B(n_76), .Y(n_117) );
AND2x2_ASAP7_75t_L g689 ( .A(n_57), .B(n_142), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g897 ( .A1(n_58), .A2(n_74), .B1(n_898), .B2(n_899), .Y(n_897) );
INVx1_ASAP7_75t_L g899 ( .A(n_58), .Y(n_899) );
INVx1_ASAP7_75t_L g933 ( .A(n_59), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_60), .B(n_259), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_61), .B(n_149), .Y(n_165) );
NAND2x1_ASAP7_75t_L g582 ( .A(n_62), .B(n_216), .Y(n_582) );
INVx1_ASAP7_75t_L g300 ( .A(n_63), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_64), .B(n_657), .Y(n_656) );
CKINVDCx5p33_ASAP7_75t_R g912 ( .A(n_65), .Y(n_912) );
NAND2xp5_ASAP7_75t_SL g603 ( .A(n_66), .B(n_219), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_67), .B(n_306), .Y(n_638) );
INVx2_ASAP7_75t_L g114 ( .A(n_68), .Y(n_114) );
AND3x2_ASAP7_75t_L g928 ( .A(n_68), .B(n_124), .C(n_929), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_69), .B(n_234), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_70), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g328 ( .A(n_71), .B(n_242), .Y(n_328) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_72), .B(n_242), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_73), .B(n_202), .Y(n_621) );
CKINVDCx5p33_ASAP7_75t_R g898 ( .A(n_74), .Y(n_898) );
NAND2xp5_ASAP7_75t_SL g688 ( .A(n_77), .B(n_222), .Y(n_688) );
CKINVDCx5p33_ASAP7_75t_R g580 ( .A(n_78), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_79), .B(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_80), .B(n_154), .Y(n_578) );
NAND2xp33_ASAP7_75t_SL g640 ( .A(n_81), .B(n_155), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_82), .B(n_335), .Y(n_637) );
INVx1_ASAP7_75t_L g184 ( .A(n_83), .Y(n_184) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_84), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_85), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_86), .B(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g160 ( .A(n_88), .Y(n_160) );
INVx1_ASAP7_75t_L g200 ( .A(n_88), .Y(n_200) );
BUFx3_ASAP7_75t_L g276 ( .A(n_88), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g619 ( .A(n_89), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_90), .B(n_196), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_91), .B(n_234), .Y(n_329) );
INVx1_ASAP7_75t_L g284 ( .A(n_92), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_93), .B(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_94), .B(n_142), .Y(n_226) );
NAND2xp33_ASAP7_75t_L g653 ( .A(n_95), .B(n_164), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_96), .B(n_163), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_97), .Y(n_279) );
INVx1_ASAP7_75t_L g274 ( .A(n_98), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_99), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g918 ( .A(n_100), .Y(n_918) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_101), .B(n_335), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_102), .B(n_149), .Y(n_148) );
OR2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_900), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_118), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g913 ( .A1(n_107), .A2(n_914), .B(n_916), .Y(n_913) );
NOR2xp67_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
CKINVDCx8_ASAP7_75t_R g907 ( .A(n_109), .Y(n_907) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx3_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
NOR2x1p5_ASAP7_75t_L g112 ( .A(n_113), .B(n_115), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
BUFx2_ASAP7_75t_L g125 ( .A(n_114), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
BUFx2_ASAP7_75t_L g566 ( .A(n_116), .Y(n_566) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_117), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_128), .Y(n_118) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OR2x6_ASAP7_75t_L g122 ( .A(n_123), .B(n_126), .Y(n_122) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
INVx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx6f_ASAP7_75t_L g903 ( .A(n_127), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_127), .B(n_922), .Y(n_921) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
XNOR2x1_ASAP7_75t_L g129 ( .A(n_130), .B(n_897), .Y(n_129) );
OAI22x1_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_563), .B1(n_567), .B2(n_896), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_500), .Y(n_131) );
NOR3xp33_ASAP7_75t_L g132 ( .A(n_133), .B(n_393), .C(n_471), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g133 ( .A(n_134), .B(n_354), .Y(n_133) );
AOI21xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_246), .B(n_308), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_176), .Y(n_136) );
AND2x2_ASAP7_75t_L g310 ( .A(n_137), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g423 ( .A(n_137), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g444 ( .A(n_137), .B(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g512 ( .A(n_137), .B(n_363), .Y(n_512) );
OR2x2_ASAP7_75t_L g515 ( .A(n_137), .B(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OR2x2_ASAP7_75t_L g352 ( .A(n_138), .B(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g375 ( .A(n_138), .Y(n_375) );
AND2x2_ASAP7_75t_L g407 ( .A(n_138), .B(n_378), .Y(n_407) );
BUFx2_ASAP7_75t_L g416 ( .A(n_138), .Y(n_416) );
INVx1_ASAP7_75t_L g449 ( .A(n_138), .Y(n_449) );
AND2x4_ASAP7_75t_L g468 ( .A(n_138), .B(n_426), .Y(n_468) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NAND2x1_ASAP7_75t_L g139 ( .A(n_140), .B(n_146), .Y(n_139) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_141), .Y(n_230) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_144), .Y(n_170) );
BUFx2_ASAP7_75t_L g293 ( .A(n_144), .Y(n_293) );
INVxp33_ASAP7_75t_L g645 ( .A(n_144), .Y(n_645) );
INVx1_ASAP7_75t_L g206 ( .A(n_145), .Y(n_206) );
OAI21x1_ASAP7_75t_SL g146 ( .A1(n_147), .A2(n_161), .B(n_168), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_153), .B(n_158), .Y(n_147) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_149), .A2(n_283), .B1(n_285), .B2(n_287), .Y(n_282) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_150), .B(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g196 ( .A(n_151), .Y(n_196) );
INVx1_ASAP7_75t_L g306 ( .A(n_151), .Y(n_306) );
INVx2_ASAP7_75t_L g632 ( .A(n_151), .Y(n_632) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_152), .Y(n_183) );
INVx2_ASAP7_75t_L g243 ( .A(n_152), .Y(n_243) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g164 ( .A(n_156), .Y(n_164) );
INVx2_ASAP7_75t_L g194 ( .A(n_156), .Y(n_194) );
INVx2_ASAP7_75t_L g335 ( .A(n_156), .Y(n_335) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g188 ( .A(n_157), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_158), .Y(n_189) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g281 ( .A(n_159), .Y(n_281) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
BUFx3_ASAP7_75t_L g167 ( .A(n_160), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_165), .B(n_166), .Y(n_161) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g682 ( .A1(n_166), .A2(n_683), .B(n_684), .Y(n_682) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_167), .A2(n_213), .B(n_215), .Y(n_212) );
O2A1O1Ixp5_ASAP7_75t_L g579 ( .A1(n_167), .A2(n_580), .B(n_581), .C(n_582), .Y(n_579) );
NAND3xp33_ASAP7_75t_L g630 ( .A(n_167), .B(n_264), .C(n_269), .Y(n_630) );
NOR2x1_ASAP7_75t_SL g168 ( .A(n_169), .B(n_171), .Y(n_168) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_169), .Y(n_210) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g380 ( .A(n_170), .Y(n_380) );
INVxp67_ASAP7_75t_SL g588 ( .A(n_170), .Y(n_588) );
NOR2xp67_ASAP7_75t_SL g680 ( .A(n_170), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_172), .B(n_203), .Y(n_615) );
INVx2_ASAP7_75t_SL g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g244 ( .A(n_173), .Y(n_244) );
INVx1_ASAP7_75t_L g583 ( .A(n_173), .Y(n_583) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g207 ( .A(n_174), .Y(n_207) );
BUFx6f_ASAP7_75t_SL g225 ( .A(n_174), .Y(n_225) );
INVx3_ASAP7_75t_L g277 ( .A(n_174), .Y(n_277) );
INVx1_ASAP7_75t_L g681 ( .A(n_174), .Y(n_681) );
INVx2_ASAP7_75t_L g392 ( .A(n_176), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_176), .A2(n_536), .B1(n_551), .B2(n_552), .Y(n_550) );
AND2x2_ASAP7_75t_L g176 ( .A(n_177), .B(n_208), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_L g311 ( .A(n_178), .B(n_312), .Y(n_311) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_178), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_178), .B(n_426), .Y(n_425) );
AND2x4_ASAP7_75t_L g432 ( .A(n_178), .B(n_209), .Y(n_432) );
AND2x2_ASAP7_75t_L g445 ( .A(n_178), .B(n_378), .Y(n_445) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g364 ( .A(n_179), .Y(n_364) );
OAI21x1_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_190), .B(n_201), .Y(n_179) );
AOI21x1_ASAP7_75t_SL g180 ( .A1(n_181), .A2(n_185), .B(n_189), .Y(n_180) );
OR2x2_ASAP7_75t_L g181 ( .A(n_182), .B(n_184), .Y(n_181) );
INVx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g214 ( .A(n_183), .Y(n_214) );
INVx2_ASAP7_75t_L g234 ( .A(n_183), .Y(n_234) );
INVx3_ASAP7_75t_L g253 ( .A(n_183), .Y(n_253) );
INVx2_ASAP7_75t_L g259 ( .A(n_183), .Y(n_259) );
INVx2_ASAP7_75t_L g333 ( .A(n_183), .Y(n_333) );
INVx2_ASAP7_75t_L g657 ( .A(n_183), .Y(n_657) );
HB1xp67_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g216 ( .A(n_187), .Y(n_216) );
INVx2_ASAP7_75t_L g219 ( .A(n_187), .Y(n_219) );
INVx2_ASAP7_75t_L g236 ( .A(n_187), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_187), .B(n_619), .Y(n_618) );
INVx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_188), .Y(n_222) );
AOI22x1_ASAP7_75t_L g250 ( .A1(n_189), .A2(n_199), .B1(n_251), .B2(n_257), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_191), .B(n_192), .Y(n_190) );
OAI21xp33_ASAP7_75t_L g201 ( .A1(n_191), .A2(n_202), .B(n_207), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_193), .A2(n_258), .B1(n_260), .B2(n_261), .Y(n_257) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AOI21x1_ASAP7_75t_L g232 ( .A1(n_199), .A2(n_233), .B(n_235), .Y(n_232) );
BUFx3_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g224 ( .A(n_200), .Y(n_224) );
INVxp67_ASAP7_75t_L g262 ( .A(n_202), .Y(n_262) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_203), .B(n_625), .Y(n_624) );
AO21x2_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_206), .Y(n_203) );
AOI21x1_ASAP7_75t_L g270 ( .A1(n_204), .A2(n_205), .B(n_206), .Y(n_270) );
INVx1_ASAP7_75t_L g264 ( .A(n_207), .Y(n_264) );
AND2x2_ASAP7_75t_L g399 ( .A(n_208), .B(n_400), .Y(n_399) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_208), .Y(n_443) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_227), .Y(n_208) );
AND2x4_ASAP7_75t_L g462 ( .A(n_209), .B(n_415), .Y(n_462) );
AND2x4_ASAP7_75t_L g475 ( .A(n_209), .B(n_468), .Y(n_475) );
OR2x2_ASAP7_75t_L g505 ( .A(n_209), .B(n_377), .Y(n_505) );
OAI21x1_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_226), .Y(n_209) );
OAI21x1_ASAP7_75t_L g313 ( .A1(n_210), .A2(n_211), .B(n_226), .Y(n_313) );
OAI21x1_ASAP7_75t_L g341 ( .A1(n_210), .A2(n_250), .B(n_342), .Y(n_341) );
OAI21x1_ASAP7_75t_L g574 ( .A1(n_210), .A2(n_575), .B(n_584), .Y(n_574) );
OAI21xp5_ASAP7_75t_L g597 ( .A1(n_210), .A2(n_598), .B(n_605), .Y(n_597) );
OAI21x1_ASAP7_75t_L g709 ( .A1(n_210), .A2(n_598), .B(n_605), .Y(n_709) );
OAI21x1_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_217), .B(n_225), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_220), .B(n_223), .Y(n_217) );
INVx2_ASAP7_75t_L g255 ( .A(n_219), .Y(n_255) );
INVxp67_ASAP7_75t_L g240 ( .A(n_221), .Y(n_240) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_222), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g287 ( .A(n_222), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_222), .B(n_614), .Y(n_613) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_223), .A2(n_304), .B(n_305), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_223), .A2(n_328), .B(n_329), .Y(n_327) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_223), .A2(n_577), .B(n_578), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g594 ( .A1(n_223), .A2(n_595), .B(n_596), .Y(n_594) );
AOI21xp5_ASAP7_75t_L g602 ( .A1(n_223), .A2(n_603), .B(n_604), .Y(n_602) );
AO21x1_ASAP7_75t_L g636 ( .A1(n_223), .A2(n_637), .B(n_638), .Y(n_636) );
BUFx10_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g239 ( .A(n_224), .Y(n_239) );
OAI21x1_ASAP7_75t_L g294 ( .A1(n_225), .A2(n_295), .B(n_303), .Y(n_294) );
AOI21xp5_ASAP7_75t_L g587 ( .A1(n_225), .A2(n_588), .B(n_589), .Y(n_587) );
OAI21x1_ASAP7_75t_L g598 ( .A1(n_225), .A2(n_599), .B(n_602), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g646 ( .A1(n_225), .A2(n_643), .B(n_647), .Y(n_646) );
OAI21x1_ASAP7_75t_L g650 ( .A1(n_225), .A2(n_651), .B(n_655), .Y(n_650) );
OR2x6_ASAP7_75t_L g363 ( .A(n_227), .B(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVxp67_ASAP7_75t_SL g353 ( .A(n_228), .Y(n_353) );
INVx2_ASAP7_75t_L g426 ( .A(n_228), .Y(n_426) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
OAI21x1_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_245), .Y(n_229) );
OA21x2_ASAP7_75t_L g378 ( .A1(n_231), .A2(n_245), .B(n_379), .Y(n_378) );
OAI21x1_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_237), .B(n_244), .Y(n_231) );
OAI21xp5_ASAP7_75t_L g591 ( .A1(n_236), .A2(n_592), .B(n_593), .Y(n_591) );
OAI21xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_240), .B(n_241), .Y(n_237) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g302 ( .A(n_243), .Y(n_302) );
INVx2_ASAP7_75t_L g659 ( .A(n_243), .Y(n_659) );
OAI21xp5_ASAP7_75t_L g326 ( .A1(n_244), .A2(n_327), .B(n_330), .Y(n_326) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_266), .Y(n_246) );
OR2x2_ASAP7_75t_L g391 ( .A(n_247), .B(n_360), .Y(n_391) );
INVx1_ASAP7_75t_L g491 ( .A(n_247), .Y(n_491) );
OR2x2_ASAP7_75t_L g547 ( .A(n_247), .B(n_344), .Y(n_547) );
BUFx3_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g435 ( .A(n_248), .Y(n_435) );
AO31x2_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_262), .A3(n_263), .B(n_265), .Y(n_248) );
AO31x2_ASAP7_75t_L g318 ( .A1(n_249), .A2(n_262), .A3(n_263), .B(n_265), .Y(n_318) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
OAI22x1_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_254), .B1(n_255), .B2(n_256), .Y(n_251) );
INVxp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVxp67_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVxp67_ASAP7_75t_L g296 ( .A(n_259), .Y(n_296) );
BUFx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND3xp33_ASAP7_75t_L g627 ( .A(n_264), .B(n_269), .C(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g342 ( .A(n_265), .Y(n_342) );
AND2x2_ASAP7_75t_L g463 ( .A(n_266), .B(n_358), .Y(n_463) );
AND2x2_ASAP7_75t_L g477 ( .A(n_266), .B(n_435), .Y(n_477) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_266), .Y(n_497) );
AND2x2_ASAP7_75t_L g557 ( .A(n_266), .B(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_290), .Y(n_266) );
INVx3_ASAP7_75t_L g346 ( .A(n_267), .Y(n_346) );
AO21x2_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_271), .B(n_288), .Y(n_267) );
AO21x1_ASAP7_75t_L g323 ( .A1(n_268), .A2(n_271), .B(n_288), .Y(n_323) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NOR2xp33_ASAP7_75t_SL g288 ( .A(n_269), .B(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_282), .Y(n_271) );
AOI22xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_275), .B1(n_278), .B2(n_280), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
NOR3xp33_ASAP7_75t_L g283 ( .A(n_276), .B(n_277), .C(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g301 ( .A(n_276), .Y(n_301) );
INVx2_ASAP7_75t_L g336 ( .A(n_276), .Y(n_336) );
AOI211x1_ASAP7_75t_L g590 ( .A1(n_276), .A2(n_589), .B(n_591), .C(n_594), .Y(n_590) );
INVx1_ASAP7_75t_L g654 ( .A(n_276), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_277), .B(n_281), .Y(n_280) );
NOR3xp33_ASAP7_75t_L g285 ( .A(n_277), .B(n_281), .C(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g628 ( .A(n_281), .Y(n_628) );
INVx3_ASAP7_75t_L g319 ( .A(n_290), .Y(n_319) );
AND2x2_ASAP7_75t_L g340 ( .A(n_290), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g361 ( .A(n_290), .Y(n_361) );
INVx2_ASAP7_75t_L g387 ( .A(n_290), .Y(n_387) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_290), .Y(n_398) );
AND2x2_ASAP7_75t_L g404 ( .A(n_290), .B(n_346), .Y(n_404) );
INVx1_ASAP7_75t_L g516 ( .A(n_290), .Y(n_516) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OAI21x1_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_294), .B(n_307), .Y(n_291) );
OAI21x1_ASAP7_75t_L g325 ( .A1(n_292), .A2(n_326), .B(n_337), .Y(n_325) );
OAI21x1_ASAP7_75t_L g649 ( .A1(n_292), .A2(n_650), .B(n_660), .Y(n_649) );
BUFx3_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g647 ( .A(n_293), .Y(n_647) );
OAI21xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_297), .B(n_298), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_302), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx1_ASAP7_75t_L g620 ( .A(n_301), .Y(n_620) );
INVx2_ASAP7_75t_L g581 ( .A(n_306), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_314), .B1(n_338), .B2(n_347), .Y(n_308) );
NAND2xp33_ASAP7_75t_L g456 ( .A(n_309), .B(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g383 ( .A(n_311), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_311), .B(n_468), .Y(n_545) );
BUFx3_ASAP7_75t_L g350 ( .A(n_312), .Y(n_350) );
AND2x2_ASAP7_75t_L g374 ( .A(n_312), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g499 ( .A(n_312), .Y(n_499) );
AND2x4_ASAP7_75t_L g539 ( .A(n_312), .B(n_415), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_312), .B(n_535), .Y(n_542) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_313), .Y(n_420) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AOI22xp33_ASAP7_75t_SL g560 ( .A1(n_315), .A2(n_450), .B1(n_466), .B2(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_320), .Y(n_315) );
INVx2_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g417 ( .A(n_317), .B(n_344), .Y(n_417) );
OR2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx1_ASAP7_75t_L g369 ( .A(n_318), .Y(n_369) );
OR2x2_ASAP7_75t_L g554 ( .A(n_318), .B(n_345), .Y(n_554) );
INVx2_ASAP7_75t_L g371 ( .A(n_319), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_319), .B(n_455), .Y(n_470) );
AND2x2_ASAP7_75t_L g522 ( .A(n_320), .B(n_523), .Y(n_522) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g411 ( .A(n_321), .Y(n_411) );
INVx1_ASAP7_75t_L g495 ( .A(n_321), .Y(n_495) );
AND2x2_ASAP7_75t_L g536 ( .A(n_321), .B(n_435), .Y(n_536) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g386 ( .A(n_323), .B(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_323), .B(n_453), .Y(n_452) );
INVx3_ASAP7_75t_L g345 ( .A(n_324), .Y(n_345) );
INVx1_ASAP7_75t_L g368 ( .A(n_324), .Y(n_368) );
INVx2_ASAP7_75t_L g455 ( .A(n_324), .Y(n_455) );
AND2x2_ASAP7_75t_L g558 ( .A(n_324), .B(n_341), .Y(n_558) );
INVx3_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
O2A1O1Ixp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_332), .B(n_334), .C(n_336), .Y(n_330) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AOI21xp5_ASAP7_75t_L g599 ( .A1(n_336), .A2(n_600), .B(n_601), .Y(n_599) );
AO21x1_ASAP7_75t_L g639 ( .A1(n_336), .A2(n_640), .B(n_641), .Y(n_639) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_340), .B(n_343), .Y(n_339) );
INVx1_ASAP7_75t_L g410 ( .A(n_340), .Y(n_410) );
AND2x4_ASAP7_75t_L g358 ( .A(n_341), .B(n_345), .Y(n_358) );
INVx1_ASAP7_75t_L g453 ( .A(n_341), .Y(n_453) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_346), .B(n_361), .Y(n_360) );
NOR2x1_ASAP7_75t_L g519 ( .A(n_346), .B(n_455), .Y(n_519) );
BUFx2_ASAP7_75t_L g553 ( .A(n_346), .Y(n_553) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_351), .Y(n_348) );
OR2x2_ASAP7_75t_L g405 ( .A(n_349), .B(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g362 ( .A(n_350), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_350), .B(n_421), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_350), .B(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_350), .B(n_445), .Y(n_521) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g382 ( .A(n_352), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g466 ( .A(n_352), .Y(n_466) );
OR2x2_ASAP7_75t_L g559 ( .A(n_352), .B(n_446), .Y(n_559) );
AND2x2_ASAP7_75t_L g421 ( .A(n_353), .B(n_375), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_355), .B(n_381), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_362), .B1(n_365), .B2(n_372), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_358), .B(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g440 ( .A(n_358), .Y(n_440) );
AOI322xp5_ASAP7_75t_L g513 ( .A1(n_358), .A2(n_376), .A3(n_514), .B1(n_517), .B2(n_520), .C1(n_522), .C2(n_524), .Y(n_513) );
INVxp67_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_SL g509 ( .A(n_362), .Y(n_509) );
OR2x2_ASAP7_75t_L g457 ( .A(n_363), .B(n_416), .Y(n_457) );
OR2x2_ASAP7_75t_SL g377 ( .A(n_364), .B(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g415 ( .A(n_364), .Y(n_415) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_370), .Y(n_366) );
AND2x2_ASAP7_75t_L g527 ( .A(n_367), .B(n_516), .Y(n_527) );
AND2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx1_ASAP7_75t_L g390 ( .A(n_368), .Y(n_390) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_368), .Y(n_403) );
INVx1_ASAP7_75t_L g492 ( .A(n_370), .Y(n_492) );
BUFx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NOR2xp67_ASAP7_75t_L g454 ( .A(n_371), .B(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g532 ( .A(n_371), .B(n_411), .Y(n_532) );
INVxp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_376), .Y(n_373) );
INVx1_ASAP7_75t_L g431 ( .A(n_375), .Y(n_431) );
BUFx2_ASAP7_75t_L g489 ( .A(n_375), .Y(n_489) );
INVx2_ASAP7_75t_SL g408 ( .A(n_376), .Y(n_408) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g447 ( .A(n_377), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
OAI32xp33_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_384), .A3(n_388), .B1(n_391), .B2(n_392), .Y(n_381) );
AND2x2_ASAP7_75t_L g427 ( .A(n_384), .B(n_389), .Y(n_427) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g439 ( .A(n_386), .Y(n_439) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_390), .B(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g479 ( .A(n_391), .Y(n_479) );
NAND4xp25_ASAP7_75t_L g393 ( .A(n_394), .B(n_418), .C(n_436), .D(n_458), .Y(n_393) );
AOI211x1_ASAP7_75t_SL g394 ( .A1(n_395), .A2(n_399), .B(n_401), .C(n_412), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g482 ( .A(n_397), .B(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_397), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_399), .B(n_489), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_405), .B1(n_408), .B2(n_409), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_404), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g506 ( .A(n_404), .Y(n_506) );
OR2x2_ASAP7_75t_L g460 ( .A(n_406), .B(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g538 ( .A(n_407), .B(n_539), .Y(n_538) );
AOI21xp33_ASAP7_75t_SL g412 ( .A1(n_408), .A2(n_413), .B(n_417), .Y(n_412) );
OR2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_414), .B(n_416), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_415), .Y(n_465) );
O2A1O1Ixp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_422), .B(n_427), .C(n_428), .Y(n_418) );
AOI32xp33_ASAP7_75t_L g525 ( .A1(n_419), .A2(n_459), .A3(n_506), .B1(n_526), .B2(n_527), .Y(n_525) );
AND2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
INVx1_ASAP7_75t_L g461 ( .A(n_420), .Y(n_461) );
AND2x4_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g498 ( .A(n_425), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g535 ( .A(n_426), .Y(n_535) );
AOI21xp33_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_430), .B(n_433), .Y(n_428) );
INVx2_ASAP7_75t_SL g530 ( .A(n_429), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_431), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_431), .B(n_504), .Y(n_503) );
OR2x2_ASAP7_75t_L g541 ( .A(n_431), .B(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g446 ( .A(n_432), .Y(n_446) );
INVx1_ASAP7_75t_L g476 ( .A(n_432), .Y(n_476) );
AND2x2_ASAP7_75t_L g533 ( .A(n_432), .B(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OR2x6_ASAP7_75t_L g494 ( .A(n_435), .B(n_495), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_441), .B1(n_450), .B2(n_456), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_437), .A2(n_463), .B1(n_538), .B2(n_540), .Y(n_537) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
INVx1_ASAP7_75t_L g526 ( .A(n_440), .Y(n_526) );
NAND4xp25_ASAP7_75t_L g441 ( .A(n_442), .B(n_444), .C(n_446), .D(n_447), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g551 ( .A(n_445), .B(n_448), .Y(n_551) );
INVx1_ASAP7_75t_L g480 ( .A(n_447), .Y(n_480) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_454), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_451), .B(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g469 ( .A(n_452), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g484 ( .A(n_455), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_462), .B(n_463), .C(n_464), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g524 ( .A(n_462), .B(n_489), .Y(n_524) );
O2A1O1Ixp33_ASAP7_75t_SL g464 ( .A1(n_465), .A2(n_466), .B(n_467), .C(n_469), .Y(n_464) );
INVx1_ASAP7_75t_L g478 ( .A(n_466), .Y(n_478) );
INVx1_ASAP7_75t_L g508 ( .A(n_469), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_486), .Y(n_471) );
AOI322xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_477), .A3(n_478), .B1(n_479), .B2(n_480), .C1(n_481), .C2(n_485), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_476), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
AOI31xp33_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_490), .A3(n_492), .B(n_493), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_496), .B(n_498), .Y(n_493) );
INVx1_ASAP7_75t_L g510 ( .A(n_496), .Y(n_510) );
NOR2xp67_ASAP7_75t_L g500 ( .A(n_501), .B(n_528), .Y(n_500) );
NAND4xp25_ASAP7_75t_L g501 ( .A(n_502), .B(n_507), .C(n_513), .D(n_525), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_506), .Y(n_502) );
INVx3_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B1(n_510), .B2(n_511), .Y(n_507) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_SL g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g523 ( .A(n_516), .Y(n_523) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
NAND5xp2_ASAP7_75t_L g528 ( .A(n_529), .B(n_537), .C(n_543), .D(n_548), .E(n_560), .Y(n_528) );
AOI22xp33_ASAP7_75t_SL g529 ( .A1(n_530), .A2(n_531), .B1(n_533), .B2(n_536), .Y(n_529) );
INVx1_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OAI21xp5_ASAP7_75t_L g543 ( .A1(n_540), .A2(n_544), .B(n_546), .Y(n_543) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_542), .Y(n_562) );
INVxp67_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_549), .B(n_555), .Y(n_548) );
INVxp67_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
NOR2x1_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_556), .B(n_559), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVxp67_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
CKINVDCx10_ASAP7_75t_R g563 ( .A(n_564), .Y(n_563) );
BUFx6f_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
BUFx8_ASAP7_75t_L g896 ( .A(n_565), .Y(n_896) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x4_ASAP7_75t_L g929 ( .A(n_566), .B(n_930), .Y(n_929) );
XNOR2xp5_ASAP7_75t_L g908 ( .A(n_567), .B(n_909), .Y(n_908) );
AND2x4_ASAP7_75t_L g567 ( .A(n_568), .B(n_804), .Y(n_567) );
NOR3xp33_ASAP7_75t_L g568 ( .A(n_569), .B(n_736), .C(n_772), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_703), .Y(n_569) );
AOI221xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_606), .B1(n_661), .B2(n_672), .C(n_675), .Y(n_570) );
INVx1_ASAP7_75t_L g731 ( .A(n_571), .Y(n_731) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_585), .Y(n_571) );
AND2x2_ASAP7_75t_L g837 ( .A(n_572), .B(n_775), .Y(n_837) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_573), .B(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g782 ( .A(n_573), .B(n_725), .Y(n_782) );
AND2x2_ASAP7_75t_L g819 ( .A(n_573), .B(n_708), .Y(n_819) );
INVx1_ASAP7_75t_L g841 ( .A(n_573), .Y(n_841) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g700 ( .A(n_574), .Y(n_700) );
INVx1_ASAP7_75t_L g707 ( .A(n_574), .Y(n_707) );
OAI21xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_579), .B(n_583), .Y(n_575) );
NAND2x1_ASAP7_75t_L g888 ( .A(n_585), .B(n_797), .Y(n_888) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_597), .Y(n_585) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_586), .Y(n_674) );
BUFx2_ASAP7_75t_L g696 ( .A(n_586), .Y(n_696) );
INVx2_ASAP7_75t_L g712 ( .A(n_586), .Y(n_712) );
AND2x2_ASAP7_75t_L g756 ( .A(n_586), .B(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g776 ( .A(n_586), .Y(n_776) );
INVx2_ASAP7_75t_L g786 ( .A(n_586), .Y(n_786) );
INVx1_ASAP7_75t_L g834 ( .A(n_586), .Y(n_834) );
AND2x2_ASAP7_75t_L g851 ( .A(n_586), .B(n_711), .Y(n_851) );
OR2x6_ASAP7_75t_L g586 ( .A(n_587), .B(n_590), .Y(n_586) );
INVx1_ASAP7_75t_L g698 ( .A(n_597), .Y(n_698) );
AND2x2_ASAP7_75t_L g755 ( .A(n_597), .B(n_711), .Y(n_755) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OAI221xp5_ASAP7_75t_L g716 ( .A1(n_607), .A2(n_710), .B1(n_717), .B2(n_720), .C(n_723), .Y(n_716) );
OR2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_633), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g728 ( .A(n_609), .B(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_622), .Y(n_609) );
INVx2_ASAP7_75t_L g693 ( .A(n_610), .Y(n_693) );
OR2x2_ASAP7_75t_L g722 ( .A(n_610), .B(n_635), .Y(n_722) );
AND2x2_ASAP7_75t_L g813 ( .A(n_610), .B(n_623), .Y(n_813) );
AND2x2_ASAP7_75t_L g830 ( .A(n_610), .B(n_635), .Y(n_830) );
NAND2x1p5_ASAP7_75t_L g610 ( .A(n_611), .B(n_616), .Y(n_610) );
NAND2x1p5_ASAP7_75t_L g665 ( .A(n_611), .B(n_616), .Y(n_665) );
OR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_615), .Y(n_611) );
OA21x2_ASAP7_75t_L g616 ( .A1(n_615), .A2(n_617), .B(n_621), .Y(n_616) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_620), .A2(n_656), .B(n_658), .Y(n_655) );
INVx1_ASAP7_75t_L g739 ( .A(n_622), .Y(n_739) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g669 ( .A(n_623), .Y(n_669) );
AND2x2_ASAP7_75t_L g715 ( .A(n_623), .B(n_694), .Y(n_715) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_623), .Y(n_752) );
AND2x2_ASAP7_75t_L g759 ( .A(n_623), .B(n_649), .Y(n_759) );
INVx1_ASAP7_75t_L g803 ( .A(n_623), .Y(n_803) );
INVxp67_ASAP7_75t_L g895 ( .A(n_623), .Y(n_895) );
OR2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_629), .B1(n_630), .B2(n_631), .Y(n_626) );
OR2x2_ASAP7_75t_L g831 ( .A(n_633), .B(n_663), .Y(n_831) );
OR2x2_ASAP7_75t_L g881 ( .A(n_633), .B(n_751), .Y(n_881) );
INVx3_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g702 ( .A(n_634), .B(n_663), .Y(n_702) );
AND2x2_ASAP7_75t_L g802 ( .A(n_634), .B(n_803), .Y(n_802) );
AND2x2_ASAP7_75t_L g812 ( .A(n_634), .B(n_813), .Y(n_812) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_648), .Y(n_634) );
INVx2_ASAP7_75t_L g668 ( .A(n_635), .Y(n_668) );
AND2x2_ASAP7_75t_L g729 ( .A(n_635), .B(n_649), .Y(n_729) );
AND2x2_ASAP7_75t_L g740 ( .A(n_635), .B(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g771 ( .A(n_635), .Y(n_771) );
AO31x2_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_639), .A3(n_642), .B(n_646), .Y(n_635) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g671 ( .A(n_649), .Y(n_671) );
INVx1_ASAP7_75t_L g694 ( .A(n_649), .Y(n_694) );
AND2x2_ASAP7_75t_L g780 ( .A(n_649), .B(n_669), .Y(n_780) );
AND2x2_ASAP7_75t_L g795 ( .A(n_649), .B(n_693), .Y(n_795) );
AOI21xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B(n_654), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_654), .A2(n_687), .B(n_688), .Y(n_686) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NAND2x1p5_ASAP7_75t_L g662 ( .A(n_663), .B(n_666), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
HB1xp67_ASAP7_75t_L g768 ( .A(n_664), .Y(n_768) );
AND2x2_ASAP7_75t_L g779 ( .A(n_664), .B(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g714 ( .A(n_665), .B(n_668), .Y(n_714) );
INVx1_ASAP7_75t_L g741 ( .A(n_665), .Y(n_741) );
BUFx2_ASAP7_75t_L g753 ( .A(n_665), .Y(n_753) );
AND2x2_ASAP7_75t_L g761 ( .A(n_665), .B(n_712), .Y(n_761) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_665), .Y(n_844) );
AOI22xp5_ASAP7_75t_L g861 ( .A1(n_666), .A2(n_743), .B1(n_802), .B2(n_862), .Y(n_861) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_670), .Y(n_666) );
AND2x2_ASAP7_75t_L g691 ( .A(n_667), .B(n_692), .Y(n_691) );
AND2x4_ASAP7_75t_L g794 ( .A(n_667), .B(n_795), .Y(n_794) );
AND2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
INVx1_ASAP7_75t_L g791 ( .A(n_668), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_670), .B(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g811 ( .A(n_670), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g836 ( .A(n_670), .B(n_829), .Y(n_836) );
NOR2xp33_ASAP7_75t_L g854 ( .A(n_670), .B(n_722), .Y(n_854) );
BUFx3_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_671), .B(n_771), .Y(n_770) );
INVxp67_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_690), .B1(n_695), .B2(n_701), .Y(n_675) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g719 ( .A(n_677), .Y(n_719) );
OR2x2_ASAP7_75t_L g788 ( .A(n_677), .B(n_764), .Y(n_788) );
INVx2_ASAP7_75t_L g711 ( .A(n_678), .Y(n_711) );
OR2x2_ASAP7_75t_L g727 ( .A(n_678), .B(n_709), .Y(n_727) );
AND2x2_ASAP7_75t_L g735 ( .A(n_678), .B(n_708), .Y(n_735) );
AND2x4_ASAP7_75t_L g775 ( .A(n_678), .B(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g798 ( .A(n_678), .Y(n_798) );
AND2x4_ASAP7_75t_L g678 ( .A(n_679), .B(n_685), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_682), .Y(n_679) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_680), .A2(n_686), .B(n_689), .Y(n_685) );
AOI21xp33_ASAP7_75t_SL g730 ( .A1(n_690), .A2(n_731), .B(n_732), .Y(n_730) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
INVx1_ASAP7_75t_L g733 ( .A(n_696), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_696), .B(n_726), .Y(n_748) );
INVx1_ASAP7_75t_L g853 ( .A(n_696), .Y(n_853) );
INVx2_ASAP7_75t_L g877 ( .A(n_697), .Y(n_877) );
AND2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
INVx1_ASAP7_75t_L g718 ( .A(n_698), .Y(n_718) );
INVx2_ASAP7_75t_L g745 ( .A(n_699), .Y(n_745) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g757 ( .A(n_700), .Y(n_757) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AOI211xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_713), .B(n_716), .C(n_730), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
OR2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_710), .Y(n_705) );
INVx2_ASAP7_75t_L g799 ( .A(n_706), .Y(n_799) );
INVx1_ASAP7_75t_L g848 ( .A(n_706), .Y(n_848) );
INVx2_ASAP7_75t_SL g893 ( .A(n_706), .Y(n_893) );
OR2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
INVx1_ASAP7_75t_L g725 ( .A(n_708), .Y(n_725) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g809 ( .A(n_710), .Y(n_809) );
OR2x2_ASAP7_75t_L g866 ( .A(n_710), .B(n_745), .Y(n_866) );
NAND2xp33_ASAP7_75t_L g892 ( .A(n_710), .B(n_893), .Y(n_892) );
OR2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
AND2x4_ASAP7_75t_SL g785 ( .A(n_711), .B(n_786), .Y(n_785) );
AND2x2_ASAP7_75t_L g724 ( .A(n_712), .B(n_725), .Y(n_724) );
BUFx3_ASAP7_75t_L g764 ( .A(n_712), .Y(n_764) );
AND2x4_ASAP7_75t_SL g713 ( .A(n_714), .B(n_715), .Y(n_713) );
AND2x2_ASAP7_75t_L g824 ( .A(n_714), .B(n_825), .Y(n_824) );
AND2x2_ASAP7_75t_L g878 ( .A(n_714), .B(n_759), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_714), .B(n_895), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_718), .B(n_775), .Y(n_863) );
INVx1_ASAP7_75t_L g873 ( .A(n_718), .Y(n_873) );
INVx1_ASAP7_75t_L g810 ( .A(n_721), .Y(n_810) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OR2x2_ASAP7_75t_L g815 ( .A(n_722), .B(n_816), .Y(n_815) );
OAI21xp33_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_726), .B(n_728), .Y(n_723) );
AND2x4_ASAP7_75t_L g743 ( .A(n_726), .B(n_744), .Y(n_743) );
AOI322xp5_ASAP7_75t_L g806 ( .A1(n_726), .A2(n_807), .A3(n_810), .B1(n_811), .B2(n_812), .C1(n_814), .C2(n_817), .Y(n_806) );
NAND3xp33_ASAP7_75t_L g822 ( .A(n_726), .B(n_744), .C(n_823), .Y(n_822) );
INVx4_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OAI33xp33_ASAP7_75t_L g750 ( .A1(n_727), .A2(n_751), .A3(n_753), .B1(n_754), .B2(n_758), .B3(n_760), .Y(n_750) );
NOR2x1_ASAP7_75t_L g846 ( .A(n_727), .B(n_833), .Y(n_846) );
OR2x2_ASAP7_75t_L g860 ( .A(n_727), .B(n_841), .Y(n_860) );
AND2x2_ASAP7_75t_L g867 ( .A(n_729), .B(n_813), .Y(n_867) );
OR2x2_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .Y(n_732) );
OR2x2_ASAP7_75t_L g871 ( .A(n_734), .B(n_745), .Y(n_871) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g763 ( .A(n_735), .B(n_764), .Y(n_763) );
OAI211xp5_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_742), .B(n_746), .C(n_762), .Y(n_736) );
INVx1_ASAP7_75t_L g749 ( .A(n_737), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_740), .Y(n_737) );
OR2x2_ASAP7_75t_L g828 ( .A(n_738), .B(n_829), .Y(n_828) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_740), .B(n_759), .Y(n_869) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_745), .B(n_755), .Y(n_766) );
AND2x2_ASAP7_75t_L g793 ( .A(n_745), .B(n_785), .Y(n_793) );
OR2x2_ASAP7_75t_L g890 ( .A(n_745), .B(n_891), .Y(n_890) );
AOI21xp5_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_749), .B(n_750), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
NAND4xp25_ASAP7_75t_L g883 ( .A(n_748), .B(n_884), .C(n_887), .D(n_888), .Y(n_883) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g839 ( .A(n_753), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
AND2x2_ASAP7_75t_L g840 ( .A(n_755), .B(n_841), .Y(n_840) );
AND2x2_ASAP7_75t_L g852 ( .A(n_755), .B(n_853), .Y(n_852) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_757), .Y(n_777) );
OR2x2_ASAP7_75t_L g833 ( .A(n_757), .B(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g816 ( .A(n_759), .Y(n_816) );
AND2x2_ASAP7_75t_L g838 ( .A(n_759), .B(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
OAI21xp33_ASAP7_75t_SL g762 ( .A1(n_763), .A2(n_765), .B(n_767), .Y(n_762) );
INVx2_ASAP7_75t_L g823 ( .A(n_764), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_764), .B(n_848), .Y(n_847) );
HB1xp67_ASAP7_75t_L g858 ( .A(n_764), .Y(n_858) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
OAI32xp33_ASAP7_75t_L g879 ( .A1(n_766), .A2(n_816), .A3(n_830), .B1(n_880), .B2(n_881), .Y(n_879) );
NOR2x1p5_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
BUFx3_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
OAI211xp5_ASAP7_75t_SL g772 ( .A1(n_773), .A2(n_778), .B(n_781), .C(n_792), .Y(n_772) );
NAND3xp33_ASAP7_75t_SL g876 ( .A(n_773), .B(n_788), .C(n_877), .Y(n_876) );
INVx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
AND2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_777), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_775), .B(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_780), .B(n_791), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_780), .B(n_844), .Y(n_843) );
A2O1A1Ixp33_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_783), .B(n_787), .C(n_789), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_782), .B(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g891 ( .A(n_785), .Y(n_891) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
AOI22xp33_ASAP7_75t_SL g792 ( .A1(n_793), .A2(n_794), .B1(n_796), .B2(n_800), .Y(n_792) );
INVx2_ASAP7_75t_L g874 ( .A(n_794), .Y(n_874) );
AND2x4_ASAP7_75t_SL g796 ( .A(n_797), .B(n_799), .Y(n_796) );
OR2x2_ASAP7_75t_L g832 ( .A(n_797), .B(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g885 ( .A(n_797), .Y(n_885) );
INVx4_ASAP7_75t_R g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g887 ( .A(n_799), .Y(n_887) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx2_ASAP7_75t_L g825 ( .A(n_803), .Y(n_825) );
NOR2x1_ASAP7_75t_L g804 ( .A(n_805), .B(n_855), .Y(n_804) );
NAND3xp33_ASAP7_75t_L g805 ( .A(n_806), .B(n_820), .C(n_826), .Y(n_805) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
O2A1O1Ixp33_ASAP7_75t_L g872 ( .A1(n_809), .A2(n_871), .B(n_873), .C(n_874), .Y(n_872) );
AOI21xp5_ASAP7_75t_L g882 ( .A1(n_814), .A2(n_883), .B(n_889), .Y(n_882) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
NAND2xp5_ASAP7_75t_SL g820 ( .A(n_821), .B(n_824), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
NOR2xp33_ASAP7_75t_L g826 ( .A(n_827), .B(n_842), .Y(n_826) );
A2O1A1Ixp33_ASAP7_75t_L g827 ( .A1(n_828), .A2(n_831), .B(n_832), .C(n_835), .Y(n_827) );
OAI221xp5_ASAP7_75t_L g842 ( .A1(n_828), .A2(n_843), .B1(n_845), .B2(n_847), .C(n_849), .Y(n_842) );
OA21x2_ASAP7_75t_L g856 ( .A1(n_829), .A2(n_857), .B(n_861), .Y(n_856) );
INVx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_836), .A2(n_837), .B1(n_838), .B2(n_840), .Y(n_835) );
AND2x2_ASAP7_75t_L g850 ( .A(n_841), .B(n_851), .Y(n_850) );
HB1xp67_ASAP7_75t_L g886 ( .A(n_841), .Y(n_886) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
OAI21xp33_ASAP7_75t_L g849 ( .A1(n_850), .A2(n_852), .B(n_854), .Y(n_849) );
INVx1_ASAP7_75t_L g880 ( .A(n_850), .Y(n_880) );
NAND4xp75_ASAP7_75t_L g855 ( .A(n_856), .B(n_864), .C(n_875), .D(n_882), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_858), .B(n_859), .Y(n_857) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
AOI221xp5_ASAP7_75t_L g864 ( .A1(n_865), .A2(n_867), .B1(n_868), .B2(n_870), .C(n_872), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
AOI21xp5_ASAP7_75t_L g875 ( .A1(n_876), .A2(n_878), .B(n_879), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_885), .B(n_886), .Y(n_884) );
AOI21xp33_ASAP7_75t_L g889 ( .A1(n_890), .A2(n_892), .B(n_894), .Y(n_889) );
NAND2xp5_ASAP7_75t_SL g900 ( .A(n_901), .B(n_923), .Y(n_900) );
AOI21xp5_ASAP7_75t_L g901 ( .A1(n_902), .A2(n_904), .B(n_917), .Y(n_901) );
CKINVDCx11_ASAP7_75t_R g902 ( .A(n_903), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_906), .B(n_908), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
NOR2xp33_ASAP7_75t_R g914 ( .A(n_907), .B(n_915), .Y(n_914) );
INVx1_ASAP7_75t_L g916 ( .A(n_908), .Y(n_916) );
CKINVDCx5p33_ASAP7_75t_R g909 ( .A(n_910), .Y(n_909) );
NOR2xp33_ASAP7_75t_R g917 ( .A(n_918), .B(n_919), .Y(n_917) );
BUFx6f_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
BUFx6f_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
CKINVDCx5p33_ASAP7_75t_R g924 ( .A(n_925), .Y(n_924) );
CKINVDCx5p33_ASAP7_75t_R g925 ( .A(n_926), .Y(n_925) );
BUFx6f_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
BUFx6f_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
BUFx6f_ASAP7_75t_L g935 ( .A(n_928), .Y(n_935) );
INVx1_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
CKINVDCx5p33_ASAP7_75t_R g934 ( .A(n_935), .Y(n_934) );
endmodule