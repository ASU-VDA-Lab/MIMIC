module fake_jpeg_17213_n_88 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_88);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_88;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx8_ASAP7_75t_SL g10 ( 
.A(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_1),
.B(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_0),
.C(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_20),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_2),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_21),
.B(n_22),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_16),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_13),
.B(n_16),
.C(n_15),
.Y(n_29)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_31),
.Y(n_33)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_19),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_18),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_35),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_31),
.A2(n_18),
.B1(n_12),
.B2(n_11),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_9),
.C(n_15),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_12),
.B1(n_11),
.B2(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_40),
.B(n_30),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_12),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_26),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_SL g53 ( 
.A(n_44),
.B(n_33),
.C(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_28),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_47),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_40),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_52),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_37),
.B(n_30),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_26),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_55),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_33),
.B(n_32),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_61),
.B(n_42),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_36),
.C(n_32),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_50),
.C(n_45),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_60),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_63),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_56),
.C(n_59),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_57),
.B(n_67),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_57),
.B1(n_14),
.B2(n_13),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_71),
.A2(n_73),
.B1(n_2),
.B2(n_3),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_62),
.C(n_63),
.Y(n_74)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_66),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_77),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_9),
.C(n_27),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_72),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_13),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_76),
.B(n_69),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_79),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_80),
.A2(n_3),
.B(n_4),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_81),
.A2(n_82),
.B(n_6),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_80),
.A2(n_5),
.B(n_6),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_83),
.B(n_5),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_85),
.C(n_6),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_27),
.B1(n_8),
.B2(n_7),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_7),
.Y(n_88)
);


endmodule