module fake_jpeg_14261_n_186 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_186);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_122;
wire n_75;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_19),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_8),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_5),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_51),
.Y(n_72)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_25),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_43),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_6),
.B(n_0),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_49),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_52),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_13),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_39),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_2),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

CKINVDCx9p33_ASAP7_75t_R g85 ( 
.A(n_58),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_1),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_89),
.Y(n_96)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_1),
.Y(n_89)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_64),
.Y(n_97)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_92),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_55),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_72),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_64),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_90),
.A2(n_57),
.B1(n_80),
.B2(n_65),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_103),
.A2(n_105),
.B1(n_67),
.B2(n_83),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_70),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_104),
.B(n_106),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_91),
.A2(n_57),
.B1(n_80),
.B2(n_65),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_81),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_79),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_107),
.B(n_59),
.Y(n_129)
);

HAxp5_ASAP7_75t_SL g108 ( 
.A(n_88),
.B(n_64),
.CON(n_108),
.SN(n_108)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_71),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_95),
.A2(n_84),
.B1(n_83),
.B2(n_62),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_131),
.B1(n_26),
.B2(n_47),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_110),
.A2(n_119),
.B(n_120),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_113),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_98),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_118),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_96),
.B(n_66),
.Y(n_115)
);

NAND3xp33_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_121),
.C(n_130),
.Y(n_146)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_108),
.A2(n_63),
.B(n_73),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_73),
.B(n_68),
.Y(n_120)
);

NAND2x1_ASAP7_75t_SL g121 ( 
.A(n_100),
.B(n_84),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_122),
.A2(n_125),
.B1(n_60),
.B2(n_4),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_75),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_126),
.Y(n_136)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_101),
.A2(n_67),
.B1(n_76),
.B2(n_74),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_54),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_128),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_78),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_3),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_2),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_103),
.A2(n_60),
.B1(n_4),
.B2(n_5),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_137),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_123),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_140),
.B(n_151),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_SL g141 ( 
.A1(n_120),
.A2(n_24),
.B(n_46),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_141),
.A2(n_149),
.B(n_37),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_110),
.A2(n_23),
.B1(n_44),
.B2(n_42),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_142),
.A2(n_144),
.B1(n_145),
.B2(n_147),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_122),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_119),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_15),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_18),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_152),
.B(n_28),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_20),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_156),
.B(n_160),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_159),
.Y(n_174)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_29),
.C(n_31),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_32),
.B(n_33),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_161),
.A2(n_166),
.B1(n_142),
.B2(n_141),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_36),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_162),
.A2(n_132),
.B1(n_146),
.B2(n_167),
.Y(n_171)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_164),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_139),
.B(n_148),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_165),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_133),
.A2(n_38),
.B1(n_48),
.B2(n_138),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_168),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_171),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_172),
.A2(n_154),
.B1(n_157),
.B2(n_166),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_173),
.C(n_169),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_178),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_177),
.A2(n_154),
.B(n_171),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_174),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_181),
.A2(n_155),
.B(n_162),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_175),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_170),
.C(n_160),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_146),
.B(n_179),
.Y(n_185)
);

XNOR2x2_ASAP7_75t_SL g186 ( 
.A(n_185),
.B(n_163),
.Y(n_186)
);


endmodule