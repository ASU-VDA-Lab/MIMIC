module fake_jpeg_30576_n_70 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_70);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_70;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_51;
wire n_47;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_32;
wire n_66;

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_13),
.A2(n_9),
.B(n_19),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_12),
.B(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_36),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g33 ( 
.A(n_25),
.Y(n_33)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_29),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_34),
.B(n_38),
.Y(n_41)
);

OA21x2_ASAP7_75t_L g35 ( 
.A1(n_27),
.A2(n_0),
.B(n_1),
.Y(n_35)
);

OAI22x1_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_20),
.B1(n_14),
.B2(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_24),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_27),
.A2(n_23),
.B1(n_22),
.B2(n_21),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_46),
.B1(n_41),
.B2(n_42),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_16),
.C(n_15),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_35),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_44),
.A2(n_37),
.B1(n_35),
.B2(n_8),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_50),
.B1(n_53),
.B2(n_10),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_6),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_46),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_10),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_11),
.Y(n_57)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_55),
.Y(n_60)
);

OAI211xp5_ASAP7_75t_L g63 ( 
.A1(n_56),
.A2(n_53),
.B(n_48),
.C(n_57),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_57),
.B(n_58),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_47),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_52),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_64),
.B(n_65),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_63),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_59),
.B(n_11),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_62),
.Y(n_68)
);

OA21x2_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_67),
.B(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_69),
.B(n_60),
.Y(n_70)
);


endmodule