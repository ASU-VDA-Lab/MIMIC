module fake_jpeg_919_n_199 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_199);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx4f_ASAP7_75t_SL g55 ( 
.A(n_23),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_13),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_3),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_2),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

BUFx4f_ASAP7_75t_SL g60 ( 
.A(n_45),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_47),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_7),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_19),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_74),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_0),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_1),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_55),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_52),
.Y(n_79)
);

INVx4_ASAP7_75t_SL g81 ( 
.A(n_79),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_53),
.B1(n_69),
.B2(n_50),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_82),
.A2(n_91),
.B1(n_78),
.B2(n_64),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_79),
.A2(n_52),
.B1(n_53),
.B2(n_58),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_84),
.A2(n_79),
.B1(n_78),
.B2(n_60),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_55),
.B1(n_60),
.B2(n_56),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_87),
.B1(n_81),
.B2(n_94),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_86),
.B(n_90),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_77),
.A2(n_55),
.B1(n_60),
.B2(n_57),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_62),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_76),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_66),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_80),
.A2(n_72),
.B1(n_70),
.B2(n_67),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_79),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_95),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_96),
.B(n_100),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_73),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_105),
.Y(n_119)
);

AND2x4_ASAP7_75t_SL g99 ( 
.A(n_92),
.B(n_80),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_99),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_83),
.B(n_51),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_81),
.Y(n_102)
);

INVxp67_ASAP7_75t_SL g113 ( 
.A(n_102),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_54),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_103),
.B(n_110),
.Y(n_131)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_71),
.C(n_61),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_111),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_5),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_81),
.A2(n_64),
.B1(n_68),
.B2(n_4),
.Y(n_109)
);

AOI22x1_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_64),
.B1(n_68),
.B2(n_93),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_1),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_89),
.B(n_2),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_116),
.A2(n_132),
.B1(n_15),
.B2(n_16),
.Y(n_149)
);

NOR2x1_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_68),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_117),
.A2(n_95),
.B(n_99),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_30),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_6),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_126),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_7),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_8),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_130),
.Y(n_138)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

FAx1_ASAP7_75t_SL g129 ( 
.A(n_99),
.B(n_9),
.CI(n_10),
.CON(n_129),
.SN(n_129)
);

A2O1A1O1Ixp25_ASAP7_75t_L g141 ( 
.A1(n_129),
.A2(n_11),
.B(n_12),
.C(n_13),
.D(n_14),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_26),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_136),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_137),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_104),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_105),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_139),
.B(n_144),
.Y(n_164)
);

NAND3xp33_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_155),
.C(n_18),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_112),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_142),
.Y(n_161)
);

OA21x2_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_28),
.B(n_44),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_121),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_147),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_118),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_146),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_116),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_119),
.B(n_14),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_148),
.B(n_152),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_149),
.A2(n_18),
.B1(n_24),
.B2(n_25),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_15),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_150),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_114),
.A2(n_31),
.B1(n_40),
.B2(n_39),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_151),
.A2(n_33),
.B(n_22),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_16),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_132),
.A2(n_27),
.B1(n_38),
.B2(n_20),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_153),
.A2(n_114),
.B1(n_129),
.B2(n_17),
.Y(n_157)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_140),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_129),
.B(n_17),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_157),
.A2(n_165),
.B1(n_142),
.B2(n_133),
.Y(n_181)
);

NOR3xp33_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_171),
.C(n_143),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_169),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_146),
.A2(n_34),
.B(n_35),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_170),
.A2(n_141),
.B(n_151),
.Y(n_175)
);

NAND3xp33_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_37),
.C(n_49),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_135),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_172),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_178),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_181),
.C(n_162),
.Y(n_185)
);

BUFx24_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_176),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_156),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_167),
.A2(n_143),
.B1(n_137),
.B2(n_153),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_179),
.B(n_180),
.Y(n_186)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

XOR2x2_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_158),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_184),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_164),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_187),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_166),
.C(n_159),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_186),
.A2(n_188),
.B(n_183),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_176),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_163),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_162),
.Y(n_193)
);

AOI21x1_ASAP7_75t_L g195 ( 
.A1(n_193),
.A2(n_194),
.B(n_190),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_195),
.A2(n_191),
.B(n_173),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_196),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_168),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_171),
.Y(n_199)
);


endmodule