module fake_jpeg_25241_n_141 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_141);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx5_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_19),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_43),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_30),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_36),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_4),
.B(n_12),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_35),
.Y(n_61)
);

INVx8_ASAP7_75t_SL g62 ( 
.A(n_9),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_33),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_0),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_71),
.Y(n_77)
);

BUFx4f_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_72),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_0),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_56),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_73),
.A2(n_46),
.B1(n_59),
.B2(n_69),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_74),
.A2(n_76),
.B1(n_85),
.B2(n_87),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_69),
.A2(n_59),
.B1(n_66),
.B2(n_55),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_67),
.B(n_66),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_3),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_49),
.C(n_64),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_78),
.B(n_81),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_70),
.A2(n_64),
.B1(n_50),
.B2(n_52),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVxp67_ASAP7_75t_SL g93 ( 
.A(n_84),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_72),
.A2(n_65),
.B1(n_63),
.B2(n_61),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_1),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_68),
.A2(n_47),
.B1(n_48),
.B2(n_53),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_77),
.A2(n_50),
.B(n_52),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_77),
.A2(n_57),
.B1(n_54),
.B2(n_60),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_89),
.B(n_91),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_20),
.B(n_41),
.Y(n_91)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_83),
.Y(n_94)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_96),
.B(n_97),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_84),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_99),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_81),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_5),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_4),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_80),
.C(n_75),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_6),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_108),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_110),
.B(n_5),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_103),
.A2(n_95),
.B1(n_90),
.B2(n_96),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_111),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_126)
);

AO21x1_ASAP7_75t_L g112 ( 
.A1(n_109),
.A2(n_91),
.B(n_93),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_115),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_109),
.A2(n_94),
.B1(n_101),
.B2(n_23),
.Y(n_113)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_116),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_6),
.C(n_8),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_112),
.A2(n_107),
.B(n_105),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_123),
.C(n_124),
.Y(n_129)
);

AO22x1_ASAP7_75t_SL g122 ( 
.A1(n_111),
.A2(n_102),
.B1(n_8),
.B2(n_10),
.Y(n_122)
);

BUFx4f_ASAP7_75t_SL g131 ( 
.A(n_122),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_117),
.C(n_113),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_126),
.A2(n_11),
.B(n_116),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_128),
.A2(n_120),
.B1(n_125),
.B2(n_122),
.Y(n_133)
);

NOR3xp33_ASAP7_75t_SL g130 ( 
.A(n_125),
.B(n_13),
.C(n_14),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_15),
.C(n_18),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_132),
.A2(n_133),
.B1(n_129),
.B2(n_131),
.Y(n_134)
);

OAI21x1_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_127),
.B(n_22),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_21),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_136),
.B(n_24),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_26),
.B(n_29),
.Y(n_138)
);

FAx1_ASAP7_75t_SL g139 ( 
.A(n_138),
.B(n_32),
.CI(n_37),
.CON(n_139),
.SN(n_139)
);

AOI322xp5_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_38),
.A3(n_39),
.B1(n_40),
.B2(n_44),
.C1(n_114),
.C2(n_121),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_139),
.Y(n_141)
);


endmodule