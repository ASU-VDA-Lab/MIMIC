module fake_jpeg_18960_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_26),
.B(n_16),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_12),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g38 ( 
.A(n_27),
.B(n_15),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_46),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_33),
.A2(n_25),
.B1(n_23),
.B2(n_21),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_44),
.B1(n_45),
.B2(n_22),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_31),
.A2(n_15),
.B1(n_23),
.B2(n_21),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_L g45 ( 
.A1(n_32),
.A2(n_15),
.B1(n_25),
.B2(n_16),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_48),
.B1(n_49),
.B2(n_17),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_46),
.A2(n_32),
.B1(n_27),
.B2(n_33),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_12),
.B1(n_14),
.B2(n_20),
.Y(n_49)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_12),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_18),
.B1(n_17),
.B2(n_20),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_59),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_29),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_58),
.C(n_29),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_22),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_39),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_30),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_45),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_30),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_61),
.A2(n_65),
.B(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_72),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_28),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_58),
.B(n_57),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_42),
.B1(n_43),
.B2(n_18),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_29),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_73),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_35),
.Y(n_68)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_30),
.C(n_39),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_74),
.A2(n_65),
.B(n_61),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_76),
.A2(n_58),
.B(n_71),
.Y(n_97)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_50),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_82),
.B(n_83),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_63),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_62),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_86),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_61),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_87),
.B(n_92),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_90),
.B(n_94),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_67),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_65),
.C(n_58),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_85),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_80),
.Y(n_95)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

AOI221xp5_ASAP7_75t_L g99 ( 
.A1(n_97),
.A2(n_77),
.B1(n_71),
.B2(n_86),
.C(n_78),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_99),
.B(n_100),
.Y(n_112)
);

AOI322xp5_ASAP7_75t_L g100 ( 
.A1(n_89),
.A2(n_84),
.A3(n_49),
.B1(n_47),
.B2(n_48),
.C1(n_80),
.C2(n_69),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_105),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_84),
.B(n_69),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_103),
.A2(n_90),
.B(n_93),
.Y(n_110)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_106),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_105),
.A2(n_96),
.B1(n_97),
.B2(n_94),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_111),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_110),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_107),
.A2(n_98),
.B1(n_51),
.B2(n_55),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_103),
.A2(n_51),
.B1(n_43),
.B2(n_34),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_115),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_104),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_114),
.A2(n_102),
.B1(n_108),
.B2(n_106),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_121),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_34),
.C(n_35),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_35),
.C(n_28),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_115),
.Y(n_125)
);

OA21x2_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_116),
.B(n_110),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_126),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_125),
.A2(n_9),
.B(n_3),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_117),
.A2(n_109),
.B(n_113),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_118),
.B(n_11),
.Y(n_127)
);

OAI221xp5_ASAP7_75t_L g129 ( 
.A1(n_127),
.A2(n_10),
.B1(n_9),
.B2(n_121),
.C(n_40),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_130),
.Y(n_132)
);

OAI221xp5_ASAP7_75t_L g131 ( 
.A1(n_123),
.A2(n_28),
.B1(n_4),
.B2(n_5),
.C(n_7),
.Y(n_131)
);

OAI321xp33_ASAP7_75t_L g133 ( 
.A1(n_131),
.A2(n_2),
.A3(n_5),
.B1(n_7),
.B2(n_8),
.C(n_128),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_132),
.A2(n_2),
.B(n_5),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_8),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_135),
.Y(n_137)
);


endmodule