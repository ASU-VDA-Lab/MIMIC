module real_aes_1651_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_841, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_841;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_551;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_504;
wire n_119;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_733;
wire n_552;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
NAND2xp5_ASAP7_75t_L g219 ( .A(n_0), .B(n_156), .Y(n_219) );
CKINVDCx5p33_ASAP7_75t_R g793 ( .A(n_1), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_2), .B(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g128 ( .A(n_3), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_4), .B(n_132), .Y(n_177) );
NAND2xp33_ASAP7_75t_SL g239 ( .A(n_5), .B(n_138), .Y(n_239) );
INVx1_ASAP7_75t_L g231 ( .A(n_6), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_7), .B(n_182), .Y(n_455) );
INVx1_ASAP7_75t_L g499 ( .A(n_8), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g809 ( .A(n_9), .Y(n_809) );
AND2x2_ASAP7_75t_L g175 ( .A(n_10), .B(n_161), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g491 ( .A(n_11), .Y(n_491) );
INVx2_ASAP7_75t_L g120 ( .A(n_12), .Y(n_120) );
CKINVDCx16_ASAP7_75t_R g440 ( .A(n_13), .Y(n_440) );
INVx1_ASAP7_75t_L g464 ( .A(n_14), .Y(n_464) );
AOI221x1_ASAP7_75t_L g234 ( .A1(n_15), .A2(n_140), .B1(n_235), .B2(n_237), .C(n_238), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_16), .B(n_132), .Y(n_199) );
INVx1_ASAP7_75t_L g444 ( .A(n_17), .Y(n_444) );
INVx1_ASAP7_75t_L g462 ( .A(n_18), .Y(n_462) );
INVx1_ASAP7_75t_SL g558 ( .A(n_19), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_20), .B(n_133), .Y(n_532) );
AOI33xp33_ASAP7_75t_L g508 ( .A1(n_21), .A2(n_53), .A3(n_125), .B1(n_145), .B2(n_509), .B3(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_22), .A2(n_140), .B(n_179), .Y(n_178) );
AOI221xp5_ASAP7_75t_SL g208 ( .A1(n_23), .A2(n_40), .B1(n_132), .B2(n_140), .C(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_24), .B(n_156), .Y(n_180) );
INVx1_ASAP7_75t_L g485 ( .A(n_25), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g828 ( .A(n_26), .Y(n_828) );
OAI22x1_ASAP7_75t_R g105 ( .A1(n_27), .A2(n_51), .B1(n_106), .B2(n_107), .Y(n_105) );
INVx1_ASAP7_75t_L g107 ( .A(n_27), .Y(n_107) );
OA21x2_ASAP7_75t_L g119 ( .A1(n_28), .A2(n_90), .B(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g162 ( .A(n_28), .B(n_90), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_29), .B(n_154), .Y(n_203) );
INVxp67_ASAP7_75t_L g233 ( .A(n_30), .Y(n_233) );
AND2x2_ASAP7_75t_L g172 ( .A(n_31), .B(n_160), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_32), .B(n_123), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_33), .A2(n_140), .B(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_34), .B(n_154), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g823 ( .A1(n_35), .A2(n_52), .B1(n_644), .B2(n_824), .Y(n_823) );
CKINVDCx20_ASAP7_75t_R g824 ( .A(n_35), .Y(n_824) );
AND2x2_ASAP7_75t_L g130 ( .A(n_36), .B(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g138 ( .A(n_36), .B(n_128), .Y(n_138) );
INVx1_ASAP7_75t_L g144 ( .A(n_36), .Y(n_144) );
OR2x6_ASAP7_75t_L g442 ( .A(n_37), .B(n_443), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_38), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_39), .B(n_123), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_41), .A2(n_182), .B1(n_215), .B2(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_42), .B(n_534), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g139 ( .A1(n_43), .A2(n_82), .B1(n_140), .B2(n_142), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_44), .B(n_133), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_45), .B(n_156), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_46), .B(n_118), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_47), .B(n_133), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g529 ( .A(n_48), .Y(n_529) );
AND2x2_ASAP7_75t_L g222 ( .A(n_49), .B(n_160), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_50), .B(n_160), .Y(n_212) );
INVx1_ASAP7_75t_L g106 ( .A(n_51), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g644 ( .A(n_52), .Y(n_644) );
HB1xp67_ASAP7_75t_SL g715 ( .A(n_52), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_54), .B(n_133), .Y(n_477) );
AOI222xp33_ASAP7_75t_L g101 ( .A1(n_55), .A2(n_102), .B1(n_802), .B2(n_813), .C1(n_829), .C2(n_833), .Y(n_101) );
OAI22x1_ASAP7_75t_R g822 ( .A1(n_55), .A2(n_823), .B1(n_825), .B2(n_826), .Y(n_822) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_55), .Y(n_826) );
INVx1_ASAP7_75t_L g126 ( .A(n_56), .Y(n_126) );
INVx1_ASAP7_75t_L g135 ( .A(n_56), .Y(n_135) );
AND2x2_ASAP7_75t_L g478 ( .A(n_57), .B(n_160), .Y(n_478) );
AOI221xp5_ASAP7_75t_L g497 ( .A1(n_58), .A2(n_75), .B1(n_123), .B2(n_142), .C(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_59), .B(n_123), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_60), .B(n_132), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_61), .B(n_215), .Y(n_493) );
AOI21xp5_ASAP7_75t_SL g518 ( .A1(n_62), .A2(n_142), .B(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g163 ( .A(n_63), .B(n_160), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_64), .B(n_154), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_65), .B(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_SL g204 ( .A(n_66), .B(n_161), .Y(n_204) );
INVx1_ASAP7_75t_L g458 ( .A(n_67), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_68), .A2(n_140), .B(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g476 ( .A(n_69), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_70), .B(n_154), .Y(n_181) );
AND2x2_ASAP7_75t_SL g147 ( .A(n_71), .B(n_118), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_72), .A2(n_142), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g131 ( .A(n_73), .Y(n_131) );
INVx1_ASAP7_75t_L g137 ( .A(n_73), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_74), .B(n_123), .Y(n_511) );
AND2x2_ASAP7_75t_L g560 ( .A(n_76), .B(n_237), .Y(n_560) );
INVx1_ASAP7_75t_L g460 ( .A(n_77), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_78), .A2(n_142), .B(n_557), .Y(n_556) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_79), .A2(n_117), .B(n_142), .C(n_531), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g122 ( .A1(n_80), .A2(n_85), .B1(n_123), .B2(n_132), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_81), .B(n_132), .Y(n_158) );
INVx1_ASAP7_75t_L g445 ( .A(n_83), .Y(n_445) );
AND2x2_ASAP7_75t_SL g516 ( .A(n_84), .B(n_237), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_86), .A2(n_142), .B1(n_506), .B2(n_507), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_87), .B(n_156), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_88), .B(n_156), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_89), .A2(n_140), .B(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g520 ( .A(n_91), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_92), .B(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_L g512 ( .A(n_93), .B(n_237), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_94), .A2(n_483), .B(n_484), .C(n_486), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_95), .B(n_132), .Y(n_221) );
INVxp67_ASAP7_75t_L g236 ( .A(n_96), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_97), .B(n_154), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_98), .A2(n_140), .B(n_201), .Y(n_200) );
BUFx2_ASAP7_75t_L g810 ( .A(n_99), .Y(n_810) );
BUFx2_ASAP7_75t_SL g837 ( .A(n_99), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_100), .B(n_133), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_103), .B(n_797), .Y(n_102) );
AOI21xp33_ASAP7_75t_SL g103 ( .A1(n_104), .A2(n_108), .B(n_792), .Y(n_103) );
CKINVDCx16_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
NAND2xp33_ASAP7_75t_L g797 ( .A(n_105), .B(n_798), .Y(n_797) );
OAI22x1_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_439), .B1(n_446), .B2(n_788), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OAI22xp5_ASAP7_75t_SL g798 ( .A1(n_110), .A2(n_447), .B1(n_799), .B2(n_800), .Y(n_798) );
AND3x4_ASAP7_75t_L g110 ( .A(n_111), .B(n_310), .C(n_384), .Y(n_110) );
NOR3xp33_ASAP7_75t_L g111 ( .A(n_112), .B(n_252), .C(n_283), .Y(n_111) );
A2O1A1Ixp33_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_185), .B(n_194), .C(n_223), .Y(n_112) );
AOI21x1_ASAP7_75t_SL g113 ( .A1(n_114), .A2(n_164), .B(n_183), .Y(n_113) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_114), .A2(n_286), .B1(n_292), .B2(n_295), .Y(n_285) );
AND2x2_ASAP7_75t_L g419 ( .A(n_114), .B(n_187), .Y(n_419) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_148), .Y(n_114) );
BUFx2_ASAP7_75t_L g190 ( .A(n_115), .Y(n_190) );
AND2x2_ASAP7_75t_L g278 ( .A(n_115), .B(n_149), .Y(n_278) );
AND2x2_ASAP7_75t_L g349 ( .A(n_115), .B(n_193), .Y(n_349) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_116), .Y(n_243) );
AOI21x1_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_121), .B(n_147), .Y(n_116) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_117), .A2(n_504), .B(n_512), .Y(n_503) );
AO21x2_ASAP7_75t_L g575 ( .A1(n_117), .A2(n_504), .B(n_512), .Y(n_575) );
INVx2_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_118), .A2(n_199), .B(n_200), .Y(n_198) );
OA21x2_ASAP7_75t_L g496 ( .A1(n_118), .A2(n_497), .B(n_501), .Y(n_496) );
BUFx4f_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx3_ASAP7_75t_L g215 ( .A(n_119), .Y(n_215) );
AND2x2_ASAP7_75t_SL g161 ( .A(n_120), .B(n_162), .Y(n_161) );
AND2x4_ASAP7_75t_L g182 ( .A(n_120), .B(n_162), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_139), .Y(n_121) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_123), .A2(n_142), .B1(n_230), .B2(n_232), .Y(n_229) );
INVx1_ASAP7_75t_L g494 ( .A(n_123), .Y(n_494) );
AND2x4_ASAP7_75t_L g123 ( .A(n_124), .B(n_129), .Y(n_123) );
INVx1_ASAP7_75t_L g527 ( .A(n_124), .Y(n_527) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_127), .Y(n_124) );
OR2x6_ASAP7_75t_L g459 ( .A(n_125), .B(n_146), .Y(n_459) );
INVxp33_ASAP7_75t_L g509 ( .A(n_125), .Y(n_509) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g141 ( .A(n_126), .B(n_128), .Y(n_141) );
AND2x4_ASAP7_75t_L g154 ( .A(n_126), .B(n_136), .Y(n_154) );
HB1xp67_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g528 ( .A(n_129), .Y(n_528) );
BUFx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x6_ASAP7_75t_L g140 ( .A(n_130), .B(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g146 ( .A(n_131), .Y(n_146) );
AND2x6_ASAP7_75t_L g156 ( .A(n_131), .B(n_134), .Y(n_156) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_138), .Y(n_132) );
INVx1_ASAP7_75t_L g240 ( .A(n_133), .Y(n_240) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_136), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx5_ASAP7_75t_L g157 ( .A(n_138), .Y(n_157) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_138), .Y(n_486) );
AND2x4_ASAP7_75t_L g142 ( .A(n_141), .B(n_143), .Y(n_142) );
INVxp67_ASAP7_75t_L g492 ( .A(n_142), .Y(n_492) );
NOR2x1p5_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
INVx1_ASAP7_75t_L g510 ( .A(n_145), .Y(n_510) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x4_ASAP7_75t_L g242 ( .A(n_148), .B(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g184 ( .A(n_149), .B(n_174), .Y(n_184) );
OR2x2_ASAP7_75t_L g192 ( .A(n_149), .B(n_193), .Y(n_192) );
AND2x4_ASAP7_75t_L g247 ( .A(n_149), .B(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g294 ( .A(n_149), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_149), .B(n_193), .Y(n_302) );
AND2x2_ASAP7_75t_L g339 ( .A(n_149), .B(n_243), .Y(n_339) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_149), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_149), .B(n_173), .Y(n_380) );
AO21x2_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_159), .B(n_163), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_158), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_155), .B(n_157), .Y(n_152) );
INVxp67_ASAP7_75t_L g465 ( .A(n_154), .Y(n_465) );
INVxp67_ASAP7_75t_L g463 ( .A(n_156), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_157), .A2(n_169), .B(n_170), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_157), .A2(n_180), .B(n_181), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_157), .A2(n_202), .B(n_203), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_157), .A2(n_210), .B(n_211), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_157), .A2(n_219), .B(n_220), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_157), .B(n_182), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_157), .A2(n_459), .B(n_476), .C(n_477), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_SL g498 ( .A1(n_157), .A2(n_459), .B(n_499), .C(n_500), .Y(n_498) );
INVx1_ASAP7_75t_L g506 ( .A(n_157), .Y(n_506) );
O2A1O1Ixp33_ASAP7_75t_L g519 ( .A1(n_157), .A2(n_459), .B(n_520), .C(n_521), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_157), .A2(n_532), .B(n_533), .Y(n_531) );
O2A1O1Ixp33_ASAP7_75t_SL g557 ( .A1(n_157), .A2(n_459), .B(n_558), .C(n_559), .Y(n_557) );
AO21x2_ASAP7_75t_L g165 ( .A1(n_159), .A2(n_166), .B(n_172), .Y(n_165) );
AO21x2_ASAP7_75t_L g193 ( .A1(n_159), .A2(n_166), .B(n_172), .Y(n_193) );
AO21x2_ASAP7_75t_L g553 ( .A1(n_159), .A2(n_554), .B(n_560), .Y(n_553) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_160), .Y(n_159) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_160), .A2(n_208), .B(n_212), .Y(n_207) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g281 ( .A(n_164), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_164), .B(n_242), .Y(n_337) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_164), .Y(n_438) );
AND2x4_ASAP7_75t_L g164 ( .A(n_165), .B(n_173), .Y(n_164) );
AND2x2_ASAP7_75t_L g183 ( .A(n_165), .B(n_184), .Y(n_183) );
OR2x2_ASAP7_75t_L g263 ( .A(n_165), .B(n_174), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_165), .B(n_294), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_167), .B(n_171), .Y(n_166) );
AND2x2_ASAP7_75t_L g330 ( .A(n_173), .B(n_247), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_173), .B(n_242), .Y(n_386) );
INVx5_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g188 ( .A(n_174), .Y(n_188) );
AND2x2_ASAP7_75t_L g257 ( .A(n_174), .B(n_248), .Y(n_257) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_174), .Y(n_277) );
AND2x4_ASAP7_75t_L g284 ( .A(n_174), .B(n_193), .Y(n_284) );
AND2x2_ASAP7_75t_SL g431 ( .A(n_174), .B(n_243), .Y(n_431) );
OR2x6_ASAP7_75t_L g174 ( .A(n_175), .B(n_176), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_182), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_182), .B(n_231), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_182), .B(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_182), .B(n_236), .Y(n_235) );
NOR3xp33_ASAP7_75t_L g238 ( .A(n_182), .B(n_239), .C(n_240), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_182), .A2(n_518), .B(n_522), .Y(n_517) );
INVx1_ASAP7_75t_L g410 ( .A(n_183), .Y(n_410) );
INVx1_ASAP7_75t_L g352 ( .A(n_184), .Y(n_352) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_189), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
OR2x2_ASAP7_75t_L g274 ( .A(n_188), .B(n_192), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_188), .B(n_243), .Y(n_367) );
AND2x2_ASAP7_75t_L g369 ( .A(n_188), .B(n_191), .Y(n_369) );
AOI32xp33_ASAP7_75t_L g435 ( .A1(n_188), .A2(n_251), .A3(n_406), .B1(n_436), .B2(n_438), .Y(n_435) );
AND2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
AND2x2_ASAP7_75t_L g261 ( .A(n_190), .B(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g379 ( .A(n_190), .B(n_380), .Y(n_379) );
OR2x2_ASAP7_75t_L g402 ( .A(n_190), .B(n_263), .Y(n_402) );
AND2x2_ASAP7_75t_L g429 ( .A(n_190), .B(n_330), .Y(n_429) );
AND2x2_ASAP7_75t_L g355 ( .A(n_191), .B(n_243), .Y(n_355) );
AND2x2_ASAP7_75t_L g430 ( .A(n_191), .B(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g248 ( .A(n_193), .Y(n_248) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_205), .Y(n_195) );
NOR2x1p5_ASAP7_75t_L g288 ( .A(n_196), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g306 ( .A(n_196), .Y(n_306) );
OR2x2_ASAP7_75t_L g334 ( .A(n_196), .B(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x4_ASAP7_75t_SL g251 ( .A(n_197), .B(n_228), .Y(n_251) );
AND2x4_ASAP7_75t_L g267 ( .A(n_197), .B(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g270 ( .A(n_197), .B(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g298 ( .A(n_197), .B(n_207), .Y(n_298) );
OR2x2_ASAP7_75t_L g323 ( .A(n_197), .B(n_272), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_197), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_197), .B(n_207), .Y(n_358) );
INVx2_ASAP7_75t_L g374 ( .A(n_197), .Y(n_374) );
AND2x2_ASAP7_75t_L g389 ( .A(n_197), .B(n_227), .Y(n_389) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_197), .Y(n_413) );
INVx1_ASAP7_75t_L g418 ( .A(n_197), .Y(n_418) );
OR2x6_ASAP7_75t_L g197 ( .A(n_198), .B(n_204), .Y(n_197) );
AND2x2_ASAP7_75t_L g282 ( .A(n_205), .B(n_267), .Y(n_282) );
AND2x2_ASAP7_75t_L g303 ( .A(n_205), .B(n_251), .Y(n_303) );
INVx1_ASAP7_75t_L g335 ( .A(n_205), .Y(n_335) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_213), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g226 ( .A(n_207), .Y(n_226) );
INVx2_ASAP7_75t_L g272 ( .A(n_207), .Y(n_272) );
BUFx3_ASAP7_75t_L g289 ( .A(n_207), .Y(n_289) );
AND2x2_ASAP7_75t_L g328 ( .A(n_207), .B(n_213), .Y(n_328) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_207), .Y(n_426) );
INVx2_ASAP7_75t_L g241 ( .A(n_213), .Y(n_241) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_213), .Y(n_250) );
INVx1_ASAP7_75t_L g266 ( .A(n_213), .Y(n_266) );
OR2x2_ASAP7_75t_L g271 ( .A(n_213), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g291 ( .A(n_213), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_213), .B(n_268), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_213), .B(n_374), .Y(n_373) );
INVx3_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AOI21x1_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B(n_222), .Y(n_214) );
INVx4_ASAP7_75t_L g237 ( .A(n_215), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_215), .B(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_217), .B(n_221), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_242), .B(n_244), .Y(n_223) );
AND2x2_ASAP7_75t_SL g224 ( .A(n_225), .B(n_227), .Y(n_224) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_225), .Y(n_434) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVxp67_ASAP7_75t_SL g260 ( .A(n_226), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_226), .B(n_266), .Y(n_308) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_226), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_227), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g313 ( .A(n_227), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g364 ( .A(n_227), .Y(n_364) );
AOI221xp5_ASAP7_75t_L g368 ( .A1(n_227), .A2(n_369), .B1(n_370), .B2(n_375), .C(n_378), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_227), .B(n_418), .Y(n_417) );
AND2x4_ASAP7_75t_L g227 ( .A(n_228), .B(n_241), .Y(n_227) );
INVx3_ASAP7_75t_L g268 ( .A(n_228), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_228), .B(n_272), .Y(n_372) );
AND2x2_ASAP7_75t_L g401 ( .A(n_228), .B(n_374), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_228), .B(n_433), .Y(n_432) );
AND2x4_ASAP7_75t_L g228 ( .A(n_229), .B(n_234), .Y(n_228) );
INVx3_ASAP7_75t_L g471 ( .A(n_237), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_237), .A2(n_471), .B1(n_482), .B2(n_487), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_240), .A2(n_458), .B1(n_459), .B2(n_460), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_240), .B(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g309 ( .A(n_242), .B(n_284), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g345 ( .A1(n_242), .A2(n_262), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g246 ( .A(n_243), .B(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g255 ( .A(n_243), .Y(n_255) );
OR2x2_ASAP7_75t_L g301 ( .A(n_243), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_243), .B(n_284), .Y(n_393) );
OR2x2_ASAP7_75t_L g425 ( .A(n_243), .B(n_426), .Y(n_425) );
OR2x2_ASAP7_75t_L g437 ( .A(n_243), .B(n_343), .Y(n_437) );
INVxp67_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_249), .Y(n_245) );
INVx2_ASAP7_75t_L g315 ( .A(n_246), .Y(n_315) );
INVx3_ASAP7_75t_SL g381 ( .A(n_247), .Y(n_381) );
INVxp67_ASAP7_75t_L g331 ( .A(n_249), .Y(n_331) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
AOI322xp5_ASAP7_75t_L g253 ( .A1(n_251), .A2(n_254), .A3(n_258), .B1(n_261), .B2(n_264), .C1(n_269), .C2(n_273), .Y(n_253) );
INVx1_ASAP7_75t_SL g342 ( .A(n_251), .Y(n_342) );
AND2x4_ASAP7_75t_L g427 ( .A(n_251), .B(n_314), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_275), .Y(n_252) );
NOR2x1_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
OR2x2_ASAP7_75t_L g280 ( .A(n_255), .B(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g376 ( .A(n_255), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g404 ( .A(n_255), .B(n_257), .Y(n_404) );
AOI32xp33_ASAP7_75t_L g405 ( .A1(n_255), .A2(n_256), .A3(n_406), .B1(n_408), .B2(n_411), .Y(n_405) );
OR2x2_ASAP7_75t_L g409 ( .A(n_255), .B(n_302), .Y(n_409) );
NAND3xp33_ASAP7_75t_L g365 ( .A(n_256), .B(n_281), .C(n_366), .Y(n_365) );
OAI22xp33_ASAP7_75t_SL g385 ( .A1(n_256), .A2(n_322), .B1(n_386), .B2(n_387), .Y(n_385) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVxp67_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g388 ( .A(n_259), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_263), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
OAI322xp33_ASAP7_75t_L g311 ( .A1(n_267), .A2(n_271), .A3(n_280), .B1(n_312), .B2(n_315), .C1(n_316), .C2(n_317), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_267), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_267), .B(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g290 ( .A(n_268), .B(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g322 ( .A(n_268), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_268), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g383 ( .A(n_271), .Y(n_383) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_272), .Y(n_314) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OAI21xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_279), .B(n_282), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_278), .B(n_326), .Y(n_325) );
AOI322xp5_ASAP7_75t_SL g420 ( .A1(n_278), .A2(n_284), .A3(n_401), .B1(n_419), .B2(n_421), .C1(n_424), .C2(n_427), .Y(n_420) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OAI21xp33_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_285), .B(n_299), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_284), .B(n_294), .Y(n_316) );
INVx2_ASAP7_75t_SL g326 ( .A(n_284), .Y(n_326) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
INVx1_ASAP7_75t_SL g351 ( .A(n_290), .Y(n_351) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_291), .Y(n_321) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g396 ( .A(n_297), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g350 ( .A(n_298), .B(n_351), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_303), .B1(n_304), .B2(n_309), .Y(n_299) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NOR4xp75_ASAP7_75t_L g310 ( .A(n_311), .B(n_324), .C(n_344), .D(n_360), .Y(n_310) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
INVxp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_SL g318 ( .A(n_319), .B(n_322), .Y(n_318) );
INVxp67_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_322), .A2(n_399), .B1(n_402), .B2(n_403), .Y(n_398) );
OR2x2_ASAP7_75t_L g363 ( .A(n_323), .B(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g407 ( .A(n_323), .Y(n_407) );
OAI221xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_327), .B1(n_329), .B2(n_331), .C(n_332), .Y(n_324) );
INVx2_ASAP7_75t_L g343 ( .A(n_328), .Y(n_343) );
AND2x2_ASAP7_75t_L g400 ( .A(n_328), .B(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AOI22xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_336), .B1(n_338), .B2(n_340), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g395 ( .A(n_339), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_340), .A2(n_346), .B1(n_362), .B2(n_365), .Y(n_361) );
INVx1_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
OAI221xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_350), .B1(n_352), .B2(n_353), .C(n_841), .Y(n_344) );
AND2x2_ASAP7_75t_SL g346 ( .A(n_347), .B(n_349), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g412 ( .A(n_351), .B(n_413), .Y(n_412) );
INVxp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx1_ASAP7_75t_L g397 ( .A(n_359), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_368), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
AOI21xp33_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_381), .B(n_382), .Y(n_378) );
NOR3xp33_ASAP7_75t_SL g384 ( .A(n_385), .B(n_390), .C(n_414), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_391), .B(n_405), .Y(n_390) );
O2A1O1Ixp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_394), .B(n_396), .C(n_398), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AND2x4_ASAP7_75t_L g406 ( .A(n_397), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g403 ( .A(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_SL g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
NAND4xp25_ASAP7_75t_SL g414 ( .A(n_415), .B(n_420), .C(n_428), .D(n_435), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_416), .B(n_419), .Y(n_415) );
INVx1_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
INVxp67_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
OAI21xp5_ASAP7_75t_SL g428 ( .A1(n_429), .A2(n_430), .B(n_432), .Y(n_428) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx3_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
CKINVDCx11_ASAP7_75t_R g801 ( .A(n_439), .Y(n_801) );
OR2x6_ASAP7_75t_SL g439 ( .A(n_440), .B(n_441), .Y(n_439) );
AND2x6_ASAP7_75t_SL g791 ( .A(n_440), .B(n_442), .Y(n_791) );
OR2x2_ASAP7_75t_L g796 ( .A(n_440), .B(n_442), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_440), .B(n_441), .Y(n_812) );
CKINVDCx5p33_ASAP7_75t_R g441 ( .A(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AOI211x1_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_644), .B(n_645), .C(n_785), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AND4x1_ASAP7_75t_L g785 ( .A(n_449), .B(n_646), .C(n_786), .D(n_787), .Y(n_785) );
NAND3x1_ASAP7_75t_L g820 ( .A(n_449), .B(n_646), .C(n_821), .Y(n_820) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_612), .Y(n_449) );
AOI211xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_535), .B(n_547), .C(n_588), .Y(n_450) );
OAI21xp33_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_467), .B(n_513), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
A2O1A1Ixp33_ASAP7_75t_SL g535 ( .A1(n_453), .A2(n_536), .B(n_541), .C(n_546), .Y(n_535) );
NAND2x1_ASAP7_75t_L g665 ( .A(n_453), .B(n_666), .Y(n_665) );
NOR2x1_ASAP7_75t_L g756 ( .A(n_453), .B(n_685), .Y(n_756) );
AND2x2_ASAP7_75t_L g775 ( .A(n_453), .B(n_515), .Y(n_775) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx3_ASAP7_75t_L g552 ( .A(n_454), .Y(n_552) );
AND2x2_ASAP7_75t_L g623 ( .A(n_454), .B(n_553), .Y(n_623) );
AND2x2_ASAP7_75t_L g628 ( .A(n_454), .B(n_524), .Y(n_628) );
NOR2x1_ASAP7_75t_SL g744 ( .A(n_454), .B(n_515), .Y(n_744) );
AND2x4_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
OAI21xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_461), .B(n_466), .Y(n_456) );
INVxp67_ASAP7_75t_L g483 ( .A(n_459), .Y(n_483) );
INVx2_ASAP7_75t_L g534 ( .A(n_459), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_463), .B1(n_464), .B2(n_465), .Y(n_461) );
INVx1_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_495), .Y(n_468) );
NAND2x1p5_ASAP7_75t_L g659 ( .A(n_469), .B(n_593), .Y(n_659) );
AND2x2_ASAP7_75t_L g776 ( .A(n_469), .B(n_617), .Y(n_776) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_479), .Y(n_469) );
NOR2x1_ASAP7_75t_L g544 ( .A(n_470), .B(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g565 ( .A(n_470), .Y(n_565) );
AND2x2_ASAP7_75t_L g573 ( .A(n_470), .B(n_574), .Y(n_573) );
NOR2xp67_ASAP7_75t_L g711 ( .A(n_470), .B(n_479), .Y(n_711) );
AO21x2_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B(n_478), .Y(n_470) );
AO21x2_ASAP7_75t_L g596 ( .A1(n_471), .A2(n_472), .B(n_478), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
AND2x2_ASAP7_75t_L g663 ( .A(n_479), .B(n_503), .Y(n_663) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x4_ASAP7_75t_L g539 ( .A(n_480), .B(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g543 ( .A(n_480), .Y(n_543) );
INVx1_ASAP7_75t_L g563 ( .A(n_480), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_480), .B(n_596), .Y(n_620) );
AND2x2_ASAP7_75t_L g669 ( .A(n_480), .B(n_496), .Y(n_669) );
OR2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_488), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_492), .B1(n_493), .B2(n_494), .Y(n_488) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g624 ( .A(n_495), .B(n_619), .Y(n_624) );
AND2x2_ASAP7_75t_L g680 ( .A(n_495), .B(n_563), .Y(n_680) );
AND2x2_ASAP7_75t_L g695 ( .A(n_495), .B(n_609), .Y(n_695) );
AND2x2_ASAP7_75t_L g732 ( .A(n_495), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g748 ( .A(n_495), .Y(n_748) );
AND2x4_ASAP7_75t_L g495 ( .A(n_496), .B(n_502), .Y(n_495) );
INVx2_ASAP7_75t_L g540 ( .A(n_496), .Y(n_540) );
INVx1_ASAP7_75t_L g545 ( .A(n_496), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_496), .B(n_575), .Y(n_578) );
INVx1_ASAP7_75t_L g592 ( .A(n_496), .Y(n_592) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_496), .Y(n_602) );
INVxp67_ASAP7_75t_L g618 ( .A(n_496), .Y(n_618) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g537 ( .A(n_503), .Y(n_537) );
AND2x4_ASAP7_75t_L g564 ( .A(n_503), .B(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_505), .B(n_511), .Y(n_504) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g546 ( .A(n_513), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_513), .B(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_SL g567 ( .A(n_514), .B(n_568), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_514), .B(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_514), .B(n_581), .Y(n_724) );
HB1xp67_ASAP7_75t_L g762 ( .A(n_514), .Y(n_762) );
AND2x4_ASAP7_75t_L g514 ( .A(n_515), .B(n_523), .Y(n_514) );
INVx2_ASAP7_75t_L g587 ( .A(n_515), .Y(n_587) );
AND2x2_ASAP7_75t_L g598 ( .A(n_515), .B(n_524), .Y(n_598) );
INVx4_ASAP7_75t_L g606 ( .A(n_515), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_515), .B(n_582), .Y(n_642) );
BUFx6f_ASAP7_75t_L g655 ( .A(n_515), .Y(n_655) );
OR2x6_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
AND2x4_ASAP7_75t_L g633 ( .A(n_523), .B(n_606), .Y(n_633) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x4_ASAP7_75t_L g584 ( .A(n_524), .B(n_552), .Y(n_584) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_524), .Y(n_605) );
INVx2_ASAP7_75t_L g654 ( .A(n_524), .Y(n_654) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_530), .Y(n_524) );
NOR3xp33_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .C(n_529), .Y(n_526) );
OR2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_537), .B(n_542), .Y(n_643) );
NAND2x1_ASAP7_75t_SL g757 ( .A(n_537), .B(n_539), .Y(n_757) );
OR2x2_ASAP7_75t_L g636 ( .A(n_538), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g739 ( .A(n_538), .Y(n_739) );
INVx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g629 ( .A(n_539), .B(n_564), .Y(n_629) );
AND2x2_ASAP7_75t_L g745 ( .A(n_539), .B(n_738), .Y(n_745) );
OAI221xp5_ASAP7_75t_L g753 ( .A1(n_541), .A2(n_754), .B1(n_757), .B2(n_758), .C(n_760), .Y(n_753) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_542), .A2(n_698), .B1(n_700), .B2(n_702), .Y(n_697) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_543), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_SL g611 ( .A(n_543), .Y(n_611) );
BUFx2_ASAP7_75t_L g692 ( .A(n_543), .Y(n_692) );
AND2x2_ASAP7_75t_L g662 ( .A(n_544), .B(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_548), .B(n_566), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_561), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_SL g635 ( .A(n_551), .Y(n_635) );
NAND4xp25_ASAP7_75t_L g760 ( .A(n_551), .B(n_761), .C(n_762), .D(n_763), .Y(n_760) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
INVx1_ASAP7_75t_L g570 ( .A(n_552), .Y(n_570) );
AND2x2_ASAP7_75t_L g653 ( .A(n_552), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g569 ( .A(n_553), .Y(n_569) );
INVx2_ASAP7_75t_L g583 ( .A(n_553), .Y(n_583) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_553), .Y(n_610) );
INVx1_ASAP7_75t_L g627 ( .A(n_553), .Y(n_627) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_553), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
INVx1_ASAP7_75t_L g774 ( .A(n_562), .Y(n_774) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g572 ( .A(n_563), .Y(n_572) );
AND2x2_ASAP7_75t_L g668 ( .A(n_564), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g768 ( .A(n_564), .B(n_769), .Y(n_768) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_571), .B1(n_576), .B2(n_579), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_568), .B(n_633), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_568), .B(n_732), .Y(n_731) );
AND2x4_ASAP7_75t_L g749 ( .A(n_568), .B(n_727), .Y(n_749) );
AOI21xp5_ASAP7_75t_L g779 ( .A1(n_568), .A2(n_604), .B(n_726), .Y(n_779) );
AND2x4_ASAP7_75t_SL g568 ( .A(n_569), .B(n_570), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_569), .B(n_653), .Y(n_690) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_569), .Y(n_706) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
AND2x2_ASAP7_75t_L g576 ( .A(n_572), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g593 ( .A(n_574), .Y(n_593) );
AND2x2_ASAP7_75t_L g617 ( .A(n_574), .B(n_618), .Y(n_617) );
AND2x4_ASAP7_75t_L g738 ( .A(n_574), .B(n_595), .Y(n_738) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_575), .B(n_596), .Y(n_637) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g713 ( .A(n_578), .B(n_620), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_585), .Y(n_579) );
INVx1_ASAP7_75t_L g694 ( .A(n_580), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_584), .Y(n_580) );
NOR3xp33_ASAP7_75t_L g589 ( .A(n_581), .B(n_590), .C(n_594), .Y(n_589) );
AND2x2_ASAP7_75t_L g632 ( .A(n_581), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g661 ( .A(n_581), .B(n_604), .Y(n_661) );
AND2x2_ASAP7_75t_L g743 ( .A(n_581), .B(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g769 ( .A(n_581), .Y(n_769) );
INVx1_ASAP7_75t_L g783 ( .A(n_581), .Y(n_783) );
INVx3_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g586 ( .A(n_584), .B(n_587), .Y(n_586) );
INVx4_ASAP7_75t_L g742 ( .A(n_584), .Y(n_742) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g782 ( .A(n_586), .B(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g685 ( .A(n_587), .Y(n_685) );
AO22x1_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_597), .B1(n_599), .B2(n_607), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
NAND2x1p5_ASAP7_75t_L g675 ( .A(n_591), .B(n_595), .Y(n_675) );
INVx3_ASAP7_75t_L g709 ( .A(n_591), .Y(n_709) );
BUFx3_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx3_ASAP7_75t_L g609 ( .A(n_595), .Y(n_609) );
INVx3_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g687 ( .A(n_596), .B(n_602), .Y(n_687) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_596), .Y(n_734) );
AOI31xp33_ASAP7_75t_L g638 ( .A1(n_597), .A2(n_639), .A3(n_641), .B(n_643), .Y(n_638) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AOI22xp33_ASAP7_75t_SL g614 ( .A1(n_598), .A2(n_615), .B1(n_621), .B2(n_624), .Y(n_614) );
AND2x2_ASAP7_75t_L g698 ( .A(n_598), .B(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g705 ( .A(n_598), .B(n_706), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_600), .B(n_603), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx2_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_604), .B(n_759), .Y(n_758) );
AND2x4_ASAP7_75t_SL g604 ( .A(n_605), .B(n_606), .Y(n_604) );
OR2x2_ASAP7_75t_L g634 ( .A(n_606), .B(n_635), .Y(n_634) );
HB1xp67_ASAP7_75t_L g767 ( .A(n_606), .Y(n_767) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_611), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
AND2x2_ASAP7_75t_L g729 ( .A(n_609), .B(n_669), .Y(n_729) );
INVx1_ASAP7_75t_L g764 ( .A(n_609), .Y(n_764) );
AND2x2_ASAP7_75t_L g714 ( .A(n_610), .B(n_653), .Y(n_714) );
BUFx2_ASAP7_75t_L g759 ( .A(n_610), .Y(n_759) );
AND2x2_ASAP7_75t_L g702 ( .A(n_611), .B(n_703), .Y(n_702) );
NOR3xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_630), .C(n_638), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g613 ( .A(n_614), .B(n_625), .Y(n_613) );
INVx3_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NAND2x1p5_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .Y(n_616) );
AND2x2_ASAP7_75t_L g691 ( .A(n_617), .B(n_692), .Y(n_691) );
INVx2_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_623), .B(n_633), .Y(n_656) );
AND2x2_ASAP7_75t_L g678 ( .A(n_623), .B(n_655), .Y(n_678) );
AND2x2_ASAP7_75t_SL g726 ( .A(n_623), .B(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_626), .B(n_629), .Y(n_625) );
AND2x2_ASAP7_75t_L g781 ( .A(n_626), .B(n_655), .Y(n_781) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
AND2x2_ASAP7_75t_L g755 ( .A(n_627), .B(n_756), .Y(n_755) );
INVx2_ASAP7_75t_L g672 ( .A(n_628), .Y(n_672) );
AND2x2_ASAP7_75t_L g772 ( .A(n_628), .B(n_655), .Y(n_772) );
AOI21xp33_ASAP7_75t_R g630 ( .A1(n_631), .A2(n_634), .B(n_636), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_632), .B(n_736), .Y(n_735) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_633), .Y(n_640) );
INVx1_ASAP7_75t_L g703 ( .A(n_637), .Y(n_703) );
OAI22xp33_ASAP7_75t_L g670 ( .A1(n_639), .A2(n_657), .B1(n_671), .B2(n_673), .Y(n_670) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g671 ( .A(n_642), .B(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_644), .B(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_644), .B(n_751), .Y(n_750) );
NOR2xp67_ASAP7_75t_SL g786 ( .A(n_644), .B(n_717), .Y(n_786) );
OAI211xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_715), .B(n_716), .C(n_750), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_681), .Y(n_646) );
NOR3xp33_ASAP7_75t_L g647 ( .A(n_648), .B(n_670), .C(n_676), .Y(n_647) );
OAI21xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_657), .B(n_660), .Y(n_648) );
INVxp67_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_656), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_652), .A2(n_691), .B1(n_694), .B2(n_695), .Y(n_693) );
AND2x2_ASAP7_75t_SL g652 ( .A(n_653), .B(n_655), .Y(n_652) );
INVx1_ASAP7_75t_L g728 ( .A(n_654), .Y(n_728) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OR2x2_ASAP7_75t_L g720 ( .A(n_659), .B(n_709), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_662), .B1(n_664), .B2(n_668), .Y(n_660) );
INVx1_ASAP7_75t_L g674 ( .A(n_663), .Y(n_674) );
AND2x4_ASAP7_75t_L g686 ( .A(n_663), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g722 ( .A(n_665), .Y(n_722) );
INVx1_ASAP7_75t_L g699 ( .A(n_666), .Y(n_699) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_668), .A2(n_678), .B1(n_726), .B2(n_729), .Y(n_725) );
INVxp67_ASAP7_75t_L g770 ( .A(n_669), .Y(n_770) );
NOR2x1_ASAP7_75t_L g684 ( .A(n_672), .B(n_685), .Y(n_684) );
OR2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
INVxp33_ASAP7_75t_L g784 ( .A(n_675), .Y(n_784) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_677), .B(n_679), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_682), .B(n_696), .Y(n_681) );
NAND2xp5_ASAP7_75t_SL g682 ( .A(n_683), .B(n_693), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_686), .B1(n_688), .B2(n_691), .Y(n_683) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
BUFx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_697), .B(n_704), .Y(n_696) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_707), .B1(n_712), .B2(n_714), .Y(n_704) );
NOR2xp33_ASAP7_75t_SL g707 ( .A(n_708), .B(n_710), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g761 ( .A(n_709), .Y(n_761) );
INVxp67_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g821 ( .A(n_718), .B(n_752), .Y(n_821) );
NOR2x1_ASAP7_75t_L g718 ( .A(n_719), .B(n_730), .Y(n_718) );
OAI21xp5_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_721), .B(n_725), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NAND4xp25_ASAP7_75t_SL g730 ( .A(n_731), .B(n_735), .C(n_740), .D(n_746), .Y(n_730) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_737), .B(n_739), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
AND2x2_ASAP7_75t_L g773 ( .A(n_738), .B(n_774), .Y(n_773) );
OAI21xp5_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_743), .B(n_745), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_749), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g787 ( .A(n_751), .Y(n_787) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
NOR3x1_ASAP7_75t_L g752 ( .A(n_753), .B(n_765), .C(n_777), .Y(n_752) );
INVx1_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
OAI21xp5_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_770), .B(n_771), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_767), .B(n_768), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_773), .B1(n_775), .B2(n_776), .Y(n_771) );
INVx1_ASAP7_75t_L g778 ( .A(n_776), .Y(n_778) );
OAI21xp5_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_779), .B(n_780), .Y(n_777) );
OAI21xp5_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_782), .B(n_784), .Y(n_780) );
CKINVDCx11_ASAP7_75t_R g788 ( .A(n_789), .Y(n_788) );
CKINVDCx6p67_ASAP7_75t_R g799 ( .A(n_789), .Y(n_799) );
INVx3_ASAP7_75t_SL g789 ( .A(n_790), .Y(n_789) );
CKINVDCx5p33_ASAP7_75t_R g790 ( .A(n_791), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g792 ( .A(n_793), .B(n_794), .Y(n_792) );
CKINVDCx5p33_ASAP7_75t_R g794 ( .A(n_795), .Y(n_794) );
INVx3_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_SL g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
AND2x2_ASAP7_75t_L g804 ( .A(n_805), .B(n_811), .Y(n_804) );
INVxp67_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
NAND2xp5_ASAP7_75t_SL g806 ( .A(n_807), .B(n_810), .Y(n_806) );
INVx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
OR2x2_ASAP7_75t_SL g832 ( .A(n_808), .B(n_810), .Y(n_832) );
AOI21xp5_ASAP7_75t_L g834 ( .A1(n_808), .A2(n_835), .B(n_838), .Y(n_834) );
NOR2xp33_ASAP7_75t_SL g827 ( .A(n_811), .B(n_828), .Y(n_827) );
BUFx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
BUFx3_ASAP7_75t_L g817 ( .A(n_812), .Y(n_817) );
BUFx2_ASAP7_75t_L g839 ( .A(n_812), .Y(n_839) );
INVxp67_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
AOI21xp5_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_818), .B(n_827), .Y(n_814) );
CKINVDCx11_ASAP7_75t_R g815 ( .A(n_816), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_817), .Y(n_816) );
INVx2_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
XNOR2xp5_ASAP7_75t_L g819 ( .A(n_820), .B(n_822), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g825 ( .A(n_823), .Y(n_825) );
INVx1_ASAP7_75t_SL g829 ( .A(n_830), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_SL g833 ( .A(n_834), .Y(n_833) );
CKINVDCx11_ASAP7_75t_R g835 ( .A(n_836), .Y(n_835) );
CKINVDCx8_ASAP7_75t_R g836 ( .A(n_837), .Y(n_836) );
INVx2_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
endmodule