module real_aes_1755_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_693;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g233 ( .A(n_0), .B(n_154), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_1), .B(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_2), .B(n_138), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_3), .B(n_156), .Y(n_510) );
INVx1_ASAP7_75t_L g145 ( .A(n_4), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_5), .B(n_138), .Y(n_137) );
NAND2xp33_ASAP7_75t_SL g224 ( .A(n_6), .B(n_144), .Y(n_224) );
INVx1_ASAP7_75t_L g205 ( .A(n_7), .Y(n_205) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_8), .Y(n_115) );
AND2x2_ASAP7_75t_L g132 ( .A(n_9), .B(n_133), .Y(n_132) );
XNOR2xp5_ASAP7_75t_L g123 ( .A(n_10), .B(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g520 ( .A(n_10), .B(n_221), .Y(n_520) );
AND2x2_ASAP7_75t_L g512 ( .A(n_11), .B(n_195), .Y(n_512) );
INVx2_ASAP7_75t_L g134 ( .A(n_12), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_13), .B(n_156), .Y(n_529) );
XNOR2xp5_ASAP7_75t_L g481 ( .A(n_14), .B(n_482), .Y(n_481) );
NOR3xp33_ASAP7_75t_L g113 ( .A(n_15), .B(n_114), .C(n_116), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g471 ( .A(n_15), .Y(n_471) );
AOI221x1_ASAP7_75t_L g218 ( .A1(n_16), .A2(n_147), .B1(n_219), .B2(n_221), .C(n_223), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_17), .B(n_138), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_18), .B(n_138), .Y(n_543) );
INVx1_ASAP7_75t_L g111 ( .A(n_19), .Y(n_111) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_20), .A2(n_91), .B1(n_138), .B2(n_206), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_21), .A2(n_147), .B(n_152), .Y(n_146) );
AOI221xp5_ASAP7_75t_SL g182 ( .A1(n_22), .A2(n_35), .B1(n_138), .B2(n_147), .C(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_23), .B(n_154), .Y(n_153) );
OR2x2_ASAP7_75t_L g135 ( .A(n_24), .B(n_90), .Y(n_135) );
OA21x2_ASAP7_75t_L g196 ( .A1(n_24), .A2(n_90), .B(n_134), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_25), .B(n_156), .Y(n_194) );
INVxp67_ASAP7_75t_L g217 ( .A(n_26), .Y(n_217) );
AND2x2_ASAP7_75t_L g178 ( .A(n_27), .B(n_168), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_28), .A2(n_147), .B(n_232), .Y(n_231) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_29), .A2(n_221), .B(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_30), .B(n_156), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_31), .A2(n_147), .B(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_32), .B(n_156), .Y(n_538) );
AND2x2_ASAP7_75t_L g144 ( .A(n_33), .B(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g148 ( .A(n_33), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g213 ( .A(n_33), .Y(n_213) );
INVxp67_ASAP7_75t_L g116 ( .A(n_34), .Y(n_116) );
OR2x6_ASAP7_75t_L g473 ( .A(n_34), .B(n_110), .Y(n_473) );
XOR2xp5_ASAP7_75t_L g480 ( .A(n_36), .B(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_37), .B(n_138), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g248 ( .A1(n_38), .A2(n_83), .B1(n_147), .B2(n_211), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_39), .B(n_156), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_40), .A2(n_75), .B1(n_463), .B2(n_464), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_40), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_41), .B(n_138), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_42), .B(n_154), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_43), .Y(n_796) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_44), .A2(n_147), .B(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_45), .B(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g236 ( .A(n_46), .B(n_168), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_47), .B(n_154), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_48), .B(n_168), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_49), .B(n_138), .Y(n_526) );
OAI22xp5_ASAP7_75t_SL g460 ( .A1(n_50), .A2(n_461), .B1(n_462), .B2(n_465), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_50), .Y(n_465) );
INVx1_ASAP7_75t_L g141 ( .A(n_51), .Y(n_141) );
INVx1_ASAP7_75t_L g151 ( .A(n_51), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_52), .B(n_156), .Y(n_518) );
AND2x2_ASAP7_75t_L g554 ( .A(n_53), .B(n_168), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_54), .B(n_138), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_55), .B(n_154), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_56), .B(n_154), .Y(n_537) );
AND2x2_ASAP7_75t_L g169 ( .A(n_57), .B(n_168), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_58), .B(n_138), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_59), .B(n_156), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_60), .B(n_138), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_61), .A2(n_147), .B(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_62), .B(n_154), .Y(n_165) );
AND2x2_ASAP7_75t_SL g197 ( .A(n_63), .B(n_133), .Y(n_197) );
AND2x2_ASAP7_75t_L g549 ( .A(n_64), .B(n_133), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_65), .A2(n_147), .B(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_66), .B(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_SL g249 ( .A(n_67), .B(n_195), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_68), .B(n_154), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_69), .B(n_154), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_70), .A2(n_94), .B1(n_147), .B2(n_211), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_71), .B(n_156), .Y(n_546) );
INVx1_ASAP7_75t_L g143 ( .A(n_72), .Y(n_143) );
INVx1_ASAP7_75t_L g149 ( .A(n_72), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_73), .B(n_154), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_74), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_75), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_76), .A2(n_147), .B(n_558), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_77), .A2(n_147), .B(n_500), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_78), .A2(n_147), .B(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g540 ( .A(n_79), .B(n_133), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_80), .B(n_168), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_81), .B(n_138), .Y(n_166) );
AOI22xp5_ASAP7_75t_L g247 ( .A1(n_82), .A2(n_85), .B1(n_138), .B2(n_206), .Y(n_247) );
INVx1_ASAP7_75t_L g112 ( .A(n_84), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_86), .B(n_154), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_87), .B(n_154), .Y(n_185) );
AND2x2_ASAP7_75t_L g503 ( .A(n_88), .B(n_195), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_89), .A2(n_147), .B(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_92), .B(n_156), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_93), .A2(n_147), .B(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_95), .B(n_156), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_96), .A2(n_103), .B1(n_483), .B2(n_484), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_96), .Y(n_483) );
INVxp67_ASAP7_75t_L g220 ( .A(n_97), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_98), .B(n_138), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_99), .B(n_156), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_100), .A2(n_147), .B(n_192), .Y(n_191) );
BUFx2_ASAP7_75t_L g548 ( .A(n_101), .Y(n_548) );
BUFx2_ASAP7_75t_L g121 ( .A(n_102), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_102), .B(n_474), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_103), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_117), .B(n_799), .Y(n_104) );
BUFx3_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_107), .Y(n_801) );
INVx2_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_SL g108 ( .A(n_109), .B(n_113), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
OA22x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_122), .B1(n_478), .B2(n_479), .Y(n_117) );
CKINVDCx11_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_120), .Y(n_119) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI21xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_466), .B(n_474), .Y(n_122) );
OAI22x1_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_126), .B1(n_459), .B2(n_460), .Y(n_124) );
OAI22x1_ASAP7_75t_L g793 ( .A1(n_125), .A2(n_486), .B1(n_791), .B2(n_794), .Y(n_793) );
INVx4_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_126), .A2(n_486), .B1(n_490), .B2(n_789), .Y(n_485) );
AND2x4_ASAP7_75t_L g126 ( .A(n_127), .B(n_370), .Y(n_126) );
NOR3xp33_ASAP7_75t_L g127 ( .A(n_128), .B(n_292), .C(n_342), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_259), .Y(n_128) );
AOI221xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_179), .B1(n_198), .B2(n_241), .C(n_251), .Y(n_129) );
INVx1_ASAP7_75t_SL g341 ( .A(n_130), .Y(n_341) );
AND2x4_ASAP7_75t_SL g130 ( .A(n_131), .B(n_159), .Y(n_130) );
INVx2_ASAP7_75t_L g263 ( .A(n_131), .Y(n_263) );
OR2x2_ASAP7_75t_L g285 ( .A(n_131), .B(n_276), .Y(n_285) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_131), .Y(n_300) );
INVx5_ASAP7_75t_L g307 ( .A(n_131), .Y(n_307) );
AND2x4_ASAP7_75t_L g313 ( .A(n_131), .B(n_171), .Y(n_313) );
AND2x2_ASAP7_75t_SL g316 ( .A(n_131), .B(n_243), .Y(n_316) );
OR2x2_ASAP7_75t_L g325 ( .A(n_131), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g332 ( .A(n_131), .B(n_160), .Y(n_332) );
AND2x2_ASAP7_75t_L g433 ( .A(n_131), .B(n_170), .Y(n_433) );
OR2x6_ASAP7_75t_L g131 ( .A(n_132), .B(n_136), .Y(n_131) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_133), .Y(n_168) );
AND2x2_ASAP7_75t_SL g133 ( .A(n_134), .B(n_135), .Y(n_133) );
AND2x4_ASAP7_75t_L g158 ( .A(n_134), .B(n_135), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_146), .B(n_158), .Y(n_136) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_144), .Y(n_138) );
INVx1_ASAP7_75t_L g225 ( .A(n_139), .Y(n_225) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
AND2x6_ASAP7_75t_L g154 ( .A(n_140), .B(n_149), .Y(n_154) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x4_ASAP7_75t_L g156 ( .A(n_142), .B(n_151), .Y(n_156) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx5_ASAP7_75t_L g157 ( .A(n_144), .Y(n_157) );
AND2x2_ASAP7_75t_L g150 ( .A(n_145), .B(n_151), .Y(n_150) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_145), .Y(n_209) );
AND2x6_ASAP7_75t_L g147 ( .A(n_148), .B(n_150), .Y(n_147) );
BUFx3_ASAP7_75t_L g210 ( .A(n_148), .Y(n_210) );
INVx2_ASAP7_75t_L g215 ( .A(n_149), .Y(n_215) );
AND2x4_ASAP7_75t_L g211 ( .A(n_150), .B(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g208 ( .A(n_151), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_155), .B(n_157), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_154), .B(n_548), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_157), .A2(n_164), .B(n_165), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_157), .A2(n_175), .B(n_176), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_157), .A2(n_184), .B(n_185), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_157), .A2(n_193), .B(n_194), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_157), .A2(n_233), .B(n_234), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_157), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_157), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_157), .A2(n_517), .B(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_157), .A2(n_529), .B(n_530), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_157), .A2(n_537), .B(n_538), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_157), .A2(n_546), .B(n_547), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_157), .A2(n_559), .B(n_560), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_158), .B(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_158), .B(n_217), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_158), .B(n_220), .Y(n_219) );
NOR3xp33_ASAP7_75t_L g223 ( .A(n_158), .B(n_224), .C(n_225), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_158), .A2(n_526), .B(n_527), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_158), .A2(n_556), .B(n_557), .Y(n_555) );
INVx3_ASAP7_75t_SL g284 ( .A(n_159), .Y(n_284) );
AND2x2_ASAP7_75t_L g328 ( .A(n_159), .B(n_243), .Y(n_328) );
OAI21xp5_ASAP7_75t_L g331 ( .A1(n_159), .A2(n_332), .B(n_333), .Y(n_331) );
AND2x2_ASAP7_75t_L g369 ( .A(n_159), .B(n_307), .Y(n_369) );
AND2x4_ASAP7_75t_L g159 ( .A(n_160), .B(n_170), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_160), .B(n_171), .Y(n_250) );
OR2x2_ASAP7_75t_L g254 ( .A(n_160), .B(n_171), .Y(n_254) );
INVx1_ASAP7_75t_L g262 ( .A(n_160), .Y(n_262) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_160), .Y(n_274) );
INVx2_ASAP7_75t_L g282 ( .A(n_160), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_160), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g391 ( .A(n_160), .B(n_276), .Y(n_391) );
AND2x2_ASAP7_75t_L g406 ( .A(n_160), .B(n_243), .Y(n_406) );
AO21x2_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_167), .B(n_169), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_162), .B(n_166), .Y(n_161) );
AO21x2_ASAP7_75t_L g171 ( .A1(n_167), .A2(n_172), .B(n_178), .Y(n_171) );
AO21x2_ASAP7_75t_L g326 ( .A1(n_167), .A2(n_172), .B(n_178), .Y(n_326) );
AOI21x1_ASAP7_75t_L g505 ( .A1(n_167), .A2(n_506), .B(n_512), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_168), .Y(n_167) );
OA21x2_ASAP7_75t_L g181 ( .A1(n_168), .A2(n_182), .B(n_186), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_168), .A2(n_498), .B(n_499), .Y(n_497) );
AO21x2_ASAP7_75t_L g580 ( .A1(n_168), .A2(n_581), .B(n_582), .Y(n_580) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g275 ( .A(n_171), .B(n_276), .Y(n_275) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_171), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_173), .B(n_177), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_179), .B(n_399), .Y(n_398) );
NOR2x1p5_ASAP7_75t_L g179 ( .A(n_180), .B(n_187), .Y(n_179) );
BUFx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g227 ( .A(n_181), .B(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_181), .B(n_188), .Y(n_257) );
INVx1_ASAP7_75t_L g267 ( .A(n_181), .Y(n_267) );
INVx2_ASAP7_75t_L g290 ( .A(n_181), .Y(n_290) );
INVx2_ASAP7_75t_L g296 ( .A(n_181), .Y(n_296) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_181), .Y(n_366) );
OR2x2_ASAP7_75t_L g397 ( .A(n_181), .B(n_188), .Y(n_397) );
OR2x2_ASAP7_75t_L g413 ( .A(n_187), .B(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x4_ASAP7_75t_SL g201 ( .A(n_188), .B(n_202), .Y(n_201) );
AND2x4_ASAP7_75t_L g239 ( .A(n_188), .B(n_240), .Y(n_239) );
OR2x2_ASAP7_75t_L g277 ( .A(n_188), .B(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g289 ( .A(n_188), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g302 ( .A(n_188), .B(n_268), .Y(n_302) );
OR2x2_ASAP7_75t_L g310 ( .A(n_188), .B(n_202), .Y(n_310) );
INVx2_ASAP7_75t_L g337 ( .A(n_188), .Y(n_337) );
INVx1_ASAP7_75t_L g355 ( .A(n_188), .Y(n_355) );
NOR2xp33_ASAP7_75t_R g388 ( .A(n_188), .B(n_228), .Y(n_388) );
OR2x6_ASAP7_75t_L g188 ( .A(n_189), .B(n_197), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_195), .Y(n_189) );
INVx2_ASAP7_75t_SL g245 ( .A(n_195), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_195), .A2(n_543), .B(n_544), .Y(n_542) );
BUFx4f_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx3_ASAP7_75t_L g222 ( .A(n_196), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_199), .B(n_237), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g279 ( .A1(n_199), .A2(n_280), .B1(n_283), .B2(n_286), .Y(n_279) );
OR2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_226), .Y(n_199) );
INVx1_ASAP7_75t_SL g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g294 ( .A(n_201), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g329 ( .A(n_201), .B(n_330), .Y(n_329) );
AND2x4_ASAP7_75t_L g408 ( .A(n_201), .B(n_386), .Y(n_408) );
INVx3_ASAP7_75t_L g240 ( .A(n_202), .Y(n_240) );
AND2x4_ASAP7_75t_L g268 ( .A(n_202), .B(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_202), .B(n_228), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_202), .B(n_290), .Y(n_335) );
AND2x2_ASAP7_75t_L g340 ( .A(n_202), .B(n_337), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_202), .B(n_227), .Y(n_377) );
INVx1_ASAP7_75t_L g447 ( .A(n_202), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_202), .B(n_365), .Y(n_458) );
AND2x4_ASAP7_75t_L g202 ( .A(n_203), .B(n_218), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_206), .B1(n_211), .B2(n_216), .Y(n_203) );
AND2x4_ASAP7_75t_L g206 ( .A(n_207), .B(n_210), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
NOR2x1p5_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
INVx3_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx3_ASAP7_75t_L g533 ( .A(n_221), .Y(n_533) );
INVx4_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AOI21x1_ASAP7_75t_L g229 ( .A1(n_222), .A2(n_230), .B(n_236), .Y(n_229) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_222), .A2(n_514), .B(n_520), .Y(n_513) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g238 ( .A(n_228), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_228), .B(n_240), .Y(n_258) );
INVx2_ASAP7_75t_L g269 ( .A(n_228), .Y(n_269) );
AND2x2_ASAP7_75t_L g295 ( .A(n_228), .B(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g311 ( .A(n_228), .B(n_290), .Y(n_311) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_228), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_228), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g400 ( .A(n_228), .Y(n_400) );
INVx3_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_235), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_238), .B(n_267), .Y(n_278) );
AOI221x1_ASAP7_75t_SL g372 ( .A1(n_239), .A2(n_373), .B1(n_376), .B2(n_378), .C(n_382), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_239), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g430 ( .A(n_239), .B(n_295), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_239), .B(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g361 ( .A(n_240), .B(n_289), .Y(n_361) );
AND2x2_ASAP7_75t_L g399 ( .A(n_240), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g241 ( .A(n_242), .Y(n_241) );
OR2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_250), .Y(n_242) );
AND2x2_ASAP7_75t_L g252 ( .A(n_243), .B(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g347 ( .A(n_243), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_243), .B(n_263), .Y(n_352) );
AND2x4_ASAP7_75t_L g381 ( .A(n_243), .B(n_282), .Y(n_381) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_243), .B(n_313), .Y(n_417) );
OR2x2_ASAP7_75t_L g435 ( .A(n_243), .B(n_366), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_243), .B(n_326), .Y(n_445) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g276 ( .A(n_244), .Y(n_276) );
AOI21x1_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_246), .B(n_249), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
INVx1_ASAP7_75t_L g301 ( .A(n_250), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g308 ( .A1(n_250), .A2(n_309), .B1(n_312), .B2(n_314), .Y(n_308) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_255), .Y(n_251) );
INVx2_ASAP7_75t_L g264 ( .A(n_252), .Y(n_264) );
AND2x2_ASAP7_75t_L g403 ( .A(n_253), .B(n_263), .Y(n_403) );
AND2x2_ASAP7_75t_L g449 ( .A(n_253), .B(n_316), .Y(n_449) );
AND2x2_ASAP7_75t_L g454 ( .A(n_253), .B(n_305), .Y(n_454) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AOI32xp33_ASAP7_75t_L g423 ( .A1(n_255), .A2(n_325), .A3(n_405), .B1(n_424), .B2(n_426), .Y(n_423) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
INVx1_ASAP7_75t_L g291 ( .A(n_258), .Y(n_291) );
AOI211xp5_ASAP7_75t_SL g259 ( .A1(n_260), .A2(n_265), .B(n_270), .C(n_279), .Y(n_259) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_263), .B(n_264), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_262), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_263), .B(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g443 ( .A(n_263), .Y(n_443) );
AND2x2_ASAP7_75t_L g353 ( .A(n_265), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_SL g265 ( .A(n_266), .B(n_268), .Y(n_265) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_266), .Y(n_453) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVxp67_ASAP7_75t_SL g322 ( .A(n_267), .Y(n_322) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_267), .Y(n_422) );
INVx1_ASAP7_75t_L g319 ( .A(n_268), .Y(n_319) );
AND2x2_ASAP7_75t_L g385 ( .A(n_268), .B(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_268), .B(n_396), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_271), .B(n_277), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OAI21xp33_ASAP7_75t_L g351 ( .A1(n_272), .A2(n_352), .B(n_353), .Y(n_351) );
AND2x2_ASAP7_75t_SL g272 ( .A(n_273), .B(n_275), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g281 ( .A(n_276), .B(n_282), .Y(n_281) );
BUFx2_ASAP7_75t_L g305 ( .A(n_276), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_281), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g412 ( .A(n_281), .Y(n_412) );
AND2x2_ASAP7_75t_L g442 ( .A(n_281), .B(n_443), .Y(n_442) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_282), .Y(n_419) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_284), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_SL g359 ( .A(n_285), .Y(n_359) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x4_ASAP7_75t_L g287 ( .A(n_288), .B(n_291), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g318 ( .A(n_289), .B(n_319), .Y(n_318) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_290), .Y(n_386) );
AND2x2_ASAP7_75t_L g395 ( .A(n_291), .B(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_315), .Y(n_292) );
AOI221xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_297), .B1(n_302), .B2(n_303), .C(n_308), .Y(n_293) );
INVx1_ASAP7_75t_L g414 ( .A(n_295), .Y(n_414) );
INVxp33_ASAP7_75t_SL g446 ( .A(n_295), .Y(n_446) );
AOI21xp5_ASAP7_75t_L g392 ( .A1(n_297), .A2(n_393), .B(n_401), .Y(n_392) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_299), .B(n_301), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_301), .B(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g314 ( .A(n_302), .Y(n_314) );
AND2x2_ASAP7_75t_L g349 ( .A(n_302), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g368 ( .A(n_302), .B(n_369), .Y(n_368) );
AOI22xp33_ASAP7_75t_SL g429 ( .A1(n_302), .A2(n_430), .B1(n_431), .B2(n_434), .Y(n_429) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
OR2x2_ASAP7_75t_L g324 ( .A(n_305), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_305), .B(n_313), .Y(n_363) );
AND2x4_ASAP7_75t_L g380 ( .A(n_307), .B(n_326), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_307), .B(n_381), .Y(n_427) );
AND2x2_ASAP7_75t_L g439 ( .A(n_307), .B(n_391), .Y(n_439) );
NAND2xp33_ASAP7_75t_L g424 ( .A(n_309), .B(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_SL g367 ( .A(n_310), .Y(n_367) );
INVx1_ASAP7_75t_L g438 ( .A(n_311), .Y(n_438) );
INVx2_ASAP7_75t_SL g390 ( .A(n_313), .Y(n_390) );
AOI211xp5_ASAP7_75t_SL g315 ( .A1(n_316), .A2(n_317), .B(n_320), .C(n_338), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OAI211xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_324), .B(n_327), .C(n_331), .Y(n_320) );
OR2x6_ASAP7_75t_SL g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g350 ( .A(n_322), .Y(n_350) );
INVx1_ASAP7_75t_SL g375 ( .A(n_325), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_325), .B(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_330), .B(n_340), .Y(n_339) );
INVx2_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
OAI22xp33_ASAP7_75t_L g416 ( .A1(n_334), .A2(n_417), .B1(n_418), .B2(n_420), .Y(n_416) );
OR2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
OAI211xp5_ASAP7_75t_SL g342 ( .A1(n_343), .A2(n_348), .B(n_351), .C(n_356), .Y(n_342) );
INVxp67_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_345), .B(n_347), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AOI221xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_360), .B1(n_362), .B2(n_364), .C(n_368), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_367), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AOI222xp33_ASAP7_75t_L g448 ( .A1(n_367), .A2(n_449), .B1(n_450), .B2(n_454), .C1(n_455), .C2(n_457), .Y(n_448) );
INVx2_ASAP7_75t_L g383 ( .A(n_369), .Y(n_383) );
NOR3xp33_ASAP7_75t_L g370 ( .A(n_371), .B(n_409), .C(n_428), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_392), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVxp67_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_380), .B(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_381), .B(n_443), .Y(n_456) );
OAI22xp33_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_384), .B1(n_387), .B2(n_389), .Y(n_382) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
INVxp33_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_390), .B(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_398), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_398), .A2(n_402), .B1(n_404), .B2(n_407), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
BUFx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
CKINVDCx16_ASAP7_75t_R g407 ( .A(n_408), .Y(n_407) );
OAI211xp5_ASAP7_75t_SL g409 ( .A1(n_410), .A2(n_413), .B(n_415), .C(n_423), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVxp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NAND3xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_436), .C(n_448), .Y(n_428) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OAI21xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_440), .B(n_447), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
AOI21xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_444), .B(n_446), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVxp33_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_462), .Y(n_461) );
CKINVDCx11_ASAP7_75t_R g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
BUFx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx3_ASAP7_75t_L g477 ( .A(n_470), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
AND2x6_ASAP7_75t_SL g489 ( .A(n_471), .B(n_473), .Y(n_489) );
OR2x6_ASAP7_75t_SL g791 ( .A(n_471), .B(n_472), .Y(n_791) );
OR2x2_ASAP7_75t_L g798 ( .A(n_471), .B(n_473), .Y(n_798) );
CKINVDCx5p33_ASAP7_75t_R g472 ( .A(n_473), .Y(n_472) );
BUFx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_477), .Y(n_476) );
AO221x1_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_485), .B1(n_792), .B2(n_793), .C(n_795), .Y(n_479) );
INVx1_ASAP7_75t_L g792 ( .A(n_480), .Y(n_792) );
CKINVDCx11_ASAP7_75t_R g486 ( .A(n_487), .Y(n_486) );
INVx3_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
CKINVDCx5p33_ASAP7_75t_R g488 ( .A(n_489), .Y(n_488) );
INVx5_ASAP7_75t_L g794 ( .A(n_490), .Y(n_794) );
AND2x4_ASAP7_75t_L g490 ( .A(n_491), .B(n_693), .Y(n_490) );
NOR3xp33_ASAP7_75t_L g491 ( .A(n_492), .B(n_618), .C(n_654), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_592), .Y(n_492) );
AOI211xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_521), .B(n_550), .C(n_575), .Y(n_493) );
AND2x2_ASAP7_75t_L g683 ( .A(n_494), .B(n_552), .Y(n_683) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_504), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_495), .B(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g716 ( .A(n_495), .B(n_598), .Y(n_716) );
AND2x2_ASAP7_75t_L g732 ( .A(n_495), .B(n_567), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_495), .B(n_742), .Y(n_741) );
NAND2x1p5_ASAP7_75t_L g765 ( .A(n_495), .B(n_766), .Y(n_765) );
INVx4_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x4_ASAP7_75t_SL g562 ( .A(n_496), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g587 ( .A(n_496), .Y(n_587) );
AND2x2_ASAP7_75t_L g634 ( .A(n_496), .B(n_577), .Y(n_634) );
AND2x2_ASAP7_75t_L g653 ( .A(n_496), .B(n_504), .Y(n_653) );
BUFx2_ASAP7_75t_L g658 ( .A(n_496), .Y(n_658) );
AND2x2_ASAP7_75t_L g702 ( .A(n_496), .B(n_513), .Y(n_702) );
AND2x4_ASAP7_75t_L g774 ( .A(n_496), .B(n_775), .Y(n_774) );
NOR2x1_ASAP7_75t_L g786 ( .A(n_496), .B(n_566), .Y(n_786) );
OR2x6_ASAP7_75t_L g496 ( .A(n_497), .B(n_503), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_504), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g705 ( .A(n_504), .Y(n_705) );
BUFx2_ASAP7_75t_L g754 ( .A(n_504), .Y(n_754) );
INVx1_ASAP7_75t_L g776 ( .A(n_504), .Y(n_776) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_513), .Y(n_504) );
INVx3_ASAP7_75t_L g563 ( .A(n_505), .Y(n_563) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_505), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_511), .Y(n_506) );
INVx2_ASAP7_75t_L g566 ( .A(n_513), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_513), .B(n_563), .Y(n_567) );
INVx2_ASAP7_75t_L g642 ( .A(n_513), .Y(n_642) );
OR2x2_ASAP7_75t_L g649 ( .A(n_513), .B(n_598), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_519), .Y(n_514) );
AND2x2_ASAP7_75t_L g604 ( .A(n_521), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g638 ( .A(n_521), .B(n_601), .Y(n_638) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_531), .Y(n_521) );
AND2x2_ASAP7_75t_L g674 ( .A(n_522), .B(n_573), .Y(n_674) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g631 ( .A(n_523), .B(n_532), .Y(n_631) );
AND2x2_ASAP7_75t_L g750 ( .A(n_523), .B(n_541), .Y(n_750) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g572 ( .A(n_524), .Y(n_572) );
INVx1_ASAP7_75t_L g590 ( .A(n_524), .Y(n_590) );
AND2x2_ASAP7_75t_L g646 ( .A(n_524), .B(n_532), .Y(n_646) );
AND2x2_ASAP7_75t_L g651 ( .A(n_524), .B(n_553), .Y(n_651) );
OR2x2_ASAP7_75t_L g714 ( .A(n_524), .B(n_541), .Y(n_714) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_524), .Y(n_723) );
AND2x2_ASAP7_75t_L g552 ( .A(n_531), .B(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g591 ( .A(n_531), .Y(n_591) );
NOR2x1_ASAP7_75t_SL g531 ( .A(n_532), .B(n_541), .Y(n_531) );
AO21x1_ASAP7_75t_SL g532 ( .A1(n_533), .A2(n_534), .B(n_540), .Y(n_532) );
AO21x2_ASAP7_75t_L g574 ( .A1(n_533), .A2(n_534), .B(n_540), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_539), .Y(n_534) );
AND2x2_ASAP7_75t_L g569 ( .A(n_541), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_SL g617 ( .A(n_541), .Y(n_617) );
NAND2x1_ASAP7_75t_L g627 ( .A(n_541), .B(n_553), .Y(n_627) );
OR2x2_ASAP7_75t_L g632 ( .A(n_541), .B(n_570), .Y(n_632) );
BUFx2_ASAP7_75t_L g688 ( .A(n_541), .Y(n_688) );
AND2x2_ASAP7_75t_L g724 ( .A(n_541), .B(n_603), .Y(n_724) );
AND2x2_ASAP7_75t_L g735 ( .A(n_541), .B(n_573), .Y(n_735) );
OR2x6_ASAP7_75t_L g541 ( .A(n_542), .B(n_549), .Y(n_541) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_561), .B1(n_567), .B2(n_568), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g781 ( .A1(n_552), .A2(n_732), .B1(n_782), .B2(n_787), .Y(n_781) );
INVx4_ASAP7_75t_L g570 ( .A(n_553), .Y(n_570) );
INVx2_ASAP7_75t_L g601 ( .A(n_553), .Y(n_601) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_553), .Y(n_672) );
OR2x2_ASAP7_75t_L g687 ( .A(n_553), .B(n_573), .Y(n_687) );
OR2x2_ASAP7_75t_SL g713 ( .A(n_553), .B(n_714), .Y(n_713) );
OR2x6_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
AND2x2_ASAP7_75t_SL g561 ( .A(n_562), .B(n_564), .Y(n_561) );
INVx2_ASAP7_75t_SL g594 ( .A(n_562), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_562), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g662 ( .A(n_562), .B(n_610), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_562), .B(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g584 ( .A(n_563), .Y(n_584) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_563), .Y(n_609) );
AND2x2_ASAP7_75t_L g665 ( .A(n_563), .B(n_642), .Y(n_665) );
INVx1_ASAP7_75t_L g775 ( .A(n_563), .Y(n_775) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_565), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_565), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g583 ( .A(n_566), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_567), .B(n_716), .Y(n_715) );
AOI321xp33_ASAP7_75t_L g737 ( .A1(n_568), .A2(n_639), .A3(n_707), .B1(n_738), .B2(n_739), .C(n_743), .Y(n_737) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
INVxp67_ASAP7_75t_SL g636 ( .A(n_569), .Y(n_636) );
AND2x2_ASAP7_75t_L g661 ( .A(n_569), .B(n_590), .Y(n_661) );
AND2x2_ASAP7_75t_L g736 ( .A(n_569), .B(n_646), .Y(n_736) );
INVx1_ASAP7_75t_L g605 ( .A(n_570), .Y(n_605) );
BUFx2_ASAP7_75t_L g615 ( .A(n_570), .Y(n_615) );
NOR2xp67_ASAP7_75t_L g722 ( .A(n_570), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_SL g660 ( .A(n_571), .Y(n_660) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
BUFx2_ASAP7_75t_L g667 ( .A(n_572), .Y(n_667) );
INVx2_ASAP7_75t_L g603 ( .A(n_573), .Y(n_603) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_573), .Y(n_626) );
INVx3_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AOI21xp33_ASAP7_75t_SL g575 ( .A1(n_576), .A2(n_585), .B(n_588), .Y(n_575) );
NOR2xp67_ASAP7_75t_L g719 ( .A(n_576), .B(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_583), .Y(n_577) );
INVx3_ASAP7_75t_L g610 ( .A(n_578), .Y(n_610) );
AND2x2_ASAP7_75t_L g641 ( .A(n_578), .B(n_642), .Y(n_641) );
AND2x4_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
AND2x4_ASAP7_75t_L g598 ( .A(n_579), .B(n_580), .Y(n_598) );
INVx1_ASAP7_75t_L g681 ( .A(n_583), .Y(n_681) );
INVx1_ASAP7_75t_SL g766 ( .A(n_584), .Y(n_766) );
INVxp33_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_587), .B(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g692 ( .A(n_587), .B(n_649), .Y(n_692) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_591), .Y(n_588) );
AND2x2_ASAP7_75t_L g696 ( .A(n_589), .B(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_589), .B(n_711), .Y(n_710) );
INVx3_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_590), .B(n_627), .Y(n_682) );
NOR4xp25_ASAP7_75t_L g777 ( .A(n_590), .B(n_621), .C(n_778), .D(n_779), .Y(n_777) );
OR2x2_ASAP7_75t_L g745 ( .A(n_591), .B(n_746), .Y(n_745) );
AOI221xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_599), .B1(n_604), .B2(n_606), .C(n_611), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
AND2x2_ASAP7_75t_L g620 ( .A(n_595), .B(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g657 ( .A(n_596), .B(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g677 ( .A(n_597), .Y(n_677) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
BUFx3_ASAP7_75t_L g700 ( .A(n_598), .Y(n_700) );
AND2x2_ASAP7_75t_L g707 ( .A(n_598), .B(n_708), .Y(n_707) );
INVxp67_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
OR2x2_ASAP7_75t_L g644 ( .A(n_601), .B(n_645), .Y(n_644) );
INVxp67_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_603), .B(n_617), .Y(n_616) );
INVxp67_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_610), .Y(n_607) );
INVx2_ASAP7_75t_L g621 ( .A(n_608), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_608), .B(n_691), .Y(n_690) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g613 ( .A(n_610), .Y(n_613) );
OAI321xp33_ASAP7_75t_L g725 ( .A1(n_610), .A2(n_718), .A3(n_726), .B1(n_731), .B2(n_733), .C(n_737), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
OR2x2_ASAP7_75t_L g680 ( .A(n_613), .B(n_681), .Y(n_680) );
OR2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
INVx1_ASAP7_75t_L g780 ( .A(n_616), .Y(n_780) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_617), .B(n_660), .Y(n_659) );
NAND2xp33_ASAP7_75t_SL g760 ( .A(n_617), .B(n_631), .Y(n_760) );
OAI211xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_622), .B(n_633), .C(n_637), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NOR2x1_ASAP7_75t_L g622 ( .A(n_623), .B(n_628), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g729 ( .A(n_626), .Y(n_729) );
INVx3_ASAP7_75t_L g668 ( .A(n_627), .Y(n_668) );
OR2x2_ASAP7_75t_L g771 ( .A(n_627), .B(n_645), .Y(n_771) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_629), .A2(n_713), .B1(n_715), .B2(n_717), .Y(n_712) );
OR2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_SL g711 ( .A(n_632), .Y(n_711) );
OR2x2_ASAP7_75t_L g788 ( .A(n_632), .B(n_645), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AOI21xp5_ASAP7_75t_SL g637 ( .A1(n_638), .A2(n_639), .B(n_643), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_641), .B(n_658), .Y(n_757) );
AND2x2_ASAP7_75t_L g763 ( .A(n_641), .B(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g708 ( .A(n_642), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_647), .B1(n_650), .B2(n_652), .Y(n_643) );
A2O1A1Ixp33_ASAP7_75t_L g689 ( .A1(n_645), .A2(n_688), .B(n_690), .C(n_692), .Y(n_689) );
INVx2_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_648), .B(n_718), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_648), .B(n_740), .Y(n_762) );
INVx2_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g734 ( .A(n_651), .B(n_735), .Y(n_734) );
INVx2_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
A2O1A1Ixp33_ASAP7_75t_L g684 ( .A1(n_653), .A2(n_685), .B(n_688), .C(n_689), .Y(n_684) );
NAND3xp33_ASAP7_75t_SL g654 ( .A(n_655), .B(n_669), .C(n_684), .Y(n_654) );
AOI222xp33_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_659), .B1(n_661), .B2(n_662), .C1(n_663), .C2(n_666), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g718 ( .A(n_658), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_658), .B(n_691), .Y(n_744) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_SL g678 ( .A(n_665), .Y(n_678) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
OR2x2_ASAP7_75t_L g783 ( .A(n_667), .B(n_700), .Y(n_783) );
AOI22xp5_ASAP7_75t_L g758 ( .A1(n_668), .A2(n_759), .B1(n_761), .B2(n_763), .Y(n_758) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_675), .B1(n_679), .B2(n_682), .C(n_683), .Y(n_669) );
INVx2_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
OR2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AOI21xp5_ASAP7_75t_SL g743 ( .A1(n_676), .A2(n_744), .B(n_745), .Y(n_743) );
OR2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
INVx2_ASAP7_75t_L g691 ( .A(n_677), .Y(n_691) );
AND2x2_ASAP7_75t_L g785 ( .A(n_677), .B(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g769 ( .A(n_681), .Y(n_769) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
OR2x2_ASAP7_75t_L g698 ( .A(n_687), .B(n_688), .Y(n_698) );
INVx1_ASAP7_75t_L g751 ( .A(n_687), .Y(n_751) );
NOR3xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_725), .C(n_747), .Y(n_693) );
OAI211xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_699), .B(n_701), .C(n_706), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
OAI21xp33_ASAP7_75t_L g701 ( .A1(n_696), .A2(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AOI211xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_709), .B(n_712), .C(n_719), .Y(n_706) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g730 ( .A(n_713), .Y(n_730) );
INVxp67_ASAP7_75t_SL g755 ( .A(n_714), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_716), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g778 ( .A(n_716), .Y(n_778) );
AND2x2_ASAP7_75t_L g768 ( .A(n_718), .B(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g738 ( .A(n_720), .Y(n_738) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_724), .Y(n_721) );
INVx1_ASAP7_75t_L g746 ( .A(n_722), .Y(n_746) );
INVx2_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
AND2x4_ASAP7_75t_L g727 ( .A(n_728), .B(n_730), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_736), .Y(n_733) );
AOI221xp5_ASAP7_75t_L g767 ( .A1(n_734), .A2(n_768), .B1(n_770), .B2(n_772), .C(n_777), .Y(n_767) );
OAI21xp33_ASAP7_75t_SL g782 ( .A1(n_739), .A2(n_783), .B(n_784), .Y(n_782) );
INVx2_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
NAND4xp25_ASAP7_75t_L g747 ( .A(n_748), .B(n_758), .C(n_767), .D(n_781), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_752), .B1(n_755), .B2(n_756), .Y(n_748) );
AND2x4_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVxp67_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_773), .B(n_776), .Y(n_772) );
INVx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_SL g789 ( .A(n_790), .Y(n_789) );
CKINVDCx11_ASAP7_75t_R g790 ( .A(n_791), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .Y(n_795) );
BUFx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
NOR2xp33_ASAP7_75t_L g799 ( .A(n_800), .B(n_801), .Y(n_799) );
endmodule