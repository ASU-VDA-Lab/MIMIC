module fake_jpeg_27160_n_271 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_271);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_271;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_15),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_21),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_38),
.B(n_18),
.C(n_20),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_0),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_35),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_44),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_0),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_57),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_45),
.A2(n_24),
.B1(n_32),
.B2(n_18),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_65),
.B1(n_39),
.B2(n_46),
.Y(n_75)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_37),
.B1(n_38),
.B2(n_32),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_51),
.A2(n_52),
.B1(n_57),
.B2(n_42),
.Y(n_81)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_26),
.B(n_24),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_19),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_20),
.B1(n_34),
.B2(n_33),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_46),
.B1(n_40),
.B2(n_39),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_28),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_37),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_36),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_66),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_35),
.B1(n_34),
.B2(n_33),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_31),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_73),
.A2(n_76),
.B1(n_78),
.B2(n_86),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_85),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_75),
.A2(n_84),
.B1(n_61),
.B2(n_68),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_62),
.A2(n_43),
.B1(n_28),
.B2(n_34),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_28),
.B1(n_22),
.B2(n_33),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_81),
.B(n_91),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_55),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_53),
.A2(n_43),
.B1(n_42),
.B2(n_27),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_52),
.B(n_2),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_27),
.B1(n_22),
.B2(n_19),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_59),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_89),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_59),
.A2(n_26),
.B1(n_27),
.B2(n_22),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_88),
.Y(n_108)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_69),
.B(n_66),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_31),
.B1(n_3),
.B2(n_4),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_61),
.B1(n_55),
.B2(n_64),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_49),
.Y(n_102)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g118 ( 
.A1(n_94),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_56),
.C(n_47),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_100),
.Y(n_130)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_99),
.B(n_102),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_100),
.A2(n_79),
.B(n_71),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_101),
.A2(n_106),
.B1(n_94),
.B2(n_80),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_49),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_107),
.Y(n_134)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_111),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_93),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_105),
.Y(n_131)
);

AO21x2_ASAP7_75t_L g106 ( 
.A1(n_73),
.A2(n_61),
.B(n_50),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_49),
.Y(n_107)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_2),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_112),
.Y(n_136)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_117),
.Y(n_137)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_115),
.A2(n_94),
.B1(n_80),
.B2(n_71),
.Y(n_127)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

OA21x2_ASAP7_75t_L g125 ( 
.A1(n_118),
.A2(n_92),
.B(n_79),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_4),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_95),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_117),
.A2(n_91),
.B1(n_88),
.B2(n_87),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_126),
.B1(n_140),
.B2(n_106),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_SL g146 ( 
.A1(n_125),
.A2(n_108),
.B(n_106),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_113),
.A2(n_91),
.B1(n_78),
.B2(n_80),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_127),
.A2(n_141),
.B1(n_106),
.B2(n_111),
.Y(n_147)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_133),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_129),
.A2(n_118),
.B(n_72),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_138),
.Y(n_169)
);

NOR2x1_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_103),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_139),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_95),
.B(n_6),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_97),
.A2(n_72),
.B1(n_83),
.B2(n_8),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_105),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_131),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_98),
.B(n_72),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_144),
.Y(n_165)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_145),
.A2(n_157),
.B1(n_164),
.B2(n_167),
.Y(n_185)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_147),
.B(n_168),
.Y(n_190)
);

XOR2x2_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_106),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_L g179 ( 
.A1(n_148),
.A2(n_162),
.B(n_136),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_133),
.A2(n_108),
.B(n_104),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_149),
.A2(n_155),
.B(n_158),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_96),
.C(n_99),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_152),
.C(n_170),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_96),
.C(n_110),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_154),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_132),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_119),
.B(n_118),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_140),
.A2(n_97),
.B1(n_115),
.B2(n_118),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_118),
.B(n_114),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_124),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_142),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_161),
.B(n_163),
.Y(n_188)
);

XOR2x2_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_6),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_114),
.B1(n_109),
.B2(n_8),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_137),
.A2(n_109),
.B(n_7),
.Y(n_166)
);

MAJx2_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_136),
.C(n_125),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_126),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_137),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_16),
.C(n_10),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_123),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_174),
.Y(n_201)
);

INVxp67_ASAP7_75t_SL g175 ( 
.A(n_151),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_187),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_123),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_181),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_151),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_178),
.Y(n_213)
);

XNOR2x1_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_193),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_128),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_182),
.B(n_183),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_166),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_135),
.C(n_132),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_169),
.Y(n_202)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_156),
.Y(n_189)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_189),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_149),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_191),
.A2(n_125),
.B(n_127),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_120),
.Y(n_192)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_188),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_204),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_197),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_185),
.A2(n_147),
.B1(n_145),
.B2(n_157),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_198),
.A2(n_200),
.B1(n_190),
.B2(n_171),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_185),
.A2(n_162),
.B1(n_158),
.B2(n_159),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_206),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_187),
.A2(n_156),
.B1(n_141),
.B2(n_155),
.Y(n_204)
);

NOR2x1_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_167),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_205),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_150),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_207),
.A2(n_186),
.B(n_191),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_152),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_173),
.C(n_193),
.Y(n_214)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_212),
.B(n_172),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_225),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_221),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_218),
.B(n_219),
.Y(n_232)
);

BUFx12_ASAP7_75t_L g219 ( 
.A(n_209),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_196),
.B(n_181),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_224),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_200),
.A2(n_186),
.B(n_191),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_229),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_223),
.A2(n_228),
.B1(n_227),
.B2(n_221),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_201),
.B(n_208),
.Y(n_224)
);

AOI221xp5_ASAP7_75t_L g225 ( 
.A1(n_209),
.A2(n_183),
.B1(n_193),
.B2(n_178),
.C(n_171),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_198),
.A2(n_190),
.B1(n_182),
.B2(n_189),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_211),
.B(n_170),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_226),
.C(n_217),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_237),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_217),
.A2(n_204),
.B1(n_213),
.B2(n_206),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_9),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_202),
.C(n_173),
.Y(n_237)
);

AOI21x1_ASAP7_75t_SL g238 ( 
.A1(n_227),
.A2(n_205),
.B(n_199),
.Y(n_238)
);

XOR2x1_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_219),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_210),
.C(n_194),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_240),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_203),
.C(n_120),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_241),
.A2(n_223),
.B1(n_228),
.B2(n_215),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_242),
.A2(n_234),
.B1(n_240),
.B2(n_232),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_243),
.Y(n_253)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_235),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_238),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_222),
.C(n_219),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_246),
.B(n_248),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_125),
.C(n_138),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_233),
.B(n_144),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_15),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_250),
.A2(n_231),
.B(n_10),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_255),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_254),
.Y(n_259)
);

BUFx24_ASAP7_75t_SL g255 ( 
.A(n_247),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_257),
.C(n_249),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_257),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_261),
.Y(n_266)
);

NOR2xp67_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_243),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_260),
.A2(n_253),
.B(n_244),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_262),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_263),
.A2(n_259),
.B1(n_13),
.B2(n_14),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_265),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_259),
.A2(n_9),
.B(n_12),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_13),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_266),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_267),
.Y(n_271)
);


endmodule