module real_aes_7413_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_725;
wire n_119;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_505;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g177 ( .A1(n_0), .A2(n_178), .B(n_181), .C(n_185), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_1), .B(n_169), .Y(n_188) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_2), .B(n_109), .C(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g450 ( .A(n_2), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_3), .B(n_179), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_4), .A2(n_138), .B(n_499), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_5), .A2(n_143), .B(n_146), .C(n_526), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_6), .A2(n_138), .B(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_7), .B(n_169), .Y(n_505) );
AO21x2_ASAP7_75t_L g245 ( .A1(n_8), .A2(n_171), .B(n_246), .Y(n_245) );
AND2x6_ASAP7_75t_L g143 ( .A(n_9), .B(n_144), .Y(n_143) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_10), .A2(n_143), .B(n_146), .C(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g539 ( .A(n_11), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_12), .B(n_41), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_13), .B(n_184), .Y(n_528) );
INVx1_ASAP7_75t_L g164 ( .A(n_14), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_15), .B(n_179), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_L g558 ( .A1(n_16), .A2(n_180), .B(n_559), .C(n_561), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_17), .B(n_169), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_18), .B(n_158), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_L g145 ( .A1(n_19), .A2(n_146), .B(n_149), .C(n_157), .Y(n_145) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_20), .A2(n_183), .B(n_239), .C(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_21), .B(n_184), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_22), .A2(n_40), .B1(n_728), .B2(n_729), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_22), .Y(n_729) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_23), .B(n_184), .Y(n_513) );
CKINVDCx16_ASAP7_75t_R g473 ( .A(n_24), .Y(n_473) );
INVx1_ASAP7_75t_L g512 ( .A(n_25), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_26), .A2(n_146), .B(n_157), .C(n_249), .Y(n_248) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_27), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_28), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_29), .A2(n_78), .B1(n_126), .B2(n_127), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_29), .Y(n_127) );
INVx1_ASAP7_75t_L g490 ( .A(n_30), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_31), .A2(n_138), .B(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g141 ( .A(n_32), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_33), .A2(n_197), .B(n_198), .C(n_202), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_34), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_35), .A2(n_183), .B(n_502), .C(n_504), .Y(n_501) );
INVxp67_ASAP7_75t_L g491 ( .A(n_36), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_37), .B(n_251), .Y(n_250) );
CKINVDCx14_ASAP7_75t_R g500 ( .A(n_38), .Y(n_500) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_39), .A2(n_146), .B(n_157), .C(n_511), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_40), .Y(n_728) );
A2O1A1Ixp33_ASAP7_75t_L g536 ( .A1(n_42), .A2(n_185), .B(n_537), .C(n_538), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_43), .B(n_137), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_44), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_45), .B(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_46), .B(n_179), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_47), .B(n_138), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_48), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_49), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_50), .A2(n_197), .B(n_202), .C(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g182 ( .A(n_51), .Y(n_182) );
INVx1_ASAP7_75t_L g225 ( .A(n_52), .Y(n_225) );
INVx1_ASAP7_75t_L g545 ( .A(n_53), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_54), .B(n_138), .Y(n_222) );
AOI222xp33_ASAP7_75t_L g456 ( .A1(n_55), .A2(n_457), .B1(n_723), .B2(n_724), .C1(n_730), .C2(n_735), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_56), .Y(n_166) );
CKINVDCx14_ASAP7_75t_R g535 ( .A(n_57), .Y(n_535) );
INVx1_ASAP7_75t_L g144 ( .A(n_58), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_59), .B(n_138), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_60), .B(n_169), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_61), .A2(n_156), .B(n_212), .C(n_214), .Y(n_211) );
INVx1_ASAP7_75t_L g163 ( .A(n_62), .Y(n_163) );
INVx1_ASAP7_75t_SL g503 ( .A(n_63), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_64), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_65), .B(n_179), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_66), .B(n_169), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_67), .B(n_180), .Y(n_236) );
INVx1_ASAP7_75t_L g476 ( .A(n_68), .Y(n_476) );
CKINVDCx16_ASAP7_75t_R g175 ( .A(n_69), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_70), .B(n_151), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_71), .A2(n_146), .B(n_202), .C(n_265), .Y(n_264) );
CKINVDCx16_ASAP7_75t_R g210 ( .A(n_72), .Y(n_210) );
INVx1_ASAP7_75t_L g112 ( .A(n_73), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_74), .A2(n_138), .B(n_534), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_75), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_76), .A2(n_138), .B(n_556), .Y(n_555) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_77), .A2(n_124), .B1(n_125), .B2(n_128), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_77), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_78), .Y(n_126) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_79), .A2(n_137), .B(n_486), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g509 ( .A(n_80), .Y(n_509) );
INVx1_ASAP7_75t_L g557 ( .A(n_81), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_82), .B(n_154), .Y(n_153) );
AOI22xp5_ASAP7_75t_L g724 ( .A1(n_83), .A2(n_725), .B1(n_726), .B2(n_727), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_83), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_84), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_85), .A2(n_138), .B(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g560 ( .A(n_86), .Y(n_560) );
INVx2_ASAP7_75t_L g161 ( .A(n_87), .Y(n_161) );
INVx1_ASAP7_75t_L g527 ( .A(n_88), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_89), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_90), .B(n_184), .Y(n_237) );
INVx2_ASAP7_75t_L g109 ( .A(n_91), .Y(n_109) );
OR2x2_ASAP7_75t_L g447 ( .A(n_91), .B(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_L g460 ( .A(n_91), .B(n_449), .Y(n_460) );
A2O1A1Ixp33_ASAP7_75t_L g474 ( .A1(n_92), .A2(n_146), .B(n_202), .C(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_93), .B(n_138), .Y(n_195) );
INVx1_ASAP7_75t_L g199 ( .A(n_94), .Y(n_199) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_95), .A2(n_104), .B1(n_105), .B2(n_115), .Y(n_103) );
INVxp67_ASAP7_75t_L g215 ( .A(n_96), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_97), .B(n_171), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_98), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g232 ( .A(n_99), .Y(n_232) );
INVx1_ASAP7_75t_L g266 ( .A(n_100), .Y(n_266) );
INVx2_ASAP7_75t_L g548 ( .A(n_101), .Y(n_548) );
AND2x2_ASAP7_75t_L g227 ( .A(n_102), .B(n_160), .Y(n_227) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
OR2x2_ASAP7_75t_SL g107 ( .A(n_108), .B(n_113), .Y(n_107) );
OR2x2_ASAP7_75t_L g461 ( .A(n_109), .B(n_449), .Y(n_461) );
NOR2x2_ASAP7_75t_L g737 ( .A(n_109), .B(n_448), .Y(n_737) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
INVxp67_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x2_ASAP7_75t_L g449 ( .A(n_114), .B(n_450), .Y(n_449) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_455), .Y(n_115) );
BUFx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
NAND3xp33_ASAP7_75t_L g455 ( .A(n_117), .B(n_451), .C(n_456), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_444), .B(n_451), .Y(n_121) );
AOI22xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_129), .B1(n_442), .B2(n_443), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_123), .Y(n_442) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g443 ( .A(n_129), .Y(n_443) );
OAI22xp5_ASAP7_75t_SL g730 ( .A1(n_129), .A2(n_731), .B1(n_732), .B2(n_733), .Y(n_730) );
AND2x2_ASAP7_75t_SL g129 ( .A(n_130), .B(n_378), .Y(n_129) );
NOR5xp2_ASAP7_75t_L g130 ( .A(n_131), .B(n_309), .C(n_338), .D(n_358), .E(n_365), .Y(n_130) );
OAI211xp5_ASAP7_75t_SL g131 ( .A1(n_132), .A2(n_189), .B(n_253), .C(n_296), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_133), .A2(n_381), .B1(n_383), .B2(n_384), .Y(n_380) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_168), .Y(n_133) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_134), .Y(n_256) );
AND2x4_ASAP7_75t_L g289 ( .A(n_134), .B(n_290), .Y(n_289) );
INVx5_ASAP7_75t_L g307 ( .A(n_134), .Y(n_307) );
AND2x2_ASAP7_75t_L g316 ( .A(n_134), .B(n_308), .Y(n_316) );
AND2x2_ASAP7_75t_L g328 ( .A(n_134), .B(n_193), .Y(n_328) );
AND2x2_ASAP7_75t_L g424 ( .A(n_134), .B(n_292), .Y(n_424) );
OR2x6_ASAP7_75t_L g134 ( .A(n_135), .B(n_165), .Y(n_134) );
AOI21xp5_ASAP7_75t_SL g135 ( .A1(n_136), .A2(n_145), .B(n_158), .Y(n_135) );
BUFx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_143), .Y(n_138) );
NAND2x1p5_ASAP7_75t_L g233 ( .A(n_139), .B(n_143), .Y(n_233) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
INVx1_ASAP7_75t_L g156 ( .A(n_140), .Y(n_156) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g147 ( .A(n_141), .Y(n_147) );
INVx1_ASAP7_75t_L g240 ( .A(n_141), .Y(n_240) );
INVx1_ASAP7_75t_L g148 ( .A(n_142), .Y(n_148) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_142), .Y(n_152) );
INVx3_ASAP7_75t_L g180 ( .A(n_142), .Y(n_180) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_142), .Y(n_184) );
INVx1_ASAP7_75t_L g251 ( .A(n_142), .Y(n_251) );
BUFx3_ASAP7_75t_L g157 ( .A(n_143), .Y(n_157) );
INVx4_ASAP7_75t_SL g187 ( .A(n_143), .Y(n_187) );
INVx5_ASAP7_75t_L g176 ( .A(n_146), .Y(n_176) );
AND2x6_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
BUFx3_ASAP7_75t_L g186 ( .A(n_147), .Y(n_186) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_147), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_153), .B(n_155), .Y(n_149) );
INVx2_ASAP7_75t_L g154 ( .A(n_151), .Y(n_154) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx4_ASAP7_75t_L g213 ( .A(n_152), .Y(n_213) );
O2A1O1Ixp33_ASAP7_75t_L g198 ( .A1(n_154), .A2(n_199), .B(n_200), .C(n_201), .Y(n_198) );
O2A1O1Ixp33_ASAP7_75t_L g224 ( .A1(n_154), .A2(n_201), .B(n_225), .C(n_226), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_154), .A2(n_476), .B(n_477), .C(n_478), .Y(n_475) );
O2A1O1Ixp5_ASAP7_75t_L g526 ( .A1(n_154), .A2(n_478), .B(n_527), .C(n_528), .Y(n_526) );
O2A1O1Ixp33_ASAP7_75t_L g511 ( .A1(n_155), .A2(n_179), .B(n_512), .C(n_513), .Y(n_511) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_156), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_159), .B(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g167 ( .A(n_160), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_160), .A2(n_195), .B(n_196), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_160), .A2(n_222), .B(n_223), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_160), .A2(n_233), .B(n_509), .C(n_510), .Y(n_508) );
OA21x2_ASAP7_75t_L g532 ( .A1(n_160), .A2(n_533), .B(n_540), .Y(n_532) );
AND2x2_ASAP7_75t_SL g160 ( .A(n_161), .B(n_162), .Y(n_160) );
AND2x2_ASAP7_75t_L g172 ( .A(n_161), .B(n_162), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
AO21x2_ASAP7_75t_L g522 ( .A1(n_167), .A2(n_523), .B(n_529), .Y(n_522) );
INVx2_ASAP7_75t_L g290 ( .A(n_168), .Y(n_290) );
AND2x2_ASAP7_75t_L g308 ( .A(n_168), .B(n_262), .Y(n_308) );
AND2x2_ASAP7_75t_L g327 ( .A(n_168), .B(n_261), .Y(n_327) );
AND2x2_ASAP7_75t_L g367 ( .A(n_168), .B(n_307), .Y(n_367) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_173), .B(n_188), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_170), .B(n_204), .Y(n_203) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_170), .A2(n_231), .B(n_241), .Y(n_230) );
AO21x2_ASAP7_75t_L g262 ( .A1(n_170), .A2(n_263), .B(n_271), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_170), .B(n_272), .Y(n_271) );
AO21x2_ASAP7_75t_L g471 ( .A1(n_170), .A2(n_472), .B(n_479), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_170), .B(n_515), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_170), .B(n_530), .Y(n_529) );
INVx4_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_171), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_171), .A2(n_247), .B(n_248), .Y(n_246) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g243 ( .A(n_172), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_SL g174 ( .A1(n_175), .A2(n_176), .B(n_177), .C(n_187), .Y(n_174) );
INVx2_ASAP7_75t_L g197 ( .A(n_176), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_L g209 ( .A1(n_176), .A2(n_187), .B(n_210), .C(n_211), .Y(n_209) );
O2A1O1Ixp33_ASAP7_75t_SL g486 ( .A1(n_176), .A2(n_187), .B(n_487), .C(n_488), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_L g499 ( .A1(n_176), .A2(n_187), .B(n_500), .C(n_501), .Y(n_499) );
O2A1O1Ixp33_ASAP7_75t_SL g534 ( .A1(n_176), .A2(n_187), .B(n_535), .C(n_536), .Y(n_534) );
O2A1O1Ixp33_ASAP7_75t_SL g544 ( .A1(n_176), .A2(n_187), .B(n_545), .C(n_546), .Y(n_544) );
O2A1O1Ixp33_ASAP7_75t_SL g556 ( .A1(n_176), .A2(n_187), .B(n_557), .C(n_558), .Y(n_556) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_179), .B(n_215), .Y(n_214) );
OAI22xp33_ASAP7_75t_L g489 ( .A1(n_179), .A2(n_213), .B1(n_490), .B2(n_491), .Y(n_489) );
INVx5_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_180), .B(n_539), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_183), .B(n_503), .Y(n_502) );
INVx4_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g537 ( .A(n_184), .Y(n_537) );
INVx2_ASAP7_75t_L g478 ( .A(n_185), .Y(n_478) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_186), .Y(n_201) );
INVx1_ASAP7_75t_L g561 ( .A(n_186), .Y(n_561) );
INVx1_ASAP7_75t_L g202 ( .A(n_187), .Y(n_202) );
INVxp67_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_191), .B(n_217), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AOI322xp5_ASAP7_75t_L g426 ( .A1(n_192), .A2(n_228), .A3(n_281), .B1(n_289), .B2(n_343), .C1(n_427), .C2(n_430), .Y(n_426) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_205), .Y(n_192) );
INVx5_ASAP7_75t_L g258 ( .A(n_193), .Y(n_258) );
AND2x2_ASAP7_75t_L g275 ( .A(n_193), .B(n_260), .Y(n_275) );
BUFx2_ASAP7_75t_L g353 ( .A(n_193), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_193), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g430 ( .A(n_193), .B(n_337), .Y(n_430) );
OR2x6_ASAP7_75t_L g193 ( .A(n_194), .B(n_203), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_205), .B(n_219), .Y(n_284) );
INVx1_ASAP7_75t_L g311 ( .A(n_205), .Y(n_311) );
AND2x2_ASAP7_75t_L g324 ( .A(n_205), .B(n_244), .Y(n_324) );
AND2x2_ASAP7_75t_L g425 ( .A(n_205), .B(n_343), .Y(n_425) );
INVx3_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
OR2x2_ASAP7_75t_L g279 ( .A(n_206), .B(n_219), .Y(n_279) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_206), .Y(n_287) );
OR2x2_ASAP7_75t_L g294 ( .A(n_206), .B(n_244), .Y(n_294) );
AND2x2_ASAP7_75t_L g304 ( .A(n_206), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_206), .B(n_230), .Y(n_333) );
INVxp67_ASAP7_75t_L g357 ( .A(n_206), .Y(n_357) );
AND2x2_ASAP7_75t_L g364 ( .A(n_206), .B(n_228), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_206), .B(n_244), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_206), .B(n_229), .Y(n_390) );
OA21x2_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B(n_216), .Y(n_206) );
OA21x2_ASAP7_75t_L g497 ( .A1(n_207), .A2(n_498), .B(n_505), .Y(n_497) );
OA21x2_ASAP7_75t_L g542 ( .A1(n_207), .A2(n_543), .B(n_549), .Y(n_542) );
OA21x2_ASAP7_75t_L g554 ( .A1(n_207), .A2(n_555), .B(n_562), .Y(n_554) );
O2A1O1Ixp33_ASAP7_75t_L g265 ( .A1(n_212), .A2(n_266), .B(n_267), .C(n_268), .Y(n_265) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_213), .B(n_548), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_213), .B(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_228), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_219), .B(n_245), .Y(n_334) );
OR2x2_ASAP7_75t_L g356 ( .A(n_219), .B(n_229), .Y(n_356) );
AND2x2_ASAP7_75t_L g369 ( .A(n_219), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_219), .B(n_324), .Y(n_375) );
OAI211xp5_ASAP7_75t_SL g379 ( .A1(n_219), .A2(n_380), .B(n_385), .C(n_394), .Y(n_379) );
AND2x2_ASAP7_75t_L g440 ( .A(n_219), .B(n_244), .Y(n_440) );
INVx5_ASAP7_75t_SL g219 ( .A(n_220), .Y(n_219) );
OR2x2_ASAP7_75t_L g293 ( .A(n_220), .B(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_220), .B(n_299), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_220), .B(n_288), .Y(n_300) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_220), .Y(n_302) );
OR2x2_ASAP7_75t_L g313 ( .A(n_220), .B(n_229), .Y(n_313) );
AND2x2_ASAP7_75t_SL g318 ( .A(n_220), .B(n_304), .Y(n_318) );
AND2x2_ASAP7_75t_L g343 ( .A(n_220), .B(n_229), .Y(n_343) );
AND2x2_ASAP7_75t_L g363 ( .A(n_220), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g401 ( .A(n_220), .B(n_228), .Y(n_401) );
OR2x2_ASAP7_75t_L g404 ( .A(n_220), .B(n_390), .Y(n_404) );
OR2x6_ASAP7_75t_L g220 ( .A(n_221), .B(n_227), .Y(n_220) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_244), .Y(n_228) );
A2O1A1Ixp33_ASAP7_75t_L g347 ( .A1(n_229), .A2(n_348), .B(n_351), .C(n_357), .Y(n_347) );
INVx5_ASAP7_75t_SL g229 ( .A(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_230), .B(n_244), .Y(n_278) );
AND2x2_ASAP7_75t_L g282 ( .A(n_230), .B(n_245), .Y(n_282) );
OR2x2_ASAP7_75t_L g288 ( .A(n_230), .B(n_244), .Y(n_288) );
OAI21xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_234), .Y(n_231) );
OAI21xp5_ASAP7_75t_L g472 ( .A1(n_233), .A2(n_473), .B(n_474), .Y(n_472) );
OAI21xp5_ASAP7_75t_L g523 ( .A1(n_233), .A2(n_524), .B(n_525), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B(n_238), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_238), .A2(n_250), .B(n_252), .Y(n_249) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
INVx2_ASAP7_75t_L g483 ( .A(n_243), .Y(n_483) );
INVx1_ASAP7_75t_SL g305 ( .A(n_244), .Y(n_305) );
OR2x2_ASAP7_75t_L g433 ( .A(n_244), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_273), .B(n_276), .C(n_285), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AOI31xp33_ASAP7_75t_L g358 ( .A1(n_255), .A2(n_359), .A3(n_361), .B(n_362), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_256), .B(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_257), .B(n_289), .Y(n_295) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_258), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g315 ( .A(n_258), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g320 ( .A(n_258), .B(n_290), .Y(n_320) );
AND2x2_ASAP7_75t_L g330 ( .A(n_258), .B(n_289), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_258), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g350 ( .A(n_258), .B(n_307), .Y(n_350) );
AND2x2_ASAP7_75t_L g355 ( .A(n_258), .B(n_327), .Y(n_355) );
OR2x2_ASAP7_75t_L g374 ( .A(n_258), .B(n_260), .Y(n_374) );
OR2x2_ASAP7_75t_L g376 ( .A(n_258), .B(n_377), .Y(n_376) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_258), .Y(n_423) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g323 ( .A(n_260), .B(n_290), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_260), .B(n_307), .Y(n_346) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
BUFx2_ASAP7_75t_L g292 ( .A(n_262), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_270), .Y(n_263) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx3_ASAP7_75t_L g504 ( .A(n_269), .Y(n_504) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g383 ( .A(n_275), .B(n_307), .Y(n_383) );
AOI322xp5_ASAP7_75t_L g385 ( .A1(n_275), .A2(n_289), .A3(n_327), .B1(n_386), .B2(n_387), .C1(n_388), .C2(n_391), .Y(n_385) );
INVx1_ASAP7_75t_L g393 ( .A(n_275), .Y(n_393) );
NAND2xp33_ASAP7_75t_L g276 ( .A(n_277), .B(n_280), .Y(n_276) );
INVx1_ASAP7_75t_SL g387 ( .A(n_277), .Y(n_387) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
OR2x2_ASAP7_75t_L g339 ( .A(n_278), .B(n_284), .Y(n_339) );
INVx1_ASAP7_75t_L g370 ( .A(n_278), .Y(n_370) );
INVx2_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
AND2x4_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OAI32xp33_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_289), .A3(n_291), .B1(n_293), .B2(n_295), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
AOI21xp33_ASAP7_75t_SL g325 ( .A1(n_288), .A2(n_303), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g340 ( .A(n_289), .Y(n_340) );
AND2x4_ASAP7_75t_L g337 ( .A(n_290), .B(n_307), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_290), .B(n_373), .Y(n_372) );
AOI322xp5_ASAP7_75t_L g402 ( .A1(n_291), .A2(n_318), .A3(n_337), .B1(n_370), .B2(n_403), .C1(n_405), .C2(n_406), .Y(n_402) );
OAI221xp5_ASAP7_75t_L g431 ( .A1(n_291), .A2(n_368), .B1(n_432), .B2(n_433), .C(n_435), .Y(n_431) );
AND2x2_ASAP7_75t_L g319 ( .A(n_292), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_SL g299 ( .A(n_294), .Y(n_299) );
OR2x2_ASAP7_75t_L g371 ( .A(n_294), .B(n_356), .Y(n_371) );
OAI31xp33_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_300), .A3(n_301), .B(n_306), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_297), .A2(n_330), .B1(n_331), .B2(n_335), .Y(n_329) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g342 ( .A(n_299), .B(n_343), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_301), .A2(n_342), .B1(n_395), .B2(n_398), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g384 ( .A(n_304), .B(n_353), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_304), .B(n_343), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_305), .B(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g418 ( .A(n_305), .B(n_356), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_306), .A2(n_401), .B1(n_414), .B2(n_417), .Y(n_413) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx2_ASAP7_75t_L g322 ( .A(n_307), .Y(n_322) );
AND2x2_ASAP7_75t_L g405 ( .A(n_307), .B(n_327), .Y(n_405) );
OR2x2_ASAP7_75t_L g407 ( .A(n_307), .B(n_374), .Y(n_407) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_307), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_308), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_308), .B(n_353), .Y(n_361) );
OAI211xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_314), .B(n_317), .C(n_329), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AOI221xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_319), .B1(n_321), .B2(n_324), .C(n_325), .Y(n_317) );
INVxp67_ASAP7_75t_L g429 ( .A(n_320), .Y(n_429) );
INVx1_ASAP7_75t_L g396 ( .A(n_321), .Y(n_396) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
AND2x2_ASAP7_75t_L g360 ( .A(n_322), .B(n_327), .Y(n_360) );
INVx1_ASAP7_75t_L g377 ( .A(n_323), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_323), .B(n_350), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
INVx1_ASAP7_75t_L g392 ( .A(n_327), .Y(n_392) );
AND2x2_ASAP7_75t_L g398 ( .A(n_327), .B(n_353), .Y(n_398) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx1_ASAP7_75t_SL g386 ( .A(n_334), .Y(n_386) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_337), .B(n_373), .Y(n_397) );
OAI221xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_340), .B1(n_341), .B2(n_344), .C(n_347), .Y(n_338) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g434 ( .A(n_343), .Y(n_434) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g352 ( .A(n_346), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_350), .B(n_409), .Y(n_408) );
AOI21xp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_354), .B(n_356), .Y(n_351) );
OAI211xp5_ASAP7_75t_SL g399 ( .A1(n_354), .A2(n_400), .B(n_402), .C(n_408), .Y(n_399) );
INVx1_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g411 ( .A(n_356), .Y(n_411) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI222xp33_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_368), .B1(n_371), .B2(n_372), .C1(n_375), .C2(n_376), .Y(n_365) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g441 ( .A(n_372), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_373), .B(n_416), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_373), .A2(n_420), .B1(n_422), .B2(n_425), .Y(n_419) );
INVx2_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
NOR4xp25_ASAP7_75t_L g378 ( .A(n_379), .B(n_399), .C(n_412), .D(n_431), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_381), .B(n_411), .Y(n_421) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g388 ( .A(n_386), .B(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_389), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_396), .B(n_397), .Y(n_395) );
INVx1_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NAND3xp33_ASAP7_75t_L g412 ( .A(n_413), .B(n_419), .C(n_426), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
INVx2_ASAP7_75t_L g428 ( .A(n_424), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
OAI21xp5_ASAP7_75t_SL g435 ( .A1(n_436), .A2(n_438), .B(n_441), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_443), .A2(n_458), .B1(n_461), .B2(n_462), .Y(n_457) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g454 ( .A(n_447), .Y(n_454) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g731 ( .A(n_459), .Y(n_731) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g734 ( .A(n_461), .Y(n_734) );
INVx2_ASAP7_75t_L g732 ( .A(n_462), .Y(n_732) );
OR2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_657), .Y(n_462) );
NAND5xp2_ASAP7_75t_L g463 ( .A(n_464), .B(n_586), .C(n_616), .D(n_637), .E(n_643), .Y(n_463) );
AOI221xp5_ASAP7_75t_SL g464 ( .A1(n_465), .A2(n_519), .B1(n_550), .B2(n_552), .C(n_563), .Y(n_464) );
INVxp67_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_516), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_468), .B(n_494), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_SL g637 ( .A1(n_469), .A2(n_506), .B(n_638), .C(n_641), .Y(n_637) );
AND2x2_ASAP7_75t_L g707 ( .A(n_469), .B(n_507), .Y(n_707) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_481), .Y(n_469) );
AND2x2_ASAP7_75t_L g565 ( .A(n_470), .B(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g569 ( .A(n_470), .B(n_566), .Y(n_569) );
OR2x2_ASAP7_75t_L g595 ( .A(n_470), .B(n_507), .Y(n_595) );
AND2x2_ASAP7_75t_L g597 ( .A(n_470), .B(n_497), .Y(n_597) );
AND2x2_ASAP7_75t_L g615 ( .A(n_470), .B(n_496), .Y(n_615) );
INVx1_ASAP7_75t_L g648 ( .A(n_470), .Y(n_648) );
INVx2_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g518 ( .A(n_471), .Y(n_518) );
AND2x2_ASAP7_75t_L g551 ( .A(n_471), .B(n_497), .Y(n_551) );
AND2x2_ASAP7_75t_L g704 ( .A(n_471), .B(n_507), .Y(n_704) );
AND2x2_ASAP7_75t_L g585 ( .A(n_481), .B(n_495), .Y(n_585) );
OR2x2_ASAP7_75t_L g589 ( .A(n_481), .B(n_507), .Y(n_589) );
AND2x2_ASAP7_75t_L g614 ( .A(n_481), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_SL g661 ( .A(n_481), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_481), .B(n_623), .Y(n_709) );
AO21x2_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_484), .B(n_492), .Y(n_481) );
INVx1_ASAP7_75t_L g567 ( .A(n_482), .Y(n_567) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OA21x2_ASAP7_75t_L g566 ( .A1(n_485), .A2(n_493), .B(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
OAI322xp33_ASAP7_75t_L g710 ( .A1(n_494), .A2(n_646), .A3(n_669), .B1(n_690), .B2(n_711), .C1(n_713), .C2(n_714), .Y(n_710) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_495), .B(n_566), .Y(n_713) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_506), .Y(n_495) );
AND2x2_ASAP7_75t_L g517 ( .A(n_496), .B(n_518), .Y(n_517) );
AND2x4_ASAP7_75t_L g582 ( .A(n_496), .B(n_507), .Y(n_582) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g623 ( .A(n_497), .B(n_507), .Y(n_623) );
AND2x2_ASAP7_75t_L g667 ( .A(n_497), .B(n_506), .Y(n_667) );
AND2x2_ASAP7_75t_L g550 ( .A(n_506), .B(n_551), .Y(n_550) );
OR2x2_ASAP7_75t_L g568 ( .A(n_506), .B(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_506), .B(n_597), .Y(n_721) );
INVx3_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g516 ( .A(n_507), .B(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_507), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g635 ( .A(n_507), .B(n_566), .Y(n_635) );
AND2x2_ASAP7_75t_L g662 ( .A(n_507), .B(n_597), .Y(n_662) );
OR2x2_ASAP7_75t_L g718 ( .A(n_507), .B(n_569), .Y(n_718) );
OR2x6_ASAP7_75t_L g507 ( .A(n_508), .B(n_514), .Y(n_507) );
INVx1_ASAP7_75t_SL g604 ( .A(n_516), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_517), .B(n_635), .Y(n_636) );
AND2x2_ASAP7_75t_L g670 ( .A(n_517), .B(n_660), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_517), .B(n_593), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_517), .B(n_715), .Y(n_714) );
OAI31xp33_ASAP7_75t_L g688 ( .A1(n_519), .A2(n_550), .A3(n_689), .B(n_691), .Y(n_688) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_531), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g655 ( .A(n_520), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g671 ( .A(n_520), .B(n_606), .Y(n_671) );
OR2x2_ASAP7_75t_L g678 ( .A(n_520), .B(n_679), .Y(n_678) );
OR2x2_ASAP7_75t_L g690 ( .A(n_520), .B(n_579), .Y(n_690) );
CKINVDCx16_ASAP7_75t_R g520 ( .A(n_521), .Y(n_520) );
OR2x2_ASAP7_75t_L g624 ( .A(n_521), .B(n_625), .Y(n_624) );
BUFx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g552 ( .A(n_522), .B(n_553), .Y(n_552) );
INVx4_ASAP7_75t_L g573 ( .A(n_522), .Y(n_573) );
AND2x2_ASAP7_75t_L g610 ( .A(n_522), .B(n_554), .Y(n_610) );
AND2x2_ASAP7_75t_L g609 ( .A(n_531), .B(n_610), .Y(n_609) );
INVx1_ASAP7_75t_SL g679 ( .A(n_531), .Y(n_679) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_541), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_532), .B(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g579 ( .A(n_532), .B(n_542), .Y(n_579) );
INVx2_ASAP7_75t_L g599 ( .A(n_532), .Y(n_599) );
AND2x2_ASAP7_75t_L g613 ( .A(n_532), .B(n_542), .Y(n_613) );
AND2x2_ASAP7_75t_L g620 ( .A(n_532), .B(n_576), .Y(n_620) );
BUFx3_ASAP7_75t_L g630 ( .A(n_532), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_532), .B(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g575 ( .A(n_541), .Y(n_575) );
AND2x2_ASAP7_75t_L g583 ( .A(n_541), .B(n_573), .Y(n_583) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g553 ( .A(n_542), .B(n_554), .Y(n_553) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_542), .Y(n_607) );
INVx2_ASAP7_75t_SL g590 ( .A(n_551), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_551), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_551), .B(n_660), .Y(n_681) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_552), .B(n_630), .Y(n_683) );
INVx1_ASAP7_75t_SL g717 ( .A(n_552), .Y(n_717) );
INVx1_ASAP7_75t_SL g625 ( .A(n_553), .Y(n_625) );
INVx1_ASAP7_75t_SL g576 ( .A(n_554), .Y(n_576) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_554), .Y(n_587) );
OR2x2_ASAP7_75t_L g598 ( .A(n_554), .B(n_573), .Y(n_598) );
AND2x2_ASAP7_75t_L g612 ( .A(n_554), .B(n_573), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_554), .B(n_602), .Y(n_664) );
A2O1A1Ixp33_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_568), .B(n_570), .C(n_581), .Y(n_563) );
AOI31xp33_ASAP7_75t_L g680 ( .A1(n_564), .A2(n_681), .A3(n_682), .B(n_683), .Y(n_680) );
AND2x2_ASAP7_75t_L g653 ( .A(n_565), .B(n_582), .Y(n_653) );
BUFx3_ASAP7_75t_L g593 ( .A(n_566), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_566), .B(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g629 ( .A(n_566), .B(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_566), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_SL g584 ( .A(n_569), .Y(n_584) );
OAI222xp33_ASAP7_75t_L g693 ( .A1(n_569), .A2(n_694), .B1(n_697), .B2(n_698), .C1(n_699), .C2(n_700), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_571), .B(n_577), .Y(n_570) );
INVx1_ASAP7_75t_L g699 ( .A(n_571), .Y(n_699) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_573), .B(n_576), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_573), .B(n_599), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_573), .B(n_574), .Y(n_669) );
INVx1_ASAP7_75t_L g720 ( .A(n_573), .Y(n_720) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_574), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g722 ( .A(n_574), .Y(n_722) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
INVx2_ASAP7_75t_L g602 ( .A(n_575), .Y(n_602) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_576), .Y(n_645) );
AOI32xp33_ASAP7_75t_L g581 ( .A1(n_577), .A2(n_582), .A3(n_583), .B1(n_584), .B2(n_585), .Y(n_581) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_579), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g656 ( .A(n_579), .Y(n_656) );
OR2x2_ASAP7_75t_L g697 ( .A(n_579), .B(n_598), .Y(n_697) );
INVx1_ASAP7_75t_L g633 ( .A(n_580), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_582), .B(n_593), .Y(n_618) );
INVx3_ASAP7_75t_L g627 ( .A(n_582), .Y(n_627) );
AOI322xp5_ASAP7_75t_L g643 ( .A1(n_582), .A2(n_627), .A3(n_644), .B1(n_646), .B2(n_649), .C1(n_653), .C2(n_654), .Y(n_643) );
AND2x2_ASAP7_75t_L g619 ( .A(n_583), .B(n_620), .Y(n_619) );
INVxp67_ASAP7_75t_L g696 ( .A(n_583), .Y(n_696) );
A2O1A1O1Ixp25_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_588), .B(n_591), .C(n_599), .D(n_600), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_587), .B(n_630), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
OAI221xp5_ASAP7_75t_L g600 ( .A1(n_589), .A2(n_601), .B1(n_604), .B2(n_605), .C(n_608), .Y(n_600) );
INVx1_ASAP7_75t_SL g715 ( .A(n_589), .Y(n_715) );
AOI21xp33_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_596), .B(n_598), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g703 ( .A(n_593), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OAI221xp5_ASAP7_75t_SL g685 ( .A1(n_595), .A2(n_679), .B1(n_686), .B2(n_687), .C(n_688), .Y(n_685) );
OAI222xp33_ASAP7_75t_L g716 ( .A1(n_596), .A2(n_717), .B1(n_718), .B2(n_719), .C1(n_721), .C2(n_722), .Y(n_716) );
AND2x2_ASAP7_75t_L g674 ( .A(n_597), .B(n_660), .Y(n_674) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_597), .A2(n_612), .B(n_659), .Y(n_686) );
INVx1_ASAP7_75t_L g700 ( .A(n_597), .Y(n_700) );
INVx2_ASAP7_75t_SL g603 ( .A(n_598), .Y(n_603) );
AND2x2_ASAP7_75t_L g606 ( .A(n_599), .B(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
INVx1_ASAP7_75t_SL g640 ( .A(n_602), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_602), .B(n_612), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_603), .B(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_603), .B(n_613), .Y(n_642) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OAI21xp5_ASAP7_75t_SL g608 ( .A1(n_609), .A2(n_611), .B(n_614), .Y(n_608) );
INVx1_ASAP7_75t_SL g626 ( .A(n_610), .Y(n_626) );
AND2x2_ASAP7_75t_L g673 ( .A(n_610), .B(n_656), .Y(n_673) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
AND2x2_ASAP7_75t_L g712 ( .A(n_612), .B(n_630), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_613), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_SL g698 ( .A(n_614), .Y(n_698) );
AOI221xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_619), .B1(n_621), .B2(n_628), .C(n_631), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_624), .B1(n_626), .B2(n_627), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OAI22xp33_ASAP7_75t_L g631 ( .A1(n_625), .A2(n_632), .B1(n_634), .B2(n_636), .Y(n_631) );
OR2x2_ASAP7_75t_L g702 ( .A(n_626), .B(n_630), .Y(n_702) );
OR2x2_ASAP7_75t_L g705 ( .A(n_626), .B(n_640), .Y(n_705) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OAI221xp5_ASAP7_75t_L g701 ( .A1(n_647), .A2(n_702), .B1(n_703), .B2(n_705), .C(n_706), .Y(n_701) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVxp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND3xp33_ASAP7_75t_SL g657 ( .A(n_658), .B(n_672), .C(n_684), .Y(n_657) );
AOI222xp33_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_663), .B1(n_665), .B2(n_668), .C1(n_670), .C2(n_671), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_662), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_660), .B(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g682 ( .A(n_662), .Y(n_682) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVxp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_674), .B1(n_675), .B2(n_677), .C(n_680), .Y(n_672) );
INVx1_ASAP7_75t_L g687 ( .A(n_673), .Y(n_687) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OAI21xp33_ASAP7_75t_L g706 ( .A1(n_677), .A2(n_707), .B(n_708), .Y(n_706) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
NOR5xp2_ASAP7_75t_L g684 ( .A(n_685), .B(n_693), .C(n_701), .D(n_710), .E(n_716), .Y(n_684) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
INVxp67_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx3_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
endmodule