module fake_netlist_5_483_n_2590 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_74, n_515, n_57, n_353, n_351, n_367, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_590, n_4, n_378, n_551, n_17, n_581, n_382, n_554, n_254, n_33, n_23, n_583, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_559, n_275, n_252, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_584, n_591, n_145, n_48, n_521, n_50, n_337, n_430, n_313, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_502, n_239, n_466, n_420, n_489, n_55, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_480, n_237, n_425, n_513, n_407, n_527, n_180, n_560, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_572, n_113, n_246, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_541, n_391, n_434, n_539, n_175, n_538, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_2590);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_590;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_382;
input n_554;
input n_254;
input n_33;
input n_23;
input n_583;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_559;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_584;
input n_591;
input n_145;
input n_48;
input n_521;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_480;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_560;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_541;
input n_391;
input n_434;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_2590;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_785;
wire n_2200;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_1007;
wire n_2369;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_956;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_800;
wire n_1347;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2396;
wire n_2069;
wire n_1580;
wire n_674;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_1118;
wire n_755;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_1107;
wire n_1728;
wire n_2031;
wire n_2076;
wire n_2482;
wire n_1230;
wire n_668;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_2584;
wire n_1257;
wire n_1182;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_2323;
wire n_2203;
wire n_1243;
wire n_1016;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_2515;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2276;
wire n_1547;
wire n_1070;
wire n_777;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_1561;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_845;
wire n_663;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_2300;
wire n_1796;
wire n_2551;
wire n_680;
wire n_1473;
wire n_1587;
wire n_901;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_2506;
wire n_675;
wire n_888;
wire n_1880;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_1585;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_2258;
wire n_748;
wire n_1058;
wire n_1667;
wire n_838;
wire n_1053;
wire n_1224;
wire n_2557;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2324;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_857;
wire n_832;
wire n_2305;
wire n_2450;
wire n_1319;
wire n_2379;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2331;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_702;
wire n_1276;
wire n_2548;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_1884;
wire n_2434;
wire n_1038;
wire n_1369;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_868;
wire n_2454;
wire n_639;
wire n_914;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_2518;
wire n_1415;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_1829;
wire n_1464;
wire n_649;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_604;
wire n_2007;
wire n_949;
wire n_2539;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_2577;
wire n_1760;
wire n_936;
wire n_1500;
wire n_1090;
wire n_757;
wire n_2342;
wire n_633;
wire n_1832;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_1964;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_1586;
wire n_959;
wire n_2459;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_2481;
wire n_2171;
wire n_978;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2320;
wire n_2038;
wire n_2339;
wire n_2473;
wire n_2137;
wire n_603;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_2540;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_2168;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_1574;
wire n_2399;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_1800;
wire n_1548;
wire n_614;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_2565;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2418;
wire n_829;
wire n_2519;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_1237;
wire n_700;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_2277;
wire n_761;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_1823;
wire n_874;
wire n_2464;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_860;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_628;
wire n_1849;
wire n_2410;
wire n_1131;
wire n_729;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_2467;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_1552;
wire n_2508;
wire n_602;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_623;
wire n_2088;
wire n_824;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_1821;
wire n_1381;
wire n_2555;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_716;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2534;
wire n_2092;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_803;
wire n_1092;
wire n_1776;
wire n_2198;
wire n_2572;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_1811;
wire n_2443;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_2465;
wire n_968;
wire n_912;
wire n_619;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_2541;
wire n_1139;
wire n_2333;
wire n_885;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_1283;
wire n_762;
wire n_1644;
wire n_2334;
wire n_690;
wire n_1974;
wire n_2463;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_2475;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2556;
wire n_2269;
wire n_2309;
wire n_2415;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_2533;
wire n_618;
wire n_896;
wire n_2310;
wire n_2287;
wire n_2291;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2318;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_669;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_2471;
wire n_1807;
wire n_1149;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2325;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_2588;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_849;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_2282;
wire n_2371;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_749;
wire n_1895;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_2361;
wire n_1088;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_836;
wire n_990;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_1465;
wire n_778;
wire n_1122;
wire n_770;
wire n_1375;
wire n_2494;
wire n_1102;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_1174;
wire n_2431;
wire n_2558;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_726;
wire n_982;
wire n_2575;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2437;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_1584;
wire n_1726;
wire n_665;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_2093;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_2547;
wire n_708;
wire n_1812;
wire n_735;
wire n_2501;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_1067;
wire n_1720;
wire n_2401;
wire n_2003;
wire n_1457;
wire n_766;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_872;
wire n_2012;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_2213;
wire n_2023;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_2421;
wire n_2286;
wire n_664;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_2363;
wire n_2430;
wire n_916;
wire n_1081;
wire n_2549;
wire n_2332;
wire n_1235;
wire n_980;
wire n_698;
wire n_1115;
wire n_703;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_2528;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_825;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_1489;
wire n_733;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_792;
wire n_1429;
wire n_756;
wire n_1238;
wire n_2448;
wire n_812;
wire n_2104;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_1675;
wire n_1924;
wire n_2573;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2497;
wire n_2006;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2172;
wire n_1973;
wire n_1083;
wire n_786;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2456;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_2451;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_2567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_685;
wire n_598;
wire n_928;
wire n_1367;
wire n_608;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_2531;
wire n_1589;
wire n_1086;
wire n_2570;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_1546;
wire n_595;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_2112;
wire n_1739;
wire n_616;
wire n_2278;
wire n_2394;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2569;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_2027;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_2525;
wire n_2513;
wire n_1764;
wire n_712;
wire n_2414;
wire n_1583;
wire n_2426;
wire n_1042;
wire n_1402;
wire n_2049;
wire n_2273;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_2044;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_2524;
wire n_1271;
wire n_1542;
wire n_1251;
wire n_2268;

CKINVDCx16_ASAP7_75t_R g595 ( 
.A(n_481),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_574),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_32),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_589),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_180),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_416),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_507),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_548),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_149),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_348),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_316),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_386),
.Y(n_606)
);

INVx1_ASAP7_75t_SL g607 ( 
.A(n_533),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_234),
.Y(n_608)
);

INVx1_ASAP7_75t_SL g609 ( 
.A(n_257),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_583),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_198),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_211),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_190),
.Y(n_613)
);

BUFx10_ASAP7_75t_L g614 ( 
.A(n_418),
.Y(n_614)
);

CKINVDCx16_ASAP7_75t_R g615 ( 
.A(n_4),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_128),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_244),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_308),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_254),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_464),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_177),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_105),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_539),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_30),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_239),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_258),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_448),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_79),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_552),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_38),
.Y(n_630)
);

BUFx2_ASAP7_75t_L g631 ( 
.A(n_84),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_221),
.Y(n_632)
);

CKINVDCx16_ASAP7_75t_R g633 ( 
.A(n_239),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_593),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_398),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_582),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_509),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_368),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_36),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_102),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_428),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_540),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_571),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_508),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_541),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_476),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_274),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_78),
.Y(n_648)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_377),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_273),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_528),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_447),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_24),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_413),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_47),
.Y(n_655)
);

INVxp67_ASAP7_75t_L g656 ( 
.A(n_354),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_258),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_62),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_201),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_203),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_35),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_323),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_536),
.Y(n_663)
);

BUFx10_ASAP7_75t_L g664 ( 
.A(n_130),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_393),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_248),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_14),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_160),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_521),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_438),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_300),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_500),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_337),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_14),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_275),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_579),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_91),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_61),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_128),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_372),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_51),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_80),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_236),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_104),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_255),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_58),
.Y(n_686)
);

BUFx10_ASAP7_75t_L g687 ( 
.A(n_293),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_371),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_575),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_576),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_457),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_562),
.Y(n_692)
);

INVx1_ASAP7_75t_SL g693 ( 
.A(n_6),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_477),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_445),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_471),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_335),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_68),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_189),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_185),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_178),
.Y(n_701)
);

BUFx2_ASAP7_75t_L g702 ( 
.A(n_231),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_212),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_166),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_33),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_279),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_106),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_526),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_268),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_26),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_75),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_307),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_373),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_279),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_299),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_559),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_149),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_524),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_20),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_87),
.Y(n_720)
);

CKINVDCx14_ASAP7_75t_R g721 ( 
.A(n_229),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_567),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_72),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_208),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_159),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_489),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_350),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_75),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_15),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_158),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_210),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_276),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_50),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_473),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_323),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_544),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_49),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_459),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_396),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_8),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_333),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_266),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_63),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_205),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_470),
.Y(n_745)
);

CKINVDCx20_ASAP7_75t_R g746 ( 
.A(n_490),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_150),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_177),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_550),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_12),
.Y(n_750)
);

CKINVDCx20_ASAP7_75t_R g751 ( 
.A(n_448),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_569),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_378),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_300),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_510),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_306),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_504),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_45),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_27),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_429),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_12),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_184),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_235),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_335),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_502),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_413),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_565),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_88),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_285),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_1),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_591),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_449),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_367),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_248),
.Y(n_774)
);

CKINVDCx20_ASAP7_75t_R g775 ( 
.A(n_307),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_344),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_124),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_54),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_250),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_82),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_285),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_453),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_302),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_98),
.Y(n_784)
);

BUFx5_ASAP7_75t_L g785 ( 
.A(n_196),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_70),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_42),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_112),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_250),
.Y(n_789)
);

BUFx3_ASAP7_75t_L g790 ( 
.A(n_212),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_13),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_523),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_77),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_512),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_450),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_236),
.Y(n_796)
);

CKINVDCx20_ASAP7_75t_R g797 ( 
.A(n_133),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_0),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_211),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_263),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_483),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_288),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_269),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_414),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_372),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_594),
.Y(n_806)
);

CKINVDCx20_ASAP7_75t_R g807 ( 
.A(n_87),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_377),
.Y(n_808)
);

INVx1_ASAP7_75t_SL g809 ( 
.A(n_527),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_459),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_458),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_70),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_407),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_442),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_136),
.Y(n_815)
);

BUFx10_ASAP7_75t_L g816 ( 
.A(n_256),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_122),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_292),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_331),
.Y(n_819)
);

BUFx2_ASAP7_75t_L g820 ( 
.A(n_203),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_312),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_133),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_257),
.Y(n_823)
);

CKINVDCx14_ASAP7_75t_R g824 ( 
.A(n_385),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_160),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_240),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_59),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_734),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_785),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_785),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_785),
.Y(n_831)
);

INVxp33_ASAP7_75t_L g832 ( 
.A(n_698),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_785),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_734),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_721),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_785),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_824),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_785),
.Y(n_838)
);

INVxp67_ASAP7_75t_SL g839 ( 
.A(n_759),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_785),
.Y(n_840)
);

INVxp67_ASAP7_75t_SL g841 ( 
.A(n_759),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_759),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_611),
.Y(n_843)
);

INVxp67_ASAP7_75t_SL g844 ( 
.A(n_625),
.Y(n_844)
);

INVxp67_ASAP7_75t_SL g845 ( 
.A(n_625),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_615),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_611),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_625),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_625),
.Y(n_849)
);

INVxp33_ASAP7_75t_SL g850 ( 
.A(n_613),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_684),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_622),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_684),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_771),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_684),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_684),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_787),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_787),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_787),
.Y(n_859)
);

BUFx2_ASAP7_75t_L g860 ( 
.A(n_631),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_622),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_638),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_638),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_653),
.Y(n_864)
);

CKINVDCx20_ASAP7_75t_R g865 ( 
.A(n_621),
.Y(n_865)
);

CKINVDCx16_ASAP7_75t_R g866 ( 
.A(n_633),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_653),
.Y(n_867)
);

INVxp67_ASAP7_75t_L g868 ( 
.A(n_702),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_820),
.Y(n_869)
);

CKINVDCx20_ASAP7_75t_R g870 ( 
.A(n_621),
.Y(n_870)
);

INVxp67_ASAP7_75t_L g871 ( 
.A(n_614),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_771),
.Y(n_872)
);

INVxp33_ASAP7_75t_L g873 ( 
.A(n_597),
.Y(n_873)
);

BUFx2_ASAP7_75t_SL g874 ( 
.A(n_718),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_688),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_758),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_758),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_784),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_784),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_790),
.Y(n_880)
);

BUFx2_ASAP7_75t_SL g881 ( 
.A(n_718),
.Y(n_881)
);

INVxp33_ASAP7_75t_SL g882 ( 
.A(n_613),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_787),
.Y(n_883)
);

INVxp33_ASAP7_75t_SL g884 ( 
.A(n_617),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_796),
.Y(n_885)
);

CKINVDCx20_ASAP7_75t_R g886 ( 
.A(n_640),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_796),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_669),
.B(n_801),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_796),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_796),
.Y(n_890)
);

INVx1_ASAP7_75t_SL g891 ( 
.A(n_614),
.Y(n_891)
);

INVxp67_ASAP7_75t_SL g892 ( 
.A(n_819),
.Y(n_892)
);

INVxp67_ASAP7_75t_SL g893 ( 
.A(n_819),
.Y(n_893)
);

CKINVDCx20_ASAP7_75t_R g894 ( 
.A(n_640),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_819),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_819),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_600),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_606),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_616),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_801),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_628),
.Y(n_901)
);

INVxp67_ASAP7_75t_SL g902 ( 
.A(n_596),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_632),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_650),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_639),
.Y(n_905)
);

INVxp67_ASAP7_75t_SL g906 ( 
.A(n_598),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_641),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_652),
.Y(n_908)
);

INVxp33_ASAP7_75t_L g909 ( 
.A(n_655),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_699),
.Y(n_910)
);

CKINVDCx20_ASAP7_75t_R g911 ( 
.A(n_650),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_658),
.Y(n_912)
);

CKINVDCx20_ASAP7_75t_R g913 ( 
.A(n_658),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_667),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_599),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_671),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_603),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_617),
.Y(n_918)
);

BUFx2_ASAP7_75t_SL g919 ( 
.A(n_746),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_618),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_604),
.Y(n_921)
);

CKINVDCx16_ASAP7_75t_R g922 ( 
.A(n_595),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_844),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_845),
.B(n_601),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_828),
.B(n_610),
.Y(n_925)
);

OR2x2_ASAP7_75t_L g926 ( 
.A(n_891),
.B(n_609),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_854),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_854),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_834),
.Y(n_929)
);

BUFx8_ASAP7_75t_SL g930 ( 
.A(n_865),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_854),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_888),
.B(n_902),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_848),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_854),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_906),
.B(n_607),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_834),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_848),
.Y(n_937)
);

BUFx2_ASAP7_75t_L g938 ( 
.A(n_846),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_854),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_872),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_850),
.B(n_882),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_SL g942 ( 
.A(n_922),
.B(n_746),
.Y(n_942)
);

INVx4_ASAP7_75t_L g943 ( 
.A(n_834),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_828),
.B(n_629),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_839),
.B(n_841),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_872),
.Y(n_946)
);

BUFx8_ASAP7_75t_SL g947 ( 
.A(n_865),
.Y(n_947)
);

INVx2_ASAP7_75t_SL g948 ( 
.A(n_915),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_892),
.B(n_634),
.Y(n_949)
);

BUFx12f_ASAP7_75t_L g950 ( 
.A(n_835),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_SL g951 ( 
.A(n_866),
.B(n_752),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_872),
.Y(n_952)
);

BUFx3_ASAP7_75t_L g953 ( 
.A(n_834),
.Y(n_953)
);

HB1xp67_ASAP7_75t_L g954 ( 
.A(n_918),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_850),
.B(n_623),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_920),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_835),
.B(n_637),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_893),
.B(n_645),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_872),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_834),
.B(n_672),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_842),
.B(n_690),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_868),
.B(n_692),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_849),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_849),
.Y(n_964)
);

BUFx12f_ASAP7_75t_L g965 ( 
.A(n_837),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_851),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_843),
.B(n_694),
.Y(n_967)
);

CKINVDCx20_ASAP7_75t_R g968 ( 
.A(n_870),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_851),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_900),
.B(n_889),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_889),
.B(n_696),
.Y(n_971)
);

BUFx8_ASAP7_75t_L g972 ( 
.A(n_860),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_900),
.B(n_736),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_900),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_853),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_853),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_855),
.B(n_749),
.Y(n_977)
);

AND2x6_ASAP7_75t_L g978 ( 
.A(n_831),
.B(n_767),
.Y(n_978)
);

INVx5_ASAP7_75t_L g979 ( 
.A(n_831),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_855),
.B(n_809),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_847),
.B(n_825),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_852),
.B(n_602),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_856),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_915),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_970),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_971),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_927),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_955),
.B(n_837),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_961),
.B(n_910),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_933),
.Y(n_990)
);

CKINVDCx11_ASAP7_75t_R g991 ( 
.A(n_968),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_927),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_955),
.B(n_917),
.Y(n_993)
);

AND2x6_ASAP7_75t_L g994 ( 
.A(n_924),
.B(n_699),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_971),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_945),
.B(n_882),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_935),
.B(n_856),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_971),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_927),
.Y(n_999)
);

INVx4_ASAP7_75t_L g1000 ( 
.A(n_979),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_927),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_933),
.Y(n_1002)
);

AND2x4_ASAP7_75t_L g1003 ( 
.A(n_961),
.B(n_977),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_937),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_926),
.Y(n_1005)
);

INVx5_ASAP7_75t_L g1006 ( 
.A(n_978),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_937),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_935),
.B(n_857),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_963),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_963),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_950),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_960),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_963),
.Y(n_1013)
);

INVxp67_ASAP7_75t_L g1014 ( 
.A(n_941),
.Y(n_1014)
);

OA21x2_ASAP7_75t_L g1015 ( 
.A1(n_973),
.A2(n_830),
.B(n_829),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_928),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_963),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_928),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_928),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_923),
.B(n_884),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_964),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_932),
.B(n_857),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_977),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_977),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_964),
.Y(n_1025)
);

CKINVDCx11_ASAP7_75t_R g1026 ( 
.A(n_968),
.Y(n_1026)
);

HB1xp67_ASAP7_75t_L g1027 ( 
.A(n_957),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_954),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_929),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_929),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_928),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_931),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_931),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_936),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_931),
.Y(n_1035)
);

INVx1_ASAP7_75t_SL g1036 ( 
.A(n_930),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_954),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_936),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_953),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_932),
.B(n_858),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_931),
.Y(n_1041)
);

AND2x6_ASAP7_75t_L g1042 ( 
.A(n_924),
.B(n_782),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_953),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_956),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_982),
.B(n_884),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_924),
.B(n_858),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_964),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_934),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_964),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_934),
.Y(n_1050)
);

INVxp67_ASAP7_75t_L g1051 ( 
.A(n_941),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_966),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_966),
.Y(n_1053)
);

HB1xp67_ASAP7_75t_L g1054 ( 
.A(n_956),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_961),
.B(n_910),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_966),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_965),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_934),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_966),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_969),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_969),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_967),
.B(n_833),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_969),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_967),
.B(n_861),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_925),
.B(n_836),
.Y(n_1065)
);

HB1xp67_ASAP7_75t_L g1066 ( 
.A(n_938),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_969),
.Y(n_1067)
);

INVx4_ASAP7_75t_L g1068 ( 
.A(n_979),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_943),
.B(n_859),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_975),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_934),
.Y(n_1071)
);

INVxp33_ASAP7_75t_L g1072 ( 
.A(n_1005),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_1003),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_990),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_1065),
.Y(n_1075)
);

NOR3xp33_ASAP7_75t_L g1076 ( 
.A(n_988),
.B(n_984),
.C(n_948),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_990),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_986),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_1002),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1012),
.B(n_980),
.Y(n_1080)
);

OAI22xp33_ASAP7_75t_L g1081 ( 
.A1(n_1027),
.A2(n_942),
.B1(n_951),
.B2(n_917),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_1065),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_1028),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_986),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1002),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_1004),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_1004),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_996),
.B(n_980),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_1045),
.B(n_980),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_995),
.Y(n_1090)
);

NOR2x1p5_ASAP7_75t_L g1091 ( 
.A(n_1011),
.B(n_965),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_991),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_1020),
.B(n_1014),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_995),
.Y(n_1094)
);

INVx8_ASAP7_75t_L g1095 ( 
.A(n_994),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_998),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1007),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_998),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_989),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_989),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_1051),
.B(n_993),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1007),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_1003),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1023),
.Y(n_1104)
);

AO21x2_ASAP7_75t_L g1105 ( 
.A1(n_1012),
.A2(n_958),
.B(n_949),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_SL g1106 ( 
.A(n_1065),
.Y(n_1106)
);

INVx5_ASAP7_75t_L g1107 ( 
.A(n_994),
.Y(n_1107)
);

OR2x2_ASAP7_75t_L g1108 ( 
.A(n_1028),
.B(n_874),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_1003),
.B(n_921),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_1022),
.B(n_874),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_1055),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_994),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1055),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1029),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_997),
.B(n_921),
.Y(n_1115)
);

INVx3_ASAP7_75t_L g1116 ( 
.A(n_1009),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_1008),
.B(n_1065),
.Y(n_1117)
);

CKINVDCx6p67_ASAP7_75t_R g1118 ( 
.A(n_1026),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_985),
.B(n_1023),
.Y(n_1119)
);

AO22x1_ASAP7_75t_L g1120 ( 
.A1(n_994),
.A2(n_962),
.B1(n_832),
.B2(n_944),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1029),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_1062),
.B(n_925),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1030),
.Y(n_1123)
);

INVx5_ASAP7_75t_L g1124 ( 
.A(n_994),
.Y(n_1124)
);

NAND2xp33_ASAP7_75t_L g1125 ( 
.A(n_994),
.B(n_978),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1030),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1024),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_985),
.B(n_944),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1024),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_1037),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_1062),
.B(n_962),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1034),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_1062),
.B(n_620),
.Y(n_1133)
);

INVx2_ASAP7_75t_SL g1134 ( 
.A(n_1064),
.Y(n_1134)
);

AOI22x1_ASAP7_75t_L g1135 ( 
.A1(n_1064),
.A2(n_860),
.B1(n_869),
.B2(n_981),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_1062),
.B(n_620),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_1009),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1046),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1034),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_1040),
.B(n_881),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_994),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_1037),
.B(n_722),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_1054),
.B(n_881),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1038),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1039),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1044),
.B(n_981),
.Y(n_1146)
);

AOI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1069),
.A2(n_840),
.B(n_838),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_1044),
.B(n_722),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1039),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1043),
.Y(n_1150)
);

BUFx4f_ASAP7_75t_L g1151 ( 
.A(n_1042),
.Y(n_1151)
);

NAND3xp33_ASAP7_75t_L g1152 ( 
.A(n_1066),
.B(n_869),
.C(n_871),
.Y(n_1152)
);

BUFx10_ASAP7_75t_L g1153 ( 
.A(n_1011),
.Y(n_1153)
);

AO21x2_ASAP7_75t_L g1154 ( 
.A1(n_1070),
.A2(n_859),
.B(n_883),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1015),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1042),
.B(n_1070),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1015),
.Y(n_1157)
);

AOI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1015),
.A2(n_887),
.B(n_885),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_1006),
.B(n_726),
.Y(n_1159)
);

BUFx10_ASAP7_75t_L g1160 ( 
.A(n_1057),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1015),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_1053),
.B(n_919),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1071),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_1057),
.Y(n_1164)
);

INVx4_ASAP7_75t_L g1165 ( 
.A(n_1042),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1010),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_1006),
.B(n_726),
.Y(n_1167)
);

INVx1_ASAP7_75t_SL g1168 ( 
.A(n_1036),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1042),
.B(n_862),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1013),
.Y(n_1170)
);

AO21x2_ASAP7_75t_L g1171 ( 
.A1(n_1053),
.A2(n_895),
.B(n_890),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1013),
.Y(n_1172)
);

BUFx3_ASAP7_75t_L g1173 ( 
.A(n_1042),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1017),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1017),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1021),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_1006),
.B(n_792),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1042),
.B(n_978),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1021),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_SL g1180 ( 
.A(n_1042),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_1025),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1025),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1047),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1056),
.B(n_978),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1047),
.Y(n_1185)
);

INVx8_ASAP7_75t_L g1186 ( 
.A(n_1006),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1049),
.Y(n_1187)
);

INVx3_ASAP7_75t_L g1188 ( 
.A(n_1049),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1052),
.B(n_863),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1052),
.Y(n_1190)
);

NAND2xp33_ASAP7_75t_L g1191 ( 
.A(n_1006),
.B(n_978),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1059),
.B(n_864),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1059),
.Y(n_1193)
);

OR2x6_ASAP7_75t_L g1194 ( 
.A(n_1060),
.B(n_919),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1060),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_1063),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1006),
.B(n_792),
.Y(n_1197)
);

INVx8_ASAP7_75t_L g1198 ( 
.A(n_987),
.Y(n_1198)
);

NAND2xp33_ASAP7_75t_SL g1199 ( 
.A(n_1063),
.B(n_715),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1061),
.B(n_975),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_1075),
.B(n_897),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1104),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1104),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1127),
.Y(n_1204)
);

OR2x6_ASAP7_75t_L g1205 ( 
.A(n_1083),
.B(n_825),
.Y(n_1205)
);

INVx1_ASAP7_75t_SL g1206 ( 
.A(n_1083),
.Y(n_1206)
);

XNOR2x2_ASAP7_75t_L g1207 ( 
.A(n_1093),
.B(n_657),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1129),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1078),
.Y(n_1209)
);

NAND2xp33_ASAP7_75t_SL g1210 ( 
.A(n_1180),
.B(n_715),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1088),
.B(n_720),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1117),
.A2(n_1067),
.B(n_1031),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1074),
.Y(n_1213)
);

CKINVDCx20_ASAP7_75t_R g1214 ( 
.A(n_1118),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1084),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_1089),
.B(n_720),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_1118),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1090),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1094),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1138),
.B(n_1018),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1077),
.Y(n_1221)
);

XOR2x2_ASAP7_75t_L g1222 ( 
.A(n_1076),
.B(n_930),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1096),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1098),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1101),
.B(n_748),
.Y(n_1225)
);

CKINVDCx20_ASAP7_75t_R g1226 ( 
.A(n_1092),
.Y(n_1226)
);

CKINVDCx20_ASAP7_75t_R g1227 ( 
.A(n_1092),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1181),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1181),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1114),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1114),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1121),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1121),
.Y(n_1233)
);

XNOR2xp5_ASAP7_75t_L g1234 ( 
.A(n_1164),
.B(n_870),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1123),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1110),
.B(n_748),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1077),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1123),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1079),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1126),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1126),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1140),
.B(n_751),
.Y(n_1242)
);

XOR2xp5_ASAP7_75t_L g1243 ( 
.A(n_1164),
.B(n_886),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1119),
.B(n_1018),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_1153),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1079),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1132),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_SL g1248 ( 
.A(n_1153),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1075),
.B(n_1082),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1146),
.B(n_886),
.Y(n_1250)
);

XNOR2xp5_ASAP7_75t_L g1251 ( 
.A(n_1091),
.B(n_894),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1139),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1139),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1085),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1145),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1085),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1145),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1144),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1144),
.Y(n_1259)
);

XOR2xp5_ASAP7_75t_L g1260 ( 
.A(n_1108),
.B(n_894),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1086),
.Y(n_1261)
);

XNOR2xp5_ASAP7_75t_L g1262 ( 
.A(n_1168),
.B(n_904),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1130),
.Y(n_1263)
);

NAND2xp33_ASAP7_75t_R g1264 ( 
.A(n_1108),
.B(n_947),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1082),
.B(n_898),
.Y(n_1265)
);

NOR2xp67_ASAP7_75t_L g1266 ( 
.A(n_1152),
.B(n_867),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1086),
.Y(n_1267)
);

INVxp67_ASAP7_75t_L g1268 ( 
.A(n_1080),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1087),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1097),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1097),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1102),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1102),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1111),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1111),
.Y(n_1275)
);

NAND2x1p5_ASAP7_75t_L g1276 ( 
.A(n_1151),
.B(n_1018),
.Y(n_1276)
);

INVxp33_ASAP7_75t_SL g1277 ( 
.A(n_1143),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1146),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1115),
.B(n_751),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1081),
.B(n_773),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1189),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1189),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1073),
.Y(n_1283)
);

CKINVDCx20_ASAP7_75t_R g1284 ( 
.A(n_1199),
.Y(n_1284)
);

CKINVDCx20_ASAP7_75t_R g1285 ( 
.A(n_1153),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1072),
.B(n_911),
.Y(n_1286)
);

XOR2xp5_ASAP7_75t_L g1287 ( 
.A(n_1072),
.B(n_911),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1192),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1099),
.B(n_912),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_1073),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1100),
.B(n_912),
.Y(n_1291)
);

XNOR2xp5_ASAP7_75t_L g1292 ( 
.A(n_1109),
.B(n_913),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1192),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1149),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_SL g1295 ( 
.A(n_1107),
.B(n_987),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1150),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1113),
.Y(n_1297)
);

OR2x2_ASAP7_75t_L g1298 ( 
.A(n_1134),
.B(n_1142),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1073),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1134),
.B(n_913),
.Y(n_1300)
);

INVxp33_ASAP7_75t_L g1301 ( 
.A(n_1148),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1103),
.Y(n_1302)
);

NOR2x1p5_ASAP7_75t_L g1303 ( 
.A(n_1128),
.B(n_1103),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1176),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1105),
.B(n_1031),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1176),
.Y(n_1306)
);

XNOR2xp5_ASAP7_75t_L g1307 ( 
.A(n_1135),
.B(n_947),
.Y(n_1307)
);

INVx4_ASAP7_75t_L g1308 ( 
.A(n_1106),
.Y(n_1308)
);

XNOR2xp5_ASAP7_75t_L g1309 ( 
.A(n_1135),
.B(n_1194),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1166),
.Y(n_1310)
);

CKINVDCx16_ASAP7_75t_R g1311 ( 
.A(n_1160),
.Y(n_1311)
);

BUFx5_ASAP7_75t_L g1312 ( 
.A(n_1173),
.Y(n_1312)
);

AOI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1158),
.A2(n_896),
.B(n_876),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1166),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1172),
.Y(n_1315)
);

INVxp33_ASAP7_75t_L g1316 ( 
.A(n_1131),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1172),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1174),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1174),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1105),
.B(n_1031),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1175),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1175),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1179),
.Y(n_1323)
);

XOR2xp5_ASAP7_75t_L g1324 ( 
.A(n_1120),
.B(n_773),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1179),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1183),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1183),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1190),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1196),
.B(n_775),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1190),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_L g1331 ( 
.A(n_1196),
.B(n_775),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1160),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1105),
.B(n_1155),
.Y(n_1333)
);

XOR2xp5_ASAP7_75t_L g1334 ( 
.A(n_1120),
.B(n_797),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_SL g1335 ( 
.A(n_1180),
.B(n_797),
.Y(n_1335)
);

OR2x2_ASAP7_75t_L g1336 ( 
.A(n_1199),
.B(n_875),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1195),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1162),
.B(n_798),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1155),
.B(n_1041),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1157),
.B(n_1041),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1116),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1170),
.Y(n_1342)
);

XOR2xp5_ASAP7_75t_L g1343 ( 
.A(n_1133),
.B(n_798),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1182),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1194),
.B(n_877),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1116),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1185),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_1160),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1187),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1193),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1163),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1116),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1137),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1137),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1137),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1188),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1188),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1188),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1200),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1194),
.B(n_878),
.Y(n_1360)
);

INVx1_ASAP7_75t_SL g1361 ( 
.A(n_1194),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1169),
.B(n_879),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1169),
.B(n_880),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1154),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1154),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1171),
.Y(n_1366)
);

INVxp67_ASAP7_75t_SL g1367 ( 
.A(n_1157),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1171),
.Y(n_1368)
);

INVxp67_ASAP7_75t_L g1369 ( 
.A(n_1136),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1171),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1122),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1184),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1106),
.B(n_807),
.Y(n_1373)
);

INVxp67_ASAP7_75t_L g1374 ( 
.A(n_1106),
.Y(n_1374)
);

OAI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1161),
.A2(n_1058),
.B(n_1041),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1161),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_1198),
.Y(n_1377)
);

XNOR2x2_ASAP7_75t_L g1378 ( 
.A(n_1156),
.B(n_693),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1158),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1147),
.Y(n_1380)
);

XOR2x2_ASAP7_75t_L g1381 ( 
.A(n_1159),
.B(n_972),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1147),
.Y(n_1382)
);

XNOR2xp5_ASAP7_75t_L g1383 ( 
.A(n_1167),
.B(n_807),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1268),
.B(n_1173),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1367),
.A2(n_1151),
.B1(n_1165),
.B2(n_1180),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1268),
.B(n_1112),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_1377),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1202),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1367),
.B(n_1165),
.Y(n_1389)
);

AND2x6_ASAP7_75t_SL g1390 ( 
.A(n_1280),
.B(n_680),
.Y(n_1390)
);

BUFx6f_ASAP7_75t_L g1391 ( 
.A(n_1283),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1203),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1249),
.B(n_1112),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_SL g1394 ( 
.A(n_1335),
.B(n_1316),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_SL g1395 ( 
.A(n_1335),
.B(n_1107),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1261),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1267),
.Y(n_1397)
);

AND2x6_ASAP7_75t_SL g1398 ( 
.A(n_1280),
.B(n_681),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1269),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1277),
.B(n_972),
.Y(n_1400)
);

INVx2_ASAP7_75t_SL g1401 ( 
.A(n_1206),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_SL g1402 ( 
.A(n_1316),
.B(n_1107),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_SL g1403 ( 
.A(n_1278),
.B(n_1369),
.Y(n_1403)
);

NOR2xp33_ASAP7_75t_L g1404 ( 
.A(n_1236),
.B(n_1197),
.Y(n_1404)
);

BUFx3_ASAP7_75t_L g1405 ( 
.A(n_1263),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1281),
.B(n_1112),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1206),
.B(n_873),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1282),
.B(n_1112),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1288),
.B(n_1141),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1293),
.B(n_1141),
.Y(n_1410)
);

INVxp33_ASAP7_75t_L g1411 ( 
.A(n_1286),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1270),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1236),
.B(n_909),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1300),
.Y(n_1414)
);

NOR2xp67_ASAP7_75t_L g1415 ( 
.A(n_1369),
.B(n_1177),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_SL g1416 ( 
.A(n_1298),
.B(n_1124),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_SL g1417 ( 
.A(n_1283),
.B(n_1290),
.Y(n_1417)
);

OR2x2_ASAP7_75t_L g1418 ( 
.A(n_1250),
.B(n_1242),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_L g1419 ( 
.A(n_1242),
.B(n_1141),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1271),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1338),
.B(n_1141),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1338),
.B(n_1095),
.Y(n_1422)
);

AOI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1211),
.A2(n_1095),
.B1(n_1125),
.B2(n_1178),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1228),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1308),
.B(n_1124),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_SL g1426 ( 
.A(n_1226),
.B(n_1095),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1272),
.Y(n_1427)
);

O2A1O1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1211),
.A2(n_656),
.B(n_649),
.C(n_682),
.Y(n_1428)
);

O2A1O1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1216),
.A2(n_686),
.B(n_701),
.C(n_697),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1204),
.B(n_1095),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1329),
.B(n_724),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1329),
.B(n_605),
.Y(n_1432)
);

AO22x1_ASAP7_75t_L g1433 ( 
.A1(n_1279),
.A2(n_618),
.B1(n_624),
.B2(n_619),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1331),
.B(n_608),
.Y(n_1434)
);

AOI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1216),
.A2(n_1279),
.B1(n_1210),
.B2(n_1303),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1324),
.A2(n_1334),
.B1(n_1259),
.B2(n_1258),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1208),
.B(n_1198),
.Y(n_1437)
);

INVx5_ASAP7_75t_L g1438 ( 
.A(n_1290),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1209),
.B(n_1198),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1215),
.B(n_1198),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1218),
.B(n_1041),
.Y(n_1441)
);

OAI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1301),
.A2(n_619),
.B1(n_626),
.B2(n_624),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_1308),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1219),
.B(n_1058),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_SL g1445 ( 
.A(n_1309),
.B(n_794),
.Y(n_1445)
);

INVxp67_ASAP7_75t_L g1446 ( 
.A(n_1289),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1331),
.B(n_612),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1273),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1359),
.B(n_1058),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1376),
.B(n_1058),
.Y(n_1450)
);

INVxp67_ASAP7_75t_L g1451 ( 
.A(n_1291),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_SL g1452 ( 
.A(n_1371),
.B(n_636),
.Y(n_1452)
);

NOR2xp67_ASAP7_75t_SL g1453 ( 
.A(n_1311),
.B(n_642),
.Y(n_1453)
);

AO22x1_ASAP7_75t_L g1454 ( 
.A1(n_1225),
.A2(n_630),
.B1(n_710),
.B2(n_626),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1223),
.B(n_1125),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1330),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_SL g1457 ( 
.A(n_1361),
.B(n_643),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1260),
.B(n_899),
.Y(n_1458)
);

BUFx8_ASAP7_75t_L g1459 ( 
.A(n_1248),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1230),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_1201),
.Y(n_1461)
);

AOI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1210),
.A2(n_644),
.B1(n_651),
.B2(n_646),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1225),
.B(n_1301),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_L g1464 ( 
.A(n_1343),
.B(n_635),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1362),
.A2(n_676),
.B1(n_689),
.B2(n_663),
.Y(n_1465)
);

NOR3xp33_ASAP7_75t_L g1466 ( 
.A(n_1373),
.B(n_903),
.C(n_901),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1229),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1361),
.B(n_708),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1244),
.A2(n_1186),
.B(n_1191),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1287),
.B(n_647),
.Y(n_1470)
);

INVx3_ASAP7_75t_L g1471 ( 
.A(n_1276),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_SL g1472 ( 
.A(n_1274),
.B(n_716),
.Y(n_1472)
);

A2O1A1Ixp33_ASAP7_75t_L g1473 ( 
.A1(n_1224),
.A2(n_1191),
.B(n_705),
.C(n_707),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1275),
.B(n_745),
.Y(n_1474)
);

AND2x6_ASAP7_75t_SL g1475 ( 
.A(n_1373),
.B(n_704),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1363),
.B(n_755),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_SL g1477 ( 
.A1(n_1243),
.A2(n_630),
.B1(n_710),
.B2(n_627),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1383),
.B(n_648),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1284),
.B(n_654),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1297),
.B(n_757),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1294),
.B(n_765),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_1201),
.B(n_806),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1296),
.B(n_987),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_SL g1484 ( 
.A(n_1265),
.B(n_987),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1378),
.A2(n_789),
.B1(n_804),
.B2(n_782),
.Y(n_1485)
);

AND2x2_ASAP7_75t_SL g1486 ( 
.A(n_1336),
.B(n_789),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_SL g1487 ( 
.A(n_1265),
.B(n_987),
.Y(n_1487)
);

BUFx6f_ASAP7_75t_L g1488 ( 
.A(n_1299),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1284),
.B(n_659),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1231),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_L g1491 ( 
.A(n_1234),
.B(n_660),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1232),
.B(n_992),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1233),
.B(n_992),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_SL g1494 ( 
.A(n_1226),
.B(n_664),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1235),
.B(n_1238),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1292),
.B(n_661),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1240),
.B(n_992),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1241),
.B(n_999),
.Y(n_1498)
);

BUFx6f_ASAP7_75t_SL g1499 ( 
.A(n_1205),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1247),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1262),
.B(n_662),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1252),
.B(n_999),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1253),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1255),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1257),
.B(n_999),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1213),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1207),
.B(n_665),
.Y(n_1507)
);

INVx2_ASAP7_75t_SL g1508 ( 
.A(n_1205),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_SL g1509 ( 
.A(n_1312),
.B(n_1001),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_SL g1510 ( 
.A(n_1345),
.B(n_1001),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_SL g1511 ( 
.A(n_1360),
.B(n_1016),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1220),
.B(n_1016),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1304),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1306),
.Y(n_1514)
);

BUFx3_ASAP7_75t_L g1515 ( 
.A(n_1227),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_1227),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1372),
.B(n_1016),
.Y(n_1517)
);

O2A1O1Ixp33_ASAP7_75t_L g1518 ( 
.A1(n_1342),
.A2(n_712),
.B(n_713),
.C(n_711),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1333),
.A2(n_804),
.B1(n_714),
.B2(n_725),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1205),
.B(n_666),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1344),
.B(n_1019),
.Y(n_1521)
);

BUFx12f_ASAP7_75t_L g1522 ( 
.A(n_1245),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1374),
.B(n_668),
.Y(n_1523)
);

INVxp67_ASAP7_75t_L g1524 ( 
.A(n_1266),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1347),
.B(n_1019),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1349),
.B(n_1032),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1374),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_L g1528 ( 
.A(n_1332),
.B(n_670),
.Y(n_1528)
);

OR2x6_ASAP7_75t_L g1529 ( 
.A(n_1302),
.B(n_1186),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1221),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1237),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1350),
.B(n_1032),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1351),
.B(n_1333),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1239),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1348),
.B(n_664),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1246),
.B(n_1033),
.Y(n_1536)
);

NOR2xp33_ASAP7_75t_L g1537 ( 
.A(n_1251),
.B(n_1307),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_1341),
.B(n_1033),
.Y(n_1538)
);

AOI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1264),
.A2(n_1035),
.B1(n_1048),
.B2(n_1033),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_1214),
.Y(n_1540)
);

INVxp67_ASAP7_75t_SL g1541 ( 
.A(n_1339),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1254),
.B(n_1035),
.Y(n_1542)
);

AOI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1364),
.A2(n_1048),
.B1(n_1050),
.B2(n_1035),
.Y(n_1543)
);

AND2x6_ASAP7_75t_SL g1544 ( 
.A(n_1217),
.B(n_723),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1256),
.B(n_1035),
.Y(n_1545)
);

OAI21xp33_ASAP7_75t_L g1546 ( 
.A1(n_1222),
.A2(n_791),
.B(n_627),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1365),
.A2(n_727),
.B1(n_737),
.B2(n_729),
.Y(n_1547)
);

INVxp67_ASAP7_75t_L g1548 ( 
.A(n_1248),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1305),
.B(n_1048),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_SL g1550 ( 
.A(n_1346),
.B(n_1048),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1381),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1320),
.B(n_1050),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1320),
.B(n_1050),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1339),
.B(n_1050),
.Y(n_1554)
);

NOR2xp67_ASAP7_75t_L g1555 ( 
.A(n_1366),
.B(n_463),
.Y(n_1555)
);

INVxp33_ASAP7_75t_L g1556 ( 
.A(n_1285),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1340),
.B(n_1050),
.Y(n_1557)
);

NAND3xp33_ASAP7_75t_L g1558 ( 
.A(n_1368),
.B(n_674),
.C(n_673),
.Y(n_1558)
);

AOI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1370),
.A2(n_907),
.B1(n_908),
.B2(n_905),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_SL g1560 ( 
.A(n_1217),
.B(n_687),
.Y(n_1560)
);

INVx3_ASAP7_75t_L g1561 ( 
.A(n_1425),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_L g1562 ( 
.A(n_1463),
.B(n_1310),
.Y(n_1562)
);

OAI321xp33_ASAP7_75t_L g1563 ( 
.A1(n_1507),
.A2(n_739),
.A3(n_738),
.B1(n_754),
.B2(n_750),
.C(n_747),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_SL g1564 ( 
.A(n_1486),
.B(n_1352),
.Y(n_1564)
);

AO21x1_ASAP7_75t_L g1565 ( 
.A1(n_1404),
.A2(n_1382),
.B(n_1212),
.Y(n_1565)
);

INVx3_ASAP7_75t_L g1566 ( 
.A(n_1425),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1389),
.A2(n_1375),
.B(n_1295),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1413),
.B(n_1314),
.Y(n_1568)
);

AOI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1385),
.A2(n_1295),
.B(n_1340),
.Y(n_1569)
);

OAI21xp5_ASAP7_75t_L g1570 ( 
.A1(n_1422),
.A2(n_1212),
.B(n_1380),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1388),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1392),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1533),
.A2(n_1379),
.B1(n_1317),
.B2(n_1318),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1418),
.B(n_1407),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1419),
.B(n_1315),
.Y(n_1575)
);

AOI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1385),
.A2(n_1321),
.B(n_1319),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_SL g1577 ( 
.A(n_1401),
.B(n_1353),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_1516),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1431),
.B(n_1322),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1513),
.Y(n_1580)
);

AOI21xp5_ASAP7_75t_L g1581 ( 
.A1(n_1469),
.A2(n_1325),
.B(n_1323),
.Y(n_1581)
);

INVx3_ASAP7_75t_L g1582 ( 
.A(n_1393),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1432),
.B(n_1326),
.Y(n_1583)
);

A2O1A1Ixp33_ASAP7_75t_L g1584 ( 
.A1(n_1434),
.A2(n_1328),
.B(n_1337),
.C(n_1327),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1447),
.B(n_1354),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1435),
.B(n_1355),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1514),
.A2(n_1357),
.B1(n_1358),
.B2(n_1356),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1421),
.B(n_1313),
.Y(n_1588)
);

AOI21xp33_ASAP7_75t_L g1589 ( 
.A1(n_1429),
.A2(n_916),
.B(n_914),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_1540),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1478),
.A2(n_816),
.B1(n_687),
.B2(n_764),
.Y(n_1591)
);

AOI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1541),
.A2(n_940),
.B(n_939),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_1405),
.Y(n_1593)
);

INVxp67_ASAP7_75t_L g1594 ( 
.A(n_1424),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1414),
.B(n_756),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1461),
.B(n_1443),
.Y(n_1596)
);

BUFx6f_ASAP7_75t_L g1597 ( 
.A(n_1387),
.Y(n_1597)
);

INVx2_ASAP7_75t_SL g1598 ( 
.A(n_1387),
.Y(n_1598)
);

O2A1O1Ixp33_ASAP7_75t_L g1599 ( 
.A1(n_1428),
.A2(n_786),
.B(n_793),
.C(n_788),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_SL g1600 ( 
.A(n_1461),
.B(n_719),
.Y(n_1600)
);

INVx1_ASAP7_75t_SL g1601 ( 
.A(n_1467),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1384),
.B(n_795),
.Y(n_1602)
);

NOR2xp67_ASAP7_75t_L g1603 ( 
.A(n_1524),
.B(n_465),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1446),
.B(n_802),
.Y(n_1604)
);

O2A1O1Ixp5_ASAP7_75t_L g1605 ( 
.A1(n_1395),
.A2(n_803),
.B(n_812),
.C(n_808),
.Y(n_1605)
);

AOI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1496),
.A2(n_677),
.B1(n_678),
.B2(n_675),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_L g1607 ( 
.A(n_1411),
.B(n_679),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1451),
.B(n_813),
.Y(n_1608)
);

OAI21xp33_ASAP7_75t_L g1609 ( 
.A1(n_1464),
.A2(n_783),
.B(n_719),
.Y(n_1609)
);

NAND3xp33_ASAP7_75t_L g1610 ( 
.A(n_1501),
.B(n_685),
.C(n_683),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1476),
.B(n_817),
.Y(n_1611)
);

AOI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1491),
.A2(n_691),
.B1(n_700),
.B2(n_695),
.Y(n_1612)
);

AOI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1549),
.A2(n_1553),
.B(n_1552),
.Y(n_1613)
);

INVx1_ASAP7_75t_SL g1614 ( 
.A(n_1458),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1415),
.B(n_821),
.Y(n_1615)
);

BUFx3_ASAP7_75t_L g1616 ( 
.A(n_1522),
.Y(n_1616)
);

CKINVDCx20_ASAP7_75t_R g1617 ( 
.A(n_1459),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_SL g1618 ( 
.A(n_1461),
.B(n_783),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1456),
.Y(n_1619)
);

BUFx3_ASAP7_75t_L g1620 ( 
.A(n_1443),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1386),
.B(n_823),
.Y(n_1621)
);

BUFx2_ASAP7_75t_L g1622 ( 
.A(n_1527),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1393),
.Y(n_1623)
);

OAI321xp33_ASAP7_75t_L g1624 ( 
.A1(n_1477),
.A2(n_816),
.A3(n_687),
.B1(n_826),
.B2(n_827),
.C(n_791),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1403),
.Y(n_1625)
);

O2A1O1Ixp5_ASAP7_75t_L g1626 ( 
.A1(n_1394),
.A2(n_1000),
.B(n_1068),
.C(n_816),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1480),
.B(n_703),
.Y(n_1627)
);

AOI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1552),
.A2(n_940),
.B(n_939),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_SL g1629 ( 
.A(n_1479),
.B(n_1489),
.Y(n_1629)
);

AOI21xp5_ASAP7_75t_L g1630 ( 
.A1(n_1553),
.A2(n_952),
.B(n_946),
.Y(n_1630)
);

OR2x6_ASAP7_75t_SL g1631 ( 
.A(n_1436),
.B(n_1558),
.Y(n_1631)
);

O2A1O1Ixp33_ASAP7_75t_L g1632 ( 
.A1(n_1436),
.A2(n_709),
.B(n_717),
.C(n_706),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1445),
.B(n_728),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1547),
.B(n_730),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1406),
.B(n_826),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1466),
.B(n_731),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1408),
.B(n_827),
.Y(n_1637)
);

OAI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1554),
.A2(n_733),
.B(n_732),
.Y(n_1638)
);

OAI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1554),
.A2(n_740),
.B(n_735),
.Y(n_1639)
);

AOI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1430),
.A2(n_952),
.B(n_946),
.Y(n_1640)
);

O2A1O1Ixp5_ASAP7_75t_L g1641 ( 
.A1(n_1519),
.A2(n_1452),
.B(n_1416),
.C(n_1402),
.Y(n_1641)
);

INVx3_ASAP7_75t_L g1642 ( 
.A(n_1391),
.Y(n_1642)
);

BUFx3_ASAP7_75t_L g1643 ( 
.A(n_1443),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1409),
.B(n_741),
.Y(n_1644)
);

BUFx3_ASAP7_75t_L g1645 ( 
.A(n_1387),
.Y(n_1645)
);

OAI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1557),
.A2(n_743),
.B(n_742),
.Y(n_1646)
);

A2O1A1Ixp33_ASAP7_75t_L g1647 ( 
.A1(n_1559),
.A2(n_753),
.B(n_760),
.C(n_744),
.Y(n_1647)
);

BUFx2_ASAP7_75t_L g1648 ( 
.A(n_1515),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1410),
.B(n_761),
.Y(n_1649)
);

OAI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1557),
.A2(n_763),
.B(n_762),
.Y(n_1650)
);

OAI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1423),
.A2(n_768),
.B(n_766),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_SL g1652 ( 
.A(n_1528),
.B(n_769),
.Y(n_1652)
);

AOI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1509),
.A2(n_959),
.B(n_974),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1396),
.Y(n_1654)
);

O2A1O1Ixp5_ASAP7_75t_L g1655 ( 
.A1(n_1519),
.A2(n_1068),
.B(n_1000),
.C(n_2),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1470),
.B(n_770),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1397),
.B(n_772),
.Y(n_1657)
);

OAI21xp5_ASAP7_75t_L g1658 ( 
.A1(n_1512),
.A2(n_776),
.B(n_774),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1494),
.B(n_1535),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1399),
.B(n_777),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_SL g1661 ( 
.A(n_1426),
.B(n_778),
.Y(n_1661)
);

AOI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1455),
.A2(n_974),
.B(n_1000),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1481),
.B(n_779),
.Y(n_1663)
);

O2A1O1Ixp33_ASAP7_75t_L g1664 ( 
.A1(n_1546),
.A2(n_781),
.B(n_799),
.C(n_780),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1420),
.B(n_800),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1400),
.B(n_805),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1555),
.A2(n_976),
.B(n_975),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1427),
.B(n_810),
.Y(n_1668)
);

AOI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1537),
.A2(n_814),
.B1(n_815),
.B2(n_811),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1448),
.B(n_818),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1460),
.B(n_822),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1506),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1474),
.B(n_976),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_SL g1674 ( 
.A(n_1508),
.B(n_983),
.Y(n_1674)
);

INVx4_ASAP7_75t_L g1675 ( 
.A(n_1438),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1517),
.A2(n_983),
.B(n_467),
.Y(n_1676)
);

AOI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1437),
.A2(n_983),
.B(n_468),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1490),
.Y(n_1678)
);

AOI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1439),
.A2(n_983),
.B(n_469),
.Y(n_1679)
);

INVx3_ASAP7_75t_L g1680 ( 
.A(n_1391),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1500),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_SL g1682 ( 
.A(n_1520),
.B(n_0),
.Y(n_1682)
);

AOI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1440),
.A2(n_472),
.B(n_466),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_SL g1684 ( 
.A(n_1560),
.B(n_1488),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1503),
.B(n_1),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1504),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1495),
.A2(n_475),
.B(n_474),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1488),
.B(n_2),
.Y(n_1688)
);

INVx8_ASAP7_75t_L g1689 ( 
.A(n_1438),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1412),
.B(n_3),
.Y(n_1690)
);

AOI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1484),
.A2(n_479),
.B(n_478),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1438),
.B(n_480),
.Y(n_1692)
);

INVx3_ASAP7_75t_L g1693 ( 
.A(n_1391),
.Y(n_1693)
);

BUFx2_ASAP7_75t_SL g1694 ( 
.A(n_1438),
.Y(n_1694)
);

INVx3_ASAP7_75t_L g1695 ( 
.A(n_1529),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1433),
.B(n_3),
.Y(n_1696)
);

OAI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1449),
.A2(n_484),
.B(n_482),
.Y(n_1697)
);

INVxp67_ASAP7_75t_L g1698 ( 
.A(n_1523),
.Y(n_1698)
);

BUFx2_ASAP7_75t_L g1699 ( 
.A(n_1548),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1454),
.B(n_4),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1485),
.B(n_5),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1530),
.B(n_1534),
.Y(n_1702)
);

A2O1A1Ixp33_ASAP7_75t_L g1703 ( 
.A1(n_1473),
.A2(n_1518),
.B(n_1472),
.C(n_1462),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1531),
.B(n_5),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1465),
.B(n_6),
.Y(n_1705)
);

AOI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1487),
.A2(n_486),
.B(n_485),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1449),
.A2(n_488),
.B(n_487),
.Y(n_1707)
);

AOI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1543),
.A2(n_492),
.B(n_491),
.Y(n_1708)
);

BUFx6f_ASAP7_75t_L g1709 ( 
.A(n_1488),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_SL g1710 ( 
.A(n_1442),
.B(n_7),
.Y(n_1710)
);

AOI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1510),
.A2(n_494),
.B(n_493),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1450),
.Y(n_1712)
);

AOI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1511),
.A2(n_496),
.B(n_495),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_SL g1714 ( 
.A(n_1459),
.B(n_498),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1482),
.B(n_7),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1441),
.Y(n_1716)
);

AOI21xp5_ASAP7_75t_L g1717 ( 
.A1(n_1492),
.A2(n_499),
.B(n_497),
.Y(n_1717)
);

O2A1O1Ixp5_ASAP7_75t_L g1718 ( 
.A1(n_1457),
.A2(n_10),
.B(n_8),
.C(n_9),
.Y(n_1718)
);

INVx3_ASAP7_75t_L g1719 ( 
.A(n_1529),
.Y(n_1719)
);

AOI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1493),
.A2(n_503),
.B(n_501),
.Y(n_1720)
);

NOR2xp67_ASAP7_75t_L g1721 ( 
.A(n_1468),
.B(n_592),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1450),
.Y(n_1722)
);

AOI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1497),
.A2(n_506),
.B(n_505),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1444),
.B(n_1471),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1542),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1471),
.B(n_9),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1556),
.B(n_10),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1483),
.Y(n_1728)
);

AOI21xp33_ASAP7_75t_L g1729 ( 
.A1(n_1521),
.A2(n_1526),
.B(n_1525),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1574),
.B(n_1551),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1580),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1562),
.B(n_1390),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_SL g1733 ( 
.A(n_1698),
.B(n_1539),
.Y(n_1733)
);

INVxp67_ASAP7_75t_L g1734 ( 
.A(n_1622),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1579),
.B(n_1398),
.Y(n_1735)
);

OAI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1629),
.A2(n_1499),
.B1(n_1532),
.B2(n_1417),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1568),
.B(n_1453),
.Y(n_1737)
);

AOI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1567),
.A2(n_1502),
.B(n_1498),
.Y(n_1738)
);

AOI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1613),
.A2(n_1505),
.B(n_1542),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1656),
.B(n_1475),
.Y(n_1740)
);

O2A1O1Ixp33_ASAP7_75t_SL g1741 ( 
.A1(n_1703),
.A2(n_1550),
.B(n_1538),
.C(n_1545),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1583),
.B(n_1545),
.Y(n_1742)
);

AND2x4_ASAP7_75t_L g1743 ( 
.A(n_1596),
.B(n_1536),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1701),
.B(n_11),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1585),
.B(n_1544),
.Y(n_1745)
);

INVx5_ASAP7_75t_L g1746 ( 
.A(n_1689),
.Y(n_1746)
);

AOI221xp5_ASAP7_75t_L g1747 ( 
.A1(n_1599),
.A2(n_15),
.B1(n_11),
.B2(n_13),
.C(n_16),
.Y(n_1747)
);

BUFx12f_ASAP7_75t_L g1748 ( 
.A(n_1590),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1571),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_SL g1750 ( 
.A(n_1614),
.B(n_1625),
.Y(n_1750)
);

CKINVDCx20_ASAP7_75t_R g1751 ( 
.A(n_1617),
.Y(n_1751)
);

AOI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1666),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1619),
.Y(n_1753)
);

OAI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1601),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_1754)
);

AOI21xp5_ASAP7_75t_L g1755 ( 
.A1(n_1570),
.A2(n_513),
.B(n_511),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1631),
.B(n_514),
.Y(n_1756)
);

AOI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1569),
.A2(n_590),
.B(n_516),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1594),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_1578),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1635),
.B(n_21),
.Y(n_1760)
);

AOI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1575),
.A2(n_517),
.B(n_515),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1572),
.Y(n_1762)
);

AOI21xp5_ASAP7_75t_L g1763 ( 
.A1(n_1575),
.A2(n_519),
.B(n_518),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_SL g1764 ( 
.A(n_1563),
.B(n_1633),
.Y(n_1764)
);

AOI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1581),
.A2(n_522),
.B(n_520),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1635),
.B(n_22),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1637),
.B(n_22),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1637),
.B(n_23),
.Y(n_1768)
);

BUFx2_ASAP7_75t_L g1769 ( 
.A(n_1593),
.Y(n_1769)
);

AOI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1588),
.A2(n_588),
.B(n_525),
.Y(n_1770)
);

AOI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1584),
.A2(n_587),
.B(n_529),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1727),
.B(n_23),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1610),
.B(n_530),
.Y(n_1773)
);

A2O1A1Ixp33_ASAP7_75t_L g1774 ( 
.A1(n_1632),
.A2(n_26),
.B(n_24),
.C(n_25),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1644),
.B(n_25),
.Y(n_1775)
);

AND2x4_ASAP7_75t_L g1776 ( 
.A(n_1596),
.B(n_531),
.Y(n_1776)
);

BUFx6f_ASAP7_75t_L g1777 ( 
.A(n_1597),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1644),
.B(n_27),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_SL g1779 ( 
.A(n_1714),
.B(n_28),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1636),
.B(n_28),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1654),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1652),
.B(n_532),
.Y(n_1782)
);

OAI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1564),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_1783)
);

OAI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1591),
.A2(n_32),
.B1(n_29),
.B2(n_31),
.Y(n_1784)
);

BUFx4f_ASAP7_75t_L g1785 ( 
.A(n_1689),
.Y(n_1785)
);

AOI22xp33_ASAP7_75t_L g1786 ( 
.A1(n_1710),
.A2(n_1682),
.B1(n_1705),
.B2(n_1609),
.Y(n_1786)
);

A2O1A1Ixp33_ASAP7_75t_L g1787 ( 
.A1(n_1641),
.A2(n_35),
.B(n_33),
.C(n_34),
.Y(n_1787)
);

AOI21xp5_ASAP7_75t_L g1788 ( 
.A1(n_1573),
.A2(n_535),
.B(n_534),
.Y(n_1788)
);

OAI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1678),
.A2(n_1681),
.B1(n_1686),
.B2(n_1696),
.Y(n_1789)
);

AOI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1659),
.A2(n_1607),
.B1(n_1715),
.B2(n_1684),
.Y(n_1790)
);

BUFx12f_ASAP7_75t_L g1791 ( 
.A(n_1597),
.Y(n_1791)
);

BUFx12f_ASAP7_75t_L g1792 ( 
.A(n_1597),
.Y(n_1792)
);

OAI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1627),
.A2(n_1663),
.B1(n_1634),
.B2(n_1649),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1649),
.B(n_34),
.Y(n_1794)
);

OAI22xp5_ASAP7_75t_L g1795 ( 
.A1(n_1611),
.A2(n_1586),
.B1(n_1602),
.B2(n_1657),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_SL g1796 ( 
.A(n_1648),
.B(n_36),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1621),
.B(n_37),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_SL g1798 ( 
.A(n_1615),
.B(n_37),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1638),
.B(n_38),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_L g1800 ( 
.A(n_1624),
.B(n_537),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1638),
.B(n_39),
.Y(n_1801)
);

AOI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1721),
.A2(n_1612),
.B1(n_1606),
.B2(n_1669),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1600),
.B(n_538),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1603),
.B(n_39),
.Y(n_1804)
);

AOI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1673),
.A2(n_586),
.B(n_543),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1639),
.B(n_40),
.Y(n_1806)
);

AOI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1618),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_1807)
);

AOI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1576),
.A2(n_585),
.B(n_545),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1699),
.B(n_542),
.Y(n_1809)
);

OAI22xp5_ASAP7_75t_L g1810 ( 
.A1(n_1657),
.A2(n_44),
.B1(n_41),
.B2(n_43),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_SL g1811 ( 
.A(n_1639),
.B(n_43),
.Y(n_1811)
);

OAI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1660),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_1812)
);

AOI21xp5_ASAP7_75t_L g1813 ( 
.A1(n_1662),
.A2(n_547),
.B(n_546),
.Y(n_1813)
);

A2O1A1Ixp33_ASAP7_75t_SL g1814 ( 
.A1(n_1697),
.A2(n_1651),
.B(n_1708),
.C(n_1646),
.Y(n_1814)
);

AOI22xp33_ASAP7_75t_L g1815 ( 
.A1(n_1651),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_1815)
);

AOI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1640),
.A2(n_551),
.B(n_549),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_L g1817 ( 
.A(n_1582),
.B(n_553),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1672),
.Y(n_1818)
);

AOI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1729),
.A2(n_1679),
.B(n_1677),
.Y(n_1819)
);

OAI21xp33_ASAP7_75t_L g1820 ( 
.A1(n_1700),
.A2(n_51),
.B(n_52),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1702),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1646),
.B(n_1650),
.Y(n_1822)
);

A2O1A1Ixp33_ASAP7_75t_L g1823 ( 
.A1(n_1650),
.A2(n_54),
.B(n_52),
.C(n_53),
.Y(n_1823)
);

AOI21xp5_ASAP7_75t_L g1824 ( 
.A1(n_1729),
.A2(n_584),
.B(n_555),
.Y(n_1824)
);

OAI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1655),
.A2(n_556),
.B(n_554),
.Y(n_1825)
);

AOI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1565),
.A2(n_581),
.B(n_558),
.Y(n_1826)
);

AOI221xp5_ASAP7_75t_L g1827 ( 
.A1(n_1589),
.A2(n_56),
.B1(n_53),
.B2(n_55),
.C(n_57),
.Y(n_1827)
);

NOR2xp33_ASAP7_75t_L g1828 ( 
.A(n_1623),
.B(n_557),
.Y(n_1828)
);

OAI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1660),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_1829)
);

OAI22xp5_ASAP7_75t_L g1830 ( 
.A1(n_1665),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1595),
.B(n_60),
.Y(n_1831)
);

OAI22xp5_ASAP7_75t_L g1832 ( 
.A1(n_1665),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1620),
.B(n_560),
.Y(n_1833)
);

AOI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1676),
.A2(n_580),
.B(n_563),
.Y(n_1834)
);

AOI21xp5_ASAP7_75t_L g1835 ( 
.A1(n_1592),
.A2(n_578),
.B(n_564),
.Y(n_1835)
);

AOI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1628),
.A2(n_577),
.B(n_566),
.Y(n_1836)
);

INVx1_ASAP7_75t_SL g1837 ( 
.A(n_1709),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_L g1838 ( 
.A(n_1688),
.B(n_561),
.Y(n_1838)
);

BUFx3_ASAP7_75t_L g1839 ( 
.A(n_1645),
.Y(n_1839)
);

AOI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1630),
.A2(n_570),
.B(n_568),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1604),
.B(n_64),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1608),
.B(n_64),
.Y(n_1842)
);

O2A1O1Ixp33_ASAP7_75t_L g1843 ( 
.A1(n_1647),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_1843)
);

OAI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1668),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_1844)
);

O2A1O1Ixp33_ASAP7_75t_L g1845 ( 
.A1(n_1589),
.A2(n_71),
.B(n_68),
.C(n_69),
.Y(n_1845)
);

INVx3_ASAP7_75t_L g1846 ( 
.A(n_1689),
.Y(n_1846)
);

INVx3_ASAP7_75t_L g1847 ( 
.A(n_1709),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1658),
.B(n_69),
.Y(n_1848)
);

AOI21xp5_ASAP7_75t_L g1849 ( 
.A1(n_1667),
.A2(n_573),
.B(n_572),
.Y(n_1849)
);

A2O1A1Ixp33_ASAP7_75t_L g1850 ( 
.A1(n_1658),
.A2(n_73),
.B(n_71),
.C(n_72),
.Y(n_1850)
);

NOR2xp33_ASAP7_75t_L g1851 ( 
.A(n_1726),
.B(n_74),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_SL g1852 ( 
.A(n_1709),
.B(n_74),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1716),
.B(n_76),
.Y(n_1853)
);

AOI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1724),
.A2(n_1728),
.B(n_1687),
.Y(n_1854)
);

NOR2x1_ASAP7_75t_L g1855 ( 
.A(n_1675),
.B(n_76),
.Y(n_1855)
);

AOI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1712),
.A2(n_77),
.B(n_78),
.Y(n_1856)
);

OR2x6_ASAP7_75t_L g1857 ( 
.A(n_1695),
.B(n_79),
.Y(n_1857)
);

BUFx3_ASAP7_75t_L g1858 ( 
.A(n_1598),
.Y(n_1858)
);

NOR2xp33_ASAP7_75t_L g1859 ( 
.A(n_1668),
.B(n_80),
.Y(n_1859)
);

BUFx6f_ASAP7_75t_L g1860 ( 
.A(n_1643),
.Y(n_1860)
);

NOR2xp33_ASAP7_75t_L g1861 ( 
.A(n_1670),
.B(n_81),
.Y(n_1861)
);

OAI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1626),
.A2(n_81),
.B(n_82),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1670),
.B(n_83),
.Y(n_1863)
);

OA21x2_ASAP7_75t_L g1864 ( 
.A1(n_1653),
.A2(n_85),
.B(n_86),
.Y(n_1864)
);

OAI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1707),
.A2(n_462),
.B(n_86),
.Y(n_1865)
);

NAND2x1p5_ASAP7_75t_L g1866 ( 
.A(n_1675),
.B(n_1695),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1671),
.B(n_1722),
.Y(n_1867)
);

OAI21xp5_ASAP7_75t_L g1868 ( 
.A1(n_1605),
.A2(n_88),
.B(n_89),
.Y(n_1868)
);

NOR2xp33_ASAP7_75t_L g1869 ( 
.A(n_1671),
.B(n_89),
.Y(n_1869)
);

NOR2x1_ASAP7_75t_L g1870 ( 
.A(n_1694),
.B(n_90),
.Y(n_1870)
);

A2O1A1Ixp33_ASAP7_75t_L g1871 ( 
.A1(n_1718),
.A2(n_1664),
.B(n_1683),
.C(n_1711),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1725),
.B(n_1561),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1561),
.B(n_1566),
.Y(n_1873)
);

NOR2xp33_ASAP7_75t_L g1874 ( 
.A(n_1577),
.B(n_90),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_SL g1875 ( 
.A(n_1685),
.B(n_91),
.Y(n_1875)
);

OR2x6_ASAP7_75t_SL g1876 ( 
.A(n_1704),
.B(n_92),
.Y(n_1876)
);

INVxp67_ASAP7_75t_L g1877 ( 
.A(n_1690),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1566),
.B(n_92),
.Y(n_1878)
);

OAI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1661),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1587),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1587),
.Y(n_1881)
);

INVxp33_ASAP7_75t_SL g1882 ( 
.A(n_1616),
.Y(n_1882)
);

OAI22xp5_ASAP7_75t_L g1883 ( 
.A1(n_1674),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_1883)
);

INVxp67_ASAP7_75t_L g1884 ( 
.A(n_1642),
.Y(n_1884)
);

O2A1O1Ixp5_ASAP7_75t_L g1885 ( 
.A1(n_1822),
.A2(n_1717),
.B(n_1723),
.C(n_1720),
.Y(n_1885)
);

OAI21xp5_ASAP7_75t_L g1886 ( 
.A1(n_1814),
.A2(n_1865),
.B(n_1871),
.Y(n_1886)
);

BUFx6f_ASAP7_75t_L g1887 ( 
.A(n_1860),
.Y(n_1887)
);

INVxp67_ASAP7_75t_SL g1888 ( 
.A(n_1872),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1730),
.B(n_1719),
.Y(n_1889)
);

AOI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1740),
.A2(n_1719),
.B1(n_1692),
.B2(n_1713),
.Y(n_1890)
);

INVx1_ASAP7_75t_SL g1891 ( 
.A(n_1750),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1867),
.B(n_1680),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1749),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1762),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1742),
.B(n_1692),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1744),
.B(n_1693),
.Y(n_1896)
);

OAI21xp5_ASAP7_75t_L g1897 ( 
.A1(n_1865),
.A2(n_1764),
.B(n_1787),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1880),
.B(n_1693),
.Y(n_1898)
);

NOR2xp67_ASAP7_75t_SL g1899 ( 
.A(n_1748),
.B(n_1691),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1780),
.B(n_1706),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1737),
.B(n_1756),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1781),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1795),
.B(n_96),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1799),
.B(n_96),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1821),
.B(n_1877),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1793),
.B(n_97),
.Y(n_1906)
);

A2O1A1Ixp33_ASAP7_75t_L g1907 ( 
.A1(n_1802),
.A2(n_99),
.B(n_97),
.C(n_98),
.Y(n_1907)
);

AOI21xp5_ASAP7_75t_L g1908 ( 
.A1(n_1819),
.A2(n_99),
.B(n_100),
.Y(n_1908)
);

NOR3xp33_ASAP7_75t_L g1909 ( 
.A(n_1811),
.B(n_100),
.C(n_101),
.Y(n_1909)
);

AOI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1854),
.A2(n_101),
.B(n_102),
.Y(n_1910)
);

OAI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1825),
.A2(n_103),
.B(n_104),
.Y(n_1911)
);

BUFx2_ASAP7_75t_L g1912 ( 
.A(n_1734),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1731),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1801),
.B(n_106),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1789),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1806),
.B(n_462),
.Y(n_1916)
);

OAI21xp5_ASAP7_75t_L g1917 ( 
.A1(n_1862),
.A2(n_107),
.B(n_108),
.Y(n_1917)
);

BUFx2_ASAP7_75t_L g1918 ( 
.A(n_1847),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1848),
.B(n_109),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1790),
.B(n_109),
.Y(n_1920)
);

NOR2x1_ASAP7_75t_SL g1921 ( 
.A(n_1746),
.B(n_110),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1881),
.B(n_110),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1789),
.Y(n_1923)
);

NAND3xp33_ASAP7_75t_L g1924 ( 
.A(n_1752),
.B(n_111),
.C(n_112),
.Y(n_1924)
);

OAI21x1_ASAP7_75t_L g1925 ( 
.A1(n_1739),
.A2(n_111),
.B(n_113),
.Y(n_1925)
);

AOI21xp5_ASAP7_75t_L g1926 ( 
.A1(n_1738),
.A2(n_113),
.B(n_114),
.Y(n_1926)
);

AND2x4_ASAP7_75t_L g1927 ( 
.A(n_1846),
.B(n_114),
.Y(n_1927)
);

A2O1A1Ixp33_ASAP7_75t_L g1928 ( 
.A1(n_1859),
.A2(n_117),
.B(n_115),
.C(n_116),
.Y(n_1928)
);

AOI21xp5_ASAP7_75t_L g1929 ( 
.A1(n_1757),
.A2(n_115),
.B(n_116),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1733),
.B(n_461),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1851),
.B(n_118),
.Y(n_1931)
);

OAI21x1_ASAP7_75t_L g1932 ( 
.A1(n_1826),
.A2(n_119),
.B(n_120),
.Y(n_1932)
);

OAI21x1_ASAP7_75t_SL g1933 ( 
.A1(n_1862),
.A2(n_119),
.B(n_120),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_L g1934 ( 
.A(n_1732),
.B(n_121),
.Y(n_1934)
);

A2O1A1Ixp33_ASAP7_75t_L g1935 ( 
.A1(n_1861),
.A2(n_123),
.B(n_121),
.C(n_122),
.Y(n_1935)
);

AOI21xp5_ASAP7_75t_L g1936 ( 
.A1(n_1755),
.A2(n_125),
.B(n_126),
.Y(n_1936)
);

OAI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1771),
.A2(n_126),
.B(n_127),
.Y(n_1937)
);

CKINVDCx11_ASAP7_75t_R g1938 ( 
.A(n_1751),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1869),
.B(n_127),
.Y(n_1939)
);

AOI211x1_ASAP7_75t_L g1940 ( 
.A1(n_1758),
.A2(n_131),
.B(n_129),
.C(n_130),
.Y(n_1940)
);

OAI21x1_ASAP7_75t_L g1941 ( 
.A1(n_1765),
.A2(n_132),
.B(n_134),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1753),
.Y(n_1942)
);

OAI22xp5_ASAP7_75t_L g1943 ( 
.A1(n_1815),
.A2(n_1786),
.B1(n_1823),
.B2(n_1850),
.Y(n_1943)
);

OAI21xp5_ASAP7_75t_L g1944 ( 
.A1(n_1788),
.A2(n_135),
.B(n_136),
.Y(n_1944)
);

AND2x4_ASAP7_75t_L g1945 ( 
.A(n_1846),
.B(n_135),
.Y(n_1945)
);

BUFx3_ASAP7_75t_L g1946 ( 
.A(n_1839),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_SL g1947 ( 
.A(n_1745),
.B(n_137),
.Y(n_1947)
);

OAI21x1_ASAP7_75t_L g1948 ( 
.A1(n_1813),
.A2(n_137),
.B(n_138),
.Y(n_1948)
);

A2O1A1Ixp33_ASAP7_75t_L g1949 ( 
.A1(n_1843),
.A2(n_141),
.B(n_139),
.C(n_140),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1818),
.B(n_140),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1775),
.B(n_141),
.Y(n_1951)
);

AOI21xp5_ASAP7_75t_L g1952 ( 
.A1(n_1741),
.A2(n_142),
.B(n_143),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1778),
.B(n_461),
.Y(n_1953)
);

NAND2xp33_ASAP7_75t_L g1954 ( 
.A(n_1759),
.B(n_142),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1853),
.Y(n_1955)
);

AOI21xp5_ASAP7_75t_L g1956 ( 
.A1(n_1808),
.A2(n_144),
.B(n_145),
.Y(n_1956)
);

AOI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1779),
.A2(n_1782),
.B1(n_1773),
.B2(n_1820),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1743),
.B(n_146),
.Y(n_1958)
);

A2O1A1Ixp33_ASAP7_75t_L g1959 ( 
.A1(n_1774),
.A2(n_150),
.B(n_147),
.C(n_148),
.Y(n_1959)
);

AND2x4_ASAP7_75t_L g1960 ( 
.A(n_1746),
.B(n_148),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1794),
.B(n_151),
.Y(n_1961)
);

AOI221x1_ASAP7_75t_L g1962 ( 
.A1(n_1810),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.C(n_154),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1878),
.Y(n_1963)
);

AOI22xp5_ASAP7_75t_L g1964 ( 
.A1(n_1779),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1760),
.B(n_1766),
.Y(n_1965)
);

OAI21x1_ASAP7_75t_L g1966 ( 
.A1(n_1816),
.A2(n_155),
.B(n_156),
.Y(n_1966)
);

OAI21x1_ASAP7_75t_L g1967 ( 
.A1(n_1836),
.A2(n_155),
.B(n_156),
.Y(n_1967)
);

BUFx2_ASAP7_75t_L g1968 ( 
.A(n_1847),
.Y(n_1968)
);

OAI21xp5_ASAP7_75t_L g1969 ( 
.A1(n_1868),
.A2(n_1824),
.B(n_1763),
.Y(n_1969)
);

AOI22xp5_ASAP7_75t_L g1970 ( 
.A1(n_1803),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1772),
.B(n_157),
.Y(n_1971)
);

OAI21x1_ASAP7_75t_L g1972 ( 
.A1(n_1840),
.A2(n_161),
.B(n_162),
.Y(n_1972)
);

OAI21x1_ASAP7_75t_L g1973 ( 
.A1(n_1834),
.A2(n_161),
.B(n_162),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1767),
.B(n_460),
.Y(n_1974)
);

OAI21x1_ASAP7_75t_L g1975 ( 
.A1(n_1835),
.A2(n_163),
.B(n_164),
.Y(n_1975)
);

OAI21x1_ASAP7_75t_L g1976 ( 
.A1(n_1849),
.A2(n_163),
.B(n_164),
.Y(n_1976)
);

INVx3_ASAP7_75t_L g1977 ( 
.A(n_1785),
.Y(n_1977)
);

AOI21xp5_ASAP7_75t_SL g1978 ( 
.A1(n_1868),
.A2(n_165),
.B(n_166),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1864),
.Y(n_1979)
);

AOI21xp5_ASAP7_75t_L g1980 ( 
.A1(n_1770),
.A2(n_165),
.B(n_167),
.Y(n_1980)
);

OAI21x1_ASAP7_75t_L g1981 ( 
.A1(n_1761),
.A2(n_167),
.B(n_168),
.Y(n_1981)
);

AOI21xp5_ASAP7_75t_L g1982 ( 
.A1(n_1805),
.A2(n_1828),
.B(n_1817),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_SL g1983 ( 
.A(n_1736),
.B(n_168),
.Y(n_1983)
);

NAND2x1_ASAP7_75t_L g1984 ( 
.A(n_1743),
.B(n_1857),
.Y(n_1984)
);

BUFx2_ASAP7_75t_L g1985 ( 
.A(n_1791),
.Y(n_1985)
);

BUFx6f_ASAP7_75t_L g1986 ( 
.A(n_1860),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1768),
.B(n_1863),
.Y(n_1987)
);

A2O1A1Ixp33_ASAP7_75t_L g1988 ( 
.A1(n_1838),
.A2(n_171),
.B(n_169),
.C(n_170),
.Y(n_1988)
);

OAI21x1_ASAP7_75t_L g1989 ( 
.A1(n_1866),
.A2(n_1864),
.B(n_1873),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1893),
.Y(n_1990)
);

AOI21xp5_ASAP7_75t_L g1991 ( 
.A1(n_1886),
.A2(n_1804),
.B(n_1845),
.Y(n_1991)
);

AOI21xp5_ASAP7_75t_L g1992 ( 
.A1(n_1886),
.A2(n_1856),
.B(n_1827),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1913),
.Y(n_1993)
);

BUFx12f_ASAP7_75t_L g1994 ( 
.A(n_1938),
.Y(n_1994)
);

NOR3xp33_ASAP7_75t_L g1995 ( 
.A(n_1924),
.B(n_1784),
.C(n_1747),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1915),
.B(n_1874),
.Y(n_1996)
);

CKINVDCx20_ASAP7_75t_R g1997 ( 
.A(n_1946),
.Y(n_1997)
);

OR2x6_ASAP7_75t_L g1998 ( 
.A(n_1911),
.B(n_1857),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1923),
.B(n_1797),
.Y(n_1999)
);

BUFx3_ASAP7_75t_L g2000 ( 
.A(n_1887),
.Y(n_2000)
);

BUFx2_ASAP7_75t_SL g2001 ( 
.A(n_1887),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1888),
.B(n_1875),
.Y(n_2002)
);

AND2x4_ASAP7_75t_L g2003 ( 
.A(n_1894),
.B(n_1746),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1902),
.B(n_1841),
.Y(n_2004)
);

INVx2_ASAP7_75t_SL g2005 ( 
.A(n_1887),
.Y(n_2005)
);

INVx3_ASAP7_75t_L g2006 ( 
.A(n_1889),
.Y(n_2006)
);

NOR2xp33_ASAP7_75t_L g2007 ( 
.A(n_1957),
.B(n_1876),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1901),
.B(n_1896),
.Y(n_2008)
);

OAI22xp5_ASAP7_75t_L g2009 ( 
.A1(n_1924),
.A2(n_1807),
.B1(n_1857),
.B2(n_1829),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1942),
.Y(n_2010)
);

BUFx8_ASAP7_75t_L g2011 ( 
.A(n_1985),
.Y(n_2011)
);

BUFx6f_ASAP7_75t_L g2012 ( 
.A(n_1986),
.Y(n_2012)
);

AOI21xp5_ASAP7_75t_L g2013 ( 
.A1(n_1911),
.A2(n_1785),
.B(n_1776),
.Y(n_2013)
);

BUFx8_ASAP7_75t_SL g2014 ( 
.A(n_1912),
.Y(n_2014)
);

INVx2_ASAP7_75t_SL g2015 ( 
.A(n_1986),
.Y(n_2015)
);

BUFx2_ASAP7_75t_L g2016 ( 
.A(n_1918),
.Y(n_2016)
);

INVx3_ASAP7_75t_L g2017 ( 
.A(n_1986),
.Y(n_2017)
);

OR2x2_ASAP7_75t_SL g2018 ( 
.A(n_1906),
.B(n_1735),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1963),
.B(n_1842),
.Y(n_2019)
);

BUFx2_ASAP7_75t_L g2020 ( 
.A(n_1968),
.Y(n_2020)
);

AND2x4_ASAP7_75t_L g2021 ( 
.A(n_1891),
.B(n_1837),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1891),
.B(n_1831),
.Y(n_2022)
);

BUFx3_ASAP7_75t_L g2023 ( 
.A(n_1977),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1898),
.Y(n_2024)
);

BUFx3_ASAP7_75t_L g2025 ( 
.A(n_1977),
.Y(n_2025)
);

AOI21xp5_ASAP7_75t_L g2026 ( 
.A1(n_1969),
.A2(n_1982),
.B(n_1917),
.Y(n_2026)
);

INVx2_ASAP7_75t_SL g2027 ( 
.A(n_1905),
.Y(n_2027)
);

OR2x2_ASAP7_75t_L g2028 ( 
.A(n_1955),
.B(n_1798),
.Y(n_2028)
);

INVx3_ASAP7_75t_L g2029 ( 
.A(n_1984),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1904),
.B(n_1809),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1898),
.Y(n_2031)
);

BUFx6f_ASAP7_75t_L g2032 ( 
.A(n_1892),
.Y(n_2032)
);

INVx5_ASAP7_75t_L g2033 ( 
.A(n_1960),
.Y(n_2033)
);

OAI22xp5_ASAP7_75t_L g2034 ( 
.A1(n_1907),
.A2(n_1812),
.B1(n_1832),
.B2(n_1830),
.Y(n_2034)
);

INVx1_ASAP7_75t_SL g2035 ( 
.A(n_1965),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1914),
.B(n_1971),
.Y(n_2036)
);

BUFx3_ASAP7_75t_L g2037 ( 
.A(n_1927),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1979),
.Y(n_2038)
);

OAI22xp5_ASAP7_75t_L g2039 ( 
.A1(n_1964),
.A2(n_1844),
.B1(n_1754),
.B2(n_1783),
.Y(n_2039)
);

OAI22xp5_ASAP7_75t_L g2040 ( 
.A1(n_1970),
.A2(n_1800),
.B1(n_1883),
.B2(n_1879),
.Y(n_2040)
);

AOI21xp5_ASAP7_75t_L g2041 ( 
.A1(n_1917),
.A2(n_1776),
.B(n_1852),
.Y(n_2041)
);

OAI21xp5_ASAP7_75t_L g2042 ( 
.A1(n_1936),
.A2(n_1855),
.B(n_1870),
.Y(n_2042)
);

AOI21xp5_ASAP7_75t_L g2043 ( 
.A1(n_1937),
.A2(n_1833),
.B(n_1796),
.Y(n_2043)
);

NAND2x2_ASAP7_75t_L g2044 ( 
.A(n_1903),
.B(n_1858),
.Y(n_2044)
);

BUFx3_ASAP7_75t_L g2045 ( 
.A(n_1927),
.Y(n_2045)
);

AOI21xp5_ASAP7_75t_L g2046 ( 
.A1(n_1937),
.A2(n_1833),
.B(n_1884),
.Y(n_2046)
);

INVx5_ASAP7_75t_L g2047 ( 
.A(n_1960),
.Y(n_2047)
);

INVx6_ASAP7_75t_L g2048 ( 
.A(n_1945),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_SL g2049 ( 
.A(n_1897),
.B(n_1769),
.Y(n_2049)
);

BUFx3_ASAP7_75t_L g2050 ( 
.A(n_1945),
.Y(n_2050)
);

O2A1O1Ixp33_ASAP7_75t_L g2051 ( 
.A1(n_1928),
.A2(n_1882),
.B(n_171),
.C(n_169),
.Y(n_2051)
);

CKINVDCx16_ASAP7_75t_R g2052 ( 
.A(n_1931),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_SL g2053 ( 
.A(n_1890),
.B(n_1860),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_SL g2054 ( 
.A(n_1897),
.B(n_1777),
.Y(n_2054)
);

OR2x2_ASAP7_75t_SL g2055 ( 
.A(n_1987),
.B(n_1777),
.Y(n_2055)
);

BUFx6f_ASAP7_75t_L g2056 ( 
.A(n_2012),
.Y(n_2056)
);

INVx3_ASAP7_75t_L g2057 ( 
.A(n_2029),
.Y(n_2057)
);

CKINVDCx20_ASAP7_75t_R g2058 ( 
.A(n_1997),
.Y(n_2058)
);

BUFx12f_ASAP7_75t_L g2059 ( 
.A(n_1994),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_2006),
.B(n_1989),
.Y(n_2060)
);

AOI22xp33_ASAP7_75t_L g2061 ( 
.A1(n_1995),
.A2(n_1943),
.B1(n_1909),
.B2(n_1944),
.Y(n_2061)
);

CKINVDCx6p67_ASAP7_75t_R g2062 ( 
.A(n_2033),
.Y(n_2062)
);

INVx6_ASAP7_75t_L g2063 ( 
.A(n_2011),
.Y(n_2063)
);

BUFx12f_ASAP7_75t_L g2064 ( 
.A(n_2011),
.Y(n_2064)
);

BUFx3_ASAP7_75t_L g2065 ( 
.A(n_2014),
.Y(n_2065)
);

AOI22xp33_ASAP7_75t_SL g2066 ( 
.A1(n_2009),
.A2(n_1943),
.B1(n_1944),
.B2(n_1954),
.Y(n_2066)
);

BUFx10_ASAP7_75t_L g2067 ( 
.A(n_2012),
.Y(n_2067)
);

CKINVDCx11_ASAP7_75t_R g2068 ( 
.A(n_2044),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1990),
.Y(n_2069)
);

AOI22xp33_ASAP7_75t_SL g2070 ( 
.A1(n_2009),
.A2(n_1933),
.B1(n_1920),
.B2(n_1921),
.Y(n_2070)
);

CKINVDCx20_ASAP7_75t_R g2071 ( 
.A(n_2052),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_2027),
.B(n_1895),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_2038),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1993),
.Y(n_2074)
);

CKINVDCx11_ASAP7_75t_R g2075 ( 
.A(n_2012),
.Y(n_2075)
);

AOI22xp33_ASAP7_75t_L g2076 ( 
.A1(n_1995),
.A2(n_1983),
.B1(n_1934),
.B2(n_1900),
.Y(n_2076)
);

INVx6_ASAP7_75t_L g2077 ( 
.A(n_2033),
.Y(n_2077)
);

OAI22xp5_ASAP7_75t_L g2078 ( 
.A1(n_1998),
.A2(n_1935),
.B1(n_1988),
.B2(n_1959),
.Y(n_2078)
);

BUFx3_ASAP7_75t_L g2079 ( 
.A(n_2016),
.Y(n_2079)
);

BUFx2_ASAP7_75t_SL g2080 ( 
.A(n_2033),
.Y(n_2080)
);

AOI22xp33_ASAP7_75t_L g2081 ( 
.A1(n_1998),
.A2(n_1939),
.B1(n_1980),
.B2(n_1947),
.Y(n_2081)
);

AOI22xp33_ASAP7_75t_L g2082 ( 
.A1(n_1998),
.A2(n_1956),
.B1(n_1908),
.B2(n_1929),
.Y(n_2082)
);

BUFx12f_ASAP7_75t_L g2083 ( 
.A(n_2005),
.Y(n_2083)
);

CKINVDCx5p33_ASAP7_75t_R g2084 ( 
.A(n_2000),
.Y(n_2084)
);

AOI22xp33_ASAP7_75t_L g2085 ( 
.A1(n_2040),
.A2(n_1910),
.B1(n_1916),
.B2(n_1919),
.Y(n_2085)
);

AOI22xp33_ASAP7_75t_L g2086 ( 
.A1(n_2040),
.A2(n_1926),
.B1(n_1952),
.B2(n_1899),
.Y(n_2086)
);

AOI22xp33_ASAP7_75t_L g2087 ( 
.A1(n_2007),
.A2(n_1930),
.B1(n_1981),
.B2(n_1953),
.Y(n_2087)
);

AOI22xp33_ASAP7_75t_SL g2088 ( 
.A1(n_2007),
.A2(n_2034),
.B1(n_2013),
.B2(n_2026),
.Y(n_2088)
);

AOI22xp33_ASAP7_75t_L g2089 ( 
.A1(n_2034),
.A2(n_1961),
.B1(n_1951),
.B2(n_1974),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_2010),
.Y(n_2090)
);

OAI22xp33_ASAP7_75t_R g2091 ( 
.A1(n_2035),
.A2(n_1978),
.B1(n_1962),
.B2(n_173),
.Y(n_2091)
);

INVx1_ASAP7_75t_SL g2092 ( 
.A(n_2008),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2024),
.Y(n_2093)
);

CKINVDCx11_ASAP7_75t_R g2094 ( 
.A(n_2023),
.Y(n_2094)
);

CKINVDCx11_ASAP7_75t_R g2095 ( 
.A(n_2025),
.Y(n_2095)
);

AOI22xp33_ASAP7_75t_SL g2096 ( 
.A1(n_2013),
.A2(n_1932),
.B1(n_1941),
.B2(n_1973),
.Y(n_2096)
);

BUFx2_ASAP7_75t_L g2097 ( 
.A(n_2020),
.Y(n_2097)
);

BUFx12f_ASAP7_75t_L g2098 ( 
.A(n_2015),
.Y(n_2098)
);

INVx3_ASAP7_75t_L g2099 ( 
.A(n_2029),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2031),
.Y(n_2100)
);

OAI22xp33_ASAP7_75t_SL g2101 ( 
.A1(n_2049),
.A2(n_1922),
.B1(n_1958),
.B2(n_1895),
.Y(n_2101)
);

BUFx3_ASAP7_75t_L g2102 ( 
.A(n_2017),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2073),
.Y(n_2103)
);

OAI22xp5_ASAP7_75t_L g2104 ( 
.A1(n_2066),
.A2(n_2051),
.B1(n_1949),
.B2(n_2055),
.Y(n_2104)
);

OR2x6_ASAP7_75t_L g2105 ( 
.A(n_2080),
.B(n_2026),
.Y(n_2105)
);

O2A1O1Ixp33_ASAP7_75t_L g2106 ( 
.A1(n_2078),
.A2(n_2051),
.B(n_2061),
.C(n_2049),
.Y(n_2106)
);

OAI22xp5_ASAP7_75t_L g2107 ( 
.A1(n_2088),
.A2(n_2076),
.B1(n_2086),
.B2(n_2081),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_2072),
.B(n_2006),
.Y(n_2108)
);

OAI22xp5_ASAP7_75t_L g2109 ( 
.A1(n_2085),
.A2(n_2043),
.B1(n_2018),
.B2(n_2041),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_2097),
.B(n_2079),
.Y(n_2110)
);

AOI21xp5_ASAP7_75t_L g2111 ( 
.A1(n_2091),
.A2(n_1992),
.B(n_1991),
.Y(n_2111)
);

OR2x2_ASAP7_75t_L g2112 ( 
.A(n_2092),
.B(n_2032),
.Y(n_2112)
);

BUFx8_ASAP7_75t_SL g2113 ( 
.A(n_2064),
.Y(n_2113)
);

HB1xp67_ASAP7_75t_L g2114 ( 
.A(n_2060),
.Y(n_2114)
);

OR2x2_ASAP7_75t_L g2115 ( 
.A(n_2060),
.B(n_2032),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_2073),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2079),
.B(n_2036),
.Y(n_2117)
);

BUFx6f_ASAP7_75t_L g2118 ( 
.A(n_2064),
.Y(n_2118)
);

OAI22xp5_ASAP7_75t_L g2119 ( 
.A1(n_2070),
.A2(n_2043),
.B1(n_2041),
.B2(n_2039),
.Y(n_2119)
);

BUFx3_ASAP7_75t_L g2120 ( 
.A(n_2063),
.Y(n_2120)
);

O2A1O1Ixp33_ASAP7_75t_L g2121 ( 
.A1(n_2101),
.A2(n_2042),
.B(n_1991),
.C(n_2039),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_2057),
.B(n_2099),
.Y(n_2122)
);

AOI21xp5_ASAP7_75t_SL g2123 ( 
.A1(n_2065),
.A2(n_2046),
.B(n_2054),
.Y(n_2123)
);

AND2x4_ASAP7_75t_L g2124 ( 
.A(n_2057),
.B(n_2003),
.Y(n_2124)
);

A2O1A1Ixp33_ASAP7_75t_L g2125 ( 
.A1(n_2082),
.A2(n_2046),
.B(n_1992),
.C(n_2054),
.Y(n_2125)
);

NAND2xp33_ASAP7_75t_SL g2126 ( 
.A(n_2071),
.B(n_2058),
.Y(n_2126)
);

HB1xp67_ASAP7_75t_L g2127 ( 
.A(n_2090),
.Y(n_2127)
);

AOI21x1_ASAP7_75t_SL g2128 ( 
.A1(n_2068),
.A2(n_2022),
.B(n_1999),
.Y(n_2128)
);

HB1xp67_ASAP7_75t_L g2129 ( 
.A(n_2090),
.Y(n_2129)
);

INVx3_ASAP7_75t_L g2130 ( 
.A(n_2105),
.Y(n_2130)
);

INVx3_ASAP7_75t_L g2131 ( 
.A(n_2105),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_2125),
.B(n_2108),
.Y(n_2132)
);

AND2x2_ASAP7_75t_SL g2133 ( 
.A(n_2118),
.B(n_2087),
.Y(n_2133)
);

NOR2xp33_ASAP7_75t_L g2134 ( 
.A(n_2118),
.B(n_2063),
.Y(n_2134)
);

AND2x4_ASAP7_75t_SL g2135 ( 
.A(n_2118),
.B(n_2071),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2116),
.Y(n_2136)
);

INVx8_ASAP7_75t_L g2137 ( 
.A(n_2113),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_2122),
.B(n_2110),
.Y(n_2138)
);

CKINVDCx16_ASAP7_75t_R g2139 ( 
.A(n_2126),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2122),
.B(n_2057),
.Y(n_2140)
);

INVx1_ASAP7_75t_SL g2141 ( 
.A(n_2126),
.Y(n_2141)
);

INVx3_ASAP7_75t_L g2142 ( 
.A(n_2130),
.Y(n_2142)
);

NAND4xp25_ASAP7_75t_L g2143 ( 
.A(n_2141),
.B(n_2111),
.C(n_2106),
.D(n_2121),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2136),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_2130),
.B(n_2105),
.Y(n_2145)
);

BUFx3_ASAP7_75t_L g2146 ( 
.A(n_2137),
.Y(n_2146)
);

INVx4_ASAP7_75t_L g2147 ( 
.A(n_2137),
.Y(n_2147)
);

OA21x2_ASAP7_75t_L g2148 ( 
.A1(n_2136),
.A2(n_2125),
.B(n_2116),
.Y(n_2148)
);

BUFx2_ASAP7_75t_SL g2149 ( 
.A(n_2130),
.Y(n_2149)
);

OR2x2_ASAP7_75t_L g2150 ( 
.A(n_2148),
.B(n_2132),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2144),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2144),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_2145),
.B(n_2139),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_2143),
.B(n_2133),
.Y(n_2154)
);

AOI22xp33_ASAP7_75t_L g2155 ( 
.A1(n_2143),
.A2(n_2133),
.B1(n_2119),
.B2(n_2109),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_2148),
.B(n_2133),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2149),
.Y(n_2157)
);

BUFx3_ASAP7_75t_L g2158 ( 
.A(n_2146),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2149),
.Y(n_2159)
);

OAI22xp5_ASAP7_75t_L g2160 ( 
.A1(n_2155),
.A2(n_2139),
.B1(n_2141),
.B2(n_2123),
.Y(n_2160)
);

INVxp67_ASAP7_75t_L g2161 ( 
.A(n_2153),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2152),
.Y(n_2162)
);

AOI22xp5_ASAP7_75t_L g2163 ( 
.A1(n_2154),
.A2(n_2104),
.B1(n_2107),
.B2(n_2147),
.Y(n_2163)
);

OR2x2_ASAP7_75t_SL g2164 ( 
.A(n_2156),
.B(n_2063),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2158),
.B(n_2146),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_2158),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_2153),
.Y(n_2167)
);

AOI221xp5_ASAP7_75t_L g2168 ( 
.A1(n_2150),
.A2(n_2159),
.B1(n_2157),
.B2(n_2151),
.C(n_2152),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2150),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_2153),
.B(n_2146),
.Y(n_2170)
);

OR2x2_ASAP7_75t_L g2171 ( 
.A(n_2153),
.B(n_2148),
.Y(n_2171)
);

AND2x4_ASAP7_75t_L g2172 ( 
.A(n_2170),
.B(n_2147),
.Y(n_2172)
);

AND2x4_ASAP7_75t_L g2173 ( 
.A(n_2167),
.B(n_2147),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2162),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_2161),
.B(n_2147),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2169),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_2166),
.B(n_2147),
.Y(n_2177)
);

AND2x4_ASAP7_75t_SL g2178 ( 
.A(n_2163),
.B(n_2118),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_2165),
.B(n_2135),
.Y(n_2179)
);

INVx2_ASAP7_75t_SL g2180 ( 
.A(n_2171),
.Y(n_2180)
);

INVx3_ASAP7_75t_L g2181 ( 
.A(n_2172),
.Y(n_2181)
);

BUFx2_ASAP7_75t_L g2182 ( 
.A(n_2180),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_2179),
.B(n_2135),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2176),
.B(n_2168),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_2183),
.B(n_2172),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2182),
.B(n_2178),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2181),
.Y(n_2187)
);

OR2x2_ASAP7_75t_L g2188 ( 
.A(n_2184),
.B(n_2176),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_2185),
.B(n_2181),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2187),
.Y(n_2190)
);

OR2x6_ASAP7_75t_L g2191 ( 
.A(n_2186),
.B(n_2137),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_2188),
.B(n_2184),
.Y(n_2192)
);

INVxp67_ASAP7_75t_L g2193 ( 
.A(n_2186),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2187),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2190),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2189),
.B(n_2175),
.Y(n_2196)
);

AO21x2_ASAP7_75t_L g2197 ( 
.A1(n_2192),
.A2(n_2174),
.B(n_2162),
.Y(n_2197)
);

INVx1_ASAP7_75t_SL g2198 ( 
.A(n_2191),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2194),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2193),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_SL g2201 ( 
.A(n_2191),
.B(n_2160),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2190),
.Y(n_2202)
);

INVx1_ASAP7_75t_SL g2203 ( 
.A(n_2189),
.Y(n_2203)
);

INVxp67_ASAP7_75t_L g2204 ( 
.A(n_2189),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_SL g2205 ( 
.A(n_2203),
.B(n_2173),
.Y(n_2205)
);

NOR2x1_ASAP7_75t_L g2206 ( 
.A(n_2197),
.B(n_2177),
.Y(n_2206)
);

AOI22xp5_ASAP7_75t_L g2207 ( 
.A1(n_2204),
.A2(n_2173),
.B1(n_2134),
.B2(n_2135),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_2198),
.B(n_2137),
.Y(n_2208)
);

AOI22xp5_ASAP7_75t_L g2209 ( 
.A1(n_2201),
.A2(n_2137),
.B1(n_2120),
.B2(n_2142),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2197),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_2196),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2200),
.Y(n_2212)
);

AOI22xp5_ASAP7_75t_L g2213 ( 
.A1(n_2195),
.A2(n_2202),
.B1(n_2199),
.B2(n_2120),
.Y(n_2213)
);

AOI32xp33_ASAP7_75t_L g2214 ( 
.A1(n_2203),
.A2(n_2142),
.A3(n_2164),
.B1(n_2145),
.B2(n_2131),
.Y(n_2214)
);

OR2x2_ASAP7_75t_L g2215 ( 
.A(n_2203),
.B(n_2142),
.Y(n_2215)
);

AOI22xp5_ASAP7_75t_L g2216 ( 
.A1(n_2203),
.A2(n_2142),
.B1(n_2145),
.B2(n_2148),
.Y(n_2216)
);

OR2x2_ASAP7_75t_L g2217 ( 
.A(n_2203),
.B(n_2142),
.Y(n_2217)
);

AO22x1_ASAP7_75t_L g2218 ( 
.A1(n_2206),
.A2(n_2210),
.B1(n_2208),
.B2(n_2211),
.Y(n_2218)
);

INVx2_ASAP7_75t_L g2219 ( 
.A(n_2215),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2217),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_2205),
.Y(n_2221)
);

A2O1A1Ixp33_ASAP7_75t_L g2222 ( 
.A1(n_2214),
.A2(n_2065),
.B(n_2131),
.C(n_2130),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2213),
.Y(n_2223)
);

OAI22xp5_ASAP7_75t_L g2224 ( 
.A1(n_2209),
.A2(n_2059),
.B1(n_2058),
.B2(n_2148),
.Y(n_2224)
);

INVx1_ASAP7_75t_SL g2225 ( 
.A(n_2207),
.Y(n_2225)
);

INVx1_ASAP7_75t_SL g2226 ( 
.A(n_2212),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2216),
.B(n_2113),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2206),
.Y(n_2228)
);

AOI221xp5_ASAP7_75t_L g2229 ( 
.A1(n_2210),
.A2(n_2089),
.B1(n_2131),
.B2(n_1940),
.C(n_2019),
.Y(n_2229)
);

NOR4xp25_ASAP7_75t_SL g2230 ( 
.A(n_2210),
.B(n_2059),
.C(n_2084),
.D(n_2068),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_2208),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2206),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2218),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2221),
.B(n_2131),
.Y(n_2234)
);

OR2x2_ASAP7_75t_L g2235 ( 
.A(n_2231),
.B(n_2117),
.Y(n_2235)
);

AOI22xp33_ASAP7_75t_L g2236 ( 
.A1(n_2225),
.A2(n_2105),
.B1(n_2098),
.B2(n_2083),
.Y(n_2236)
);

NOR2xp33_ASAP7_75t_L g2237 ( 
.A(n_2227),
.B(n_2226),
.Y(n_2237)
);

NAND2x1_ASAP7_75t_L g2238 ( 
.A(n_2228),
.B(n_2138),
.Y(n_2238)
);

AND2x2_ASAP7_75t_L g2239 ( 
.A(n_2230),
.B(n_2219),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2232),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_2220),
.B(n_2117),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2223),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2222),
.B(n_2030),
.Y(n_2243)
);

OAI221xp5_ASAP7_75t_L g2244 ( 
.A1(n_2224),
.A2(n_2019),
.B1(n_2022),
.B2(n_2004),
.C(n_1999),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_2230),
.B(n_2138),
.Y(n_2245)
);

AOI21xp5_ASAP7_75t_L g2246 ( 
.A1(n_2229),
.A2(n_1950),
.B(n_1958),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_2239),
.B(n_2084),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2238),
.Y(n_2248)
);

NOR3xp33_ASAP7_75t_L g2249 ( 
.A(n_2237),
.B(n_2095),
.C(n_2094),
.Y(n_2249)
);

OAI321xp33_ASAP7_75t_L g2250 ( 
.A1(n_2245),
.A2(n_1922),
.A3(n_1950),
.B1(n_2004),
.B2(n_1777),
.C(n_1996),
.Y(n_2250)
);

INVx2_ASAP7_75t_SL g2251 ( 
.A(n_2235),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2241),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2234),
.Y(n_2253)
);

AOI21xp5_ASAP7_75t_L g2254 ( 
.A1(n_2233),
.A2(n_2002),
.B(n_1996),
.Y(n_2254)
);

INVx2_ASAP7_75t_L g2255 ( 
.A(n_2240),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_SL g2256 ( 
.A(n_2236),
.B(n_1792),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2242),
.Y(n_2257)
);

NOR2xp33_ASAP7_75t_L g2258 ( 
.A(n_2243),
.B(n_2094),
.Y(n_2258)
);

OAI22xp5_ASAP7_75t_L g2259 ( 
.A1(n_2246),
.A2(n_2244),
.B1(n_2140),
.B2(n_2028),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2239),
.B(n_2140),
.Y(n_2260)
);

OR2x2_ASAP7_75t_L g2261 ( 
.A(n_2238),
.B(n_2112),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_SL g2262 ( 
.A(n_2245),
.B(n_2099),
.Y(n_2262)
);

NOR2xp33_ASAP7_75t_L g2263 ( 
.A(n_2245),
.B(n_2095),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_2239),
.B(n_170),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2238),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_2239),
.B(n_172),
.Y(n_2266)
);

AOI221x1_ASAP7_75t_L g2267 ( 
.A1(n_2233),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.C(n_175),
.Y(n_2267)
);

NOR2xp33_ASAP7_75t_L g2268 ( 
.A(n_2245),
.B(n_174),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2248),
.B(n_2265),
.Y(n_2269)
);

NOR3xp33_ASAP7_75t_L g2270 ( 
.A(n_2268),
.B(n_2002),
.C(n_2075),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_2263),
.B(n_175),
.Y(n_2271)
);

OAI21xp5_ASAP7_75t_L g2272 ( 
.A1(n_2264),
.A2(n_1976),
.B(n_1975),
.Y(n_2272)
);

AOI22xp5_ASAP7_75t_L g2273 ( 
.A1(n_2249),
.A2(n_2083),
.B1(n_2098),
.B2(n_2075),
.Y(n_2273)
);

NOR2xp33_ASAP7_75t_L g2274 ( 
.A(n_2260),
.B(n_176),
.Y(n_2274)
);

AOI21xp5_ASAP7_75t_L g2275 ( 
.A1(n_2247),
.A2(n_1885),
.B(n_1966),
.Y(n_2275)
);

NOR2xp33_ASAP7_75t_L g2276 ( 
.A(n_2266),
.B(n_176),
.Y(n_2276)
);

OAI221xp5_ASAP7_75t_L g2277 ( 
.A1(n_2258),
.A2(n_2077),
.B1(n_2053),
.B2(n_2096),
.C(n_2037),
.Y(n_2277)
);

AOI22xp5_ASAP7_75t_L g2278 ( 
.A1(n_2251),
.A2(n_2077),
.B1(n_2062),
.B2(n_2099),
.Y(n_2278)
);

AO21x1_ASAP7_75t_L g2279 ( 
.A1(n_2257),
.A2(n_178),
.B(n_179),
.Y(n_2279)
);

NOR2x1_ASAP7_75t_L g2280 ( 
.A(n_2255),
.B(n_179),
.Y(n_2280)
);

NOR2xp33_ASAP7_75t_L g2281 ( 
.A(n_2262),
.B(n_180),
.Y(n_2281)
);

OAI21xp33_ASAP7_75t_SL g2282 ( 
.A1(n_2256),
.A2(n_2128),
.B(n_2114),
.Y(n_2282)
);

NOR2xp33_ASAP7_75t_L g2283 ( 
.A(n_2261),
.B(n_181),
.Y(n_2283)
);

AOI21xp5_ASAP7_75t_L g2284 ( 
.A1(n_2253),
.A2(n_2252),
.B(n_2250),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2267),
.B(n_181),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2254),
.B(n_182),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_2259),
.B(n_182),
.Y(n_2287)
);

OAI211xp5_ASAP7_75t_L g2288 ( 
.A1(n_2247),
.A2(n_185),
.B(n_183),
.C(n_184),
.Y(n_2288)
);

INVxp67_ASAP7_75t_SL g2289 ( 
.A(n_2248),
.Y(n_2289)
);

AOI211xp5_ASAP7_75t_L g2290 ( 
.A1(n_2263),
.A2(n_187),
.B(n_183),
.C(n_186),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2248),
.B(n_186),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2260),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2260),
.Y(n_2293)
);

INVx2_ASAP7_75t_L g2294 ( 
.A(n_2261),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_SL g2295 ( 
.A(n_2248),
.B(n_2056),
.Y(n_2295)
);

NOR2xp33_ASAP7_75t_L g2296 ( 
.A(n_2260),
.B(n_187),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_2248),
.B(n_188),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_2249),
.B(n_2124),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2248),
.B(n_188),
.Y(n_2299)
);

NAND3xp33_ASAP7_75t_L g2300 ( 
.A(n_2268),
.B(n_189),
.C(n_190),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2260),
.Y(n_2301)
);

O2A1O1Ixp33_ASAP7_75t_L g2302 ( 
.A1(n_2248),
.A2(n_193),
.B(n_191),
.C(n_192),
.Y(n_2302)
);

NOR2xp33_ASAP7_75t_L g2303 ( 
.A(n_2260),
.B(n_191),
.Y(n_2303)
);

NAND3xp33_ASAP7_75t_L g2304 ( 
.A(n_2268),
.B(n_192),
.C(n_193),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_SL g2305 ( 
.A(n_2248),
.B(n_2056),
.Y(n_2305)
);

OAI31xp33_ASAP7_75t_L g2306 ( 
.A1(n_2288),
.A2(n_2050),
.A3(n_2045),
.B(n_196),
.Y(n_2306)
);

NOR2xp33_ASAP7_75t_L g2307 ( 
.A(n_2294),
.B(n_194),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2279),
.Y(n_2308)
);

AOI221xp5_ASAP7_75t_L g2309 ( 
.A1(n_2289),
.A2(n_197),
.B1(n_194),
.B2(n_195),
.C(n_198),
.Y(n_2309)
);

OR2x2_ASAP7_75t_L g2310 ( 
.A(n_2285),
.B(n_195),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2280),
.Y(n_2311)
);

NAND3xp33_ASAP7_75t_L g2312 ( 
.A(n_2290),
.B(n_197),
.C(n_199),
.Y(n_2312)
);

NOR4xp25_ASAP7_75t_L g2313 ( 
.A(n_2269),
.B(n_201),
.C(n_199),
.D(n_200),
.Y(n_2313)
);

O2A1O1Ixp33_ASAP7_75t_L g2314 ( 
.A1(n_2291),
.A2(n_204),
.B(n_200),
.C(n_202),
.Y(n_2314)
);

NAND3xp33_ASAP7_75t_SL g2315 ( 
.A(n_2297),
.B(n_202),
.C(n_204),
.Y(n_2315)
);

AND4x1_ASAP7_75t_L g2316 ( 
.A(n_2274),
.B(n_207),
.C(n_205),
.D(n_206),
.Y(n_2316)
);

NAND3xp33_ASAP7_75t_SL g2317 ( 
.A(n_2299),
.B(n_2302),
.C(n_2283),
.Y(n_2317)
);

NAND3xp33_ASAP7_75t_L g2318 ( 
.A(n_2296),
.B(n_206),
.C(n_207),
.Y(n_2318)
);

OAI211xp5_ASAP7_75t_L g2319 ( 
.A1(n_2303),
.A2(n_210),
.B(n_208),
.C(n_209),
.Y(n_2319)
);

NAND4xp25_ASAP7_75t_L g2320 ( 
.A(n_2270),
.B(n_214),
.C(n_209),
.D(n_213),
.Y(n_2320)
);

NOR2xp33_ASAP7_75t_L g2321 ( 
.A(n_2300),
.B(n_2304),
.Y(n_2321)
);

NAND4xp75_ASAP7_75t_L g2322 ( 
.A(n_2284),
.B(n_215),
.C(n_213),
.D(n_214),
.Y(n_2322)
);

NOR3xp33_ASAP7_75t_SL g2323 ( 
.A(n_2287),
.B(n_215),
.C(n_216),
.Y(n_2323)
);

AOI221xp5_ASAP7_75t_L g2324 ( 
.A1(n_2295),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.C(n_219),
.Y(n_2324)
);

NOR3x1_ASAP7_75t_L g2325 ( 
.A(n_2271),
.B(n_217),
.C(n_218),
.Y(n_2325)
);

NOR4xp25_ASAP7_75t_L g2326 ( 
.A(n_2292),
.B(n_222),
.C(n_219),
.D(n_220),
.Y(n_2326)
);

OAI21xp5_ASAP7_75t_L g2327 ( 
.A1(n_2305),
.A2(n_1972),
.B(n_1967),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_L g2328 ( 
.A(n_2298),
.B(n_220),
.Y(n_2328)
);

NAND4xp25_ASAP7_75t_L g2329 ( 
.A(n_2293),
.B(n_224),
.C(n_222),
.D(n_223),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2286),
.Y(n_2330)
);

AND2x2_ASAP7_75t_L g2331 ( 
.A(n_2301),
.B(n_2124),
.Y(n_2331)
);

AND2x4_ASAP7_75t_L g2332 ( 
.A(n_2273),
.B(n_2033),
.Y(n_2332)
);

OAI211xp5_ASAP7_75t_L g2333 ( 
.A1(n_2281),
.A2(n_225),
.B(n_223),
.C(n_224),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2276),
.B(n_225),
.Y(n_2334)
);

NOR2xp33_ASAP7_75t_L g2335 ( 
.A(n_2282),
.B(n_2278),
.Y(n_2335)
);

NOR3xp33_ASAP7_75t_L g2336 ( 
.A(n_2277),
.B(n_226),
.C(n_227),
.Y(n_2336)
);

NOR2xp33_ASAP7_75t_L g2337 ( 
.A(n_2275),
.B(n_226),
.Y(n_2337)
);

NOR2xp67_ASAP7_75t_SL g2338 ( 
.A(n_2272),
.B(n_227),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_SL g2339 ( 
.A(n_2272),
.B(n_2056),
.Y(n_2339)
);

NOR2x1_ASAP7_75t_L g2340 ( 
.A(n_2308),
.B(n_228),
.Y(n_2340)
);

NOR4xp25_ASAP7_75t_L g2341 ( 
.A(n_2317),
.B(n_230),
.C(n_228),
.D(n_229),
.Y(n_2341)
);

NAND3xp33_ASAP7_75t_L g2342 ( 
.A(n_2323),
.B(n_230),
.C(n_231),
.Y(n_2342)
);

NAND3xp33_ASAP7_75t_L g2343 ( 
.A(n_2311),
.B(n_232),
.C(n_233),
.Y(n_2343)
);

NOR3xp33_ASAP7_75t_L g2344 ( 
.A(n_2328),
.B(n_232),
.C(n_233),
.Y(n_2344)
);

AOI211xp5_ASAP7_75t_L g2345 ( 
.A1(n_2313),
.A2(n_237),
.B(n_234),
.C(n_235),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2316),
.Y(n_2346)
);

NAND4xp75_ASAP7_75t_L g2347 ( 
.A(n_2325),
.B(n_240),
.C(n_237),
.D(n_238),
.Y(n_2347)
);

NAND4xp25_ASAP7_75t_L g2348 ( 
.A(n_2306),
.B(n_242),
.C(n_238),
.D(n_241),
.Y(n_2348)
);

NAND4xp25_ASAP7_75t_SL g2349 ( 
.A(n_2312),
.B(n_243),
.C(n_241),
.D(n_242),
.Y(n_2349)
);

NOR3xp33_ASAP7_75t_L g2350 ( 
.A(n_2322),
.B(n_243),
.C(n_244),
.Y(n_2350)
);

AOI211xp5_ASAP7_75t_L g2351 ( 
.A1(n_2320),
.A2(n_247),
.B(n_245),
.C(n_246),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2326),
.B(n_245),
.Y(n_2352)
);

NOR3xp33_ASAP7_75t_L g2353 ( 
.A(n_2334),
.B(n_246),
.C(n_247),
.Y(n_2353)
);

NAND4xp25_ASAP7_75t_SL g2354 ( 
.A(n_2336),
.B(n_252),
.C(n_249),
.D(n_251),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_2310),
.Y(n_2355)
);

OAI211xp5_ASAP7_75t_L g2356 ( 
.A1(n_2333),
.A2(n_253),
.B(n_251),
.C(n_252),
.Y(n_2356)
);

AOI211xp5_ASAP7_75t_L g2357 ( 
.A1(n_2315),
.A2(n_255),
.B(n_253),
.C(n_254),
.Y(n_2357)
);

NOR4xp25_ASAP7_75t_L g2358 ( 
.A(n_2330),
.B(n_260),
.C(n_256),
.D(n_259),
.Y(n_2358)
);

NAND4xp75_ASAP7_75t_L g2359 ( 
.A(n_2321),
.B(n_261),
.C(n_259),
.D(n_260),
.Y(n_2359)
);

NOR2xp67_ASAP7_75t_L g2360 ( 
.A(n_2329),
.B(n_261),
.Y(n_2360)
);

NOR3xp33_ASAP7_75t_L g2361 ( 
.A(n_2318),
.B(n_262),
.C(n_263),
.Y(n_2361)
);

OAI221xp5_ASAP7_75t_SL g2362 ( 
.A1(n_2331),
.A2(n_2062),
.B1(n_2115),
.B2(n_265),
.C(n_266),
.Y(n_2362)
);

NOR4xp25_ASAP7_75t_L g2363 ( 
.A(n_2314),
.B(n_265),
.C(n_262),
.D(n_264),
.Y(n_2363)
);

NAND5xp2_ASAP7_75t_L g2364 ( 
.A(n_2335),
.B(n_264),
.C(n_267),
.D(n_268),
.E(n_269),
.Y(n_2364)
);

AND4x1_ASAP7_75t_L g2365 ( 
.A(n_2307),
.B(n_271),
.C(n_267),
.D(n_270),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2319),
.Y(n_2366)
);

OAI21xp5_ASAP7_75t_L g2367 ( 
.A1(n_2332),
.A2(n_1948),
.B(n_1925),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_2324),
.B(n_270),
.Y(n_2368)
);

NAND3xp33_ASAP7_75t_L g2369 ( 
.A(n_2338),
.B(n_271),
.C(n_272),
.Y(n_2369)
);

AOI211xp5_ASAP7_75t_L g2370 ( 
.A1(n_2332),
.A2(n_274),
.B(n_272),
.C(n_273),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2309),
.B(n_2337),
.Y(n_2371)
);

NOR2xp33_ASAP7_75t_L g2372 ( 
.A(n_2339),
.B(n_275),
.Y(n_2372)
);

AOI21xp5_ASAP7_75t_L g2373 ( 
.A1(n_2327),
.A2(n_276),
.B(n_277),
.Y(n_2373)
);

AOI221xp5_ASAP7_75t_L g2374 ( 
.A1(n_2308),
.A2(n_277),
.B1(n_278),
.B2(n_280),
.C(n_281),
.Y(n_2374)
);

AOI221xp5_ASAP7_75t_SL g2375 ( 
.A1(n_2308),
.A2(n_278),
.B1(n_280),
.B2(n_281),
.C(n_282),
.Y(n_2375)
);

NOR2xp67_ASAP7_75t_L g2376 ( 
.A(n_2308),
.B(n_282),
.Y(n_2376)
);

INVxp67_ASAP7_75t_L g2377 ( 
.A(n_2307),
.Y(n_2377)
);

AOI221xp5_ASAP7_75t_L g2378 ( 
.A1(n_2308),
.A2(n_283),
.B1(n_284),
.B2(n_286),
.C(n_287),
.Y(n_2378)
);

NAND3xp33_ASAP7_75t_L g2379 ( 
.A(n_2308),
.B(n_283),
.C(n_284),
.Y(n_2379)
);

NOR2x1p5_ASAP7_75t_L g2380 ( 
.A(n_2322),
.B(n_286),
.Y(n_2380)
);

AOI211xp5_ASAP7_75t_L g2381 ( 
.A1(n_2313),
.A2(n_289),
.B(n_287),
.C(n_288),
.Y(n_2381)
);

OAI211xp5_ASAP7_75t_SL g2382 ( 
.A1(n_2306),
.A2(n_291),
.B(n_289),
.C(n_290),
.Y(n_2382)
);

NOR2x1_ASAP7_75t_L g2383 ( 
.A(n_2308),
.B(n_290),
.Y(n_2383)
);

AOI21xp5_ASAP7_75t_L g2384 ( 
.A1(n_2328),
.A2(n_291),
.B(n_292),
.Y(n_2384)
);

BUFx2_ASAP7_75t_L g2385 ( 
.A(n_2308),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2313),
.B(n_293),
.Y(n_2386)
);

NOR3xp33_ASAP7_75t_L g2387 ( 
.A(n_2328),
.B(n_294),
.C(n_295),
.Y(n_2387)
);

NAND3xp33_ASAP7_75t_SL g2388 ( 
.A(n_2308),
.B(n_294),
.C(n_295),
.Y(n_2388)
);

OAI211xp5_ASAP7_75t_L g2389 ( 
.A1(n_2313),
.A2(n_298),
.B(n_296),
.C(n_297),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2316),
.Y(n_2390)
);

OA211x2_ASAP7_75t_L g2391 ( 
.A1(n_2324),
.A2(n_298),
.B(n_296),
.C(n_297),
.Y(n_2391)
);

AOI221xp5_ASAP7_75t_L g2392 ( 
.A1(n_2363),
.A2(n_299),
.B1(n_301),
.B2(n_302),
.C(n_303),
.Y(n_2392)
);

OAI21xp33_ASAP7_75t_L g2393 ( 
.A1(n_2348),
.A2(n_2102),
.B(n_2124),
.Y(n_2393)
);

AOI221xp5_ASAP7_75t_L g2394 ( 
.A1(n_2385),
.A2(n_301),
.B1(n_303),
.B2(n_304),
.C(n_305),
.Y(n_2394)
);

HB1xp67_ASAP7_75t_L g2395 ( 
.A(n_2376),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2386),
.Y(n_2396)
);

HB1xp67_ASAP7_75t_L g2397 ( 
.A(n_2365),
.Y(n_2397)
);

AOI22xp5_ASAP7_75t_L g2398 ( 
.A1(n_2360),
.A2(n_2077),
.B1(n_2056),
.B2(n_2017),
.Y(n_2398)
);

AOI21xp5_ASAP7_75t_L g2399 ( 
.A1(n_2352),
.A2(n_304),
.B(n_305),
.Y(n_2399)
);

NOR2x1_ASAP7_75t_L g2400 ( 
.A(n_2340),
.B(n_306),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2383),
.Y(n_2401)
);

AOI221xp5_ASAP7_75t_SL g2402 ( 
.A1(n_2373),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.C(n_311),
.Y(n_2402)
);

NAND2xp33_ASAP7_75t_SL g2403 ( 
.A(n_2380),
.B(n_309),
.Y(n_2403)
);

INVxp67_ASAP7_75t_L g2404 ( 
.A(n_2364),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_2358),
.B(n_310),
.Y(n_2405)
);

NOR2xp33_ASAP7_75t_R g2406 ( 
.A(n_2388),
.B(n_311),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_2358),
.B(n_2341),
.Y(n_2407)
);

AOI221xp5_ASAP7_75t_L g2408 ( 
.A1(n_2382),
.A2(n_312),
.B1(n_313),
.B2(n_314),
.C(n_315),
.Y(n_2408)
);

NAND2x1_ASAP7_75t_L g2409 ( 
.A(n_2346),
.B(n_2077),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_L g2410 ( 
.A(n_2375),
.B(n_313),
.Y(n_2410)
);

INVx1_ASAP7_75t_SL g2411 ( 
.A(n_2347),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2379),
.Y(n_2412)
);

O2A1O1Ixp33_ASAP7_75t_L g2413 ( 
.A1(n_2390),
.A2(n_314),
.B(n_315),
.C(n_316),
.Y(n_2413)
);

AND2x2_ASAP7_75t_L g2414 ( 
.A(n_2350),
.B(n_2366),
.Y(n_2414)
);

OAI22xp5_ASAP7_75t_L g2415 ( 
.A1(n_2362),
.A2(n_2342),
.B1(n_2369),
.B2(n_2343),
.Y(n_2415)
);

XNOR2x1_ASAP7_75t_L g2416 ( 
.A(n_2391),
.B(n_317),
.Y(n_2416)
);

OAI211xp5_ASAP7_75t_SL g2417 ( 
.A1(n_2377),
.A2(n_317),
.B(n_318),
.C(n_319),
.Y(n_2417)
);

NAND4xp75_ASAP7_75t_L g2418 ( 
.A(n_2372),
.B(n_318),
.C(n_319),
.D(n_320),
.Y(n_2418)
);

AND2x2_ASAP7_75t_L g2419 ( 
.A(n_2351),
.B(n_2127),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2389),
.Y(n_2420)
);

NOR2xp33_ASAP7_75t_R g2421 ( 
.A(n_2354),
.B(n_320),
.Y(n_2421)
);

XNOR2xp5_ASAP7_75t_L g2422 ( 
.A(n_2345),
.B(n_321),
.Y(n_2422)
);

CKINVDCx5p33_ASAP7_75t_R g2423 ( 
.A(n_2355),
.Y(n_2423)
);

NAND4xp75_ASAP7_75t_L g2424 ( 
.A(n_2384),
.B(n_321),
.C(n_322),
.D(n_324),
.Y(n_2424)
);

AOI211xp5_ASAP7_75t_L g2425 ( 
.A1(n_2349),
.A2(n_322),
.B(n_324),
.C(n_325),
.Y(n_2425)
);

AND2x2_ASAP7_75t_L g2426 ( 
.A(n_2344),
.B(n_2129),
.Y(n_2426)
);

INVx1_ASAP7_75t_SL g2427 ( 
.A(n_2359),
.Y(n_2427)
);

NOR3xp33_ASAP7_75t_L g2428 ( 
.A(n_2371),
.B(n_325),
.C(n_326),
.Y(n_2428)
);

AOI22xp33_ASAP7_75t_L g2429 ( 
.A1(n_2361),
.A2(n_2102),
.B1(n_2001),
.B2(n_2100),
.Y(n_2429)
);

AOI211xp5_ASAP7_75t_L g2430 ( 
.A1(n_2356),
.A2(n_326),
.B(n_327),
.C(n_328),
.Y(n_2430)
);

OAI322xp33_ASAP7_75t_L g2431 ( 
.A1(n_2368),
.A2(n_327),
.A3(n_328),
.B1(n_329),
.B2(n_330),
.C1(n_331),
.C2(n_332),
.Y(n_2431)
);

NOR2xp33_ASAP7_75t_R g2432 ( 
.A(n_2381),
.B(n_329),
.Y(n_2432)
);

OAI22xp5_ASAP7_75t_L g2433 ( 
.A1(n_2357),
.A2(n_2048),
.B1(n_2047),
.B2(n_2103),
.Y(n_2433)
);

XNOR2xp5_ASAP7_75t_L g2434 ( 
.A(n_2370),
.B(n_330),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2387),
.Y(n_2435)
);

OAI211xp5_ASAP7_75t_SL g2436 ( 
.A1(n_2353),
.A2(n_332),
.B(n_333),
.C(n_334),
.Y(n_2436)
);

AO22x2_ASAP7_75t_L g2437 ( 
.A1(n_2374),
.A2(n_2378),
.B1(n_2367),
.B2(n_337),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_2376),
.B(n_334),
.Y(n_2438)
);

OAI322xp33_ASAP7_75t_L g2439 ( 
.A1(n_2366),
.A2(n_336),
.A3(n_338),
.B1(n_339),
.B2(n_340),
.C1(n_341),
.C2(n_342),
.Y(n_2439)
);

INVx1_ASAP7_75t_SL g2440 ( 
.A(n_2347),
.Y(n_2440)
);

HB1xp67_ASAP7_75t_L g2441 ( 
.A(n_2416),
.Y(n_2441)
);

XNOR2xp5_ASAP7_75t_L g2442 ( 
.A(n_2422),
.B(n_336),
.Y(n_2442)
);

XNOR2x1_ASAP7_75t_L g2443 ( 
.A(n_2424),
.B(n_338),
.Y(n_2443)
);

OAI322xp33_ASAP7_75t_L g2444 ( 
.A1(n_2404),
.A2(n_339),
.A3(n_340),
.B1(n_341),
.B2(n_342),
.C1(n_343),
.C2(n_344),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_SL g2445 ( 
.A(n_2408),
.B(n_343),
.Y(n_2445)
);

NOR2x1_ASAP7_75t_L g2446 ( 
.A(n_2400),
.B(n_345),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2392),
.B(n_345),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_2397),
.B(n_2003),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2405),
.Y(n_2449)
);

NAND4xp75_ASAP7_75t_L g2450 ( 
.A(n_2399),
.B(n_2414),
.C(n_2420),
.D(n_2438),
.Y(n_2450)
);

OAI21xp5_ASAP7_75t_SL g2451 ( 
.A1(n_2434),
.A2(n_346),
.B(n_347),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2407),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2410),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2425),
.B(n_346),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2395),
.Y(n_2455)
);

NOR2xp33_ASAP7_75t_L g2456 ( 
.A(n_2436),
.B(n_347),
.Y(n_2456)
);

AND2x4_ASAP7_75t_L g2457 ( 
.A(n_2401),
.B(n_348),
.Y(n_2457)
);

AOI22xp5_ASAP7_75t_L g2458 ( 
.A1(n_2423),
.A2(n_2048),
.B1(n_2021),
.B2(n_2067),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_2428),
.B(n_349),
.Y(n_2459)
);

AOI22xp5_ASAP7_75t_L g2460 ( 
.A1(n_2411),
.A2(n_2048),
.B1(n_2021),
.B2(n_2067),
.Y(n_2460)
);

AND2x2_ASAP7_75t_L g2461 ( 
.A(n_2440),
.B(n_2047),
.Y(n_2461)
);

NAND4xp75_ASAP7_75t_L g2462 ( 
.A(n_2412),
.B(n_2402),
.C(n_2396),
.D(n_2435),
.Y(n_2462)
);

NAND4xp75_ASAP7_75t_L g2463 ( 
.A(n_2394),
.B(n_349),
.C(n_351),
.D(n_352),
.Y(n_2463)
);

XNOR2xp5_ASAP7_75t_L g2464 ( 
.A(n_2418),
.B(n_351),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2403),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2419),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_2409),
.Y(n_2467)
);

OR2x2_ASAP7_75t_L g2468 ( 
.A(n_2427),
.B(n_352),
.Y(n_2468)
);

NOR2xp33_ASAP7_75t_L g2469 ( 
.A(n_2431),
.B(n_2417),
.Y(n_2469)
);

INVx2_ASAP7_75t_L g2470 ( 
.A(n_2437),
.Y(n_2470)
);

INVx1_ASAP7_75t_SL g2471 ( 
.A(n_2421),
.Y(n_2471)
);

XNOR2xp5_ASAP7_75t_L g2472 ( 
.A(n_2430),
.B(n_353),
.Y(n_2472)
);

INVx2_ASAP7_75t_L g2473 ( 
.A(n_2437),
.Y(n_2473)
);

NAND3x1_ASAP7_75t_L g2474 ( 
.A(n_2406),
.B(n_353),
.C(n_354),
.Y(n_2474)
);

AND2x2_ASAP7_75t_L g2475 ( 
.A(n_2426),
.B(n_2429),
.Y(n_2475)
);

NOR2x1_ASAP7_75t_L g2476 ( 
.A(n_2439),
.B(n_355),
.Y(n_2476)
);

NOR3x2_ASAP7_75t_L g2477 ( 
.A(n_2413),
.B(n_355),
.C(n_356),
.Y(n_2477)
);

NOR2x1p5_ASAP7_75t_L g2478 ( 
.A(n_2432),
.B(n_2415),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_2398),
.Y(n_2479)
);

INVxp33_ASAP7_75t_L g2480 ( 
.A(n_2433),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2468),
.Y(n_2481)
);

NOR2x1_ASAP7_75t_L g2482 ( 
.A(n_2446),
.B(n_2393),
.Y(n_2482)
);

NOR3xp33_ASAP7_75t_SL g2483 ( 
.A(n_2462),
.B(n_356),
.C(n_357),
.Y(n_2483)
);

NOR4xp75_ASAP7_75t_L g2484 ( 
.A(n_2474),
.B(n_357),
.C(n_358),
.D(n_359),
.Y(n_2484)
);

NAND4xp75_ASAP7_75t_L g2485 ( 
.A(n_2455),
.B(n_358),
.C(n_359),
.D(n_360),
.Y(n_2485)
);

NAND4xp25_ASAP7_75t_SL g2486 ( 
.A(n_2454),
.B(n_360),
.C(n_361),
.D(n_362),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2464),
.Y(n_2487)
);

NAND4xp25_ASAP7_75t_L g2488 ( 
.A(n_2469),
.B(n_361),
.C(n_362),
.D(n_363),
.Y(n_2488)
);

NOR4xp25_ASAP7_75t_L g2489 ( 
.A(n_2452),
.B(n_363),
.C(n_364),
.D(n_365),
.Y(n_2489)
);

NOR5xp2_ASAP7_75t_L g2490 ( 
.A(n_2441),
.B(n_364),
.C(n_365),
.D(n_366),
.E(n_367),
.Y(n_2490)
);

NOR3xp33_ASAP7_75t_SL g2491 ( 
.A(n_2450),
.B(n_366),
.C(n_368),
.Y(n_2491)
);

NAND2x1_ASAP7_75t_L g2492 ( 
.A(n_2467),
.B(n_369),
.Y(n_2492)
);

XNOR2x1_ASAP7_75t_L g2493 ( 
.A(n_2443),
.B(n_369),
.Y(n_2493)
);

NOR3xp33_ASAP7_75t_L g2494 ( 
.A(n_2465),
.B(n_370),
.C(n_371),
.Y(n_2494)
);

NOR3xp33_ASAP7_75t_L g2495 ( 
.A(n_2465),
.B(n_370),
.C(n_373),
.Y(n_2495)
);

NAND4xp25_ASAP7_75t_L g2496 ( 
.A(n_2456),
.B(n_374),
.C(n_375),
.D(n_376),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_2461),
.B(n_374),
.Y(n_2497)
);

NAND5xp2_ASAP7_75t_L g2498 ( 
.A(n_2466),
.B(n_375),
.C(n_376),
.D(n_378),
.E(n_379),
.Y(n_2498)
);

NOR3x2_ASAP7_75t_L g2499 ( 
.A(n_2463),
.B(n_379),
.C(n_380),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2477),
.Y(n_2500)
);

OR5x1_ASAP7_75t_L g2501 ( 
.A(n_2442),
.B(n_2480),
.C(n_2476),
.D(n_2478),
.E(n_2472),
.Y(n_2501)
);

OR5x1_ASAP7_75t_L g2502 ( 
.A(n_2471),
.B(n_2445),
.C(n_2447),
.D(n_2473),
.E(n_2470),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2448),
.Y(n_2503)
);

NOR3xp33_ASAP7_75t_SL g2504 ( 
.A(n_2451),
.B(n_2449),
.C(n_2459),
.Y(n_2504)
);

OR5x1_ASAP7_75t_L g2505 ( 
.A(n_2475),
.B(n_380),
.C(n_381),
.D(n_382),
.E(n_383),
.Y(n_2505)
);

AND2x2_ASAP7_75t_L g2506 ( 
.A(n_2479),
.B(n_2047),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_2457),
.Y(n_2507)
);

INVxp67_ASAP7_75t_L g2508 ( 
.A(n_2457),
.Y(n_2508)
);

OAI22xp5_ASAP7_75t_L g2509 ( 
.A1(n_2460),
.A2(n_2047),
.B1(n_2093),
.B2(n_2069),
.Y(n_2509)
);

CKINVDCx16_ASAP7_75t_R g2510 ( 
.A(n_2503),
.Y(n_2510)
);

NOR3xp33_ASAP7_75t_L g2511 ( 
.A(n_2508),
.B(n_2453),
.C(n_2444),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_2489),
.B(n_2458),
.Y(n_2512)
);

NAND2xp33_ASAP7_75t_L g2513 ( 
.A(n_2494),
.B(n_2495),
.Y(n_2513)
);

CKINVDCx20_ASAP7_75t_R g2514 ( 
.A(n_2483),
.Y(n_2514)
);

CKINVDCx20_ASAP7_75t_R g2515 ( 
.A(n_2504),
.Y(n_2515)
);

BUFx2_ASAP7_75t_L g2516 ( 
.A(n_2491),
.Y(n_2516)
);

CKINVDCx5p33_ASAP7_75t_R g2517 ( 
.A(n_2507),
.Y(n_2517)
);

NAND2xp33_ASAP7_75t_R g2518 ( 
.A(n_2500),
.B(n_381),
.Y(n_2518)
);

HB1xp67_ASAP7_75t_L g2519 ( 
.A(n_2484),
.Y(n_2519)
);

NOR3xp33_ASAP7_75t_L g2520 ( 
.A(n_2481),
.B(n_382),
.C(n_383),
.Y(n_2520)
);

CKINVDCx5p33_ASAP7_75t_R g2521 ( 
.A(n_2487),
.Y(n_2521)
);

NOR2x1p5_ASAP7_75t_L g2522 ( 
.A(n_2492),
.B(n_384),
.Y(n_2522)
);

BUFx2_ASAP7_75t_L g2523 ( 
.A(n_2497),
.Y(n_2523)
);

NOR4xp25_ASAP7_75t_L g2524 ( 
.A(n_2496),
.B(n_384),
.C(n_385),
.D(n_386),
.Y(n_2524)
);

AOI221xp5_ASAP7_75t_L g2525 ( 
.A1(n_2506),
.A2(n_387),
.B1(n_388),
.B2(n_389),
.C(n_390),
.Y(n_2525)
);

HB1xp67_ASAP7_75t_L g2526 ( 
.A(n_2505),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2499),
.Y(n_2527)
);

INVx1_ASAP7_75t_SL g2528 ( 
.A(n_2485),
.Y(n_2528)
);

CKINVDCx16_ASAP7_75t_R g2529 ( 
.A(n_2482),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2488),
.B(n_387),
.Y(n_2530)
);

CKINVDCx5p33_ASAP7_75t_R g2531 ( 
.A(n_2501),
.Y(n_2531)
);

AND2x4_ASAP7_75t_L g2532 ( 
.A(n_2522),
.B(n_2502),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2530),
.Y(n_2533)
);

OAI322xp33_ASAP7_75t_SL g2534 ( 
.A1(n_2531),
.A2(n_2493),
.A3(n_2490),
.B1(n_2486),
.B2(n_2509),
.C1(n_2498),
.C2(n_393),
.Y(n_2534)
);

OAI322xp33_ASAP7_75t_L g2535 ( 
.A1(n_2529),
.A2(n_388),
.A3(n_389),
.B1(n_390),
.B2(n_391),
.C1(n_392),
.C2(n_394),
.Y(n_2535)
);

OAI31xp33_ASAP7_75t_L g2536 ( 
.A1(n_2526),
.A2(n_391),
.A3(n_392),
.B(n_394),
.Y(n_2536)
);

AOI221xp5_ASAP7_75t_L g2537 ( 
.A1(n_2524),
.A2(n_2511),
.B1(n_2528),
.B2(n_2517),
.C(n_2527),
.Y(n_2537)
);

AND2x2_ASAP7_75t_L g2538 ( 
.A(n_2519),
.B(n_2074),
.Y(n_2538)
);

XNOR2xp5_ASAP7_75t_L g2539 ( 
.A(n_2515),
.B(n_395),
.Y(n_2539)
);

OAI211xp5_ASAP7_75t_L g2540 ( 
.A1(n_2516),
.A2(n_2525),
.B(n_2521),
.C(n_2523),
.Y(n_2540)
);

AOI22xp5_ASAP7_75t_L g2541 ( 
.A1(n_2510),
.A2(n_395),
.B1(n_396),
.B2(n_397),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2512),
.Y(n_2542)
);

AOI322xp5_ASAP7_75t_L g2543 ( 
.A1(n_2513),
.A2(n_397),
.A3(n_398),
.B1(n_399),
.B2(n_400),
.C1(n_401),
.C2(n_402),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2514),
.Y(n_2544)
);

OAI221xp5_ASAP7_75t_L g2545 ( 
.A1(n_2518),
.A2(n_399),
.B1(n_400),
.B2(n_401),
.C(n_402),
.Y(n_2545)
);

AOI322xp5_ASAP7_75t_L g2546 ( 
.A1(n_2520),
.A2(n_403),
.A3(n_404),
.B1(n_405),
.B2(n_406),
.C1(n_407),
.C2(n_408),
.Y(n_2546)
);

AOI322xp5_ASAP7_75t_L g2547 ( 
.A1(n_2528),
.A2(n_403),
.A3(n_404),
.B1(n_405),
.B2(n_406),
.C1(n_408),
.C2(n_409),
.Y(n_2547)
);

A2O1A1Ixp33_ASAP7_75t_L g2548 ( 
.A1(n_2511),
.A2(n_409),
.B(n_410),
.C(n_411),
.Y(n_2548)
);

A2O1A1Ixp33_ASAP7_75t_L g2549 ( 
.A1(n_2511),
.A2(n_410),
.B(n_411),
.C(n_412),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2539),
.Y(n_2550)
);

AO22x2_ASAP7_75t_L g2551 ( 
.A1(n_2532),
.A2(n_412),
.B1(n_414),
.B2(n_415),
.Y(n_2551)
);

AO22x2_ASAP7_75t_SL g2552 ( 
.A1(n_2542),
.A2(n_415),
.B1(n_416),
.B2(n_417),
.Y(n_2552)
);

AOI22xp5_ASAP7_75t_L g2553 ( 
.A1(n_2532),
.A2(n_417),
.B1(n_418),
.B2(n_419),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_2545),
.Y(n_2554)
);

AOI22xp5_ASAP7_75t_L g2555 ( 
.A1(n_2544),
.A2(n_419),
.B1(n_420),
.B2(n_421),
.Y(n_2555)
);

AOI211xp5_ASAP7_75t_L g2556 ( 
.A1(n_2548),
.A2(n_420),
.B(n_421),
.C(n_422),
.Y(n_2556)
);

AOI22xp5_ASAP7_75t_L g2557 ( 
.A1(n_2537),
.A2(n_422),
.B1(n_423),
.B2(n_424),
.Y(n_2557)
);

AO22x2_ASAP7_75t_L g2558 ( 
.A1(n_2540),
.A2(n_423),
.B1(n_424),
.B2(n_425),
.Y(n_2558)
);

AND4x2_ASAP7_75t_L g2559 ( 
.A(n_2534),
.B(n_425),
.C(n_426),
.D(n_427),
.Y(n_2559)
);

AO22x2_ASAP7_75t_L g2560 ( 
.A1(n_2533),
.A2(n_426),
.B1(n_427),
.B2(n_428),
.Y(n_2560)
);

CKINVDCx20_ASAP7_75t_R g2561 ( 
.A(n_2541),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2549),
.Y(n_2562)
);

AOI221x1_ASAP7_75t_L g2563 ( 
.A1(n_2550),
.A2(n_2538),
.B1(n_2536),
.B2(n_2546),
.C(n_2535),
.Y(n_2563)
);

AOI211xp5_ASAP7_75t_L g2564 ( 
.A1(n_2562),
.A2(n_2547),
.B(n_2543),
.C(n_431),
.Y(n_2564)
);

OAI221xp5_ASAP7_75t_L g2565 ( 
.A1(n_2556),
.A2(n_429),
.B1(n_430),
.B2(n_431),
.C(n_432),
.Y(n_2565)
);

NOR4xp25_ASAP7_75t_L g2566 ( 
.A(n_2554),
.B(n_432),
.C(n_433),
.D(n_434),
.Y(n_2566)
);

AND4x1_ASAP7_75t_L g2567 ( 
.A(n_2557),
.B(n_433),
.C(n_434),
.D(n_435),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2558),
.Y(n_2568)
);

NAND2x1p5_ASAP7_75t_L g2569 ( 
.A(n_2568),
.B(n_2553),
.Y(n_2569)
);

AOI21x1_ASAP7_75t_L g2570 ( 
.A1(n_2567),
.A2(n_2551),
.B(n_2560),
.Y(n_2570)
);

NAND3xp33_ASAP7_75t_L g2571 ( 
.A(n_2563),
.B(n_2561),
.C(n_2555),
.Y(n_2571)
);

OAI21xp5_ASAP7_75t_L g2572 ( 
.A1(n_2564),
.A2(n_2559),
.B(n_2552),
.Y(n_2572)
);

AOI21xp5_ASAP7_75t_L g2573 ( 
.A1(n_2572),
.A2(n_2565),
.B(n_2566),
.Y(n_2573)
);

BUFx2_ASAP7_75t_L g2574 ( 
.A(n_2569),
.Y(n_2574)
);

OAI21x1_ASAP7_75t_L g2575 ( 
.A1(n_2570),
.A2(n_436),
.B(n_437),
.Y(n_2575)
);

AO22x2_ASAP7_75t_L g2576 ( 
.A1(n_2571),
.A2(n_436),
.B1(n_437),
.B2(n_438),
.Y(n_2576)
);

AOI22xp5_ASAP7_75t_L g2577 ( 
.A1(n_2571),
.A2(n_439),
.B1(n_440),
.B2(n_441),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2574),
.B(n_2577),
.Y(n_2578)
);

AOI221xp5_ASAP7_75t_L g2579 ( 
.A1(n_2573),
.A2(n_439),
.B1(n_440),
.B2(n_441),
.C(n_442),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_L g2580 ( 
.A(n_2576),
.B(n_443),
.Y(n_2580)
);

AOI21xp33_ASAP7_75t_SL g2581 ( 
.A1(n_2575),
.A2(n_443),
.B(n_444),
.Y(n_2581)
);

AOI21xp5_ASAP7_75t_L g2582 ( 
.A1(n_2578),
.A2(n_444),
.B(n_445),
.Y(n_2582)
);

INVxp67_ASAP7_75t_L g2583 ( 
.A(n_2580),
.Y(n_2583)
);

AOI21xp5_ASAP7_75t_L g2584 ( 
.A1(n_2581),
.A2(n_446),
.B(n_447),
.Y(n_2584)
);

AOI22xp5_ASAP7_75t_L g2585 ( 
.A1(n_2583),
.A2(n_2579),
.B1(n_449),
.B2(n_450),
.Y(n_2585)
);

AND2x2_ASAP7_75t_L g2586 ( 
.A(n_2585),
.B(n_2584),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2586),
.Y(n_2587)
);

AOI221xp5_ASAP7_75t_L g2588 ( 
.A1(n_2587),
.A2(n_2582),
.B1(n_451),
.B2(n_452),
.C(n_453),
.Y(n_2588)
);

AOI22xp33_ASAP7_75t_L g2589 ( 
.A1(n_2588),
.A2(n_446),
.B1(n_451),
.B2(n_452),
.Y(n_2589)
);

AOI211xp5_ASAP7_75t_L g2590 ( 
.A1(n_2589),
.A2(n_454),
.B(n_455),
.C(n_456),
.Y(n_2590)
);


endmodule