module fake_jpeg_1848_n_142 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_142);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx14_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx8_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_4),
.B(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_29),
.Y(n_30)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_0),
.C(n_2),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_17),
.C(n_27),
.Y(n_49)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_16),
.B(n_5),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_16),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_28),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_46),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_59),
.C(n_40),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_60),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g55 ( 
.A1(n_33),
.A2(n_18),
.B(n_27),
.Y(n_55)
);

OR2x2_ASAP7_75t_SL g76 ( 
.A(n_55),
.B(n_63),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_30),
.B(n_22),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_25),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_31),
.B(n_25),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_26),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_57),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_78),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_70),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

CKINVDCx11_ASAP7_75t_R g70 ( 
.A(n_48),
.Y(n_70)
);

AND2x6_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_9),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_SL g97 ( 
.A(n_71),
.B(n_76),
.C(n_15),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_49),
.A2(n_38),
.B1(n_36),
.B2(n_43),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_72),
.A2(n_77),
.B1(n_47),
.B2(n_44),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_62),
.Y(n_90)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_46),
.A2(n_35),
.B1(n_18),
.B2(n_32),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_82),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_59),
.A2(n_13),
.B(n_34),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_23),
.B(n_53),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_64),
.B(n_26),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_84),
.B(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_80),
.B(n_23),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_90),
.B(n_78),
.Y(n_105)
);

O2A1O1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_53),
.B(n_63),
.C(n_56),
.Y(n_91)
);

AO22x1_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_69),
.B1(n_65),
.B2(n_81),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_92),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_94),
.A2(n_72),
.B1(n_68),
.B2(n_74),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_47),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_97),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_100),
.A2(n_103),
.B1(n_109),
.B2(n_45),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_66),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_104),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_94),
.A2(n_92),
.B1(n_90),
.B2(n_87),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_79),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_89),
.C(n_86),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_71),
.B(n_70),
.C(n_75),
.Y(n_106)
);

A2O1A1O1Ixp25_ASAP7_75t_L g110 ( 
.A1(n_106),
.A2(n_97),
.B(n_88),
.C(n_83),
.D(n_87),
.Y(n_110)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_87),
.A2(n_44),
.B1(n_68),
.B2(n_58),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_110),
.A2(n_98),
.B(n_100),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_108),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_86),
.C(n_93),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_105),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_99),
.A2(n_96),
.B(n_93),
.Y(n_114)
);

OA21x2_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_98),
.B(n_106),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_96),
.Y(n_116)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_124),
.C(n_125),
.Y(n_126)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_123),
.A2(n_111),
.B1(n_110),
.B2(n_45),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_118),
.C(n_114),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_129),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_111),
.C(n_107),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_130),
.B(n_123),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_126),
.A2(n_120),
.B(n_123),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_133),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_121),
.B(n_28),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_0),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_131),
.A2(n_21),
.B(n_15),
.C(n_3),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_137),
.Y(n_138)
);

AOI322xp5_ASAP7_75t_L g139 ( 
.A1(n_136),
.A2(n_135),
.A3(n_9),
.B1(n_12),
.B2(n_21),
.C1(n_2),
.C2(n_3),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_0),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_138),
.B(n_3),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_4),
.Y(n_142)
);


endmodule