module fake_jpeg_13623_n_339 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_43),
.Y(n_48)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_0),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_49),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_29),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_63),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_24),
.B1(n_19),
.B2(n_20),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_51),
.A2(n_57),
.B1(n_20),
.B2(n_26),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_21),
.B(n_17),
.C(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_53),
.B(n_69),
.Y(n_92)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_39),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_54),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_24),
.B1(n_19),
.B2(n_20),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_47),
.A2(n_30),
.B1(n_25),
.B2(n_33),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_60),
.A2(n_33),
.B1(n_25),
.B2(n_30),
.Y(n_93)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_27),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_27),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_28),
.Y(n_83)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_46),
.B(n_23),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_22),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_72),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_45),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_71),
.A2(n_46),
.B1(n_45),
.B2(n_24),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_75),
.A2(n_93),
.B1(n_61),
.B2(n_22),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_SL g77 ( 
.A(n_48),
.B(n_50),
.C(n_63),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_58),
.C(n_52),
.Y(n_110)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_53),
.A2(n_34),
.B1(n_25),
.B2(n_30),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_98),
.B1(n_99),
.B2(n_101),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_83),
.B(n_81),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_84),
.A2(n_96),
.B1(n_100),
.B2(n_56),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_48),
.A2(n_21),
.B(n_17),
.C(n_22),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_90),
.A2(n_83),
.B(n_85),
.C(n_92),
.Y(n_115)
);

NAND2xp33_ASAP7_75t_SL g91 ( 
.A(n_71),
.B(n_19),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_91),
.Y(n_112)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_72),
.A2(n_20),
.B1(n_33),
.B2(n_26),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_62),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_56),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_69),
.A2(n_25),
.B1(n_30),
.B2(n_34),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_62),
.A2(n_21),
.B1(n_17),
.B2(n_22),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_56),
.A2(n_26),
.B1(n_28),
.B2(n_35),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_65),
.A2(n_35),
.B1(n_26),
.B2(n_28),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_103),
.B(n_113),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_89),
.B(n_16),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_109),
.B(n_111),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_91),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_76),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_81),
.B(n_58),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_124),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_82),
.A2(n_65),
.B1(n_55),
.B2(n_67),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_116),
.A2(n_118),
.B1(n_75),
.B2(n_74),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_92),
.A2(n_65),
.B1(n_55),
.B2(n_67),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_117),
.A2(n_125),
.B1(n_128),
.B2(n_73),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_67),
.B1(n_55),
.B2(n_70),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_76),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_126),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_85),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_121),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_122),
.A2(n_74),
.B1(n_95),
.B2(n_84),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_70),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_86),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_93),
.A2(n_61),
.B1(n_54),
.B2(n_26),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_26),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_79),
.Y(n_146)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_104),
.Y(n_131)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_131),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_132),
.A2(n_158),
.B1(n_18),
.B2(n_1),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_130),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_139),
.Y(n_168)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_117),
.Y(n_172)
);

AO22x1_ASAP7_75t_SL g138 ( 
.A1(n_120),
.A2(n_78),
.B1(n_88),
.B2(n_77),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_138),
.B(n_146),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_111),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_140),
.A2(n_144),
.B1(n_160),
.B2(n_128),
.Y(n_173)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_100),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_142),
.A2(n_161),
.B(n_49),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_107),
.A2(n_96),
.B1(n_99),
.B2(n_101),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_143),
.A2(n_125),
.B1(n_119),
.B2(n_105),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_129),
.A2(n_97),
.B1(n_94),
.B2(n_87),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_80),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_152),
.C(n_123),
.Y(n_162)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_79),
.C(n_73),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_16),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_154),
.B(n_156),
.Y(n_167)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_103),
.B(n_14),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_107),
.A2(n_54),
.B1(n_56),
.B2(n_49),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_112),
.A2(n_49),
.B(n_22),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_162),
.B(n_170),
.C(n_174),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_148),
.B(n_113),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_163),
.B(n_147),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_150),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_164),
.B(n_176),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_157),
.B(n_126),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_165),
.B(n_181),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_142),
.A2(n_116),
.B1(n_115),
.B2(n_118),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_169),
.A2(n_180),
.B1(n_193),
.B2(n_160),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_121),
.C(n_112),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_172),
.B(n_18),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_173),
.A2(n_179),
.B1(n_18),
.B2(n_1),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_115),
.C(n_105),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_150),
.Y(n_176)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_178),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_142),
.A2(n_106),
.B1(n_114),
.B2(n_102),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_106),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_139),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_182),
.B(n_2),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_138),
.B(n_106),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_184),
.B(n_194),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_114),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_192),
.C(n_18),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_188),
.A2(n_191),
.B(n_153),
.Y(n_210)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_135),
.Y(n_189)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_189),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_133),
.A2(n_102),
.B1(n_22),
.B2(n_18),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_145),
.B(n_18),
.C(n_13),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_145),
.B(n_13),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_195),
.A2(n_200),
.B1(n_201),
.B2(n_191),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_179),
.A2(n_158),
.B1(n_146),
.B2(n_159),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_197),
.A2(n_199),
.B1(n_204),
.B2(n_212),
.Y(n_224)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_198),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_173),
.A2(n_159),
.B1(n_133),
.B2(n_134),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_169),
.A2(n_144),
.B1(n_140),
.B2(n_138),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_164),
.A2(n_138),
.B1(n_131),
.B2(n_151),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_202),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_203),
.B(n_214),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_190),
.A2(n_152),
.B1(n_136),
.B2(n_161),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_182),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_211),
.Y(n_225)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_210),
.A2(n_219),
.B(n_222),
.Y(n_246)
);

OAI32xp33_ASAP7_75t_L g211 ( 
.A1(n_190),
.A2(n_155),
.A3(n_141),
.B1(n_12),
.B2(n_3),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_177),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_183),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_163),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_218),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_172),
.C(n_183),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_188),
.A2(n_0),
.B(n_1),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_175),
.Y(n_220)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_175),
.Y(n_221)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_176),
.A2(n_0),
.B(n_2),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_223),
.Y(n_226)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_228),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_239),
.C(n_248),
.Y(n_264)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_230),
.Y(n_262)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_231),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_187),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_238),
.Y(n_259)
);

AND2x4_ASAP7_75t_L g235 ( 
.A(n_199),
.B(n_180),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_235),
.A2(n_5),
.B(n_6),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_197),
.A2(n_170),
.B1(n_174),
.B2(n_162),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_236),
.A2(n_240),
.B1(n_237),
.B2(n_239),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_216),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_198),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_186),
.C(n_185),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_204),
.A2(n_192),
.B1(n_186),
.B2(n_185),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_205),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_243),
.B(n_245),
.Y(n_271)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_207),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_208),
.B(n_171),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_250),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_171),
.C(n_189),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_201),
.B(n_177),
.C(n_178),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_5),
.C(n_6),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_200),
.A2(n_167),
.B1(n_3),
.B2(n_4),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_225),
.A2(n_243),
.B(n_210),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_SL g277 ( 
.A1(n_251),
.A2(n_266),
.B(n_246),
.C(n_235),
.Y(n_277)
);

NOR2xp67_ASAP7_75t_SL g252 ( 
.A(n_248),
.B(n_203),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_252),
.A2(n_247),
.B(n_249),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_255),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_256),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_217),
.Y(n_255)
);

XNOR2x1_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_195),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_244),
.A2(n_213),
.B1(n_221),
.B2(n_220),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_257),
.A2(n_263),
.B1(n_268),
.B2(n_242),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_196),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_272),
.Y(n_285)
);

MAJx2_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_209),
.C(n_202),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_265),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_225),
.A2(n_222),
.B1(n_219),
.B2(n_196),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_207),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_246),
.A2(n_2),
.B(n_3),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_227),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_234),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_273),
.A2(n_271),
.B(n_266),
.Y(n_290)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_267),
.Y(n_274)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_274),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_269),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_251),
.A2(n_224),
.B1(n_231),
.B2(n_250),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_278),
.B(n_287),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_254),
.C(n_256),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_286),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_262),
.Y(n_300)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_258),
.A2(n_228),
.B1(n_242),
.B2(n_241),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_270),
.C(n_261),
.Y(n_295)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_285),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_241),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_224),
.C(n_235),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_233),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_288),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_235),
.C(n_233),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_262),
.C(n_245),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_290),
.A2(n_303),
.B1(n_293),
.B2(n_282),
.Y(n_309)
);

A2O1A1Ixp33_ASAP7_75t_SL g291 ( 
.A1(n_277),
.A2(n_258),
.B(n_267),
.C(n_271),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_291),
.B(n_277),
.C(n_6),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_293),
.A2(n_5),
.B(n_7),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_259),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_295),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_272),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_301),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_289),
.Y(n_307)
);

NOR3xp33_ASAP7_75t_SL g303 ( 
.A(n_277),
.B(n_230),
.C(n_6),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_275),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_309),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_307),
.B(n_310),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_280),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_298),
.A2(n_282),
.B1(n_281),
.B2(n_280),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_312),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_279),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_313),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_11),
.C(n_7),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_316),
.C(n_291),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_315),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_299),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_306),
.B(n_297),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_319),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_304),
.C(n_307),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_318),
.A2(n_310),
.B(n_314),
.Y(n_327)
);

AOI322xp5_ASAP7_75t_L g322 ( 
.A1(n_313),
.A2(n_303),
.A3(n_291),
.B1(n_10),
.B2(n_11),
.C1(n_8),
.C2(n_7),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_316),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_327),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_324),
.C(n_325),
.Y(n_328)
);

AO21x1_ASAP7_75t_L g334 ( 
.A1(n_328),
.A2(n_329),
.B(n_330),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_315),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_323),
.A2(n_291),
.B1(n_8),
.B2(n_10),
.Y(n_331)
);

AOI211x1_ASAP7_75t_L g333 ( 
.A1(n_331),
.A2(n_332),
.B(n_321),
.C(n_10),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_8),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_333),
.B(n_326),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_335),
.B(n_328),
.Y(n_337)
);

XNOR2x2_ASAP7_75t_SL g338 ( 
.A(n_337),
.B(n_334),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_332),
.Y(n_339)
);


endmodule