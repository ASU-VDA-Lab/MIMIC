module fake_jpeg_25437_n_329 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_19),
.Y(n_57)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_55),
.Y(n_64)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_34),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_33),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_34),
.B1(n_18),
.B2(n_30),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_60),
.A2(n_26),
.B1(n_29),
.B2(n_21),
.Y(n_91)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_72),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_69),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_75),
.Y(n_100)
);

AO22x2_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_43),
.B1(n_42),
.B2(n_39),
.Y(n_74)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_74),
.A2(n_70),
.B1(n_82),
.B2(n_81),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_53),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_79),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_28),
.B(n_1),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_85),
.Y(n_97)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_46),
.A2(n_28),
.B1(n_26),
.B2(n_29),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_80),
.A2(n_26),
.B1(n_29),
.B2(n_33),
.Y(n_106)
);

NAND2xp33_ASAP7_75t_SL g81 ( 
.A(n_47),
.B(n_32),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_54),
.Y(n_102)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_84),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_28),
.B1(n_30),
.B2(n_18),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_83),
.A2(n_91),
.B1(n_48),
.B2(n_16),
.Y(n_110)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_28),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_87),
.Y(n_109)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_90),
.Y(n_112)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_73),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_94),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_78),
.B1(n_85),
.B2(n_49),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_93),
.A2(n_98),
.B1(n_110),
.B2(n_114),
.Y(n_127)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_74),
.A2(n_54),
.B1(n_58),
.B2(n_52),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_28),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_108),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_102),
.A2(n_38),
.B(n_32),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_67),
.B(n_21),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_103),
.B(n_25),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_106),
.A2(n_113),
.B1(n_119),
.B2(n_76),
.Y(n_123)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_64),
.B(n_23),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_65),
.B1(n_71),
.B2(n_88),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_74),
.A2(n_23),
.B1(n_19),
.B2(n_20),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_74),
.A2(n_77),
.B1(n_79),
.B2(n_87),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_84),
.A2(n_68),
.B1(n_90),
.B2(n_70),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_71),
.B1(n_88),
.B2(n_65),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_20),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_117),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_20),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_69),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_75),
.A2(n_23),
.B1(n_19),
.B2(n_20),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

OAI21xp33_ASAP7_75t_SL g121 ( 
.A1(n_99),
.A2(n_97),
.B(n_108),
.Y(n_121)
);

AO21x1_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_122),
.B(n_102),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_92),
.A2(n_66),
.B1(n_65),
.B2(n_76),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_123),
.A2(n_143),
.B1(n_110),
.B2(n_98),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_124),
.B(n_129),
.Y(n_163)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_94),
.B(n_88),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_137),
.Y(n_157)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_130),
.A2(n_141),
.B1(n_113),
.B2(n_117),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_138),
.Y(n_158)
);

OA22x2_ASAP7_75t_L g167 ( 
.A1(n_133),
.A2(n_139),
.B1(n_107),
.B2(n_111),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_134),
.A2(n_148),
.B(n_104),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_135),
.B(n_136),
.Y(n_180)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

OAI22x1_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_32),
.B1(n_31),
.B2(n_16),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_142),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_27),
.B1(n_23),
.B2(n_25),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_97),
.A2(n_27),
.B1(n_31),
.B2(n_25),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_102),
.B(n_22),
.C(n_16),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_105),
.C(n_116),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_103),
.B(n_22),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_109),
.Y(n_159)
);

AOI21xp33_ASAP7_75t_L g148 ( 
.A1(n_96),
.A2(n_22),
.B(n_15),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_149),
.A2(n_151),
.B(n_156),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_150),
.A2(n_167),
.B1(n_171),
.B2(n_0),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_111),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_96),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_152),
.B(n_155),
.Y(n_195)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_154),
.B(n_161),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_102),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_93),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_159),
.B(n_170),
.Y(n_199)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_162),
.A2(n_147),
.B1(n_144),
.B2(n_138),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_134),
.A2(n_139),
.B(n_125),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_164),
.A2(n_168),
.B(n_174),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_111),
.Y(n_165)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_165),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_169),
.Y(n_196)
);

MAJx2_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_109),
.C(n_115),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_112),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_123),
.A2(n_107),
.B1(n_106),
.B2(n_118),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_104),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_172),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_119),
.Y(n_173)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_0),
.B(n_1),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_127),
.A2(n_27),
.B1(n_31),
.B2(n_15),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_175),
.A2(n_174),
.B1(n_141),
.B2(n_156),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_27),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_178),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_127),
.B(n_14),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_130),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_181),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_124),
.B(n_14),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_182),
.A2(n_188),
.B1(n_191),
.B2(n_204),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_201),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_180),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_184),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_156),
.A2(n_165),
.B1(n_150),
.B2(n_179),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_149),
.A2(n_146),
.B(n_132),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_189),
.A2(n_149),
.B(n_151),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_190),
.A2(n_209),
.B1(n_153),
.B2(n_177),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_175),
.A2(n_144),
.B1(n_120),
.B2(n_2),
.Y(n_191)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

AOI32xp33_ASAP7_75t_L g200 ( 
.A1(n_168),
.A2(n_144),
.A3(n_13),
.B1(n_2),
.B2(n_3),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_8),
.Y(n_236)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_157),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_157),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_210),
.Y(n_225)
);

OAI32xp33_ASAP7_75t_L g203 ( 
.A1(n_169),
.A2(n_13),
.A3(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_203)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_203),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_173),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_205),
.A2(n_153),
.B1(n_154),
.B2(n_161),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_160),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_206),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_164),
.A2(n_5),
.B(n_6),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_208),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_151),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_159),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_163),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_211),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_199),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_219),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_152),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_218),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_214),
.B(n_223),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_216),
.A2(n_227),
.B1(n_229),
.B2(n_230),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_195),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_198),
.Y(n_219)
);

OAI21x1_ASAP7_75t_R g224 ( 
.A1(n_183),
.A2(n_167),
.B(n_162),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_224),
.A2(n_186),
.B(n_191),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_211),
.A2(n_167),
.B1(n_178),
.B2(n_166),
.Y(n_226)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_192),
.A2(n_167),
.B1(n_155),
.B2(n_176),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_5),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_237),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_188),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_182),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_187),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_185),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_197),
.Y(n_235)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_235),
.Y(n_247)
);

NOR3xp33_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_203),
.C(n_208),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_207),
.B(n_9),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_207),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_240),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_210),
.C(n_202),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_246),
.C(n_248),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_234),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_245),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_201),
.C(n_189),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_192),
.C(n_197),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_222),
.A2(n_194),
.B1(n_190),
.B2(n_186),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_249),
.A2(n_224),
.B1(n_215),
.B2(n_222),
.Y(n_262)
);

O2A1O1Ixp33_ASAP7_75t_L g275 ( 
.A1(n_250),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_275)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_224),
.Y(n_252)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_252),
.Y(n_274)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_253),
.B(n_255),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_194),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_9),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_223),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_216),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_193),
.C(n_209),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_229),
.C(n_230),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_257),
.Y(n_259)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_259),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_262),
.A2(n_270),
.B1(n_275),
.B2(n_250),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_244),
.Y(n_284)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_212),
.Y(n_266)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_266),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_254),
.B(n_228),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_273),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_243),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_252),
.A2(n_220),
.B1(n_231),
.B2(n_233),
.Y(n_269)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_256),
.A2(n_233),
.B1(n_217),
.B2(n_11),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_249),
.A2(n_217),
.B(n_10),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_271),
.B(n_247),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_241),
.C(n_239),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_278),
.C(n_279),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_246),
.C(n_240),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_238),
.C(n_248),
.Y(n_279)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_280),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_281),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_285),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_244),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_287),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_288),
.B(n_243),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_264),
.B(n_272),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_289),
.B(n_261),
.Y(n_291)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_291),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_290),
.A2(n_258),
.B1(n_274),
.B2(n_262),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_297),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_275),
.Y(n_297)
);

AO21x1_ASAP7_75t_L g298 ( 
.A1(n_283),
.A2(n_265),
.B(n_271),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_299),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_270),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_273),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_303),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_302),
.B(n_267),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_277),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_278),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_309),
.C(n_293),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_276),
.Y(n_307)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_307),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_279),
.C(n_282),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_282),
.Y(n_310)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_310),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_313),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_10),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_299),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_317),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_315),
.Y(n_323)
);

NOR2x1_ASAP7_75t_R g316 ( 
.A(n_312),
.B(n_300),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_316),
.B(n_309),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_295),
.C(n_292),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_318),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_324),
.Y(n_325)
);

AOI321xp33_ASAP7_75t_SL g326 ( 
.A1(n_325),
.A2(n_323),
.A3(n_322),
.B1(n_319),
.B2(n_320),
.C(n_314),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_308),
.C(n_306),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_298),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_10),
.B(n_11),
.Y(n_329)
);


endmodule