module fake_jpeg_29391_n_34 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_34);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_34;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;
wire n_15;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_12),
.Y(n_17)
);

OA22x2_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_19),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_17),
.B(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_2),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_21),
.B(n_15),
.Y(n_26)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_24),
.B1(n_26),
.B2(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_13),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_29),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_14),
.C(n_16),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_3),
.B(n_4),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_4),
.B(n_10),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_31),
.C(n_28),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_25),
.Y(n_34)
);


endmodule