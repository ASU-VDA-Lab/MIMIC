module real_jpeg_12967_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_70;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_4),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_4),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_4),
.B(n_24),
.C(n_41),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_4),
.A2(n_31),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_4),
.B(n_42),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_4),
.B(n_22),
.C(n_28),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_4),
.B(n_51),
.C(n_66),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_4),
.B(n_139),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_6),
.A2(n_51),
.B1(n_52),
.B2(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_9),
.A2(n_51),
.B1(n_52),
.B2(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_9),
.Y(n_90)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_96),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_94),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_77),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_14),
.B(n_77),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_58),
.C(n_73),
.Y(n_14)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_15),
.B(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_17),
.B1(n_44),
.B2(n_57),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_16),
.A2(n_17),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_32),
.B2(n_43),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_18),
.B(n_43),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_18),
.A2(n_19),
.B1(n_63),
.B2(n_64),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_18),
.B(n_48),
.C(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_18),
.A2(n_19),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_19),
.B(n_32),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_19),
.B(n_63),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_19),
.A2(n_63),
.B(n_116),
.C(n_121),
.Y(n_115)
);

AO21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_27),
.B(n_30),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_27),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_21)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

OA22x2_ASAP7_75t_SL g27 ( 
.A1(n_22),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

AO22x1_ASAP7_75t_L g42 ( 
.A1(n_23),
.A2(n_24),
.B1(n_40),
.B2(n_41),
.Y(n_42)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_24),
.B(n_120),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_27),
.Y(n_139)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_28),
.A2(n_29),
.B1(n_66),
.B2(n_67),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_28),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_31),
.B(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_31),
.B(n_55),
.Y(n_148)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_32),
.A2(n_43),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_37),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_35),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_47),
.Y(n_46)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_42),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_42),
.Y(n_38)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI211xp5_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_64),
.B(n_75),
.C(n_76),
.Y(n_74)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_44),
.A2(n_79),
.B(n_80),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_48),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_45),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_48),
.A2(n_49),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_48),
.A2(n_49),
.B1(n_110),
.B2(n_111),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_48),
.B(n_118),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_48),
.A2(n_49),
.B1(n_136),
.B2(n_140),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_48),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_48),
.B(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_48),
.B(n_64),
.C(n_137),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_49),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_54),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_55),
.Y(n_56)
);

AO22x1_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_52),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

INVx5_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_52),
.B(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_55),
.A2(n_56),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_55),
.A2(n_56),
.B1(n_61),
.B2(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_58),
.A2(n_73),
.B1(n_74),
.B2(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_63),
.B1(n_64),
.B2(n_72),
.Y(n_58)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_64),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_63),
.A2(n_64),
.B1(n_88),
.B2(n_91),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_63),
.A2(n_64),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_63),
.B(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_63),
.A2(n_64),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_63),
.A2(n_64),
.B1(n_133),
.B2(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_64),
.B(n_123),
.C(n_127),
.Y(n_162)
);

OA21x2_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_69),
.B(n_71),
.Y(n_64)
);

NOR2x1_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_65),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B1(n_82),
.B2(n_93),
.Y(n_77)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_86),
.B1(n_87),
.B2(n_92),
.Y(n_82)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_84),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_164),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_112),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_100),
.B(n_103),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.C(n_109),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_104),
.B(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_105),
.A2(n_106),
.B1(n_116),
.B2(n_117),
.Y(n_154)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_158),
.B(n_163),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_129),
.B(n_157),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_122),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_115),
.B(n_122),
.Y(n_157)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_153),
.B(n_156),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_141),
.B(n_152),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_135),
.Y(n_152)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_136),
.Y(n_140)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_149),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_154),
.B(n_155),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_162),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);


endmodule