module fake_netlist_5_1647_n_1772 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1772);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1772;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1726;
wire n_665;
wire n_1584;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1752;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_131),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_119),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_53),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_151),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_27),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_85),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_20),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_2),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_68),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_123),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_90),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_29),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_156),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_132),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_159),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_28),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_41),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_77),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_60),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_135),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_112),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_154),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_21),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_88),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_6),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_54),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_138),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g191 ( 
.A(n_23),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_37),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_62),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_142),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_137),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_48),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_58),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_12),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_39),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_3),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_95),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_0),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_38),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_16),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_33),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_126),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_23),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_71),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_146),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_79),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_161),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_114),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_162),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_3),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_145),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_152),
.Y(n_216)
);

BUFx8_ASAP7_75t_SL g217 ( 
.A(n_153),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_25),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_116),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_75),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_7),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_98),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_134),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_52),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_106),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_99),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_40),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_22),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_8),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_67),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_100),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_117),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_5),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_55),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_115),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_39),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_50),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_25),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_66),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_17),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_9),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_122),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_160),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_118),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_89),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_121),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_136),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_4),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_84),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_20),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_53),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_87),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_63),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_130),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_92),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_69),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_0),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_29),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_125),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_40),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_148),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_128),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_10),
.Y(n_263)
);

BUFx5_ASAP7_75t_L g264 ( 
.A(n_36),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_21),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_96),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_110),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_83),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_157),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_35),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_94),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_59),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_104),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_59),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_72),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_64),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_36),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_93),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_15),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_8),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_1),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_113),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_28),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_73),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_147),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_109),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_14),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_41),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_19),
.Y(n_289)
);

BUFx5_ASAP7_75t_L g290 ( 
.A(n_22),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_14),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_4),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_18),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_65),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_17),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_51),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_48),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_10),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_103),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_78),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_163),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_30),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_16),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_56),
.Y(n_304)
);

BUFx5_ASAP7_75t_L g305 ( 
.A(n_32),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_56),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_158),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_80),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_26),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_143),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_26),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_81),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_30),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_7),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_70),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_13),
.Y(n_316)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_144),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_129),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_45),
.Y(n_319)
);

BUFx10_ASAP7_75t_L g320 ( 
.A(n_150),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_74),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_217),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_264),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_176),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_192),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_264),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_264),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_264),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_264),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_264),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_194),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_264),
.Y(n_332)
);

NOR2xp67_ASAP7_75t_L g333 ( 
.A(n_260),
.B(n_1),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_264),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_290),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_195),
.Y(n_336)
);

NOR2xp67_ASAP7_75t_L g337 ( 
.A(n_311),
.B(n_2),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_201),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_263),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_283),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_185),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_290),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_290),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_206),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_171),
.Y(n_345)
);

INVxp33_ASAP7_75t_SL g346 ( 
.A(n_204),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_290),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_208),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_212),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_254),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_210),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_213),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_210),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_215),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_290),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_166),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_290),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_255),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_290),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_308),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_216),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_310),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_290),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_219),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_305),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_320),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_225),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_223),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_305),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_305),
.B(n_5),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_235),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_275),
.B(n_6),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_242),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_305),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_244),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_305),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_245),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_246),
.Y(n_378)
);

NOR2xp67_ASAP7_75t_L g379 ( 
.A(n_238),
.B(n_9),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_305),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_191),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_179),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_L g383 ( 
.A(n_238),
.B(n_11),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_305),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_305),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_247),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_166),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_166),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_252),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_166),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_166),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_171),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_175),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_253),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_256),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_175),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_175),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_175),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_262),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_387),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_343),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_343),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_323),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_323),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_326),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_356),
.B(n_175),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_387),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_388),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_382),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_326),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_388),
.Y(n_411)
);

AND2x4_ASAP7_75t_SL g412 ( 
.A(n_367),
.B(n_320),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_327),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_327),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_356),
.B(n_240),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_390),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_328),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_390),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_346),
.A2(n_280),
.B1(n_289),
.B2(n_170),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_328),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_356),
.B(n_211),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_329),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_351),
.B(n_211),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_391),
.B(n_240),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_391),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_393),
.B(n_240),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_393),
.B(n_285),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_396),
.Y(n_428)
);

OAI21x1_ASAP7_75t_L g429 ( 
.A1(n_370),
.A2(n_177),
.B(n_173),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_329),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_396),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_397),
.B(n_240),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_351),
.B(n_285),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_330),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_330),
.Y(n_435)
);

AND2x6_ASAP7_75t_L g436 ( 
.A(n_332),
.B(n_173),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_397),
.B(n_240),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_332),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_372),
.B(n_320),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_398),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_398),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_334),
.B(n_243),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_366),
.A2(n_234),
.B1(n_248),
.B2(n_277),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_334),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_335),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_366),
.B(n_314),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_335),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_342),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_342),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_347),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_347),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_355),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_355),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_357),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_357),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_359),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_359),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_345),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_363),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_363),
.Y(n_460)
);

CKINVDCx8_ASAP7_75t_R g461 ( 
.A(n_325),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_365),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_365),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_369),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_369),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_374),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_374),
.Y(n_467)
);

CKINVDCx6p67_ASAP7_75t_R g468 ( 
.A(n_325),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_345),
.Y(n_469)
);

INVx6_ASAP7_75t_L g470 ( 
.A(n_353),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_376),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_324),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_376),
.B(n_314),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_470),
.B(n_331),
.Y(n_474)
);

NAND3xp33_ASAP7_75t_L g475 ( 
.A(n_439),
.B(n_368),
.C(n_338),
.Y(n_475)
);

OR2x6_ASAP7_75t_L g476 ( 
.A(n_446),
.B(n_333),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_439),
.B(n_336),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_446),
.B(n_344),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g479 ( 
.A(n_472),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_445),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_401),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_470),
.B(n_348),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_409),
.B(n_349),
.Y(n_483)
);

NAND3xp33_ASAP7_75t_L g484 ( 
.A(n_409),
.B(n_354),
.C(n_352),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_445),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_423),
.B(n_353),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_470),
.B(n_361),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_455),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_419),
.A2(n_304),
.B1(n_337),
.B2(n_292),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_458),
.B(n_364),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_405),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_405),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_470),
.B(n_373),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_461),
.B(n_377),
.Y(n_494)
);

BUFx4f_ASAP7_75t_L g495 ( 
.A(n_405),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_405),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_419),
.A2(n_179),
.B1(n_182),
.B2(n_180),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_458),
.Y(n_498)
);

INVxp67_ASAP7_75t_SL g499 ( 
.A(n_444),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_401),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_469),
.B(n_378),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_401),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_455),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_457),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_401),
.Y(n_505)
);

OR2x6_ASAP7_75t_L g506 ( 
.A(n_423),
.B(n_279),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_423),
.B(n_433),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_405),
.Y(n_508)
);

NAND2xp33_ASAP7_75t_L g509 ( 
.A(n_436),
.B(n_232),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_457),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_402),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_470),
.B(n_386),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_402),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_469),
.B(n_394),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_443),
.A2(n_241),
.B1(n_182),
.B2(n_186),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_402),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_470),
.Y(n_517)
);

OAI22xp33_ASAP7_75t_L g518 ( 
.A1(n_461),
.A2(n_339),
.B1(n_340),
.B2(n_379),
.Y(n_518)
);

CKINVDCx16_ASAP7_75t_R g519 ( 
.A(n_443),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_468),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_470),
.B(n_399),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_450),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_433),
.B(n_371),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_450),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_450),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_433),
.A2(n_180),
.B1(n_272),
.B2(n_186),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_452),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_402),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_461),
.B(n_339),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_452),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_442),
.B(n_392),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_442),
.B(n_380),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_442),
.B(n_380),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_442),
.B(n_427),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_412),
.B(n_340),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_452),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_403),
.Y(n_537)
);

AND2x2_ASAP7_75t_SL g538 ( 
.A(n_442),
.B(n_177),
.Y(n_538)
);

INVxp33_ASAP7_75t_L g539 ( 
.A(n_421),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_412),
.A2(n_395),
.B1(n_389),
.B2(n_375),
.Y(n_540)
);

BUFx10_ASAP7_75t_L g541 ( 
.A(n_412),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_472),
.Y(n_542)
);

AND2x6_ASAP7_75t_L g543 ( 
.A(n_442),
.B(n_220),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_427),
.B(n_392),
.Y(n_544)
);

NAND2x1p5_ASAP7_75t_L g545 ( 
.A(n_429),
.B(n_181),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_403),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_403),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_462),
.B(n_322),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_462),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_468),
.Y(n_550)
);

INVx4_ASAP7_75t_L g551 ( 
.A(n_405),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_412),
.B(n_381),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_403),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_404),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_404),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_404),
.Y(n_556)
);

BUFx8_ASAP7_75t_SL g557 ( 
.A(n_468),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_462),
.B(n_465),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_404),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_465),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_465),
.B(n_384),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_466),
.Y(n_562)
);

NAND2x1p5_ASAP7_75t_L g563 ( 
.A(n_429),
.B(n_183),
.Y(n_563)
);

BUFx4f_ASAP7_75t_L g564 ( 
.A(n_405),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_417),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_466),
.Y(n_566)
);

NAND2xp33_ASAP7_75t_R g567 ( 
.A(n_429),
.B(n_164),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_466),
.B(n_384),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_417),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_467),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_427),
.B(n_164),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_405),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_410),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_467),
.B(n_385),
.Y(n_574)
);

BUFx10_ASAP7_75t_L g575 ( 
.A(n_421),
.Y(n_575)
);

NAND3xp33_ASAP7_75t_L g576 ( 
.A(n_427),
.B(n_383),
.C(n_198),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_410),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_467),
.Y(n_578)
);

OR2x6_ASAP7_75t_L g579 ( 
.A(n_421),
.B(n_279),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_410),
.Y(n_580)
);

OAI22xp33_ASAP7_75t_L g581 ( 
.A1(n_473),
.A2(n_197),
.B1(n_200),
.B2(n_199),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_417),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_427),
.B(n_341),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_406),
.Y(n_584)
);

NAND2xp33_ASAP7_75t_L g585 ( 
.A(n_436),
.B(n_232),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_427),
.B(n_165),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_421),
.A2(n_314),
.B1(n_168),
.B2(n_302),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_406),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_410),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_417),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_421),
.Y(n_591)
);

INVxp67_ASAP7_75t_SL g592 ( 
.A(n_444),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_410),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_410),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_420),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_415),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_444),
.B(n_385),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_420),
.Y(n_598)
);

AND2x6_ASAP7_75t_L g599 ( 
.A(n_444),
.B(n_220),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_444),
.B(n_350),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g601 ( 
.A(n_415),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_420),
.Y(n_602)
);

INVx6_ASAP7_75t_L g603 ( 
.A(n_410),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_454),
.Y(n_604)
);

NAND2xp33_ASAP7_75t_L g605 ( 
.A(n_436),
.B(n_232),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_473),
.B(n_237),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_471),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_454),
.A2(n_314),
.B1(n_302),
.B2(n_168),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_408),
.B(n_237),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_471),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_424),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_410),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_420),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_454),
.B(n_243),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_454),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_471),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_471),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_424),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_454),
.B(n_456),
.Y(n_619)
);

INVx4_ASAP7_75t_L g620 ( 
.A(n_413),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_456),
.Y(n_621)
);

NOR3xp33_ASAP7_75t_L g622 ( 
.A(n_426),
.B(n_249),
.C(n_209),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_413),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_534),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_534),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_507),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_498),
.B(n_188),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_522),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_477),
.B(n_266),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_601),
.B(n_456),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_538),
.B(n_456),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_522),
.Y(n_632)
);

AOI22x1_ASAP7_75t_L g633 ( 
.A1(n_545),
.A2(n_563),
.B1(n_588),
.B2(n_584),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_538),
.A2(n_291),
.B1(n_203),
.B2(n_196),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_601),
.B(n_456),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_611),
.B(n_464),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_575),
.Y(n_637)
);

OR2x2_ASAP7_75t_L g638 ( 
.A(n_479),
.B(n_188),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_611),
.B(n_464),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_507),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_575),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_486),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_486),
.Y(n_643)
);

INVx8_ASAP7_75t_L g644 ( 
.A(n_579),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_538),
.A2(n_288),
.B1(n_218),
.B2(n_228),
.Y(n_645)
);

NAND2xp33_ASAP7_75t_L g646 ( 
.A(n_543),
.B(n_267),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_480),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_490),
.B(n_300),
.Y(n_648)
);

NAND2x1p5_ASAP7_75t_L g649 ( 
.A(n_591),
.B(n_222),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_600),
.A2(n_362),
.B1(n_358),
.B2(n_360),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_584),
.A2(n_189),
.B1(n_287),
.B2(n_295),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_531),
.B(n_191),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_544),
.B(n_251),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_618),
.B(n_464),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_481),
.Y(n_655)
);

A2O1A1Ixp33_ASAP7_75t_L g656 ( 
.A1(n_588),
.A2(n_257),
.B(n_313),
.C(n_306),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_480),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_596),
.A2(n_273),
.B1(n_276),
.B2(n_317),
.Y(n_658)
);

BUFx6f_ASAP7_75t_SL g659 ( 
.A(n_541),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_524),
.Y(n_660)
);

INVxp67_ASAP7_75t_L g661 ( 
.A(n_501),
.Y(n_661)
);

NAND2xp33_ASAP7_75t_L g662 ( 
.A(n_543),
.B(n_269),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_485),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_618),
.B(n_464),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_606),
.Y(n_665)
);

INVx8_ASAP7_75t_L g666 ( 
.A(n_579),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_596),
.B(n_485),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_575),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_591),
.Y(n_669)
);

OAI221xp5_ASAP7_75t_L g670 ( 
.A1(n_489),
.A2(n_251),
.B1(n_273),
.B2(n_276),
.C(n_317),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_488),
.B(n_464),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_606),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_514),
.B(n_165),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_481),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_478),
.B(n_484),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_609),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_503),
.B(n_413),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_R g678 ( 
.A(n_520),
.B(n_167),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_525),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_503),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_609),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_532),
.B(n_413),
.Y(n_682)
);

NOR2xp67_ASAP7_75t_L g683 ( 
.A(n_475),
.B(n_426),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_504),
.B(n_413),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_525),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_539),
.A2(n_437),
.B(n_432),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_504),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_510),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_510),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_527),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_544),
.B(n_230),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_517),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_527),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_579),
.B(n_231),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_530),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_476),
.B(n_167),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_517),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_499),
.B(n_413),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_500),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_533),
.B(n_413),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_531),
.B(n_191),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_592),
.B(n_414),
.Y(n_702)
);

INVxp67_ASAP7_75t_L g703 ( 
.A(n_542),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_558),
.B(n_414),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_536),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_536),
.B(n_414),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_579),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_476),
.B(n_169),
.Y(n_708)
);

AO22x2_ASAP7_75t_L g709 ( 
.A1(n_540),
.A2(n_226),
.B1(n_239),
.B2(n_299),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_549),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_549),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_560),
.B(n_414),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_476),
.A2(n_226),
.B1(n_239),
.B2(n_299),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_560),
.B(n_414),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_562),
.B(n_414),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_562),
.B(n_414),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_476),
.A2(n_278),
.B1(n_286),
.B2(n_282),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_483),
.B(n_169),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_519),
.B(n_241),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_566),
.B(n_414),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_523),
.B(n_202),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_566),
.Y(n_722)
);

INVxp67_ASAP7_75t_L g723 ( 
.A(n_548),
.Y(n_723)
);

BUFx6f_ASAP7_75t_SL g724 ( 
.A(n_541),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_570),
.B(n_430),
.Y(n_725)
);

BUFx2_ASAP7_75t_L g726 ( 
.A(n_583),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_578),
.B(n_430),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_578),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_619),
.B(n_430),
.Y(n_729)
);

NOR3xp33_ASAP7_75t_L g730 ( 
.A(n_519),
.B(n_227),
.C(n_205),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_604),
.B(n_430),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_604),
.B(n_430),
.Y(n_732)
);

O2A1O1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_581),
.A2(n_586),
.B(n_571),
.C(n_561),
.Y(n_733)
);

INVxp67_ASAP7_75t_L g734 ( 
.A(n_552),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_615),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_615),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_621),
.B(n_430),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_567),
.A2(n_271),
.B1(n_174),
.B2(n_178),
.Y(n_738)
);

A2O1A1Ixp33_ASAP7_75t_L g739 ( 
.A1(n_497),
.A2(n_278),
.B(n_259),
.C(n_261),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_557),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_621),
.B(n_430),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_474),
.B(n_447),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_506),
.B(n_518),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_482),
.B(n_447),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_487),
.B(n_447),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_568),
.Y(n_746)
);

NOR3xp33_ASAP7_75t_L g747 ( 
.A(n_529),
.B(n_221),
.C(n_207),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_493),
.B(n_447),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_583),
.Y(n_749)
);

NAND2x1p5_ASAP7_75t_L g750 ( 
.A(n_494),
.B(n_268),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_599),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_506),
.B(n_526),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_506),
.B(n_172),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_576),
.A2(n_172),
.B1(n_174),
.B2(n_178),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_574),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_502),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_512),
.B(n_447),
.Y(n_757)
);

BUFx6f_ASAP7_75t_SL g758 ( 
.A(n_541),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_521),
.B(n_447),
.Y(n_759)
);

A2O1A1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_497),
.A2(n_515),
.B(n_526),
.C(n_622),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_505),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_506),
.B(n_284),
.Y(n_762)
);

A2O1A1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_515),
.A2(n_312),
.B(n_321),
.C(n_318),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_535),
.B(n_214),
.Y(n_764)
);

BUFx6f_ASAP7_75t_SL g765 ( 
.A(n_520),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_603),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_545),
.B(n_447),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_491),
.B(n_451),
.Y(n_768)
);

NAND2xp33_ASAP7_75t_L g769 ( 
.A(n_543),
.B(n_232),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_545),
.B(n_451),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_491),
.B(n_451),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_550),
.B(n_587),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_508),
.B(n_451),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_563),
.B(n_451),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_537),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_597),
.B(n_614),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_550),
.B(n_224),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_543),
.A2(n_190),
.B1(n_184),
.B2(n_315),
.Y(n_778)
);

AOI22x1_ASAP7_75t_L g779 ( 
.A1(n_563),
.A2(n_463),
.B1(n_460),
.B2(n_459),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_543),
.B(n_294),
.Y(n_780)
);

INVxp67_ASAP7_75t_L g781 ( 
.A(n_509),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_508),
.B(n_184),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_543),
.A2(n_190),
.B1(n_315),
.B2(n_307),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_537),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_508),
.B(n_451),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_572),
.B(n_451),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_628),
.Y(n_787)
);

NOR2x2_ASAP7_75t_L g788 ( 
.A(n_760),
.B(n_272),
.Y(n_788)
);

A2O1A1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_629),
.A2(n_648),
.B(n_760),
.C(n_634),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_742),
.A2(n_745),
.B(n_744),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_629),
.B(n_543),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_746),
.B(n_572),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_748),
.A2(n_564),
.B(n_495),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_628),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_632),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_668),
.B(n_669),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_755),
.B(n_572),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_668),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_669),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_757),
.A2(n_759),
.B(n_704),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_648),
.B(n_573),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_723),
.B(n_573),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_632),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_767),
.A2(n_564),
.B(n_495),
.Y(n_804)
);

AOI21x1_ASAP7_75t_L g805 ( 
.A1(n_767),
.A2(n_547),
.B(n_546),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_770),
.A2(n_564),
.B(n_495),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_680),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_680),
.B(n_667),
.Y(n_808)
);

INVx1_ASAP7_75t_SL g809 ( 
.A(n_638),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_SL g810 ( 
.A(n_765),
.B(n_703),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_661),
.B(n_274),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_626),
.B(n_573),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_626),
.B(n_577),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_634),
.A2(n_599),
.B1(n_608),
.B2(n_314),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_770),
.A2(n_551),
.B(n_496),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_660),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_673),
.B(n_647),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_673),
.B(n_577),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_657),
.B(n_577),
.Y(n_819)
);

INVx5_ASAP7_75t_L g820 ( 
.A(n_668),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_721),
.B(n_274),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_765),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_665),
.B(n_580),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_774),
.A2(n_551),
.B(n_496),
.Y(n_824)
);

NOR3xp33_ASAP7_75t_L g825 ( 
.A(n_718),
.B(n_193),
.C(n_187),
.Y(n_825)
);

O2A1O1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_763),
.A2(n_585),
.B(n_509),
.C(n_605),
.Y(n_826)
);

NOR2xp67_ASAP7_75t_L g827 ( 
.A(n_650),
.B(n_432),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_672),
.B(n_281),
.Y(n_828)
);

A2O1A1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_645),
.A2(n_763),
.B(n_752),
.C(n_739),
.Y(n_829)
);

O2A1O1Ixp33_ASAP7_75t_L g830 ( 
.A1(n_739),
.A2(n_585),
.B(n_605),
.C(n_616),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_774),
.A2(n_551),
.B(n_496),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_631),
.A2(n_590),
.B(n_546),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_663),
.B(n_580),
.Y(n_833)
);

O2A1O1Ixp5_ASAP7_75t_L g834 ( 
.A1(n_776),
.A2(n_580),
.B(n_589),
.C(n_594),
.Y(n_834)
);

OR2x2_ASAP7_75t_L g835 ( 
.A(n_719),
.B(n_281),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_645),
.A2(n_603),
.B1(n_589),
.B2(n_594),
.Y(n_836)
);

NOR3xp33_ASAP7_75t_L g837 ( 
.A(n_718),
.B(n_187),
.C(n_193),
.Y(n_837)
);

OAI22xp5_ASAP7_75t_L g838 ( 
.A1(n_631),
.A2(n_772),
.B1(n_625),
.B2(n_624),
.Y(n_838)
);

NAND2x1p5_ASAP7_75t_L g839 ( 
.A(n_668),
.B(n_594),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_776),
.A2(n_582),
.B(n_547),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_687),
.B(n_553),
.Y(n_841)
);

INVx11_ASAP7_75t_L g842 ( 
.A(n_659),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_729),
.A2(n_623),
.B(n_620),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_636),
.A2(n_617),
.B(n_616),
.Y(n_844)
);

NAND2xp33_ASAP7_75t_L g845 ( 
.A(n_692),
.B(n_599),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_688),
.B(n_553),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_652),
.B(n_701),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_L g848 ( 
.A1(n_710),
.A2(n_675),
.B1(n_640),
.B2(n_633),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_689),
.B(n_710),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_690),
.B(n_554),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_676),
.B(n_293),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_679),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_686),
.A2(n_593),
.B(n_492),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_698),
.A2(n_593),
.B(n_492),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_702),
.A2(n_593),
.B(n_492),
.Y(n_855)
);

OAI321xp33_ASAP7_75t_L g856 ( 
.A1(n_670),
.A2(n_416),
.A3(n_441),
.B1(n_440),
.B2(n_431),
.C(n_428),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_693),
.B(n_554),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_653),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_695),
.B(n_555),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_653),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_679),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_685),
.Y(n_862)
);

OAI22xp33_ASAP7_75t_L g863 ( 
.A1(n_681),
.A2(n_297),
.B1(n_319),
.B2(n_316),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_685),
.Y(n_864)
);

INVx4_ASAP7_75t_L g865 ( 
.A(n_692),
.Y(n_865)
);

O2A1O1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_656),
.A2(n_617),
.B(n_613),
.C(n_610),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_762),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_642),
.Y(n_868)
);

NOR3xp33_ASAP7_75t_L g869 ( 
.A(n_749),
.B(n_301),
.C(n_307),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_630),
.A2(n_492),
.B(n_612),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_675),
.B(n_612),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_635),
.A2(n_612),
.B(n_613),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_639),
.A2(n_555),
.B(n_610),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_711),
.B(n_556),
.Y(n_874)
);

AO21x1_ASAP7_75t_L g875 ( 
.A1(n_733),
.A2(n_598),
.B(n_556),
.Y(n_875)
);

INVx1_ASAP7_75t_SL g876 ( 
.A(n_627),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_644),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_654),
.A2(n_612),
.B(n_607),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_734),
.B(n_559),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_722),
.B(n_559),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_728),
.B(n_565),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_664),
.A2(n_700),
.B(n_682),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_683),
.B(n_565),
.Y(n_883)
);

A2O1A1Ixp33_ASAP7_75t_L g884 ( 
.A1(n_752),
.A2(n_293),
.B(n_316),
.C(n_309),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_705),
.B(n_612),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_651),
.A2(n_599),
.B1(n_436),
.B2(n_602),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_682),
.A2(n_607),
.B(n_569),
.Y(n_887)
);

OAI21xp5_ASAP7_75t_L g888 ( 
.A1(n_671),
.A2(n_590),
.B(n_602),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_643),
.B(n_582),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_743),
.B(n_595),
.Y(n_890)
);

BUFx4f_ASAP7_75t_L g891 ( 
.A(n_644),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_691),
.B(n_595),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_761),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_637),
.B(n_641),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_761),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_735),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_637),
.B(n_505),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_700),
.A2(n_511),
.B(n_528),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_691),
.B(n_513),
.Y(n_899)
);

A2O1A1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_743),
.A2(n_296),
.B(n_319),
.C(n_309),
.Y(n_900)
);

AO21x1_ASAP7_75t_L g901 ( 
.A1(n_713),
.A2(n_400),
.B(n_418),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_781),
.A2(n_516),
.B(n_528),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_692),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_736),
.B(n_599),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_775),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_641),
.A2(n_435),
.B(n_422),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_696),
.B(n_603),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_769),
.A2(n_435),
.B(n_422),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_R g909 ( 
.A(n_740),
.B(n_301),
.Y(n_909)
);

INVx4_ASAP7_75t_L g910 ( 
.A(n_692),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_649),
.B(n_451),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_696),
.B(n_603),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_655),
.Y(n_913)
);

OR2x2_ASAP7_75t_SL g914 ( 
.A(n_726),
.B(n_296),
.Y(n_914)
);

A2O1A1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_708),
.A2(n_303),
.B(n_298),
.C(n_297),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_784),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_782),
.B(n_599),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_768),
.A2(n_449),
.B(n_463),
.Y(n_918)
);

INVx4_ASAP7_75t_L g919 ( 
.A(n_697),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_651),
.A2(n_599),
.B1(n_436),
.B2(n_303),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_649),
.B(n_677),
.Y(n_921)
);

INVx4_ASAP7_75t_L g922 ( 
.A(n_697),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_708),
.A2(n_298),
.B(n_233),
.C(n_236),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_706),
.A2(n_463),
.B(n_460),
.Y(n_924)
);

AO22x1_ASAP7_75t_L g925 ( 
.A1(n_730),
.A2(n_229),
.B1(n_250),
.B2(n_258),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_684),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_674),
.Y(n_927)
);

OAI22xp5_ASAP7_75t_L g928 ( 
.A1(n_658),
.A2(n_416),
.B1(n_265),
.B2(n_270),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_771),
.A2(n_463),
.B(n_460),
.Y(n_929)
);

O2A1O1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_656),
.A2(n_460),
.B(n_459),
.C(n_453),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_773),
.A2(n_459),
.B(n_453),
.Y(n_931)
);

INVx2_ASAP7_75t_SL g932 ( 
.A(n_762),
.Y(n_932)
);

AND2x2_ASAP7_75t_SL g933 ( 
.A(n_658),
.B(n_747),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_785),
.A2(n_459),
.B(n_453),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_694),
.A2(n_436),
.B1(n_448),
.B2(n_438),
.Y(n_935)
);

NOR2xp67_ASAP7_75t_SL g936 ( 
.A(n_751),
.B(n_449),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_786),
.A2(n_449),
.B(n_448),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_782),
.B(n_449),
.Y(n_938)
);

BUFx8_ASAP7_75t_L g939 ( 
.A(n_659),
.Y(n_939)
);

AO21x1_ASAP7_75t_L g940 ( 
.A1(n_717),
.A2(n_428),
.B(n_407),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_699),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_712),
.A2(n_716),
.B(n_727),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_756),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_732),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_714),
.A2(n_448),
.B(n_438),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_715),
.A2(n_438),
.B(n_435),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_737),
.A2(n_438),
.B(n_434),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_646),
.A2(n_434),
.B(n_425),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_662),
.A2(n_434),
.B(n_425),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_720),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_644),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_738),
.B(n_11),
.Y(n_952)
);

AOI22xp33_ASAP7_75t_L g953 ( 
.A1(n_709),
.A2(n_436),
.B1(n_431),
.B2(n_428),
.Y(n_953)
);

NAND2x1p5_ASAP7_75t_L g954 ( 
.A(n_751),
.B(n_400),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_725),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_697),
.B(n_418),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_731),
.A2(n_411),
.B(n_407),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_787),
.Y(n_958)
);

NAND2x1p5_ASAP7_75t_L g959 ( 
.A(n_820),
.B(n_707),
.Y(n_959)
);

XNOR2xp5_ASAP7_75t_L g960 ( 
.A(n_914),
.B(n_777),
.Y(n_960)
);

INVx3_ASAP7_75t_L g961 ( 
.A(n_798),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_852),
.Y(n_962)
);

O2A1O1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_789),
.A2(n_750),
.B(n_741),
.C(n_400),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_798),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_798),
.Y(n_965)
);

INVx4_ASAP7_75t_L g966 ( 
.A(n_798),
.Y(n_966)
);

OAI22xp5_ASAP7_75t_L g967 ( 
.A1(n_789),
.A2(n_707),
.B1(n_778),
.B2(n_783),
.Y(n_967)
);

OR2x6_ASAP7_75t_L g968 ( 
.A(n_877),
.B(n_666),
.Y(n_968)
);

BUFx2_ASAP7_75t_L g969 ( 
.A(n_858),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_865),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_787),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_817),
.B(n_764),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_860),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_829),
.A2(n_753),
.B(n_694),
.C(n_754),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_794),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_877),
.B(n_780),
.Y(n_976)
);

AOI21x1_ASAP7_75t_L g977 ( 
.A1(n_894),
.A2(n_741),
.B(n_780),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_794),
.Y(n_978)
);

HB1xp67_ASAP7_75t_L g979 ( 
.A(n_868),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_847),
.B(n_709),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_809),
.B(n_753),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_876),
.B(n_750),
.Y(n_982)
);

O2A1O1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_829),
.A2(n_407),
.B(n_411),
.C(n_766),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_803),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_790),
.A2(n_779),
.B(n_666),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_868),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_835),
.B(n_758),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_SL g988 ( 
.A1(n_952),
.A2(n_709),
.B1(n_758),
.B2(n_724),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_865),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_808),
.B(n_666),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_890),
.B(n_678),
.Y(n_991)
);

HB1xp67_ASAP7_75t_L g992 ( 
.A(n_852),
.Y(n_992)
);

INVx4_ASAP7_75t_L g993 ( 
.A(n_820),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_811),
.B(n_724),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_821),
.B(n_12),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_890),
.B(n_436),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_803),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_800),
.A2(n_436),
.B(n_155),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_917),
.A2(n_436),
.B(n_149),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_951),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_828),
.B(n_13),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_820),
.B(n_141),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_838),
.A2(n_436),
.B(n_18),
.C(n_24),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_861),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_879),
.B(n_15),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_933),
.B(n_140),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_938),
.A2(n_139),
.B(n_133),
.Y(n_1007)
);

BUFx2_ASAP7_75t_L g1008 ( 
.A(n_788),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_951),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_861),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_933),
.B(n_127),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_791),
.A2(n_102),
.B(n_120),
.Y(n_1012)
);

INVx1_ASAP7_75t_SL g1013 ( 
.A(n_851),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_879),
.B(n_27),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_848),
.A2(n_124),
.B(n_111),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_818),
.A2(n_108),
.B(n_107),
.Y(n_1016)
);

AOI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_952),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_827),
.B(n_31),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_807),
.A2(n_912),
.B1(n_907),
.B2(n_849),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_807),
.A2(n_105),
.B1(n_101),
.B2(n_97),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_893),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_867),
.B(n_91),
.Y(n_1022)
);

INVx4_ASAP7_75t_L g1023 ( 
.A(n_910),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_795),
.Y(n_1024)
);

O2A1O1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_923),
.A2(n_34),
.B(n_35),
.C(n_38),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_825),
.B(n_86),
.Y(n_1026)
);

INVxp67_ASAP7_75t_L g1027 ( 
.A(n_802),
.Y(n_1027)
);

BUFx4f_ASAP7_75t_L g1028 ( 
.A(n_932),
.Y(n_1028)
);

OAI21xp33_ASAP7_75t_SL g1029 ( 
.A1(n_814),
.A2(n_34),
.B(n_42),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_907),
.A2(n_82),
.B1(n_76),
.B2(n_44),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_895),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_912),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_837),
.B(n_43),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_891),
.Y(n_1034)
);

BUFx10_ASAP7_75t_L g1035 ( 
.A(n_822),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_801),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_944),
.B(n_46),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_SL g1038 ( 
.A1(n_814),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_926),
.B(n_896),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_823),
.B(n_51),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_823),
.B(n_799),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_871),
.A2(n_921),
.B(n_793),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_799),
.B(n_816),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_842),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_871),
.A2(n_921),
.B(n_806),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_804),
.A2(n_52),
.B(n_54),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_923),
.B(n_55),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_891),
.Y(n_1048)
);

OAI21xp33_ASAP7_75t_L g1049 ( 
.A1(n_915),
.A2(n_57),
.B(n_58),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_900),
.A2(n_57),
.B(n_60),
.C(n_61),
.Y(n_1050)
);

A2O1A1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_882),
.A2(n_61),
.B(n_915),
.C(n_884),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_853),
.A2(n_843),
.B(n_854),
.Y(n_1052)
);

AO32x2_ASAP7_75t_L g1053 ( 
.A1(n_836),
.A2(n_928),
.A3(n_919),
.B1(n_922),
.B2(n_910),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_919),
.Y(n_1054)
);

AO22x1_ASAP7_75t_L g1055 ( 
.A1(n_869),
.A2(n_939),
.B1(n_905),
.B2(n_916),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_895),
.Y(n_1056)
);

INVx2_ASAP7_75t_SL g1057 ( 
.A(n_909),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_900),
.A2(n_884),
.B(n_889),
.C(n_892),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_810),
.B(n_899),
.Y(n_1059)
);

CKINVDCx11_ASAP7_75t_R g1060 ( 
.A(n_939),
.Y(n_1060)
);

INVx5_ASAP7_75t_L g1061 ( 
.A(n_903),
.Y(n_1061)
);

NAND2x1p5_ASAP7_75t_L g1062 ( 
.A(n_903),
.B(n_796),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_925),
.B(n_909),
.Y(n_1063)
);

BUFx3_ASAP7_75t_L g1064 ( 
.A(n_927),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_950),
.A2(n_955),
.B(n_864),
.C(n_862),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_941),
.B(n_913),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_792),
.B(n_797),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_863),
.B(n_856),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_855),
.A2(n_840),
.B(n_942),
.Y(n_1069)
);

OAI22x1_ASAP7_75t_L g1070 ( 
.A1(n_863),
.A2(n_894),
.B1(n_954),
.B2(n_935),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_841),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_846),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_839),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_834),
.A2(n_832),
.B(n_887),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_812),
.A2(n_813),
.B1(n_954),
.B2(n_883),
.Y(n_1075)
);

NAND3xp33_ASAP7_75t_L g1076 ( 
.A(n_920),
.B(n_953),
.C(n_886),
.Y(n_1076)
);

O2A1O1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_850),
.A2(n_881),
.B(n_874),
.C(n_857),
.Y(n_1077)
);

AOI21x1_ASAP7_75t_L g1078 ( 
.A1(n_897),
.A2(n_805),
.B(n_885),
.Y(n_1078)
);

OAI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_859),
.A2(n_880),
.B1(n_943),
.B2(n_819),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_833),
.B(n_953),
.Y(n_1080)
);

INVx4_ASAP7_75t_L g1081 ( 
.A(n_839),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_911),
.A2(n_924),
.B(n_946),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_920),
.Y(n_1083)
);

NAND2xp33_ASAP7_75t_L g1084 ( 
.A(n_904),
.B(n_886),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_911),
.A2(n_815),
.B(n_824),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_956),
.B(n_875),
.Y(n_1086)
);

BUFx10_ASAP7_75t_L g1087 ( 
.A(n_940),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_902),
.B(n_844),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_SL g1089 ( 
.A1(n_898),
.A2(n_873),
.B1(n_888),
.B2(n_826),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_901),
.Y(n_1090)
);

AOI221xp5_ASAP7_75t_L g1091 ( 
.A1(n_830),
.A2(n_866),
.B1(n_930),
.B2(n_957),
.C(n_885),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_897),
.Y(n_1092)
);

OR2x6_ASAP7_75t_SL g1093 ( 
.A(n_845),
.B(n_936),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_947),
.Y(n_1094)
);

OR2x6_ASAP7_75t_L g1095 ( 
.A(n_831),
.B(n_870),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_906),
.A2(n_872),
.B(n_878),
.C(n_929),
.Y(n_1096)
);

AND2x2_ASAP7_75t_SL g1097 ( 
.A(n_948),
.B(n_949),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1069),
.A2(n_908),
.B(n_918),
.Y(n_1098)
);

OAI22x1_ASAP7_75t_L g1099 ( 
.A1(n_1047),
.A2(n_931),
.B1(n_934),
.B2(n_937),
.Y(n_1099)
);

AO31x2_ASAP7_75t_L g1100 ( 
.A1(n_1042),
.A2(n_1069),
.A3(n_1045),
.B(n_1052),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_974),
.A2(n_945),
.B(n_972),
.C(n_995),
.Y(n_1101)
);

OA21x2_ASAP7_75t_L g1102 ( 
.A1(n_1074),
.A2(n_1042),
.B(n_1045),
.Y(n_1102)
);

AO31x2_ASAP7_75t_L g1103 ( 
.A1(n_1052),
.A2(n_1096),
.A3(n_1085),
.B(n_1082),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1024),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_991),
.B(n_1071),
.Y(n_1105)
);

NAND3x1_ASAP7_75t_L g1106 ( 
.A(n_1063),
.B(n_994),
.C(n_987),
.Y(n_1106)
);

AO21x1_ASAP7_75t_L g1107 ( 
.A1(n_1015),
.A2(n_1003),
.B(n_1046),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_1034),
.Y(n_1108)
);

BUFx12f_ASAP7_75t_L g1109 ( 
.A(n_1060),
.Y(n_1109)
);

OR2x2_ASAP7_75t_L g1110 ( 
.A(n_1013),
.B(n_986),
.Y(n_1110)
);

AO31x2_ASAP7_75t_L g1111 ( 
.A1(n_1085),
.A2(n_1082),
.A3(n_985),
.B(n_1019),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_979),
.Y(n_1112)
);

O2A1O1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_1033),
.A2(n_1032),
.B(n_1051),
.C(n_1068),
.Y(n_1113)
);

NAND3xp33_ASAP7_75t_L g1114 ( 
.A(n_1017),
.B(n_981),
.C(n_1025),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1097),
.A2(n_985),
.B(n_1089),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1058),
.A2(n_996),
.B(n_967),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_982),
.B(n_1064),
.Y(n_1117)
);

OAI22x1_ASAP7_75t_L g1118 ( 
.A1(n_1006),
.A2(n_1011),
.B1(n_1008),
.B2(n_1083),
.Y(n_1118)
);

AOI221xp5_ASAP7_75t_SL g1119 ( 
.A1(n_1017),
.A2(n_1049),
.B1(n_1003),
.B2(n_1025),
.C(n_1038),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_SL g1120 ( 
.A1(n_1026),
.A2(n_1002),
.B(n_1065),
.C(n_980),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_1034),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_1027),
.B(n_1059),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_1027),
.B(n_979),
.Y(n_1123)
);

INVx3_ASAP7_75t_SL g1124 ( 
.A(n_1044),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_1050),
.A2(n_1036),
.B(n_1014),
.C(n_1005),
.Y(n_1125)
);

A2O1A1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_1058),
.A2(n_1018),
.B(n_1015),
.C(n_963),
.Y(n_1126)
);

NAND3xp33_ASAP7_75t_L g1127 ( 
.A(n_1050),
.B(n_988),
.C(n_1046),
.Y(n_1127)
);

INVx4_ASAP7_75t_L g1128 ( 
.A(n_965),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_1037),
.A2(n_1040),
.B(n_1030),
.C(n_1029),
.Y(n_1129)
);

BUFx12f_ASAP7_75t_L g1130 ( 
.A(n_1035),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_SL g1131 ( 
.A1(n_1080),
.A2(n_1086),
.B(n_990),
.C(n_1041),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_SL g1132 ( 
.A(n_1035),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1066),
.Y(n_1133)
);

OAI22xp33_ASAP7_75t_L g1134 ( 
.A1(n_1057),
.A2(n_1039),
.B1(n_1028),
.B2(n_1072),
.Y(n_1134)
);

A2O1A1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_963),
.A2(n_1077),
.B(n_1090),
.C(n_1076),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_1034),
.Y(n_1136)
);

AO31x2_ASAP7_75t_L g1137 ( 
.A1(n_998),
.A2(n_1088),
.A3(n_1075),
.B(n_1070),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_960),
.B(n_969),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1097),
.A2(n_1077),
.B(n_1067),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_958),
.Y(n_1140)
);

BUFx12f_ASAP7_75t_L g1141 ( 
.A(n_1048),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_988),
.A2(n_1022),
.B1(n_1001),
.B2(n_976),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_977),
.A2(n_998),
.B(n_1094),
.Y(n_1143)
);

BUFx2_ASAP7_75t_L g1144 ( 
.A(n_973),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1022),
.B(n_976),
.Y(n_1145)
);

AO31x2_ASAP7_75t_L g1146 ( 
.A1(n_999),
.A2(n_1012),
.A3(n_1007),
.B(n_1016),
.Y(n_1146)
);

INVx2_ASAP7_75t_SL g1147 ( 
.A(n_1028),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_983),
.A2(n_999),
.B(n_1062),
.Y(n_1148)
);

INVx3_ASAP7_75t_L g1149 ( 
.A(n_993),
.Y(n_1149)
);

INVx2_ASAP7_75t_SL g1150 ( 
.A(n_1000),
.Y(n_1150)
);

NAND3x1_ASAP7_75t_L g1151 ( 
.A(n_961),
.B(n_964),
.C(n_1055),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_971),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_975),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1084),
.A2(n_1079),
.B(n_1043),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1062),
.A2(n_1091),
.B(n_1092),
.Y(n_1155)
);

BUFx10_ASAP7_75t_L g1156 ( 
.A(n_1048),
.Y(n_1156)
);

AO31x2_ASAP7_75t_L g1157 ( 
.A1(n_1012),
.A2(n_1007),
.A3(n_1016),
.B(n_1010),
.Y(n_1157)
);

AO31x2_ASAP7_75t_L g1158 ( 
.A1(n_978),
.A2(n_997),
.A3(n_984),
.B(n_1004),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_992),
.A2(n_1093),
.B1(n_959),
.B2(n_968),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1021),
.A2(n_1056),
.B(n_1031),
.Y(n_1160)
);

A2O1A1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_962),
.A2(n_1073),
.B(n_1020),
.C(n_970),
.Y(n_1161)
);

OA21x2_ASAP7_75t_L g1162 ( 
.A1(n_1087),
.A2(n_1095),
.B(n_1053),
.Y(n_1162)
);

HB1xp67_ASAP7_75t_SL g1163 ( 
.A(n_1048),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1095),
.A2(n_1073),
.B(n_1081),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_993),
.A2(n_989),
.B(n_1054),
.Y(n_1165)
);

INVx3_ASAP7_75t_L g1166 ( 
.A(n_1081),
.Y(n_1166)
);

BUFx2_ASAP7_75t_L g1167 ( 
.A(n_1009),
.Y(n_1167)
);

CKINVDCx14_ASAP7_75t_R g1168 ( 
.A(n_1009),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1054),
.A2(n_1061),
.B(n_959),
.Y(n_1169)
);

AO32x2_ASAP7_75t_L g1170 ( 
.A1(n_1087),
.A2(n_966),
.A3(n_1023),
.B1(n_1053),
.B2(n_1061),
.Y(n_1170)
);

INVx3_ASAP7_75t_L g1171 ( 
.A(n_1023),
.Y(n_1171)
);

OA21x2_ASAP7_75t_L g1172 ( 
.A1(n_1053),
.A2(n_1061),
.B(n_964),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_SL g1173 ( 
.A(n_1009),
.Y(n_1173)
);

OR2x2_ASAP7_75t_L g1174 ( 
.A(n_968),
.B(n_961),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_966),
.B(n_965),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_965),
.B(n_1061),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_968),
.B(n_1053),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_SL g1178 ( 
.A(n_1044),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1024),
.Y(n_1179)
);

AO31x2_ASAP7_75t_L g1180 ( 
.A1(n_1042),
.A2(n_875),
.A3(n_1069),
.B(n_1045),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1069),
.A2(n_1097),
.B(n_790),
.Y(n_1181)
);

AO31x2_ASAP7_75t_L g1182 ( 
.A1(n_1042),
.A2(n_875),
.A3(n_1069),
.B(n_1045),
.Y(n_1182)
);

AOI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_981),
.A2(n_629),
.B1(n_648),
.B2(n_324),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1069),
.A2(n_1097),
.B(n_790),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1069),
.A2(n_1097),
.B(n_790),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_991),
.A2(n_629),
.B(n_789),
.C(n_648),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1069),
.A2(n_1097),
.B(n_790),
.Y(n_1187)
);

CKINVDCx16_ASAP7_75t_R g1188 ( 
.A(n_1035),
.Y(n_1188)
);

O2A1O1Ixp33_ASAP7_75t_SL g1189 ( 
.A1(n_1006),
.A2(n_789),
.B(n_829),
.C(n_1011),
.Y(n_1189)
);

AO31x2_ASAP7_75t_L g1190 ( 
.A1(n_1042),
.A2(n_875),
.A3(n_1069),
.B(n_1045),
.Y(n_1190)
);

OAI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_972),
.A2(n_789),
.B(n_629),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1024),
.Y(n_1192)
);

AND2x6_ASAP7_75t_L g1193 ( 
.A(n_1090),
.B(n_965),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_972),
.B(n_629),
.Y(n_1194)
);

AOI21x1_ASAP7_75t_L g1195 ( 
.A1(n_985),
.A2(n_1082),
.B(n_1042),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1052),
.A2(n_1085),
.B(n_1078),
.Y(n_1196)
);

AOI21x1_ASAP7_75t_L g1197 ( 
.A1(n_985),
.A2(n_1082),
.B(n_1042),
.Y(n_1197)
);

AOI221x1_ASAP7_75t_L g1198 ( 
.A1(n_1015),
.A2(n_789),
.B1(n_629),
.B2(n_1049),
.C(n_1046),
.Y(n_1198)
);

BUFx12f_ASAP7_75t_L g1199 ( 
.A(n_1060),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1024),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_972),
.B(n_629),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_SL g1202 ( 
.A1(n_1083),
.A2(n_519),
.B1(n_648),
.B2(n_629),
.Y(n_1202)
);

INVx6_ASAP7_75t_SL g1203 ( 
.A(n_1035),
.Y(n_1203)
);

A2O1A1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_974),
.A2(n_629),
.B(n_789),
.C(n_648),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1069),
.A2(n_1097),
.B(n_790),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1069),
.A2(n_1097),
.B(n_790),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1069),
.A2(n_1097),
.B(n_790),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_972),
.B(n_629),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1013),
.B(n_821),
.Y(n_1209)
);

AO31x2_ASAP7_75t_L g1210 ( 
.A1(n_1042),
.A2(n_875),
.A3(n_1069),
.B(n_1045),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_SL g1211 ( 
.A1(n_974),
.A2(n_789),
.B(n_668),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1069),
.A2(n_1097),
.B(n_790),
.Y(n_1212)
);

INVx6_ASAP7_75t_SL g1213 ( 
.A(n_1035),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_974),
.A2(n_629),
.B(n_789),
.C(n_648),
.Y(n_1214)
);

OA21x2_ASAP7_75t_L g1215 ( 
.A1(n_1074),
.A2(n_1042),
.B(n_1045),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_986),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1069),
.A2(n_1097),
.B(n_790),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_991),
.B(n_661),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1083),
.A2(n_629),
.B1(n_648),
.B2(n_952),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_974),
.A2(n_629),
.B(n_789),
.C(n_648),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1069),
.A2(n_1097),
.B(n_790),
.Y(n_1221)
);

OA21x2_ASAP7_75t_L g1222 ( 
.A1(n_1074),
.A2(n_1042),
.B(n_1045),
.Y(n_1222)
);

AO31x2_ASAP7_75t_L g1223 ( 
.A1(n_1042),
.A2(n_875),
.A3(n_1069),
.B(n_1045),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_972),
.A2(n_789),
.B(n_629),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_972),
.B(n_719),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1069),
.A2(n_1097),
.B(n_790),
.Y(n_1226)
);

A2O1A1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_974),
.A2(n_629),
.B(n_789),
.C(n_648),
.Y(n_1227)
);

AO32x2_ASAP7_75t_L g1228 ( 
.A1(n_1089),
.A2(n_1038),
.A3(n_1036),
.B1(n_967),
.B2(n_848),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1052),
.A2(n_1085),
.B(n_1078),
.Y(n_1229)
);

AO21x1_ASAP7_75t_L g1230 ( 
.A1(n_1015),
.A2(n_629),
.B(n_1003),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_991),
.B(n_661),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_972),
.B(n_629),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1083),
.A2(n_629),
.B1(n_789),
.B2(n_991),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_972),
.B(n_629),
.Y(n_1234)
);

NAND2x1_ASAP7_75t_L g1235 ( 
.A(n_993),
.B(n_798),
.Y(n_1235)
);

INVxp67_ASAP7_75t_L g1236 ( 
.A(n_986),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1052),
.A2(n_1085),
.B(n_1078),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_991),
.B(n_661),
.Y(n_1238)
);

BUFx3_ASAP7_75t_L g1239 ( 
.A(n_1000),
.Y(n_1239)
);

A2O1A1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_974),
.A2(n_629),
.B(n_789),
.C(n_648),
.Y(n_1240)
);

OAI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1083),
.A2(n_519),
.B1(n_629),
.B2(n_650),
.Y(n_1241)
);

A2O1A1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_974),
.A2(n_629),
.B(n_789),
.C(n_648),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_972),
.B(n_629),
.Y(n_1243)
);

AOI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1219),
.A2(n_1183),
.B1(n_1202),
.B2(n_1241),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_1178),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1114),
.A2(n_1233),
.B1(n_1191),
.B2(n_1224),
.Y(n_1246)
);

INVx6_ASAP7_75t_L g1247 ( 
.A(n_1156),
.Y(n_1247)
);

CKINVDCx14_ASAP7_75t_R g1248 ( 
.A(n_1168),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1194),
.B(n_1201),
.Y(n_1249)
);

BUFx12f_ASAP7_75t_L g1250 ( 
.A(n_1109),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_SL g1251 ( 
.A1(n_1208),
.A2(n_1243),
.B1(n_1232),
.B2(n_1234),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1127),
.A2(n_1230),
.B1(n_1225),
.B2(n_1118),
.Y(n_1252)
);

INVx6_ASAP7_75t_L g1253 ( 
.A(n_1156),
.Y(n_1253)
);

INVx5_ASAP7_75t_L g1254 ( 
.A(n_1193),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1104),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_1124),
.Y(n_1256)
);

BUFx2_ASAP7_75t_R g1257 ( 
.A(n_1239),
.Y(n_1257)
);

OAI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1105),
.A2(n_1142),
.B1(n_1198),
.B2(n_1133),
.Y(n_1258)
);

CKINVDCx6p67_ASAP7_75t_R g1259 ( 
.A(n_1199),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1108),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1218),
.A2(n_1231),
.B1(n_1238),
.B2(n_1122),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1179),
.Y(n_1262)
);

CKINVDCx11_ASAP7_75t_R g1263 ( 
.A(n_1130),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1204),
.A2(n_1242),
.B1(n_1240),
.B2(n_1227),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1192),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_SL g1266 ( 
.A(n_1108),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1107),
.A2(n_1116),
.B1(n_1115),
.B2(n_1134),
.Y(n_1267)
);

INVx3_ASAP7_75t_L g1268 ( 
.A(n_1166),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1200),
.Y(n_1269)
);

BUFx10_ASAP7_75t_L g1270 ( 
.A(n_1173),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1209),
.B(n_1145),
.Y(n_1271)
);

BUFx12f_ASAP7_75t_L g1272 ( 
.A(n_1141),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_1167),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_SL g1274 ( 
.A1(n_1119),
.A2(n_1117),
.B1(n_1162),
.B2(n_1139),
.Y(n_1274)
);

CKINVDCx11_ASAP7_75t_R g1275 ( 
.A(n_1188),
.Y(n_1275)
);

OAI21xp33_ASAP7_75t_L g1276 ( 
.A1(n_1214),
.A2(n_1220),
.B(n_1186),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1123),
.B(n_1216),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1154),
.A2(n_1112),
.B1(n_1138),
.B2(n_1152),
.Y(n_1278)
);

BUFx2_ASAP7_75t_L g1279 ( 
.A(n_1144),
.Y(n_1279)
);

CKINVDCx16_ASAP7_75t_R g1280 ( 
.A(n_1163),
.Y(n_1280)
);

CKINVDCx11_ASAP7_75t_R g1281 ( 
.A(n_1108),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1236),
.A2(n_1135),
.B1(n_1126),
.B2(n_1106),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1140),
.A2(n_1153),
.B1(n_1187),
.B2(n_1212),
.Y(n_1283)
);

BUFx8_ASAP7_75t_L g1284 ( 
.A(n_1132),
.Y(n_1284)
);

BUFx12f_ASAP7_75t_L g1285 ( 
.A(n_1121),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_1155),
.Y(n_1286)
);

BUFx3_ASAP7_75t_L g1287 ( 
.A(n_1121),
.Y(n_1287)
);

OAI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1159),
.A2(n_1177),
.B1(n_1174),
.B2(n_1147),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1113),
.B(n_1101),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1211),
.A2(n_1125),
.B1(n_1151),
.B2(n_1129),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1181),
.A2(n_1205),
.B1(n_1185),
.B2(n_1207),
.Y(n_1291)
);

BUFx12f_ASAP7_75t_L g1292 ( 
.A(n_1136),
.Y(n_1292)
);

BUFx2_ASAP7_75t_L g1293 ( 
.A(n_1150),
.Y(n_1293)
);

INVx3_ASAP7_75t_SL g1294 ( 
.A(n_1136),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_1203),
.Y(n_1295)
);

OAI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1228),
.A2(n_1206),
.B1(n_1217),
.B2(n_1221),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1158),
.Y(n_1297)
);

INVx6_ASAP7_75t_L g1298 ( 
.A(n_1136),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1172),
.Y(n_1299)
);

BUFx12f_ASAP7_75t_L g1300 ( 
.A(n_1128),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1193),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1160),
.Y(n_1302)
);

CKINVDCx14_ASAP7_75t_R g1303 ( 
.A(n_1193),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_SL g1304 ( 
.A1(n_1164),
.A2(n_1175),
.B1(n_1176),
.B2(n_1128),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1193),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1235),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1184),
.A2(n_1226),
.B1(n_1215),
.B2(n_1102),
.Y(n_1307)
);

INVx4_ASAP7_75t_L g1308 ( 
.A(n_1171),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1102),
.A2(n_1222),
.B1(n_1215),
.B2(n_1228),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_SL g1310 ( 
.A1(n_1228),
.A2(n_1189),
.B(n_1161),
.Y(n_1310)
);

AOI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1120),
.A2(n_1131),
.B1(n_1171),
.B2(n_1149),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1203),
.A2(n_1213),
.B1(n_1162),
.B2(n_1169),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1213),
.A2(n_1172),
.B1(n_1165),
.B2(n_1222),
.Y(n_1313)
);

OAI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1099),
.A2(n_1197),
.B1(n_1195),
.B2(n_1170),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1098),
.A2(n_1170),
.B1(n_1148),
.B2(n_1146),
.Y(n_1315)
);

BUFx12f_ASAP7_75t_L g1316 ( 
.A(n_1157),
.Y(n_1316)
);

CKINVDCx6p67_ASAP7_75t_R g1317 ( 
.A(n_1157),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1143),
.A2(n_1237),
.B1(n_1229),
.B2(n_1196),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1157),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1170),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1137),
.A2(n_1111),
.B1(n_1223),
.B2(n_1182),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1100),
.B(n_1182),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1137),
.A2(n_1111),
.B1(n_1180),
.B2(n_1182),
.Y(n_1323)
);

INVx4_ASAP7_75t_L g1324 ( 
.A(n_1103),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1190),
.A2(n_1210),
.B1(n_1223),
.B2(n_1103),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1190),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1210),
.A2(n_1219),
.B1(n_1202),
.B2(n_1114),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1223),
.A2(n_1219),
.B1(n_1183),
.B2(n_629),
.Y(n_1328)
);

OAI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1183),
.A2(n_1114),
.B1(n_1083),
.B2(n_1241),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_SL g1330 ( 
.A1(n_1202),
.A2(n_1219),
.B1(n_1183),
.B2(n_519),
.Y(n_1330)
);

CKINVDCx11_ASAP7_75t_R g1331 ( 
.A(n_1109),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1219),
.A2(n_1183),
.B1(n_629),
.B2(n_1202),
.Y(n_1332)
);

NAND2x1p5_ASAP7_75t_L g1333 ( 
.A(n_1166),
.B(n_820),
.Y(n_1333)
);

BUFx10_ASAP7_75t_L g1334 ( 
.A(n_1173),
.Y(n_1334)
);

BUFx8_ASAP7_75t_L g1335 ( 
.A(n_1173),
.Y(n_1335)
);

CKINVDCx11_ASAP7_75t_R g1336 ( 
.A(n_1109),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1219),
.A2(n_1202),
.B1(n_1114),
.B2(n_1017),
.Y(n_1337)
);

BUFx10_ASAP7_75t_L g1338 ( 
.A(n_1173),
.Y(n_1338)
);

BUFx12f_ASAP7_75t_L g1339 ( 
.A(n_1109),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1219),
.A2(n_1202),
.B1(n_1114),
.B2(n_1017),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1219),
.A2(n_629),
.B(n_648),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_SL g1342 ( 
.A1(n_1114),
.A2(n_1038),
.B1(n_519),
.B2(n_1083),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1194),
.B(n_1201),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_1108),
.Y(n_1344)
);

CKINVDCx11_ASAP7_75t_R g1345 ( 
.A(n_1109),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_L g1346 ( 
.A(n_1108),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1178),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1219),
.A2(n_1202),
.B1(n_1114),
.B2(n_1017),
.Y(n_1348)
);

BUFx8_ASAP7_75t_L g1349 ( 
.A(n_1173),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1219),
.A2(n_1202),
.B1(n_1114),
.B2(n_1017),
.Y(n_1350)
);

CKINVDCx20_ASAP7_75t_R g1351 ( 
.A(n_1124),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1104),
.Y(n_1352)
);

BUFx4f_ASAP7_75t_SL g1353 ( 
.A(n_1203),
.Y(n_1353)
);

CKINVDCx20_ASAP7_75t_R g1354 ( 
.A(n_1124),
.Y(n_1354)
);

BUFx2_ASAP7_75t_L g1355 ( 
.A(n_1216),
.Y(n_1355)
);

BUFx6f_ASAP7_75t_L g1356 ( 
.A(n_1108),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1219),
.A2(n_629),
.B1(n_1183),
.B2(n_1202),
.Y(n_1357)
);

INVx3_ASAP7_75t_L g1358 ( 
.A(n_1166),
.Y(n_1358)
);

BUFx12f_ASAP7_75t_L g1359 ( 
.A(n_1109),
.Y(n_1359)
);

INVx2_ASAP7_75t_SL g1360 ( 
.A(n_1239),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1219),
.A2(n_1183),
.B1(n_629),
.B2(n_1202),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_1216),
.Y(n_1362)
);

INVx1_ASAP7_75t_SL g1363 ( 
.A(n_1110),
.Y(n_1363)
);

OAI21xp5_ASAP7_75t_SL g1364 ( 
.A1(n_1183),
.A2(n_1219),
.B(n_1202),
.Y(n_1364)
);

INVx1_ASAP7_75t_SL g1365 ( 
.A(n_1110),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1251),
.B(n_1274),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1246),
.B(n_1327),
.Y(n_1367)
);

INVxp67_ASAP7_75t_L g1368 ( 
.A(n_1255),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_1254),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1297),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1251),
.B(n_1246),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1342),
.A2(n_1337),
.B1(n_1340),
.B2(n_1348),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1326),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1277),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1315),
.A2(n_1291),
.B(n_1318),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1322),
.B(n_1319),
.Y(n_1376)
);

OAI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1341),
.A2(n_1328),
.B(n_1332),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1299),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1361),
.A2(n_1330),
.B1(n_1337),
.B2(n_1350),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1327),
.B(n_1325),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1299),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1325),
.B(n_1321),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1316),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1324),
.B(n_1302),
.Y(n_1384)
);

INVx4_ASAP7_75t_L g1385 ( 
.A(n_1301),
.Y(n_1385)
);

BUFx2_ASAP7_75t_L g1386 ( 
.A(n_1286),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1286),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1320),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1291),
.A2(n_1318),
.B(n_1307),
.Y(n_1389)
);

INVxp67_ASAP7_75t_L g1390 ( 
.A(n_1262),
.Y(n_1390)
);

OA21x2_ASAP7_75t_L g1391 ( 
.A1(n_1267),
.A2(n_1321),
.B(n_1323),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1252),
.B(n_1249),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1363),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1261),
.B(n_1365),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1355),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1265),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1317),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1269),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1323),
.B(n_1309),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1352),
.Y(n_1400)
);

INVx1_ASAP7_75t_SL g1401 ( 
.A(n_1362),
.Y(n_1401)
);

AO21x2_ASAP7_75t_L g1402 ( 
.A1(n_1314),
.A2(n_1296),
.B(n_1276),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1314),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1309),
.B(n_1252),
.Y(n_1404)
);

AOI21xp33_ASAP7_75t_L g1405 ( 
.A1(n_1329),
.A2(n_1340),
.B(n_1350),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1313),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1289),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1307),
.A2(n_1283),
.B(n_1264),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1305),
.B(n_1283),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1343),
.B(n_1258),
.Y(n_1410)
);

BUFx6f_ASAP7_75t_L g1411 ( 
.A(n_1301),
.Y(n_1411)
);

CKINVDCx20_ASAP7_75t_R g1412 ( 
.A(n_1256),
.Y(n_1412)
);

BUFx6f_ASAP7_75t_L g1413 ( 
.A(n_1301),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1310),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1296),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1311),
.Y(n_1416)
);

OAI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1357),
.A2(n_1244),
.B1(n_1364),
.B2(n_1329),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1290),
.A2(n_1312),
.B(n_1282),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1271),
.B(n_1278),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1304),
.Y(n_1420)
);

BUFx3_ASAP7_75t_L g1421 ( 
.A(n_1273),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1279),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1278),
.A2(n_1358),
.B(n_1268),
.Y(n_1423)
);

INVxp33_ASAP7_75t_L g1424 ( 
.A(n_1293),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1258),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1288),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1288),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1273),
.Y(n_1428)
);

INVx1_ASAP7_75t_SL g1429 ( 
.A(n_1294),
.Y(n_1429)
);

INVxp67_ASAP7_75t_SL g1430 ( 
.A(n_1348),
.Y(n_1430)
);

BUFx4f_ASAP7_75t_L g1431 ( 
.A(n_1333),
.Y(n_1431)
);

BUFx2_ASAP7_75t_L g1432 ( 
.A(n_1303),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1303),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1342),
.B(n_1344),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1308),
.B(n_1306),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1260),
.Y(n_1436)
);

AO21x2_ASAP7_75t_L g1437 ( 
.A1(n_1266),
.A2(n_1294),
.B(n_1344),
.Y(n_1437)
);

INVx3_ASAP7_75t_L g1438 ( 
.A(n_1260),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1260),
.Y(n_1439)
);

INVx4_ASAP7_75t_SL g1440 ( 
.A(n_1298),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1298),
.A2(n_1300),
.B(n_1292),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1399),
.B(n_1280),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1399),
.B(n_1346),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1370),
.Y(n_1444)
);

AND2x2_ASAP7_75t_SL g1445 ( 
.A(n_1391),
.B(n_1356),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_SL g1446 ( 
.A1(n_1377),
.A2(n_1372),
.B(n_1420),
.Y(n_1446)
);

AO32x1_ASAP7_75t_L g1447 ( 
.A1(n_1372),
.A2(n_1360),
.A3(n_1275),
.B1(n_1257),
.B2(n_1281),
.Y(n_1447)
);

OA21x2_ASAP7_75t_L g1448 ( 
.A1(n_1375),
.A2(n_1245),
.B(n_1347),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1403),
.B(n_1380),
.Y(n_1449)
);

AND2x2_ASAP7_75t_SL g1450 ( 
.A(n_1391),
.B(n_1248),
.Y(n_1450)
);

AOI221xp5_ASAP7_75t_L g1451 ( 
.A1(n_1417),
.A2(n_1248),
.B1(n_1295),
.B2(n_1287),
.C(n_1354),
.Y(n_1451)
);

INVxp67_ASAP7_75t_L g1452 ( 
.A(n_1374),
.Y(n_1452)
);

OA21x2_ASAP7_75t_L g1453 ( 
.A1(n_1375),
.A2(n_1285),
.B(n_1247),
.Y(n_1453)
);

AND2x4_ASAP7_75t_SL g1454 ( 
.A(n_1393),
.B(n_1351),
.Y(n_1454)
);

A2O1A1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1377),
.A2(n_1405),
.B(n_1379),
.C(n_1420),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1403),
.B(n_1334),
.Y(n_1456)
);

OR2x6_ASAP7_75t_L g1457 ( 
.A(n_1408),
.B(n_1272),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1386),
.Y(n_1458)
);

OAI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1405),
.A2(n_1284),
.B(n_1247),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1394),
.B(n_1259),
.Y(n_1460)
);

BUFx2_ASAP7_75t_L g1461 ( 
.A(n_1386),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1420),
.A2(n_1247),
.B1(n_1253),
.B2(n_1353),
.Y(n_1462)
);

INVx3_ASAP7_75t_L g1463 ( 
.A(n_1384),
.Y(n_1463)
);

NAND4xp25_ASAP7_75t_SL g1464 ( 
.A(n_1371),
.B(n_1335),
.C(n_1349),
.D(n_1284),
.Y(n_1464)
);

OAI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1430),
.A2(n_1253),
.B(n_1263),
.Y(n_1465)
);

AOI221xp5_ASAP7_75t_L g1466 ( 
.A1(n_1430),
.A2(n_1270),
.B1(n_1338),
.B2(n_1334),
.C(n_1349),
.Y(n_1466)
);

OAI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1371),
.A2(n_1253),
.B(n_1270),
.Y(n_1467)
);

AO21x2_ASAP7_75t_L g1468 ( 
.A1(n_1389),
.A2(n_1338),
.B(n_1335),
.Y(n_1468)
);

OA21x2_ASAP7_75t_L g1469 ( 
.A1(n_1375),
.A2(n_1353),
.B(n_1336),
.Y(n_1469)
);

OR2x6_ASAP7_75t_L g1470 ( 
.A(n_1408),
.B(n_1250),
.Y(n_1470)
);

OAI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1418),
.A2(n_1336),
.B(n_1345),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1373),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1380),
.B(n_1339),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1392),
.A2(n_1359),
.B1(n_1345),
.B2(n_1331),
.Y(n_1474)
);

O2A1O1Ixp33_ASAP7_75t_L g1475 ( 
.A1(n_1410),
.A2(n_1392),
.B(n_1366),
.C(n_1425),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1404),
.B(n_1376),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1404),
.B(n_1376),
.Y(n_1477)
);

OAI22xp5_ASAP7_75t_SL g1478 ( 
.A1(n_1366),
.A2(n_1410),
.B1(n_1414),
.B2(n_1425),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1373),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1396),
.B(n_1400),
.Y(n_1480)
);

O2A1O1Ixp33_ASAP7_75t_L g1481 ( 
.A1(n_1367),
.A2(n_1427),
.B(n_1426),
.C(n_1407),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1400),
.B(n_1415),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_1383),
.Y(n_1483)
);

A2O1A1Ixp33_ASAP7_75t_L g1484 ( 
.A1(n_1418),
.A2(n_1367),
.B(n_1408),
.C(n_1427),
.Y(n_1484)
);

A2O1A1Ixp33_ASAP7_75t_L g1485 ( 
.A1(n_1418),
.A2(n_1426),
.B(n_1416),
.C(n_1415),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1368),
.Y(n_1486)
);

OA21x2_ASAP7_75t_L g1487 ( 
.A1(n_1389),
.A2(n_1406),
.B(n_1423),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1378),
.B(n_1381),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1388),
.B(n_1382),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1382),
.B(n_1398),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1397),
.Y(n_1491)
);

BUFx12f_ASAP7_75t_L g1492 ( 
.A(n_1432),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1414),
.A2(n_1401),
.B1(n_1432),
.B2(n_1429),
.Y(n_1493)
);

A2O1A1Ixp33_ASAP7_75t_L g1494 ( 
.A1(n_1416),
.A2(n_1431),
.B(n_1389),
.C(n_1369),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1419),
.A2(n_1434),
.B1(n_1383),
.B2(n_1409),
.Y(n_1495)
);

OAI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1423),
.A2(n_1424),
.B(n_1441),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1444),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1472),
.Y(n_1498)
);

INVxp67_ASAP7_75t_SL g1499 ( 
.A(n_1488),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1476),
.B(n_1477),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1472),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1449),
.B(n_1490),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1479),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1463),
.B(n_1397),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1476),
.B(n_1381),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1449),
.B(n_1402),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1477),
.B(n_1387),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1458),
.B(n_1461),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1490),
.B(n_1402),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1489),
.B(n_1402),
.Y(n_1510)
);

INVx3_ASAP7_75t_L g1511 ( 
.A(n_1463),
.Y(n_1511)
);

BUFx2_ASAP7_75t_L g1512 ( 
.A(n_1463),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1488),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1489),
.B(n_1402),
.Y(n_1514)
);

BUFx2_ASAP7_75t_L g1515 ( 
.A(n_1483),
.Y(n_1515)
);

BUFx2_ASAP7_75t_L g1516 ( 
.A(n_1483),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1480),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1478),
.A2(n_1434),
.B1(n_1409),
.B2(n_1433),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1480),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1445),
.B(n_1391),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1486),
.B(n_1390),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1482),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1498),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_1515),
.Y(n_1524)
);

INVx2_ASAP7_75t_SL g1525 ( 
.A(n_1511),
.Y(n_1525)
);

NAND4xp25_ASAP7_75t_L g1526 ( 
.A(n_1518),
.B(n_1446),
.C(n_1455),
.D(n_1475),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1520),
.B(n_1453),
.Y(n_1527)
);

OR2x6_ASAP7_75t_L g1528 ( 
.A(n_1520),
.B(n_1470),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1509),
.B(n_1487),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1511),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1498),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1498),
.Y(n_1532)
);

INVx4_ASAP7_75t_L g1533 ( 
.A(n_1504),
.Y(n_1533)
);

BUFx3_ASAP7_75t_L g1534 ( 
.A(n_1515),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1499),
.B(n_1484),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1508),
.B(n_1487),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1519),
.B(n_1453),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1519),
.B(n_1453),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1501),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1501),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1503),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1509),
.B(n_1487),
.Y(n_1542)
);

OAI33xp33_ASAP7_75t_L g1543 ( 
.A1(n_1521),
.A2(n_1478),
.A3(n_1493),
.B1(n_1452),
.B2(n_1481),
.B3(n_1474),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1510),
.A2(n_1446),
.B(n_1447),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1506),
.A2(n_1450),
.B1(n_1451),
.B2(n_1495),
.Y(n_1545)
);

OAI222xp33_ASAP7_75t_L g1546 ( 
.A1(n_1506),
.A2(n_1442),
.B1(n_1447),
.B2(n_1473),
.C1(n_1470),
.C2(n_1401),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1500),
.B(n_1445),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1513),
.B(n_1505),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1500),
.B(n_1445),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1505),
.B(n_1485),
.Y(n_1550)
);

AOI221xp5_ASAP7_75t_L g1551 ( 
.A1(n_1510),
.A2(n_1471),
.B1(n_1466),
.B2(n_1459),
.C(n_1473),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1497),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1497),
.Y(n_1553)
);

INVx4_ASAP7_75t_L g1554 ( 
.A(n_1504),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1517),
.B(n_1448),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1526),
.A2(n_1450),
.B1(n_1442),
.B2(n_1470),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1527),
.B(n_1512),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1552),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1527),
.B(n_1547),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1535),
.B(n_1550),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1523),
.Y(n_1561)
);

INVx4_ASAP7_75t_L g1562 ( 
.A(n_1534),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1527),
.B(n_1512),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1543),
.B(n_1460),
.Y(n_1564)
);

INVx2_ASAP7_75t_SL g1565 ( 
.A(n_1534),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1529),
.B(n_1514),
.Y(n_1566)
);

NOR3xp33_ASAP7_75t_L g1567 ( 
.A(n_1543),
.B(n_1464),
.C(n_1465),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1547),
.B(n_1522),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1547),
.B(n_1522),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1552),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1549),
.B(n_1448),
.Y(n_1571)
);

NOR2x1_ASAP7_75t_L g1572 ( 
.A(n_1534),
.B(n_1468),
.Y(n_1572)
);

INVx1_ASAP7_75t_SL g1573 ( 
.A(n_1524),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1526),
.B(n_1454),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1553),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1529),
.B(n_1514),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1549),
.B(n_1448),
.Y(n_1577)
);

INVx1_ASAP7_75t_SL g1578 ( 
.A(n_1524),
.Y(n_1578)
);

OR2x6_ASAP7_75t_L g1579 ( 
.A(n_1528),
.B(n_1470),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1553),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1532),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1523),
.Y(n_1582)
);

NAND2x1_ASAP7_75t_L g1583 ( 
.A(n_1528),
.B(n_1469),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1523),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1549),
.B(n_1537),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1535),
.B(n_1502),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1537),
.B(n_1448),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1537),
.B(n_1517),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1531),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1532),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1550),
.B(n_1502),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1540),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1538),
.B(n_1511),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1529),
.B(n_1507),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1558),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1559),
.B(n_1533),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1589),
.Y(n_1597)
);

OR2x6_ASAP7_75t_L g1598 ( 
.A(n_1562),
.B(n_1544),
.Y(n_1598)
);

OAI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1564),
.A2(n_1544),
.B(n_1545),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1559),
.B(n_1533),
.Y(n_1600)
);

INVxp33_ASAP7_75t_L g1601 ( 
.A(n_1574),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1558),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1559),
.B(n_1533),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1564),
.B(n_1454),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1586),
.B(n_1548),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1570),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1570),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1556),
.A2(n_1560),
.B1(n_1567),
.B2(n_1545),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_L g1609 ( 
.A(n_1574),
.B(n_1492),
.Y(n_1609)
);

NOR2x1_ASAP7_75t_L g1610 ( 
.A(n_1562),
.B(n_1546),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1586),
.B(n_1591),
.Y(n_1611)
);

INVxp67_ASAP7_75t_L g1612 ( 
.A(n_1560),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1585),
.B(n_1568),
.Y(n_1613)
);

NOR2x1_ASAP7_75t_L g1614 ( 
.A(n_1562),
.B(n_1546),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1575),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1575),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1591),
.B(n_1551),
.Y(n_1617)
);

INVx2_ASAP7_75t_SL g1618 ( 
.A(n_1565),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1567),
.B(n_1551),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1580),
.Y(n_1620)
);

OAI21xp5_ASAP7_75t_SL g1621 ( 
.A1(n_1556),
.A2(n_1467),
.B(n_1462),
.Y(n_1621)
);

INVxp67_ASAP7_75t_L g1622 ( 
.A(n_1565),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1580),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1592),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1592),
.Y(n_1625)
);

A2O1A1Ixp33_ASAP7_75t_L g1626 ( 
.A1(n_1583),
.A2(n_1450),
.B(n_1494),
.C(n_1447),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1585),
.B(n_1533),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1568),
.B(n_1507),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1581),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1581),
.Y(n_1630)
);

NOR3xp33_ASAP7_75t_L g1631 ( 
.A(n_1562),
.B(n_1583),
.C(n_1572),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1590),
.Y(n_1632)
);

INVx2_ASAP7_75t_SL g1633 ( 
.A(n_1565),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1590),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1585),
.B(n_1554),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1561),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1594),
.B(n_1566),
.Y(n_1637)
);

NAND2x1p5_ASAP7_75t_L g1638 ( 
.A(n_1610),
.B(n_1562),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1613),
.B(n_1571),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1613),
.B(n_1571),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1612),
.B(n_1617),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1595),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1619),
.B(n_1568),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1608),
.B(n_1569),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1599),
.B(n_1573),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1602),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1604),
.B(n_1569),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1614),
.B(n_1571),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1604),
.B(n_1569),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1598),
.B(n_1577),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1605),
.B(n_1611),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1597),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1597),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1606),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1607),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1637),
.B(n_1566),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1624),
.B(n_1566),
.Y(n_1657)
);

INVx2_ASAP7_75t_SL g1658 ( 
.A(n_1618),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1598),
.B(n_1596),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1618),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1601),
.B(n_1573),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1625),
.B(n_1576),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1601),
.B(n_1578),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1622),
.B(n_1578),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1633),
.Y(n_1665)
);

INVx1_ASAP7_75t_SL g1666 ( 
.A(n_1633),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1598),
.B(n_1577),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_SL g1668 ( 
.A(n_1626),
.B(n_1572),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1615),
.Y(n_1669)
);

AOI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1626),
.A2(n_1447),
.B(n_1583),
.Y(n_1670)
);

OAI21xp33_ASAP7_75t_L g1671 ( 
.A1(n_1598),
.A2(n_1587),
.B(n_1456),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1609),
.B(n_1412),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1616),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_SL g1674 ( 
.A1(n_1645),
.A2(n_1644),
.B1(n_1638),
.B2(n_1648),
.Y(n_1674)
);

OAI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1645),
.A2(n_1621),
.B1(n_1528),
.B2(n_1579),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1642),
.Y(n_1676)
);

OAI211xp5_ASAP7_75t_L g1677 ( 
.A1(n_1668),
.A2(n_1631),
.B(n_1609),
.C(n_1629),
.Y(n_1677)
);

AOI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1670),
.A2(n_1579),
.B1(n_1528),
.B2(n_1577),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1643),
.B(n_1630),
.Y(n_1679)
);

INVxp67_ASAP7_75t_L g1680 ( 
.A(n_1661),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1672),
.B(n_1628),
.Y(n_1681)
);

OAI221xp5_ASAP7_75t_L g1682 ( 
.A1(n_1638),
.A2(n_1579),
.B1(n_1632),
.B2(n_1634),
.C(n_1623),
.Y(n_1682)
);

OAI322xp33_ASAP7_75t_L g1683 ( 
.A1(n_1638),
.A2(n_1620),
.A3(n_1576),
.B1(n_1542),
.B2(n_1636),
.C1(n_1594),
.C2(n_1536),
.Y(n_1683)
);

OAI21xp33_ASAP7_75t_SL g1684 ( 
.A1(n_1648),
.A2(n_1641),
.B(n_1659),
.Y(n_1684)
);

INVx1_ASAP7_75t_SL g1685 ( 
.A(n_1666),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1663),
.B(n_1492),
.Y(n_1686)
);

OAI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1664),
.A2(n_1635),
.B(n_1627),
.Y(n_1687)
);

INVx1_ASAP7_75t_SL g1688 ( 
.A(n_1666),
.Y(n_1688)
);

A2O1A1Ixp33_ASAP7_75t_SL g1689 ( 
.A1(n_1660),
.A2(n_1496),
.B(n_1456),
.C(n_1589),
.Y(n_1689)
);

AOI22xp33_ASAP7_75t_L g1690 ( 
.A1(n_1647),
.A2(n_1579),
.B1(n_1528),
.B2(n_1470),
.Y(n_1690)
);

INVx2_ASAP7_75t_SL g1691 ( 
.A(n_1658),
.Y(n_1691)
);

AOI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1649),
.A2(n_1579),
.B1(n_1528),
.B2(n_1635),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1651),
.B(n_1576),
.Y(n_1693)
);

AOI322xp5_ASAP7_75t_L g1694 ( 
.A1(n_1671),
.A2(n_1587),
.A3(n_1627),
.B1(n_1603),
.B2(n_1600),
.C1(n_1596),
.C2(n_1563),
.Y(n_1694)
);

OAI211xp5_ASAP7_75t_SL g1695 ( 
.A1(n_1671),
.A2(n_1395),
.B(n_1422),
.C(n_1429),
.Y(n_1695)
);

NAND2xp33_ASAP7_75t_L g1696 ( 
.A(n_1651),
.B(n_1600),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1659),
.A2(n_1579),
.B1(n_1457),
.B2(n_1603),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1658),
.Y(n_1698)
);

OAI21xp5_ASAP7_75t_SL g1699 ( 
.A1(n_1650),
.A2(n_1587),
.B(n_1447),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1676),
.Y(n_1700)
);

NOR4xp25_ASAP7_75t_L g1701 ( 
.A(n_1677),
.B(n_1660),
.C(n_1669),
.D(n_1655),
.Y(n_1701)
);

INVx2_ASAP7_75t_SL g1702 ( 
.A(n_1691),
.Y(n_1702)
);

OAI222xp33_ASAP7_75t_L g1703 ( 
.A1(n_1674),
.A2(n_1665),
.B1(n_1660),
.B2(n_1657),
.C1(n_1662),
.C2(n_1667),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1685),
.B(n_1656),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1688),
.Y(n_1705)
);

O2A1O1Ixp5_ASAP7_75t_SL g1706 ( 
.A1(n_1680),
.A2(n_1655),
.B(n_1646),
.C(n_1654),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1698),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1693),
.Y(n_1708)
);

AOI221xp5_ASAP7_75t_L g1709 ( 
.A1(n_1674),
.A2(n_1699),
.B1(n_1683),
.B2(n_1684),
.C(n_1675),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1679),
.Y(n_1710)
);

XNOR2xp5_ASAP7_75t_L g1711 ( 
.A(n_1692),
.B(n_1650),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1681),
.B(n_1696),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1687),
.Y(n_1713)
);

OAI211xp5_ASAP7_75t_L g1714 ( 
.A1(n_1678),
.A2(n_1682),
.B(n_1694),
.C(n_1689),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1686),
.B(n_1642),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1697),
.B(n_1667),
.Y(n_1716)
);

INVxp67_ASAP7_75t_SL g1717 ( 
.A(n_1690),
.Y(n_1717)
);

NAND3xp33_ASAP7_75t_SL g1718 ( 
.A(n_1695),
.B(n_1662),
.C(n_1657),
.Y(n_1718)
);

OAI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1695),
.A2(n_1579),
.B1(n_1656),
.B2(n_1639),
.Y(n_1719)
);

OAI32xp33_ASAP7_75t_L g1720 ( 
.A1(n_1684),
.A2(n_1673),
.A3(n_1669),
.B1(n_1646),
.B2(n_1654),
.Y(n_1720)
);

AOI221xp5_ASAP7_75t_L g1721 ( 
.A1(n_1701),
.A2(n_1673),
.B1(n_1640),
.B2(n_1639),
.C(n_1652),
.Y(n_1721)
);

O2A1O1Ixp33_ASAP7_75t_L g1722 ( 
.A1(n_1703),
.A2(n_1653),
.B(n_1652),
.C(n_1640),
.Y(n_1722)
);

O2A1O1Ixp33_ASAP7_75t_L g1723 ( 
.A1(n_1703),
.A2(n_1653),
.B(n_1652),
.C(n_1542),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1704),
.Y(n_1724)
);

OAI21xp33_ASAP7_75t_L g1725 ( 
.A1(n_1709),
.A2(n_1653),
.B(n_1483),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1702),
.B(n_1557),
.Y(n_1726)
);

OAI21xp33_ASAP7_75t_L g1727 ( 
.A1(n_1717),
.A2(n_1521),
.B(n_1443),
.Y(n_1727)
);

AOI211xp5_ASAP7_75t_L g1728 ( 
.A1(n_1714),
.A2(n_1441),
.B(n_1542),
.C(n_1555),
.Y(n_1728)
);

AOI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1718),
.A2(n_1457),
.B1(n_1469),
.B2(n_1491),
.Y(n_1729)
);

NAND2x1_ASAP7_75t_SL g1730 ( 
.A(n_1705),
.B(n_1557),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1716),
.B(n_1557),
.Y(n_1731)
);

OAI321xp33_ASAP7_75t_L g1732 ( 
.A1(n_1728),
.A2(n_1718),
.A3(n_1713),
.B1(n_1708),
.B2(n_1717),
.C(n_1712),
.Y(n_1732)
);

INVx3_ASAP7_75t_L g1733 ( 
.A(n_1724),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1725),
.B(n_1702),
.Y(n_1734)
);

AOI22xp33_ASAP7_75t_L g1735 ( 
.A1(n_1731),
.A2(n_1711),
.B1(n_1719),
.B2(n_1710),
.Y(n_1735)
);

A2O1A1Ixp33_ASAP7_75t_L g1736 ( 
.A1(n_1730),
.A2(n_1720),
.B(n_1707),
.C(n_1715),
.Y(n_1736)
);

AOI221xp5_ASAP7_75t_L g1737 ( 
.A1(n_1723),
.A2(n_1700),
.B1(n_1706),
.B2(n_1555),
.C(n_1589),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1726),
.B(n_1563),
.Y(n_1738)
);

NOR3xp33_ASAP7_75t_L g1739 ( 
.A(n_1727),
.B(n_1441),
.C(n_1491),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1721),
.B(n_1563),
.Y(n_1740)
);

NAND4xp25_ASAP7_75t_L g1741 ( 
.A(n_1735),
.B(n_1729),
.C(n_1722),
.D(n_1428),
.Y(n_1741)
);

AOI221xp5_ASAP7_75t_L g1742 ( 
.A1(n_1732),
.A2(n_1589),
.B1(n_1555),
.B2(n_1584),
.C(n_1582),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1734),
.B(n_1561),
.Y(n_1743)
);

AOI311xp33_ASAP7_75t_L g1744 ( 
.A1(n_1736),
.A2(n_1439),
.A3(n_1436),
.B(n_1539),
.C(n_1541),
.Y(n_1744)
);

OAI221xp5_ASAP7_75t_SL g1745 ( 
.A1(n_1740),
.A2(n_1457),
.B1(n_1536),
.B2(n_1508),
.C(n_1516),
.Y(n_1745)
);

AOI222xp33_ASAP7_75t_L g1746 ( 
.A1(n_1743),
.A2(n_1737),
.B1(n_1733),
.B2(n_1738),
.C1(n_1739),
.C2(n_1593),
.Y(n_1746)
);

NAND3xp33_ASAP7_75t_L g1747 ( 
.A(n_1741),
.B(n_1582),
.C(n_1561),
.Y(n_1747)
);

AOI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1742),
.A2(n_1593),
.B1(n_1468),
.B2(n_1554),
.Y(n_1748)
);

NOR3xp33_ASAP7_75t_L g1749 ( 
.A(n_1745),
.B(n_1435),
.C(n_1385),
.Y(n_1749)
);

NOR3xp33_ASAP7_75t_L g1750 ( 
.A(n_1744),
.B(n_1435),
.C(n_1385),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1743),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1751),
.Y(n_1752)
);

INVxp33_ASAP7_75t_L g1753 ( 
.A(n_1749),
.Y(n_1753)
);

OAI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1748),
.A2(n_1582),
.B1(n_1584),
.B2(n_1593),
.Y(n_1754)
);

XNOR2xp5_ASAP7_75t_L g1755 ( 
.A(n_1747),
.B(n_1469),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1750),
.B(n_1584),
.Y(n_1756)
);

AND2x4_ASAP7_75t_L g1757 ( 
.A(n_1752),
.B(n_1756),
.Y(n_1757)
);

O2A1O1Ixp33_ASAP7_75t_L g1758 ( 
.A1(n_1753),
.A2(n_1754),
.B(n_1746),
.C(n_1755),
.Y(n_1758)
);

NOR2x1_ASAP7_75t_L g1759 ( 
.A(n_1752),
.B(n_1437),
.Y(n_1759)
);

NOR2x1_ASAP7_75t_L g1760 ( 
.A(n_1757),
.B(n_1437),
.Y(n_1760)
);

AOI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1760),
.A2(n_1759),
.B1(n_1758),
.B2(n_1588),
.Y(n_1761)
);

AOI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1761),
.A2(n_1588),
.B1(n_1525),
.B2(n_1554),
.Y(n_1762)
);

INVx4_ASAP7_75t_L g1763 ( 
.A(n_1761),
.Y(n_1763)
);

NAND3xp33_ASAP7_75t_L g1764 ( 
.A(n_1763),
.B(n_1554),
.C(n_1421),
.Y(n_1764)
);

CKINVDCx20_ASAP7_75t_R g1765 ( 
.A(n_1762),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1765),
.Y(n_1766)
);

INVxp67_ASAP7_75t_L g1767 ( 
.A(n_1764),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1766),
.B(n_1588),
.Y(n_1768)
);

A2O1A1Ixp33_ASAP7_75t_SL g1769 ( 
.A1(n_1768),
.A2(n_1767),
.B(n_1530),
.C(n_1438),
.Y(n_1769)
);

AOI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1769),
.A2(n_1437),
.B1(n_1525),
.B2(n_1530),
.Y(n_1770)
);

OAI221xp5_ASAP7_75t_R g1771 ( 
.A1(n_1770),
.A2(n_1525),
.B1(n_1530),
.B2(n_1437),
.C(n_1440),
.Y(n_1771)
);

AOI211xp5_ASAP7_75t_L g1772 ( 
.A1(n_1771),
.A2(n_1413),
.B(n_1411),
.C(n_1421),
.Y(n_1772)
);


endmodule