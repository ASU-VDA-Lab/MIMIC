module real_aes_8017_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_357;
wire n_287;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_374;
wire n_379;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_462;
wire n_289;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
A2O1A1Ixp33_ASAP7_75t_L g320 ( .A1(n_0), .A2(n_231), .B(n_234), .C(n_321), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_1), .A2(n_259), .B(n_260), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_2), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g216 ( .A(n_3), .Y(n_216) );
AND2x6_ASAP7_75t_L g231 ( .A(n_3), .B(n_214), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_3), .B(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g376 ( .A(n_4), .Y(n_376) );
NAND2xp5_ASAP7_75t_SL g323 ( .A(n_5), .B(n_242), .Y(n_323) );
AO22x2_ASAP7_75t_L g103 ( .A1(n_6), .A2(n_28), .B1(n_95), .B2(n_100), .Y(n_103) );
INVx1_ASAP7_75t_L g250 ( .A(n_7), .Y(n_250) );
AOI22xp5_ASAP7_75t_L g196 ( .A1(n_8), .A2(n_41), .B1(n_197), .B2(n_198), .Y(n_196) );
INVx1_ASAP7_75t_L g198 ( .A(n_8), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_9), .Y(n_179) );
A2O1A1Ixp33_ASAP7_75t_L g331 ( .A1(n_10), .A2(n_240), .B(n_332), .C(n_334), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_11), .B(n_271), .Y(n_335) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_12), .Y(n_166) );
AO22x2_ASAP7_75t_L g105 ( .A1(n_13), .A2(n_30), .B1(n_95), .B2(n_96), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_14), .B(n_290), .Y(n_289) );
A2O1A1Ixp33_ASAP7_75t_L g340 ( .A1(n_15), .A2(n_264), .B(n_341), .C(n_343), .Y(n_340) );
INVx1_ASAP7_75t_L g539 ( .A(n_15), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_16), .B(n_242), .Y(n_301) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_17), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_18), .B(n_242), .Y(n_241) );
CKINVDCx16_ASAP7_75t_R g295 ( .A(n_19), .Y(n_295) );
INVx1_ASAP7_75t_L g238 ( .A(n_20), .Y(n_238) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_21), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g113 ( .A1(n_22), .A2(n_40), .B1(n_114), .B2(n_119), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g319 ( .A(n_23), .Y(n_319) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_24), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_25), .Y(n_153) );
INVx1_ASAP7_75t_L g285 ( .A(n_26), .Y(n_285) );
INVx2_ASAP7_75t_L g229 ( .A(n_27), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g325 ( .A(n_29), .Y(n_325) );
OAI221xp5_ASAP7_75t_L g207 ( .A1(n_30), .A2(n_45), .B1(n_54), .B2(n_208), .C(n_209), .Y(n_207) );
INVxp67_ASAP7_75t_L g210 ( .A(n_30), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g263 ( .A1(n_31), .A2(n_264), .B(n_265), .C(n_267), .Y(n_263) );
INVxp67_ASAP7_75t_L g286 ( .A(n_32), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_33), .A2(n_193), .B1(n_194), .B2(n_203), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_33), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g136 ( .A1(n_34), .A2(n_55), .B1(n_137), .B2(n_141), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g233 ( .A1(n_35), .A2(n_234), .B(n_237), .C(n_245), .Y(n_233) );
CKINVDCx14_ASAP7_75t_R g261 ( .A(n_36), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_L g373 ( .A1(n_37), .A2(n_303), .B(n_374), .C(n_375), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g252 ( .A(n_38), .Y(n_252) );
CKINVDCx20_ASAP7_75t_R g282 ( .A(n_39), .Y(n_282) );
INVx1_ASAP7_75t_L g197 ( .A(n_41), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g171 ( .A(n_42), .Y(n_171) );
INVx1_ASAP7_75t_L g339 ( .A(n_43), .Y(n_339) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_44), .Y(n_106) );
AO22x2_ASAP7_75t_L g94 ( .A1(n_45), .A2(n_65), .B1(n_95), .B2(n_96), .Y(n_94) );
INVxp67_ASAP7_75t_L g211 ( .A(n_45), .Y(n_211) );
CKINVDCx14_ASAP7_75t_R g372 ( .A(n_46), .Y(n_372) );
INVx1_ASAP7_75t_L g214 ( .A(n_47), .Y(n_214) );
INVx1_ASAP7_75t_L g249 ( .A(n_48), .Y(n_249) );
INVx1_ASAP7_75t_SL g266 ( .A(n_49), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_50), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_51), .B(n_271), .Y(n_345) );
AOI22xp5_ASAP7_75t_L g194 ( .A1(n_52), .A2(n_195), .B1(n_201), .B2(n_202), .Y(n_194) );
INVx1_ASAP7_75t_L g201 ( .A(n_52), .Y(n_201) );
INVx1_ASAP7_75t_L g298 ( .A(n_53), .Y(n_298) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_54), .A2(n_71), .B1(n_95), .B2(n_100), .Y(n_99) );
AOI21xp5_ASAP7_75t_L g370 ( .A1(n_56), .A2(n_259), .B(n_371), .Y(n_370) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_57), .Y(n_135) );
INVx1_ASAP7_75t_L g84 ( .A(n_58), .Y(n_84) );
AOI21xp5_ASAP7_75t_L g328 ( .A1(n_58), .A2(n_259), .B(n_329), .Y(n_328) );
CKINVDCx20_ASAP7_75t_R g307 ( .A(n_59), .Y(n_307) );
OAI22xp5_ASAP7_75t_SL g82 ( .A1(n_60), .A2(n_83), .B1(n_84), .B2(n_85), .Y(n_82) );
CKINVDCx20_ASAP7_75t_R g85 ( .A(n_60), .Y(n_85) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_60), .A2(n_280), .B(n_281), .Y(n_279) );
CKINVDCx16_ASAP7_75t_R g232 ( .A(n_61), .Y(n_232) );
INVx1_ASAP7_75t_L g330 ( .A(n_62), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_63), .A2(n_259), .B(n_338), .Y(n_337) );
AOI22xp5_ASAP7_75t_SL g528 ( .A1(n_63), .A2(n_86), .B1(n_191), .B2(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_63), .Y(n_529) );
INVx1_ASAP7_75t_L g333 ( .A(n_64), .Y(n_333) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_66), .Y(n_177) );
INVx2_ASAP7_75t_L g247 ( .A(n_67), .Y(n_247) );
INVx1_ASAP7_75t_L g322 ( .A(n_68), .Y(n_322) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_69), .Y(n_147) );
A2O1A1Ixp33_ASAP7_75t_L g296 ( .A1(n_70), .A2(n_234), .B(n_297), .C(n_305), .Y(n_296) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_72), .A2(n_196), .B1(n_199), .B2(n_200), .Y(n_195) );
INVx1_ASAP7_75t_L g199 ( .A(n_72), .Y(n_199) );
XNOR2xp5_ASAP7_75t_L g540 ( .A(n_73), .B(n_191), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_74), .B(n_254), .Y(n_377) );
INVx1_ASAP7_75t_L g95 ( .A(n_75), .Y(n_95) );
INVx1_ASAP7_75t_L g97 ( .A(n_75), .Y(n_97) );
INVx2_ASAP7_75t_L g342 ( .A(n_76), .Y(n_342) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_77), .Y(n_184) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_204), .B1(n_217), .B2(n_523), .C(n_527), .Y(n_78) );
XOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_192), .Y(n_79) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_81), .A2(n_82), .B1(n_86), .B2(n_191), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_82), .Y(n_81) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_84), .Y(n_83) );
INVx1_ASAP7_75t_SL g191 ( .A(n_86), .Y(n_191) );
AND2x2_ASAP7_75t_SL g86 ( .A(n_87), .B(n_145), .Y(n_86) );
NOR2xp33_ASAP7_75t_L g87 ( .A(n_88), .B(n_124), .Y(n_87) );
OAI221xp5_ASAP7_75t_SL g88 ( .A1(n_89), .A2(n_106), .B1(n_107), .B2(n_112), .C(n_113), .Y(n_88) );
INVx3_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
AND2x2_ASAP7_75t_L g91 ( .A(n_92), .B(n_101), .Y(n_91) );
AND2x6_ASAP7_75t_L g116 ( .A(n_92), .B(n_117), .Y(n_116) );
AND2x4_ASAP7_75t_L g127 ( .A(n_92), .B(n_128), .Y(n_127) );
AND2x6_ASAP7_75t_L g169 ( .A(n_92), .B(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_L g92 ( .A(n_93), .B(n_98), .Y(n_92) );
AND2x2_ASAP7_75t_L g111 ( .A(n_93), .B(n_99), .Y(n_111) );
INVx2_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_94), .B(n_99), .Y(n_123) );
AND2x2_ASAP7_75t_L g133 ( .A(n_94), .B(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g165 ( .A(n_94), .B(n_103), .Y(n_165) );
INVx1_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
INVx1_ASAP7_75t_L g100 ( .A(n_97), .Y(n_100) );
INVx1_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
INVx1_ASAP7_75t_L g134 ( .A(n_99), .Y(n_134) );
INVx1_ASAP7_75t_L g164 ( .A(n_99), .Y(n_164) );
AND2x4_ASAP7_75t_L g110 ( .A(n_101), .B(n_111), .Y(n_110) );
AND2x4_ASAP7_75t_L g121 ( .A(n_101), .B(n_122), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_101), .B(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_104), .Y(n_101) );
OR2x2_ASAP7_75t_L g118 ( .A(n_102), .B(n_105), .Y(n_118) );
AND2x2_ASAP7_75t_L g128 ( .A(n_102), .B(n_105), .Y(n_128) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_L g170 ( .A(n_103), .B(n_105), .Y(n_170) );
AND2x2_ASAP7_75t_L g163 ( .A(n_104), .B(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g183 ( .A(n_104), .Y(n_183) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g144 ( .A(n_105), .Y(n_144) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx3_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g152 ( .A(n_111), .Y(n_152) );
NAND2x1p5_ASAP7_75t_L g157 ( .A(n_111), .B(n_128), .Y(n_157) );
INVx4_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx11_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OR2x2_ASAP7_75t_L g151 ( .A(n_118), .B(n_152), .Y(n_151) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OR2x6_ASAP7_75t_L g143 ( .A(n_123), .B(n_144), .Y(n_143) );
OAI221xp5_ASAP7_75t_SL g124 ( .A1(n_125), .A2(n_129), .B1(n_130), .B2(n_135), .C(n_136), .Y(n_124) );
INVx3_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
BUFx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g140 ( .A(n_128), .B(n_133), .Y(n_140) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g190 ( .A(n_134), .Y(n_190) );
BUFx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx5_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx8_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx4f_ASAP7_75t_SL g141 ( .A(n_142), .Y(n_141) );
INVx6_ASAP7_75t_SL g142 ( .A(n_143), .Y(n_142) );
NOR3xp33_ASAP7_75t_L g145 ( .A(n_146), .B(n_158), .C(n_178), .Y(n_145) );
OAI22xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B1(n_153), .B2(n_154), .Y(n_146) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
OAI222xp33_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_166), .B1(n_167), .B2(n_171), .C1(n_172), .C2(n_177), .Y(n_158) );
INVx2_ASAP7_75t_SL g159 ( .A(n_160), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_163), .B(n_165), .Y(n_162) );
INVx1_ASAP7_75t_L g176 ( .A(n_164), .Y(n_176) );
AND2x4_ASAP7_75t_L g175 ( .A(n_165), .B(n_176), .Y(n_175) );
NAND2x1p5_ASAP7_75t_L g182 ( .A(n_165), .B(n_183), .Y(n_182) );
INVx2_ASAP7_75t_SL g167 ( .A(n_168), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g188 ( .A(n_170), .Y(n_188) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
BUFx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
OAI22xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B1(n_184), .B2(n_185), .Y(n_178) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx4_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
CKINVDCx16_ASAP7_75t_R g186 ( .A(n_187), .Y(n_186) );
OR2x6_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_194), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_195), .Y(n_202) );
INVx1_ASAP7_75t_L g200 ( .A(n_196), .Y(n_200) );
CKINVDCx16_ASAP7_75t_R g204 ( .A(n_205), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_206), .Y(n_205) );
AND3x1_ASAP7_75t_SL g206 ( .A(n_207), .B(n_212), .C(n_215), .Y(n_206) );
INVxp67_ASAP7_75t_L g533 ( .A(n_207), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
INVx1_ASAP7_75t_SL g535 ( .A(n_212), .Y(n_535) );
OAI21xp5_ASAP7_75t_L g537 ( .A1(n_212), .A2(n_525), .B(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g544 ( .A(n_212), .Y(n_544) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_213), .B(n_216), .Y(n_538) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
OR2x2_ASAP7_75t_SL g543 ( .A(n_215), .B(n_544), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_216), .Y(n_215) );
OR3x1_ASAP7_75t_L g217 ( .A(n_218), .B(n_434), .C(n_481), .Y(n_217) );
NAND3xp33_ASAP7_75t_SL g218 ( .A(n_219), .B(n_380), .C(n_405), .Y(n_218) );
AOI221xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_315), .B1(n_346), .B2(n_349), .C(n_357), .Y(n_219) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_272), .B(n_308), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_222), .B(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_222), .B(n_362), .Y(n_478) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_256), .Y(n_222) );
AND2x2_ASAP7_75t_L g348 ( .A(n_223), .B(n_314), .Y(n_348) );
AND2x2_ASAP7_75t_L g398 ( .A(n_223), .B(n_313), .Y(n_398) );
AND2x2_ASAP7_75t_L g419 ( .A(n_223), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g424 ( .A(n_223), .B(n_391), .Y(n_424) );
OR2x2_ASAP7_75t_L g432 ( .A(n_223), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g504 ( .A(n_223), .B(n_292), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_223), .B(n_453), .Y(n_518) );
INVx3_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g363 ( .A(n_224), .B(n_256), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_224), .B(n_292), .Y(n_364) );
AND2x4_ASAP7_75t_L g386 ( .A(n_224), .B(n_314), .Y(n_386) );
AND2x2_ASAP7_75t_L g416 ( .A(n_224), .B(n_274), .Y(n_416) );
AND2x2_ASAP7_75t_L g425 ( .A(n_224), .B(n_415), .Y(n_425) );
AND2x2_ASAP7_75t_L g441 ( .A(n_224), .B(n_293), .Y(n_441) );
OR2x2_ASAP7_75t_L g450 ( .A(n_224), .B(n_433), .Y(n_450) );
AND2x2_ASAP7_75t_L g456 ( .A(n_224), .B(n_391), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_224), .B(n_462), .Y(n_461) );
OR2x2_ASAP7_75t_L g470 ( .A(n_224), .B(n_310), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_224), .B(n_359), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_224), .B(n_420), .Y(n_509) );
OR2x6_ASAP7_75t_L g224 ( .A(n_225), .B(n_251), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_232), .B(n_233), .C(n_246), .Y(n_225) );
OAI21xp5_ASAP7_75t_L g294 ( .A1(n_226), .A2(n_295), .B(n_296), .Y(n_294) );
OAI21xp5_ASAP7_75t_L g318 ( .A1(n_226), .A2(n_319), .B(n_320), .Y(n_318) );
NAND2x1p5_ASAP7_75t_L g226 ( .A(n_227), .B(n_231), .Y(n_226) );
AND2x4_ASAP7_75t_L g259 ( .A(n_227), .B(n_231), .Y(n_259) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_230), .Y(n_227) );
INVx1_ASAP7_75t_L g244 ( .A(n_228), .Y(n_244) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g235 ( .A(n_229), .Y(n_235) );
INVx1_ASAP7_75t_L g344 ( .A(n_229), .Y(n_344) );
INVx1_ASAP7_75t_L g236 ( .A(n_230), .Y(n_236) );
INVx3_ASAP7_75t_L g240 ( .A(n_230), .Y(n_240) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_230), .Y(n_242) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_230), .Y(n_288) );
BUFx3_ASAP7_75t_L g245 ( .A(n_231), .Y(n_245) );
INVx4_ASAP7_75t_SL g269 ( .A(n_231), .Y(n_269) );
INVx5_ASAP7_75t_L g262 ( .A(n_234), .Y(n_262) );
AND2x6_ASAP7_75t_L g234 ( .A(n_235), .B(n_236), .Y(n_234) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_235), .Y(n_268) );
BUFx3_ASAP7_75t_L g304 ( .A(n_235), .Y(n_304) );
O2A1O1Ixp33_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B(n_241), .C(n_243), .Y(n_237) );
OAI22xp33_ASAP7_75t_L g284 ( .A1(n_239), .A2(n_285), .B1(n_286), .B2(n_287), .Y(n_284) );
INVx5_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_240), .B(n_376), .Y(n_375) );
INVx4_ASAP7_75t_L g264 ( .A(n_242), .Y(n_264) );
INVx2_ASAP7_75t_L g374 ( .A(n_242), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_243), .B(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_244), .B(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_245), .B(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g291 ( .A(n_246), .Y(n_291) );
INVx1_ASAP7_75t_L g317 ( .A(n_246), .Y(n_317) );
OA21x2_ASAP7_75t_L g369 ( .A1(n_246), .A2(n_370), .B(n_377), .Y(n_369) );
AND2x2_ASAP7_75t_SL g246 ( .A(n_247), .B(n_248), .Y(n_246) );
AND2x2_ASAP7_75t_L g255 ( .A(n_247), .B(n_248), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
INVx3_ASAP7_75t_L g271 ( .A(n_253), .Y(n_271) );
AO21x2_ASAP7_75t_L g293 ( .A1(n_253), .A2(n_294), .B(n_306), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_253), .B(n_325), .Y(n_324) );
INVx4_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_254), .Y(n_257) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g278 ( .A(n_255), .Y(n_278) );
INVx2_ASAP7_75t_L g314 ( .A(n_256), .Y(n_314) );
AND2x2_ASAP7_75t_L g415 ( .A(n_256), .B(n_292), .Y(n_415) );
AND2x2_ASAP7_75t_L g420 ( .A(n_256), .B(n_293), .Y(n_420) );
INVx1_ASAP7_75t_L g476 ( .A(n_256), .Y(n_476) );
OA21x2_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_258), .B(n_270), .Y(n_256) );
OA21x2_ASAP7_75t_L g327 ( .A1(n_257), .A2(n_328), .B(n_335), .Y(n_327) );
OA21x2_ASAP7_75t_L g336 ( .A1(n_257), .A2(n_337), .B(n_345), .Y(n_336) );
BUFx2_ASAP7_75t_L g280 ( .A(n_259), .Y(n_280) );
O2A1O1Ixp33_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_262), .B(n_263), .C(n_269), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_SL g281 ( .A1(n_262), .A2(n_269), .B(n_282), .C(n_283), .Y(n_281) );
O2A1O1Ixp33_ASAP7_75t_SL g329 ( .A1(n_262), .A2(n_269), .B(n_330), .C(n_331), .Y(n_329) );
O2A1O1Ixp33_ASAP7_75t_SL g338 ( .A1(n_262), .A2(n_269), .B(n_339), .C(n_340), .Y(n_338) );
O2A1O1Ixp33_ASAP7_75t_SL g371 ( .A1(n_262), .A2(n_269), .B(n_372), .C(n_373), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_264), .B(n_266), .Y(n_265) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g305 ( .A(n_269), .Y(n_305) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g385 ( .A(n_273), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_292), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_274), .B(n_348), .Y(n_347) );
BUFx3_ASAP7_75t_L g362 ( .A(n_274), .Y(n_362) );
OR2x2_ASAP7_75t_L g433 ( .A(n_274), .B(n_292), .Y(n_433) );
OR2x2_ASAP7_75t_L g494 ( .A(n_274), .B(n_401), .Y(n_494) );
OA21x2_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_279), .B(n_289), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AO21x2_ASAP7_75t_L g310 ( .A1(n_276), .A2(n_311), .B(n_312), .Y(n_310) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g311 ( .A(n_279), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_287), .B(n_333), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_287), .B(n_342), .Y(n_341) );
INVx4_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g300 ( .A(n_288), .Y(n_300) );
INVx1_ASAP7_75t_L g312 ( .A(n_289), .Y(n_312) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_291), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g313 ( .A(n_292), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g453 ( .A(n_292), .B(n_310), .Y(n_453) );
INVx2_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
BUFx2_ASAP7_75t_L g392 ( .A(n_293), .Y(n_392) );
O2A1O1Ixp33_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B(n_301), .C(n_302), .Y(n_297) );
O2A1O1Ixp5_ASAP7_75t_L g321 ( .A1(n_299), .A2(n_302), .B(n_322), .C(n_323), .Y(n_321) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_299), .Y(n_526) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g334 ( .A(n_304), .Y(n_334) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
AOI221xp5_ASAP7_75t_L g497 ( .A1(n_309), .A2(n_498), .B1(n_502), .B2(n_505), .C(n_506), .Y(n_497) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_313), .Y(n_309) );
INVx1_ASAP7_75t_SL g360 ( .A(n_310), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_310), .B(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g492 ( .A(n_310), .B(n_348), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_313), .B(n_362), .Y(n_484) );
AND2x2_ASAP7_75t_L g391 ( .A(n_314), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_SL g395 ( .A(n_315), .Y(n_395) );
NAND2xp5_ASAP7_75t_SL g431 ( .A(n_315), .B(n_401), .Y(n_431) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_326), .Y(n_315) );
AND2x2_ASAP7_75t_L g356 ( .A(n_316), .B(n_327), .Y(n_356) );
INVx4_ASAP7_75t_L g368 ( .A(n_316), .Y(n_368) );
BUFx3_ASAP7_75t_L g411 ( .A(n_316), .Y(n_411) );
AND3x2_ASAP7_75t_L g426 ( .A(n_316), .B(n_427), .C(n_428), .Y(n_426) );
AO21x2_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_318), .B(n_324), .Y(n_316) );
AND2x2_ASAP7_75t_L g508 ( .A(n_326), .B(n_422), .Y(n_508) );
AND2x2_ASAP7_75t_L g516 ( .A(n_326), .B(n_401), .Y(n_516) );
INVx1_ASAP7_75t_SL g521 ( .A(n_326), .Y(n_521) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_336), .Y(n_326) );
INVx1_ASAP7_75t_SL g379 ( .A(n_327), .Y(n_379) );
AND2x2_ASAP7_75t_L g402 ( .A(n_327), .B(n_368), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_327), .B(n_352), .Y(n_404) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_327), .Y(n_444) );
OR2x2_ASAP7_75t_L g449 ( .A(n_327), .B(n_368), .Y(n_449) );
INVx2_ASAP7_75t_L g354 ( .A(n_336), .Y(n_354) );
AND2x2_ASAP7_75t_L g389 ( .A(n_336), .B(n_369), .Y(n_389) );
OR2x2_ASAP7_75t_L g409 ( .A(n_336), .B(n_369), .Y(n_409) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_336), .Y(n_429) );
INVx3_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
AOI21xp33_ASAP7_75t_L g479 ( .A1(n_347), .A2(n_388), .B(n_480), .Y(n_479) );
AOI322xp5_ASAP7_75t_L g515 ( .A1(n_349), .A2(n_359), .A3(n_386), .B1(n_516), .B2(n_517), .C1(n_519), .C2(n_522), .Y(n_515) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_355), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_351), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_352), .B(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g378 ( .A(n_353), .B(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g446 ( .A(n_354), .B(n_368), .Y(n_446) );
AND2x2_ASAP7_75t_L g513 ( .A(n_354), .B(n_369), .Y(n_513) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g454 ( .A(n_356), .B(n_408), .Y(n_454) );
AOI31xp33_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_361), .A3(n_364), .B(n_365), .Y(n_357) );
AND2x2_ASAP7_75t_L g413 ( .A(n_359), .B(n_391), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_359), .B(n_383), .Y(n_495) );
AND2x2_ASAP7_75t_L g514 ( .A(n_359), .B(n_419), .Y(n_514) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_362), .B(n_391), .Y(n_403) );
NAND2x1p5_ASAP7_75t_L g437 ( .A(n_362), .B(n_420), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g440 ( .A(n_362), .B(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_362), .B(n_504), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_363), .B(n_420), .Y(n_452) );
INVx1_ASAP7_75t_L g496 ( .A(n_363), .Y(n_496) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_378), .Y(n_366) );
INVxp67_ASAP7_75t_L g448 ( .A(n_367), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_368), .B(n_379), .Y(n_384) );
INVx1_ASAP7_75t_L g490 ( .A(n_368), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_368), .B(n_467), .Y(n_501) );
BUFx3_ASAP7_75t_L g401 ( .A(n_369), .Y(n_401) );
AND2x2_ASAP7_75t_L g427 ( .A(n_369), .B(n_379), .Y(n_427) );
INVx2_ASAP7_75t_L g467 ( .A(n_369), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_378), .B(n_500), .Y(n_499) );
AOI211xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_385), .B(n_387), .C(n_396), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AOI21xp33_ASAP7_75t_L g430 ( .A1(n_382), .A2(n_431), .B(n_432), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_383), .B(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_383), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g463 ( .A(n_384), .B(n_409), .Y(n_463) );
INVx3_ASAP7_75t_L g394 ( .A(n_386), .Y(n_394) );
OAI22xp5_ASAP7_75t_SL g387 ( .A1(n_388), .A2(n_390), .B1(n_393), .B2(n_395), .Y(n_387) );
OAI21xp5_ASAP7_75t_SL g412 ( .A1(n_389), .A2(n_413), .B(n_414), .Y(n_412) );
AND2x2_ASAP7_75t_L g438 ( .A(n_389), .B(n_402), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_389), .B(n_490), .Y(n_489) );
INVxp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g393 ( .A(n_392), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g462 ( .A(n_392), .Y(n_462) );
OAI21xp5_ASAP7_75t_SL g406 ( .A1(n_393), .A2(n_407), .B(n_412), .Y(n_406) );
OAI22xp33_ASAP7_75t_SL g396 ( .A1(n_397), .A2(n_399), .B1(n_403), .B2(n_404), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_398), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
INVx1_ASAP7_75t_L g422 ( .A(n_401), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_401), .B(n_444), .Y(n_443) );
NOR3xp33_ASAP7_75t_L g405 ( .A(n_406), .B(n_417), .C(n_430), .Y(n_405) );
OAI22xp5_ASAP7_75t_SL g472 ( .A1(n_407), .A2(n_473), .B1(n_477), .B2(n_478), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g407 ( .A(n_408), .B(n_410), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g477 ( .A(n_409), .B(n_410), .Y(n_477) );
AND2x2_ASAP7_75t_L g485 ( .A(n_410), .B(n_466), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g410 ( .A(n_411), .Y(n_410) );
O2A1O1Ixp33_ASAP7_75t_SL g493 ( .A1(n_411), .A2(n_494), .B(n_495), .C(n_496), .Y(n_493) );
OR2x2_ASAP7_75t_L g520 ( .A(n_411), .B(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
OAI21xp33_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_421), .B(n_423), .Y(n_417) );
INVx1_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
O2A1O1Ixp33_ASAP7_75t_L g455 ( .A1(n_419), .A2(n_456), .B(n_457), .C(n_460), .Y(n_455) );
OAI21xp33_ASAP7_75t_SL g423 ( .A1(n_424), .A2(n_425), .B(n_426), .Y(n_423) );
AND2x2_ASAP7_75t_L g488 ( .A(n_427), .B(n_446), .Y(n_488) );
INVxp67_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g466 ( .A(n_429), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g471 ( .A(n_431), .Y(n_471) );
NAND3xp33_ASAP7_75t_SL g434 ( .A(n_435), .B(n_455), .C(n_468), .Y(n_434) );
AOI211xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_438), .B(n_439), .C(n_447), .Y(n_435) );
INVx1_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_440), .B(n_442), .Y(n_439) );
INVx1_ASAP7_75t_L g505 ( .A(n_442), .Y(n_505) );
OR2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_445), .Y(n_442) );
INVx1_ASAP7_75t_L g465 ( .A(n_444), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_444), .B(n_513), .Y(n_512) );
INVxp67_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_449), .B(n_450), .C(n_451), .Y(n_447) );
INVx2_ASAP7_75t_SL g459 ( .A(n_449), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_450), .A2(n_461), .B1(n_463), .B2(n_464), .Y(n_460) );
OAI21xp33_ASAP7_75t_SL g451 ( .A1(n_452), .A2(n_453), .B(n_454), .Y(n_451) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
AOI211xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_471), .B(n_472), .C(n_479), .Y(n_468) );
INVx1_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
INVxp33_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g522 ( .A(n_476), .Y(n_522) );
NAND4xp25_ASAP7_75t_L g481 ( .A(n_482), .B(n_497), .C(n_510), .D(n_515), .Y(n_481) );
AOI211xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_485), .B(n_486), .C(n_493), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_489), .B(n_491), .Y(n_486) );
AOI21xp33_ASAP7_75t_L g506 ( .A1(n_487), .A2(n_507), .B(n_509), .Y(n_506) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_494), .B(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_514), .Y(n_510) );
INVxp67_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
CKINVDCx16_ASAP7_75t_R g523 ( .A(n_524), .Y(n_523) );
OAI322xp33_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_530), .A3(n_534), .B1(n_536), .B2(n_539), .C1(n_540), .C2(n_541), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_531), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_532), .Y(n_531) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_537), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_542), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_543), .Y(n_542) );
endmodule