module fake_netlist_5_1227_n_2781 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_74, n_515, n_57, n_353, n_351, n_367, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_4, n_378, n_551, n_17, n_581, n_382, n_554, n_254, n_33, n_23, n_583, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_559, n_275, n_252, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_584, n_145, n_48, n_521, n_50, n_337, n_430, n_313, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_502, n_239, n_466, n_420, n_489, n_55, n_49, n_310, n_54, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_480, n_237, n_425, n_513, n_407, n_527, n_180, n_560, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_572, n_113, n_246, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_541, n_391, n_434, n_539, n_175, n_538, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_2781);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_382;
input n_554;
input n_254;
input n_33;
input n_23;
input n_583;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_559;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_584;
input n_145;
input n_48;
input n_521;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_49;
input n_310;
input n_54;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_480;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_560;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_541;
input n_391;
input n_434;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_2781;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_611;
wire n_2756;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_785;
wire n_2617;
wire n_2200;
wire n_1161;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_1007;
wire n_2369;
wire n_1528;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_956;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_800;
wire n_1347;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_1118;
wire n_755;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_1728;
wire n_1107;
wire n_2076;
wire n_2031;
wire n_2482;
wire n_2677;
wire n_1230;
wire n_668;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_2770;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1016;
wire n_1243;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_2761;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_2515;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_2715;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_2672;
wire n_775;
wire n_2651;
wire n_600;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_1414;
wire n_1216;
wire n_2693;
wire n_1040;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_926;
wire n_2249;
wire n_2180;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_1070;
wire n_777;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_1561;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_2300;
wire n_1796;
wire n_2551;
wire n_1473;
wire n_680;
wire n_1587;
wire n_2682;
wire n_901;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_1672;
wire n_2506;
wire n_675;
wire n_2699;
wire n_888;
wire n_1880;
wire n_2769;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_2615;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_2753;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_2738;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_1585;
wire n_2712;
wire n_2684;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_2713;
wire n_2644;
wire n_2700;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_736;
wire n_892;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_1581;
wire n_1463;
wire n_2100;
wire n_593;
wire n_2258;
wire n_748;
wire n_1058;
wire n_1667;
wire n_838;
wire n_1053;
wire n_1224;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2757;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_857;
wire n_832;
wire n_2305;
wire n_2636;
wire n_2450;
wire n_1319;
wire n_2379;
wire n_2616;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2331;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_2762;
wire n_1276;
wire n_702;
wire n_2548;
wire n_822;
wire n_1412;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_1038;
wire n_1369;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_2698;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_2626;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_868;
wire n_2454;
wire n_639;
wire n_914;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2690;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_2621;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_2671;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_2518;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_1829;
wire n_1464;
wire n_649;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_2631;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_604;
wire n_2007;
wire n_949;
wire n_2539;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_2736;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_2718;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_2577;
wire n_1760;
wire n_936;
wire n_1500;
wire n_1090;
wire n_757;
wire n_2342;
wire n_633;
wire n_1832;
wire n_1851;
wire n_999;
wire n_758;
wire n_2046;
wire n_2741;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_1964;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_1586;
wire n_959;
wire n_2459;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_1017;
wire n_2481;
wire n_2171;
wire n_978;
wire n_2768;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_2093;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2320;
wire n_2038;
wire n_2339;
wire n_2473;
wire n_2137;
wire n_603;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_2540;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_2168;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_614;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_2565;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2729;
wire n_2418;
wire n_829;
wire n_2519;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_700;
wire n_1237;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_2277;
wire n_761;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2604;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_2681;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_1913;
wire n_1823;
wire n_874;
wire n_2464;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_860;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_628;
wire n_1849;
wire n_2410;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_2645;
wire n_2467;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_1552;
wire n_2508;
wire n_602;
wire n_2593;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_623;
wire n_2088;
wire n_824;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_2658;
wire n_1717;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_1821;
wire n_1381;
wire n_2555;
wire n_2662;
wire n_2740;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2534;
wire n_2092;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_2647;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_2465;
wire n_2650;
wire n_912;
wire n_968;
wire n_619;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_2333;
wire n_885;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_1050;
wire n_841;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_2760;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_2637;
wire n_690;
wire n_1974;
wire n_2463;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2701;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_753;
wire n_621;
wire n_2475;
wire n_2733;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2556;
wire n_2269;
wire n_2732;
wire n_2309;
wire n_2415;
wire n_2646;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_1312;
wire n_1439;
wire n_804;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_2755;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_2533;
wire n_618;
wire n_896;
wire n_2310;
wire n_2780;
wire n_2287;
wire n_2291;
wire n_2596;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_2318;
wire n_833;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2749;
wire n_2043;
wire n_1940;
wire n_814;
wire n_2707;
wire n_2751;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_2758;
wire n_669;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_2471;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_783;
wire n_1928;
wire n_1848;
wire n_2126;
wire n_1188;
wire n_2588;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_2600;
wire n_849;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_2282;
wire n_2371;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_749;
wire n_1895;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_2638;
wire n_866;
wire n_969;
wire n_1401;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_2653;
wire n_836;
wire n_990;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_1465;
wire n_778;
wire n_1122;
wire n_2608;
wire n_2657;
wire n_770;
wire n_1375;
wire n_2494;
wire n_2649;
wire n_1102;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_2633;
wire n_1441;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_1174;
wire n_2431;
wire n_2558;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_726;
wire n_982;
wire n_2575;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_2766;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2745;
wire n_2117;
wire n_2722;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1514;
wire n_1335;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2437;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_2634;
wire n_910;
wire n_2232;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_2547;
wire n_708;
wire n_1812;
wire n_735;
wire n_2501;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_2121;
wire n_1803;
wire n_2665;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_1067;
wire n_1720;
wire n_2401;
wire n_2003;
wire n_766;
wire n_1457;
wire n_2692;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_2754;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_2213;
wire n_2023;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_855;
wire n_1178;
wire n_1461;
wire n_2697;
wire n_850;
wire n_684;
wire n_2421;
wire n_2286;
wire n_664;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_605;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_2363;
wire n_2430;
wire n_916;
wire n_1081;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_1235;
wire n_980;
wire n_703;
wire n_1115;
wire n_698;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2601;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_2686;
wire n_2528;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2773;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_2687;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_2654;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_825;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_812;
wire n_2104;
wire n_2748;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_2717;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_1675;
wire n_1924;
wire n_2573;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_1745;
wire n_2735;
wire n_769;
wire n_2497;
wire n_2006;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_2726;
wire n_2774;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2172;
wire n_1973;
wire n_1083;
wire n_786;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2456;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_771;
wire n_2778;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_2451;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_930;
wire n_1873;
wire n_1411;
wire n_1962;
wire n_622;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_682;
wire n_1567;
wire n_2567;
wire n_1247;
wire n_2709;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_2531;
wire n_1589;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2591;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_1546;
wire n_595;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_2112;
wire n_1739;
wire n_616;
wire n_2278;
wire n_2594;
wire n_2394;
wire n_1914;
wire n_2335;
wire n_2135;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2569;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2734;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1956;
wire n_1936;
wire n_1642;
wire n_2279;
wire n_2655;
wire n_2027;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_2525;
wire n_2513;
wire n_2695;
wire n_1764;
wire n_712;
wire n_2414;
wire n_1583;
wire n_2426;
wire n_1042;
wire n_1402;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2708;
wire n_2113;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_2044;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2689;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_1693;
wire n_2599;
wire n_713;
wire n_2704;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_2524;
wire n_1271;
wire n_1542;
wire n_1251;
wire n_2728;
wire n_2268;

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_418),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_243),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_410),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_408),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_546),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_311),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_89),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_439),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_195),
.Y(n_595)
);

INVxp67_ASAP7_75t_SL g596 ( 
.A(n_123),
.Y(n_596)
);

INVx1_ASAP7_75t_SL g597 ( 
.A(n_517),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_46),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g599 ( 
.A(n_473),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_255),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_338),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_182),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_231),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_420),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_492),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_320),
.Y(n_606)
);

INVx1_ASAP7_75t_SL g607 ( 
.A(n_422),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_371),
.Y(n_608)
);

INVx4_ASAP7_75t_R g609 ( 
.A(n_464),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_468),
.Y(n_610)
);

BUFx2_ASAP7_75t_L g611 ( 
.A(n_116),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_477),
.Y(n_612)
);

INVxp67_ASAP7_75t_L g613 ( 
.A(n_436),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_561),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_255),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_442),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_174),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_510),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_479),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_70),
.Y(n_620)
);

INVx1_ASAP7_75t_SL g621 ( 
.A(n_329),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_505),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_483),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_12),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_266),
.Y(n_625)
);

CKINVDCx16_ASAP7_75t_R g626 ( 
.A(n_441),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_565),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_474),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_61),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_324),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_56),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_469),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_138),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_471),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g635 ( 
.A(n_215),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_51),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_558),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_93),
.Y(n_638)
);

HB1xp67_ASAP7_75t_L g639 ( 
.A(n_278),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_376),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_476),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_95),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_205),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_182),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_503),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_107),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_499),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_560),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_340),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_554),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_211),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_163),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_10),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_468),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_125),
.Y(n_655)
);

INVx1_ASAP7_75t_SL g656 ( 
.A(n_557),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_434),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_344),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_513),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_439),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_563),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_73),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_241),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_167),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_346),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_309),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_585),
.Y(n_667)
);

INVx1_ASAP7_75t_SL g668 ( 
.A(n_519),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_120),
.Y(n_669)
);

BUFx10_ASAP7_75t_L g670 ( 
.A(n_151),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_74),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_167),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_116),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_183),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_509),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_95),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_88),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_528),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_559),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_136),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_272),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_331),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_134),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_289),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_448),
.Y(n_685)
);

CKINVDCx14_ASAP7_75t_R g686 ( 
.A(n_579),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_160),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_44),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_586),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_108),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_580),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_339),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_2),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_48),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_110),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_120),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_382),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_183),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_581),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_325),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_376),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_115),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_470),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_62),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_436),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_284),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_314),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_368),
.Y(n_708)
);

CKINVDCx20_ASAP7_75t_R g709 ( 
.A(n_257),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_455),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_539),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_205),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_536),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_107),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_357),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_408),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_440),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_404),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_571),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_91),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_92),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_472),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_50),
.Y(n_723)
);

BUFx10_ASAP7_75t_L g724 ( 
.A(n_584),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_100),
.Y(n_725)
);

BUFx10_ASAP7_75t_L g726 ( 
.A(n_115),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_289),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_80),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_288),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_9),
.Y(n_730)
);

CKINVDCx14_ASAP7_75t_R g731 ( 
.A(n_252),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_473),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_556),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_564),
.Y(n_734)
);

BUFx10_ASAP7_75t_L g735 ( 
.A(n_485),
.Y(n_735)
);

INVx1_ASAP7_75t_SL g736 ( 
.A(n_420),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_578),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_283),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_78),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_61),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_514),
.Y(n_741)
);

BUFx10_ASAP7_75t_L g742 ( 
.A(n_541),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_38),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_568),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_498),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_467),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_577),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_159),
.Y(n_748)
);

CKINVDCx16_ASAP7_75t_R g749 ( 
.A(n_301),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_394),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_555),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_339),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_493),
.Y(n_753)
);

BUFx10_ASAP7_75t_L g754 ( 
.A(n_573),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_472),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_45),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_574),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_26),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_570),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_475),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_457),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_298),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_207),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_13),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_412),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_520),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_441),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_500),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_490),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_478),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_128),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_93),
.Y(n_772)
);

BUFx10_ASAP7_75t_L g773 ( 
.A(n_575),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_334),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_535),
.Y(n_775)
);

BUFx8_ASAP7_75t_SL g776 ( 
.A(n_474),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_426),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_75),
.Y(n_778)
);

CKINVDCx20_ASAP7_75t_R g779 ( 
.A(n_567),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_168),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_211),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_254),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_258),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_346),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_31),
.Y(n_785)
);

BUFx10_ASAP7_75t_L g786 ( 
.A(n_330),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_576),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_495),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_583),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_227),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_569),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_457),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_64),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_356),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_486),
.Y(n_795)
);

INVx1_ASAP7_75t_SL g796 ( 
.A(n_34),
.Y(n_796)
);

INVxp33_ASAP7_75t_R g797 ( 
.A(n_236),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_350),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_463),
.Y(n_799)
);

INVxp67_ASAP7_75t_SL g800 ( 
.A(n_175),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_231),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_71),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_477),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_469),
.Y(n_804)
);

BUFx10_ASAP7_75t_L g805 ( 
.A(n_213),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_566),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_15),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_147),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_186),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_572),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_143),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_342),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_471),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_64),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_57),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_148),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_55),
.Y(n_817)
);

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_100),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_75),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_131),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_371),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_25),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_54),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_582),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_562),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_321),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_28),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_237),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_300),
.Y(n_829)
);

BUFx2_ASAP7_75t_L g830 ( 
.A(n_476),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_217),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_479),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_275),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_776),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_592),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_588),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_592),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_604),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_604),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_624),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_624),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_776),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_763),
.Y(n_843)
);

CKINVDCx20_ASAP7_75t_R g844 ( 
.A(n_612),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_636),
.Y(n_845)
);

INVx1_ASAP7_75t_SL g846 ( 
.A(n_611),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_763),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_636),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_731),
.Y(n_849)
);

INVxp67_ASAP7_75t_SL g850 ( 
.A(n_789),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_778),
.Y(n_851)
);

BUFx2_ASAP7_75t_L g852 ( 
.A(n_635),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_778),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_731),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_626),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_766),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_749),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_636),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_636),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_655),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_724),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_655),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_655),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_724),
.Y(n_864)
);

INVxp33_ASAP7_75t_L g865 ( 
.A(n_639),
.Y(n_865)
);

BUFx3_ASAP7_75t_L g866 ( 
.A(n_724),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_655),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_690),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_735),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_690),
.Y(n_870)
);

BUFx10_ASAP7_75t_L g871 ( 
.A(n_690),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_690),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_720),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_720),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_720),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_720),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_729),
.Y(n_877)
);

CKINVDCx16_ASAP7_75t_R g878 ( 
.A(n_686),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_729),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_729),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_729),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_813),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_587),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_813),
.Y(n_884)
);

CKINVDCx14_ASAP7_75t_R g885 ( 
.A(n_686),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_589),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_813),
.Y(n_887)
);

INVxp67_ASAP7_75t_SL g888 ( 
.A(n_675),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_813),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_590),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_594),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_593),
.Y(n_892)
);

CKINVDCx20_ASAP7_75t_R g893 ( 
.A(n_612),
.Y(n_893)
);

INVxp67_ASAP7_75t_SL g894 ( 
.A(n_605),
.Y(n_894)
);

INVx1_ASAP7_75t_SL g895 ( 
.A(n_830),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_601),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_602),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_598),
.Y(n_898)
);

CKINVDCx20_ASAP7_75t_R g899 ( 
.A(n_681),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_591),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_603),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_644),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_766),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_608),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_600),
.Y(n_905)
);

INVxp33_ASAP7_75t_SL g906 ( 
.A(n_606),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_620),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_644),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_625),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_629),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_633),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_634),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_642),
.Y(n_913)
);

CKINVDCx16_ASAP7_75t_R g914 ( 
.A(n_650),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_652),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_657),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_663),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_671),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_610),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_672),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_680),
.Y(n_921)
);

CKINVDCx20_ASAP7_75t_R g922 ( 
.A(n_681),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_682),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_684),
.Y(n_924)
);

OR2x2_ASAP7_75t_L g925 ( 
.A(n_595),
.B(n_0),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_766),
.Y(n_926)
);

CKINVDCx20_ASAP7_75t_R g927 ( 
.A(n_692),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_651),
.Y(n_928)
);

INVxp67_ASAP7_75t_SL g929 ( 
.A(n_614),
.Y(n_929)
);

INVxp67_ASAP7_75t_L g930 ( 
.A(n_670),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_615),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_685),
.Y(n_932)
);

CKINVDCx20_ASAP7_75t_R g933 ( 
.A(n_692),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_688),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_616),
.Y(n_935)
);

INVxp33_ASAP7_75t_L g936 ( 
.A(n_865),
.Y(n_936)
);

CKINVDCx20_ASAP7_75t_R g937 ( 
.A(n_844),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_859),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_860),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_900),
.Y(n_940)
);

CKINVDCx20_ASAP7_75t_R g941 ( 
.A(n_844),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_883),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_883),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_862),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_886),
.Y(n_945)
);

CKINVDCx16_ASAP7_75t_R g946 ( 
.A(n_914),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_855),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_863),
.Y(n_948)
);

CKINVDCx16_ASAP7_75t_R g949 ( 
.A(n_878),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_867),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_868),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_870),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_886),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_874),
.Y(n_954)
);

INVxp67_ASAP7_75t_SL g955 ( 
.A(n_856),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_875),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_877),
.Y(n_957)
);

CKINVDCx20_ASAP7_75t_R g958 ( 
.A(n_893),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_888),
.B(n_597),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_891),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_879),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_880),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_881),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_845),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_849),
.B(n_656),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_849),
.B(n_668),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_891),
.Y(n_967)
);

CKINVDCx20_ASAP7_75t_R g968 ( 
.A(n_893),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_882),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_898),
.Y(n_970)
);

CKINVDCx20_ASAP7_75t_R g971 ( 
.A(n_899),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_854),
.B(n_734),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_884),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_887),
.Y(n_974)
);

CKINVDCx20_ASAP7_75t_R g975 ( 
.A(n_899),
.Y(n_975)
);

CKINVDCx20_ASAP7_75t_R g976 ( 
.A(n_922),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_889),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_898),
.Y(n_978)
);

INVxp67_ASAP7_75t_L g979 ( 
.A(n_861),
.Y(n_979)
);

XNOR2xp5_ASAP7_75t_L g980 ( 
.A(n_922),
.B(n_927),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_845),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_854),
.B(n_734),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_885),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_885),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_848),
.Y(n_985)
);

CKINVDCx20_ASAP7_75t_R g986 ( 
.A(n_927),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_848),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_858),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_905),
.Y(n_989)
);

NOR2xp67_ASAP7_75t_L g990 ( 
.A(n_905),
.B(n_637),
.Y(n_990)
);

CKINVDCx20_ASAP7_75t_R g991 ( 
.A(n_933),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_858),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_873),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_873),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_876),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_876),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_894),
.B(n_689),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_872),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_856),
.Y(n_999)
);

CKINVDCx20_ASAP7_75t_R g1000 ( 
.A(n_933),
.Y(n_1000)
);

CKINVDCx20_ASAP7_75t_R g1001 ( 
.A(n_834),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_959),
.A2(n_850),
.B1(n_906),
.B2(n_925),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_955),
.B(n_929),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_990),
.B(n_872),
.Y(n_1004)
);

INVxp67_ASAP7_75t_L g1005 ( 
.A(n_972),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_999),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_999),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_964),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_999),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_983),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_964),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_998),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_965),
.A2(n_857),
.B1(n_855),
.B2(n_919),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_936),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_966),
.B(n_872),
.Y(n_1015)
);

BUFx10_ASAP7_75t_L g1016 ( 
.A(n_982),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_981),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_983),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_985),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_987),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_938),
.Y(n_1021)
);

INVx2_ASAP7_75t_SL g1022 ( 
.A(n_947),
.Y(n_1022)
);

BUFx2_ASAP7_75t_L g1023 ( 
.A(n_979),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_997),
.B(n_902),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_939),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_988),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_944),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_948),
.B(n_950),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_951),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_992),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_952),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_984),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_954),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_956),
.B(n_902),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_942),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_957),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_961),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_962),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_963),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_969),
.B(n_919),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_973),
.B(n_906),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_974),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_977),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_984),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_993),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_994),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_995),
.B(n_908),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_949),
.B(n_846),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_946),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_996),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_940),
.B(n_895),
.Y(n_1051)
);

HB1xp67_ASAP7_75t_L g1052 ( 
.A(n_943),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_945),
.A2(n_857),
.B1(n_935),
.B2(n_931),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_953),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_960),
.A2(n_836),
.B1(n_935),
.B2(n_931),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_967),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_937),
.Y(n_1057)
);

XNOR2x2_ASAP7_75t_R g1058 ( 
.A(n_980),
.B(n_797),
.Y(n_1058)
);

INVx3_ASAP7_75t_L g1059 ( 
.A(n_970),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_978),
.Y(n_1060)
);

AND2x6_ASAP7_75t_L g1061 ( 
.A(n_989),
.B(n_689),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_1001),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1001),
.B(n_926),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_937),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_941),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_1000),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1000),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_941),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_991),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_958),
.B(n_908),
.Y(n_1070)
);

BUFx8_ASAP7_75t_L g1071 ( 
.A(n_958),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_968),
.B(n_928),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_968),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_971),
.B(n_928),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_991),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_971),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_975),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_975),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_976),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_976),
.B(n_861),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_986),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_986),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_999),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_983),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_964),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_998),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_998),
.Y(n_1087)
);

AND2x2_ASAP7_75t_SL g1088 ( 
.A(n_959),
.B(n_766),
.Y(n_1088)
);

INVx4_ASAP7_75t_L g1089 ( 
.A(n_999),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_999),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_936),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1028),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_1089),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1028),
.Y(n_1094)
);

INVxp67_ASAP7_75t_L g1095 ( 
.A(n_1014),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1088),
.B(n_647),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1028),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1021),
.Y(n_1098)
);

NAND2xp33_ASAP7_75t_SL g1099 ( 
.A(n_1002),
.B(n_650),
.Y(n_1099)
);

INVx3_ASAP7_75t_L g1100 ( 
.A(n_1089),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1088),
.B(n_667),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1008),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_1089),
.Y(n_1103)
);

INVx1_ASAP7_75t_SL g1104 ( 
.A(n_1051),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1008),
.Y(n_1105)
);

INVx1_ASAP7_75t_SL g1106 ( 
.A(n_1091),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_1023),
.B(n_864),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_1005),
.A2(n_779),
.B1(n_691),
.B2(n_699),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1025),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_1006),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1027),
.Y(n_1111)
);

BUFx3_ASAP7_75t_L g1112 ( 
.A(n_1056),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1031),
.Y(n_1113)
);

INVx1_ASAP7_75t_SL g1114 ( 
.A(n_1048),
.Y(n_1114)
);

OA21x2_ASAP7_75t_L g1115 ( 
.A1(n_1011),
.A2(n_719),
.B(n_678),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_1029),
.B(n_795),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1024),
.B(n_733),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_SL g1118 ( 
.A1(n_1079),
.A2(n_709),
.B1(n_758),
.B2(n_696),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_1029),
.B(n_795),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1024),
.B(n_751),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_1006),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1085),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_1057),
.Y(n_1123)
);

AOI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1061),
.A2(n_779),
.B1(n_622),
.B2(n_623),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1085),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1033),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1047),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1036),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1037),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1038),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_SL g1131 ( 
.A(n_1062),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_1034),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1039),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1047),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1034),
.Y(n_1135)
);

INVx1_ASAP7_75t_SL g1136 ( 
.A(n_1074),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1034),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_SL g1138 ( 
.A1(n_1079),
.A2(n_709),
.B1(n_758),
.B2(n_696),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_1006),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1017),
.Y(n_1140)
);

INVxp67_ASAP7_75t_L g1141 ( 
.A(n_1074),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1017),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1019),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1019),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1020),
.Y(n_1145)
);

INVxp67_ASAP7_75t_L g1146 ( 
.A(n_1041),
.Y(n_1146)
);

AND2x6_ASAP7_75t_L g1147 ( 
.A(n_1054),
.B(n_768),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_1012),
.B(n_769),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1020),
.Y(n_1149)
);

AOI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1061),
.A2(n_627),
.B1(n_645),
.B2(n_618),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_1006),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_1007),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_SL g1153 ( 
.A1(n_1081),
.A2(n_818),
.B1(n_822),
.B2(n_771),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1026),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1022),
.B(n_1059),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1026),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1030),
.Y(n_1157)
);

INVxp67_ASAP7_75t_L g1158 ( 
.A(n_1041),
.Y(n_1158)
);

INVx4_ASAP7_75t_L g1159 ( 
.A(n_1007),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_SL g1160 ( 
.A(n_1062),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1030),
.Y(n_1161)
);

AND2x6_ASAP7_75t_L g1162 ( 
.A(n_1054),
.B(n_810),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1045),
.Y(n_1163)
);

XOR2x2_ASAP7_75t_L g1164 ( 
.A(n_1058),
.B(n_852),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_1070),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1050),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1086),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_1029),
.B(n_795),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1087),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1003),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1004),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_SL g1172 ( 
.A1(n_1081),
.A2(n_818),
.B1(n_822),
.B2(n_771),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_L g1173 ( 
.A(n_1070),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1029),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_SL g1175 ( 
.A1(n_1064),
.A2(n_826),
.B1(n_842),
.B2(n_834),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1042),
.Y(n_1176)
);

INVx8_ASAP7_75t_L g1177 ( 
.A(n_1061),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1015),
.B(n_824),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1022),
.B(n_864),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1042),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1061),
.B(n_825),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_1007),
.Y(n_1182)
);

HB1xp67_ASAP7_75t_L g1183 ( 
.A(n_1070),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1042),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1042),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1040),
.A2(n_837),
.B(n_835),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1061),
.B(n_866),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1043),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_1007),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1043),
.Y(n_1190)
);

INVxp67_ASAP7_75t_L g1191 ( 
.A(n_1080),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1046),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1043),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1046),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1043),
.Y(n_1195)
);

INVx3_ASAP7_75t_L g1196 ( 
.A(n_1009),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_1009),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1061),
.B(n_1009),
.Y(n_1198)
);

INVx1_ASAP7_75t_SL g1199 ( 
.A(n_1082),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1059),
.B(n_866),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1046),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1009),
.B(n_869),
.Y(n_1202)
);

INVx5_ASAP7_75t_L g1203 ( 
.A(n_1083),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_1072),
.B(n_890),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1046),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1083),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1083),
.B(n_1090),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_1072),
.B(n_892),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1059),
.B(n_869),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1072),
.Y(n_1210)
);

AOI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1055),
.A2(n_1013),
.B1(n_1053),
.B2(n_1063),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1083),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_SL g1213 ( 
.A(n_1016),
.B(n_795),
.Y(n_1213)
);

BUFx2_ASAP7_75t_L g1214 ( 
.A(n_1082),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1090),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1090),
.Y(n_1216)
);

OA21x2_ASAP7_75t_L g1217 ( 
.A1(n_1060),
.A2(n_839),
.B(n_838),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1090),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1016),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_1016),
.Y(n_1220)
);

INVx1_ASAP7_75t_SL g1221 ( 
.A(n_1049),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_1056),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1056),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1056),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1035),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_SL g1226 ( 
.A(n_1062),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1084),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1052),
.B(n_865),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1080),
.Y(n_1229)
);

INVx3_ASAP7_75t_L g1230 ( 
.A(n_1132),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1104),
.B(n_1066),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1135),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1137),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1102),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_1123),
.Y(n_1235)
);

AND2x6_ASAP7_75t_L g1236 ( 
.A(n_1170),
.B(n_1065),
.Y(n_1236)
);

AND2x6_ASAP7_75t_L g1237 ( 
.A(n_1112),
.B(n_1065),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1179),
.B(n_1066),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_SL g1239 ( 
.A(n_1155),
.B(n_1010),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1099),
.A2(n_746),
.B1(n_595),
.B2(n_683),
.Y(n_1240)
);

OR2x2_ASAP7_75t_SL g1241 ( 
.A(n_1227),
.B(n_1058),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1132),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1102),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1140),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1105),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1105),
.Y(n_1246)
);

INVx1_ASAP7_75t_SL g1247 ( 
.A(n_1114),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1140),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1142),
.Y(n_1249)
);

AND2x4_ASAP7_75t_L g1250 ( 
.A(n_1112),
.B(n_1065),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1146),
.B(n_1158),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1146),
.B(n_1068),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1142),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1214),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_R g1255 ( 
.A(n_1220),
.B(n_1049),
.Y(n_1255)
);

AND2x6_ASAP7_75t_L g1256 ( 
.A(n_1093),
.B(n_1068),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1122),
.Y(n_1257)
);

AND2x6_ASAP7_75t_L g1258 ( 
.A(n_1093),
.B(n_1069),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1206),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1110),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1206),
.Y(n_1261)
);

INVx1_ASAP7_75t_SL g1262 ( 
.A(n_1106),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1099),
.A2(n_746),
.B1(n_651),
.B2(n_683),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1127),
.B(n_596),
.Y(n_1264)
);

AO22x2_ASAP7_75t_L g1265 ( 
.A1(n_1108),
.A2(n_1069),
.B1(n_1073),
.B2(n_1067),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1125),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1144),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1127),
.B(n_800),
.Y(n_1268)
);

INVx2_ASAP7_75t_SL g1269 ( 
.A(n_1107),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_1110),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1144),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1145),
.Y(n_1272)
);

INVx1_ASAP7_75t_SL g1273 ( 
.A(n_1136),
.Y(n_1273)
);

OAI22x1_ASAP7_75t_L g1274 ( 
.A1(n_1211),
.A2(n_1158),
.B1(n_1073),
.B2(n_1229),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1125),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1191),
.B(n_1075),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_1222),
.B(n_1010),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1145),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1149),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_1141),
.Y(n_1280)
);

INVx6_ASAP7_75t_L g1281 ( 
.A(n_1227),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1149),
.Y(n_1282)
);

INVx1_ASAP7_75t_SL g1283 ( 
.A(n_1228),
.Y(n_1283)
);

BUFx6f_ASAP7_75t_L g1284 ( 
.A(n_1110),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1191),
.B(n_1076),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1117),
.B(n_648),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1222),
.B(n_1018),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1141),
.B(n_1077),
.Y(n_1288)
);

AND2x4_ASAP7_75t_L g1289 ( 
.A(n_1222),
.B(n_1062),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1156),
.Y(n_1290)
);

BUFx3_ASAP7_75t_L g1291 ( 
.A(n_1227),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1156),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1161),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1161),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1143),
.Y(n_1295)
);

INVx4_ASAP7_75t_L g1296 ( 
.A(n_1110),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1154),
.Y(n_1297)
);

INVxp67_ASAP7_75t_SL g1298 ( 
.A(n_1093),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1120),
.B(n_659),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1157),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1163),
.Y(n_1301)
);

BUFx2_ASAP7_75t_L g1302 ( 
.A(n_1165),
.Y(n_1302)
);

AND2x2_ASAP7_75t_SL g1303 ( 
.A(n_1227),
.B(n_1078),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1095),
.B(n_1018),
.Y(n_1304)
);

AO21x2_ASAP7_75t_L g1305 ( 
.A1(n_1181),
.A2(n_697),
.B(n_695),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1200),
.B(n_1032),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1209),
.B(n_1095),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1171),
.B(n_661),
.Y(n_1308)
);

AND2x4_ASAP7_75t_L g1309 ( 
.A(n_1223),
.B(n_896),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1220),
.B(n_1032),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1098),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1163),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1096),
.A2(n_826),
.B1(n_762),
.B2(n_811),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_1131),
.Y(n_1314)
);

INVx2_ASAP7_75t_SL g1315 ( 
.A(n_1204),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1109),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1100),
.B(n_679),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1167),
.Y(n_1318)
);

INVx4_ASAP7_75t_L g1319 ( 
.A(n_1121),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_1121),
.Y(n_1320)
);

NAND3xp33_ASAP7_75t_L g1321 ( 
.A(n_1101),
.B(n_1178),
.C(n_1113),
.Y(n_1321)
);

BUFx6f_ASAP7_75t_L g1322 ( 
.A(n_1121),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1121),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1167),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1204),
.B(n_1044),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1204),
.Y(n_1326)
);

BUFx6f_ASAP7_75t_L g1327 ( 
.A(n_1182),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1111),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1169),
.Y(n_1329)
);

INVx1_ASAP7_75t_SL g1330 ( 
.A(n_1199),
.Y(n_1330)
);

INVx1_ASAP7_75t_SL g1331 ( 
.A(n_1165),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1169),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1126),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1224),
.B(n_897),
.Y(n_1334)
);

AND2x6_ASAP7_75t_L g1335 ( 
.A(n_1198),
.B(n_1092),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1128),
.Y(n_1336)
);

AND2x6_ASAP7_75t_L g1337 ( 
.A(n_1094),
.B(n_762),
.Y(n_1337)
);

INVx3_ASAP7_75t_L g1338 ( 
.A(n_1212),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1129),
.Y(n_1339)
);

OR2x2_ASAP7_75t_L g1340 ( 
.A(n_1173),
.B(n_1044),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_1097),
.B(n_901),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1130),
.Y(n_1342)
);

AND2x2_ASAP7_75t_SL g1343 ( 
.A(n_1173),
.B(n_1071),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_1182),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1100),
.B(n_711),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1133),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1166),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_SL g1348 ( 
.A(n_1103),
.B(n_842),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1134),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1212),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_1183),
.Y(n_1351)
);

AND2x6_ASAP7_75t_L g1352 ( 
.A(n_1103),
.B(n_798),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1192),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1192),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1210),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1194),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_1131),
.Y(n_1357)
);

INVx2_ASAP7_75t_SL g1358 ( 
.A(n_1208),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1217),
.B(n_713),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1194),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1208),
.B(n_904),
.Y(n_1361)
);

BUFx6f_ASAP7_75t_L g1362 ( 
.A(n_1182),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1205),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_SL g1364 ( 
.A(n_1177),
.B(n_1221),
.Y(n_1364)
);

AND2x6_ASAP7_75t_L g1365 ( 
.A(n_1187),
.B(n_798),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1160),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1217),
.A2(n_811),
.B1(n_703),
.B2(n_704),
.Y(n_1367)
);

BUFx3_ASAP7_75t_L g1368 ( 
.A(n_1208),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1174),
.B(n_737),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1205),
.Y(n_1370)
);

AOI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1148),
.A2(n_741),
.B1(n_745),
.B2(n_744),
.Y(n_1371)
);

BUFx6f_ASAP7_75t_L g1372 ( 
.A(n_1182),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1176),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_1139),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1147),
.A2(n_706),
.B1(n_708),
.B2(n_700),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1183),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_SL g1377 ( 
.A(n_1124),
.B(n_747),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1180),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1184),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_SL g1380 ( 
.A(n_1225),
.B(n_753),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1185),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1188),
.B(n_757),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1190),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1139),
.Y(n_1384)
);

BUFx3_ASAP7_75t_L g1385 ( 
.A(n_1219),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1193),
.B(n_759),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1139),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_SL g1388 ( 
.A(n_1202),
.B(n_775),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1196),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1147),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1195),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1213),
.B(n_1147),
.Y(n_1392)
);

INVx4_ASAP7_75t_L g1393 ( 
.A(n_1196),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_1148),
.B(n_907),
.Y(n_1394)
);

INVx4_ASAP7_75t_L g1395 ( 
.A(n_1196),
.Y(n_1395)
);

BUFx6f_ASAP7_75t_L g1396 ( 
.A(n_1197),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1148),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1213),
.B(n_930),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1215),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1197),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1147),
.A2(n_716),
.B1(n_721),
.B2(n_714),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1216),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1147),
.B(n_787),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1197),
.Y(n_1404)
);

BUFx3_ASAP7_75t_L g1405 ( 
.A(n_1162),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1218),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1160),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1162),
.A2(n_760),
.B1(n_761),
.B2(n_725),
.Y(n_1408)
);

INVxp33_ASAP7_75t_L g1409 ( 
.A(n_1118),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1201),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1151),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_SL g1412 ( 
.A(n_1150),
.B(n_788),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1164),
.B(n_840),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1162),
.A2(n_1138),
.B1(n_1172),
.B2(n_1153),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1162),
.B(n_791),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_1162),
.Y(n_1416)
);

INVx2_ASAP7_75t_SL g1417 ( 
.A(n_1164),
.Y(n_1417)
);

INVxp67_ASAP7_75t_L g1418 ( 
.A(n_1226),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1151),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1152),
.Y(n_1420)
);

AND2x6_ASAP7_75t_L g1421 ( 
.A(n_1177),
.B(n_1152),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1189),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1175),
.B(n_841),
.Y(n_1423)
);

AND2x4_ASAP7_75t_L g1424 ( 
.A(n_1189),
.B(n_909),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1186),
.B(n_843),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1115),
.A2(n_780),
.B1(n_781),
.B2(n_774),
.Y(n_1426)
);

AND2x6_ASAP7_75t_L g1427 ( 
.A(n_1177),
.B(n_783),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1251),
.B(n_1159),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1244),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1248),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1298),
.B(n_1159),
.Y(n_1431)
);

O2A1O1Ixp5_ASAP7_75t_L g1432 ( 
.A1(n_1412),
.A2(n_1392),
.B(n_1377),
.C(n_1388),
.Y(n_1432)
);

A2O1A1Ixp33_ASAP7_75t_L g1433 ( 
.A1(n_1398),
.A2(n_1186),
.B(n_1207),
.C(n_1116),
.Y(n_1433)
);

AOI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1315),
.A2(n_1226),
.B1(n_806),
.B2(n_1159),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1249),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1393),
.Y(n_1436)
);

NOR2xp67_ASAP7_75t_L g1437 ( 
.A(n_1269),
.B(n_847),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1298),
.B(n_1116),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_SL g1439 ( 
.A(n_1262),
.B(n_1071),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1274),
.A2(n_1168),
.B1(n_1119),
.B2(n_742),
.Y(n_1440)
);

INVx3_ASAP7_75t_L g1441 ( 
.A(n_1393),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_SL g1442 ( 
.A(n_1307),
.B(n_1203),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1397),
.A2(n_1168),
.B1(n_1119),
.B2(n_742),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_L g1444 ( 
.A(n_1247),
.B(n_599),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_SL g1445 ( 
.A(n_1303),
.B(n_1203),
.Y(n_1445)
);

INVxp33_ASAP7_75t_L g1446 ( 
.A(n_1235),
.Y(n_1446)
);

INVx3_ASAP7_75t_L g1447 ( 
.A(n_1395),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1252),
.B(n_1203),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1247),
.B(n_607),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1273),
.B(n_621),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1263),
.A2(n_613),
.B1(n_785),
.B2(n_784),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_1254),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1283),
.B(n_851),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1264),
.B(n_1203),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1283),
.B(n_853),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1264),
.B(n_1115),
.Y(n_1456)
);

AOI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1358),
.A2(n_1115),
.B1(n_742),
.B2(n_754),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_SL g1458 ( 
.A(n_1273),
.B(n_735),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1268),
.B(n_736),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1234),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1330),
.B(n_796),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_SL g1462 ( 
.A(n_1330),
.B(n_1289),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1268),
.B(n_617),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_L g1464 ( 
.A(n_1276),
.B(n_619),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1253),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1286),
.B(n_628),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1243),
.Y(n_1467)
);

A2O1A1Ixp33_ASAP7_75t_L g1468 ( 
.A1(n_1321),
.A2(n_804),
.B(n_816),
.C(n_792),
.Y(n_1468)
);

INVx2_ASAP7_75t_SL g1469 ( 
.A(n_1231),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1299),
.B(n_630),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1347),
.A2(n_773),
.B1(n_754),
.B2(n_823),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1263),
.A2(n_829),
.B1(n_828),
.B2(n_710),
.Y(n_1472)
);

INVx3_ASAP7_75t_L g1473 ( 
.A(n_1395),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_SL g1474 ( 
.A(n_1289),
.B(n_754),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1285),
.B(n_631),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1267),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1238),
.B(n_1349),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1304),
.B(n_632),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1271),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1280),
.B(n_638),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_SL g1481 ( 
.A(n_1325),
.B(n_773),
.Y(n_1481)
);

OAI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1321),
.A2(n_911),
.B(n_910),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_L g1483 ( 
.A(n_1331),
.B(n_640),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1245),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1272),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1246),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1280),
.B(n_641),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1311),
.B(n_643),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1316),
.B(n_646),
.Y(n_1489)
);

OAI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1409),
.A2(n_710),
.B1(n_831),
.B2(n_606),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_SL g1491 ( 
.A(n_1331),
.B(n_773),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1313),
.A2(n_913),
.B1(n_915),
.B2(n_912),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_SL g1493 ( 
.A(n_1250),
.B(n_1326),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1328),
.B(n_649),
.Y(n_1494)
);

INVx8_ASAP7_75t_L g1495 ( 
.A(n_1237),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_SL g1496 ( 
.A(n_1250),
.B(n_916),
.Y(n_1496)
);

INVx2_ASAP7_75t_SL g1497 ( 
.A(n_1288),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1278),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1333),
.B(n_653),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1336),
.B(n_654),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1340),
.B(n_658),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1339),
.B(n_660),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1342),
.B(n_662),
.Y(n_1503)
);

NAND2x1p5_ASAP7_75t_L g1504 ( 
.A(n_1291),
.B(n_856),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1313),
.A2(n_918),
.B1(n_920),
.B2(n_917),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1302),
.B(n_664),
.Y(n_1506)
);

INVx8_ASAP7_75t_L g1507 ( 
.A(n_1237),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1346),
.B(n_1308),
.Y(n_1508)
);

AOI221xp5_ASAP7_75t_L g1509 ( 
.A1(n_1414),
.A2(n_833),
.B1(n_832),
.B2(n_831),
.C(n_666),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1282),
.Y(n_1510)
);

AOI221xp5_ASAP7_75t_L g1511 ( 
.A1(n_1414),
.A2(n_833),
.B1(n_832),
.B2(n_669),
.C(n_674),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_1351),
.B(n_665),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1257),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1308),
.B(n_673),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_1255),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1376),
.B(n_676),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1417),
.B(n_921),
.Y(n_1517)
);

AND2x2_ASAP7_75t_SL g1518 ( 
.A(n_1343),
.B(n_609),
.Y(n_1518)
);

A2O1A1Ixp33_ASAP7_75t_L g1519 ( 
.A1(n_1392),
.A2(n_924),
.B(n_932),
.C(n_923),
.Y(n_1519)
);

NAND3xp33_ASAP7_75t_L g1520 ( 
.A(n_1240),
.B(n_687),
.C(n_677),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_SL g1521 ( 
.A(n_1368),
.B(n_1364),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1232),
.B(n_693),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1290),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1233),
.B(n_1301),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_SL g1525 ( 
.A(n_1364),
.B(n_934),
.Y(n_1525)
);

AOI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1306),
.A2(n_694),
.B1(n_701),
.B2(n_698),
.Y(n_1526)
);

AOI221xp5_ASAP7_75t_L g1527 ( 
.A1(n_1240),
.A2(n_705),
.B1(n_712),
.B2(n_707),
.C(n_702),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1312),
.B(n_715),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1239),
.B(n_717),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1396),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1266),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_SL g1532 ( 
.A(n_1371),
.B(n_1230),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1318),
.B(n_718),
.Y(n_1533)
);

INVx2_ASAP7_75t_SL g1534 ( 
.A(n_1281),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1324),
.B(n_722),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1329),
.B(n_723),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1332),
.B(n_727),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1413),
.B(n_1355),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1295),
.B(n_728),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1394),
.A2(n_726),
.B1(n_786),
.B2(n_670),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1297),
.B(n_730),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1275),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1293),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1300),
.B(n_732),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1394),
.A2(n_726),
.B1(n_786),
.B2(n_670),
.Y(n_1545)
);

AOI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1277),
.A2(n_738),
.B1(n_740),
.B2(n_739),
.Y(n_1546)
);

AOI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1287),
.A2(n_743),
.B1(n_750),
.B2(n_748),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_SL g1548 ( 
.A(n_1371),
.B(n_752),
.Y(n_1548)
);

AOI221xp5_ASAP7_75t_L g1549 ( 
.A1(n_1265),
.A2(n_756),
.B1(n_765),
.B2(n_764),
.C(n_755),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1230),
.B(n_767),
.Y(n_1550)
);

AOI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1236),
.A2(n_770),
.B1(n_777),
.B2(n_772),
.Y(n_1551)
);

BUFx12f_ASAP7_75t_L g1552 ( 
.A(n_1314),
.Y(n_1552)
);

BUFx12f_ASAP7_75t_L g1553 ( 
.A(n_1357),
.Y(n_1553)
);

INVx2_ASAP7_75t_SL g1554 ( 
.A(n_1281),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1361),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1310),
.B(n_782),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1424),
.B(n_790),
.Y(n_1557)
);

INVx2_ASAP7_75t_SL g1558 ( 
.A(n_1385),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1396),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_L g1560 ( 
.A(n_1423),
.B(n_793),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1366),
.Y(n_1561)
);

OR2x6_ASAP7_75t_L g1562 ( 
.A(n_1418),
.B(n_856),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1348),
.B(n_1380),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1361),
.B(n_794),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1279),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1309),
.Y(n_1566)
);

INVxp67_ASAP7_75t_SL g1567 ( 
.A(n_1260),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1294),
.Y(n_1568)
);

AO22x1_ASAP7_75t_L g1569 ( 
.A1(n_1237),
.A2(n_801),
.B1(n_802),
.B2(n_799),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1292),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1309),
.B(n_803),
.Y(n_1571)
);

NAND2x1p5_ASAP7_75t_L g1572 ( 
.A(n_1296),
.B(n_1319),
.Y(n_1572)
);

INVxp67_ASAP7_75t_L g1573 ( 
.A(n_1265),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1341),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1334),
.B(n_807),
.Y(n_1575)
);

INVx2_ASAP7_75t_SL g1576 ( 
.A(n_1334),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1341),
.B(n_808),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1242),
.B(n_809),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1353),
.B(n_812),
.Y(n_1579)
);

INVx4_ASAP7_75t_L g1580 ( 
.A(n_1260),
.Y(n_1580)
);

NAND3xp33_ASAP7_75t_L g1581 ( 
.A(n_1375),
.B(n_1408),
.C(n_1401),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_SL g1582 ( 
.A(n_1260),
.B(n_814),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1354),
.B(n_815),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1418),
.B(n_817),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1350),
.Y(n_1585)
);

BUFx3_ASAP7_75t_L g1586 ( 
.A(n_1407),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_SL g1587 ( 
.A(n_1270),
.B(n_819),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1360),
.B(n_820),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1369),
.B(n_821),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1259),
.B(n_1261),
.Y(n_1590)
);

INVxp67_ASAP7_75t_SL g1591 ( 
.A(n_1270),
.Y(n_1591)
);

INVx2_ASAP7_75t_SL g1592 ( 
.A(n_1237),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_SL g1593 ( 
.A(n_1270),
.B(n_827),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1259),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1356),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1261),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1338),
.B(n_480),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1337),
.A2(n_805),
.B1(n_871),
.B2(n_903),
.Y(n_1598)
);

INVx2_ASAP7_75t_SL g1599 ( 
.A(n_1396),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_SL g1600 ( 
.A(n_1284),
.B(n_805),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1338),
.B(n_481),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1363),
.B(n_482),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1370),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1337),
.A2(n_871),
.B1(n_926),
.B2(n_903),
.Y(n_1604)
);

AND2x4_ASAP7_75t_L g1605 ( 
.A(n_1405),
.B(n_484),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1374),
.B(n_487),
.Y(n_1606)
);

INVxp67_ASAP7_75t_L g1607 ( 
.A(n_1369),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1373),
.Y(n_1608)
);

OAI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1367),
.A2(n_871),
.B(n_489),
.Y(n_1609)
);

AOI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1236),
.A2(n_926),
.B1(n_903),
.B2(n_491),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1374),
.B(n_1404),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_1416),
.Y(n_1612)
);

AOI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1236),
.A2(n_1337),
.B1(n_1386),
.B2(n_1382),
.Y(n_1613)
);

INVx8_ASAP7_75t_L g1614 ( 
.A(n_1421),
.Y(n_1614)
);

INVxp67_ASAP7_75t_L g1615 ( 
.A(n_1382),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1404),
.B(n_488),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1386),
.B(n_0),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1256),
.B(n_494),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1256),
.B(n_496),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1384),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1256),
.B(n_497),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1425),
.A2(n_926),
.B1(n_903),
.B2(n_3),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1367),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_SL g1624 ( 
.A(n_1284),
.B(n_501),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1236),
.B(n_1),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1317),
.B(n_4),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1378),
.Y(n_1627)
);

INVxp67_ASAP7_75t_L g1628 ( 
.A(n_1399),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1459),
.B(n_1317),
.Y(n_1629)
);

INVx5_ASAP7_75t_L g1630 ( 
.A(n_1495),
.Y(n_1630)
);

NOR2x1_ASAP7_75t_L g1631 ( 
.A(n_1580),
.B(n_1296),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1574),
.B(n_1379),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1460),
.Y(n_1633)
);

INVxp67_ASAP7_75t_L g1634 ( 
.A(n_1461),
.Y(n_1634)
);

INVx5_ASAP7_75t_L g1635 ( 
.A(n_1495),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1467),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1484),
.Y(n_1637)
);

INVx2_ASAP7_75t_SL g1638 ( 
.A(n_1452),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1538),
.B(n_1345),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1508),
.B(n_1256),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1469),
.B(n_1375),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_1515),
.Y(n_1642)
);

NOR2xp67_ASAP7_75t_L g1643 ( 
.A(n_1607),
.B(n_1403),
.Y(n_1643)
);

INVx2_ASAP7_75t_SL g1644 ( 
.A(n_1558),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1429),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1615),
.B(n_1258),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1464),
.B(n_1475),
.Y(n_1647)
);

BUFx2_ASAP7_75t_L g1648 ( 
.A(n_1555),
.Y(n_1648)
);

BUFx3_ASAP7_75t_L g1649 ( 
.A(n_1586),
.Y(n_1649)
);

INVxp67_ASAP7_75t_L g1650 ( 
.A(n_1444),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_SL g1651 ( 
.A(n_1497),
.B(n_1345),
.Y(n_1651)
);

OR2x6_ASAP7_75t_L g1652 ( 
.A(n_1495),
.B(n_1507),
.Y(n_1652)
);

AND2x6_ASAP7_75t_SL g1653 ( 
.A(n_1560),
.B(n_1403),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1566),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1430),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_SL g1656 ( 
.A(n_1449),
.B(n_1284),
.Y(n_1656)
);

OAI22xp33_ASAP7_75t_L g1657 ( 
.A1(n_1478),
.A2(n_1415),
.B1(n_1390),
.B2(n_1410),
.Y(n_1657)
);

BUFx3_ASAP7_75t_L g1658 ( 
.A(n_1552),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1459),
.B(n_1258),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1581),
.A2(n_1426),
.B1(n_1401),
.B2(n_1408),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1446),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1450),
.B(n_1320),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1435),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_1553),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1486),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1453),
.B(n_1381),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1477),
.B(n_1241),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1465),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1517),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1463),
.B(n_1258),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1480),
.B(n_1359),
.Y(n_1671)
);

INVx3_ASAP7_75t_L g1672 ( 
.A(n_1614),
.Y(n_1672)
);

BUFx6f_ASAP7_75t_L g1673 ( 
.A(n_1614),
.Y(n_1673)
);

INVx1_ASAP7_75t_SL g1674 ( 
.A(n_1455),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_SL g1675 ( 
.A(n_1576),
.B(n_1320),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_L g1676 ( 
.A(n_1514),
.B(n_1383),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1501),
.B(n_1391),
.Y(n_1677)
);

AND2x4_ASAP7_75t_L g1678 ( 
.A(n_1493),
.B(n_1402),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1476),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1462),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1479),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1589),
.B(n_1258),
.Y(n_1682)
);

NAND2x1p5_ASAP7_75t_L g1683 ( 
.A(n_1436),
.B(n_1319),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1483),
.B(n_1305),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1506),
.B(n_1305),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1485),
.Y(n_1686)
);

HB1xp67_ASAP7_75t_L g1687 ( 
.A(n_1573),
.Y(n_1687)
);

INVxp67_ASAP7_75t_L g1688 ( 
.A(n_1512),
.Y(n_1688)
);

NAND2x1p5_ASAP7_75t_L g1689 ( 
.A(n_1436),
.B(n_1322),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1498),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1428),
.B(n_1510),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1521),
.B(n_1406),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1523),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1543),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1568),
.Y(n_1695)
);

NAND2x1p5_ASAP7_75t_L g1696 ( 
.A(n_1441),
.B(n_1322),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1516),
.B(n_1411),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1608),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_1561),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_1612),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1627),
.Y(n_1701)
);

BUFx6f_ASAP7_75t_L g1702 ( 
.A(n_1614),
.Y(n_1702)
);

BUFx4f_ASAP7_75t_L g1703 ( 
.A(n_1518),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1524),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1595),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1487),
.B(n_1419),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1548),
.A2(n_1365),
.B1(n_1335),
.B2(n_1352),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_1439),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1466),
.B(n_1387),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1470),
.B(n_1389),
.Y(n_1710)
);

NOR2xp67_ASAP7_75t_L g1711 ( 
.A(n_1626),
.B(n_1400),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1603),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_SL g1713 ( 
.A(n_1437),
.B(n_1563),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1513),
.Y(n_1714)
);

AND2x2_ASAP7_75t_SL g1715 ( 
.A(n_1617),
.B(n_1320),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1556),
.B(n_1420),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1520),
.A2(n_1365),
.B1(n_1335),
.B2(n_1352),
.Y(n_1717)
);

BUFx3_ASAP7_75t_L g1718 ( 
.A(n_1534),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1531),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1431),
.B(n_1335),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1554),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1564),
.B(n_1422),
.Y(n_1722)
);

BUFx4f_ASAP7_75t_L g1723 ( 
.A(n_1605),
.Y(n_1723)
);

BUFx8_ASAP7_75t_L g1724 ( 
.A(n_1605),
.Y(n_1724)
);

AND2x6_ASAP7_75t_L g1725 ( 
.A(n_1441),
.B(n_1322),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1628),
.B(n_1335),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1542),
.Y(n_1727)
);

INVx2_ASAP7_75t_SL g1728 ( 
.A(n_1599),
.Y(n_1728)
);

BUFx2_ASAP7_75t_L g1729 ( 
.A(n_1562),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1579),
.B(n_1583),
.Y(n_1730)
);

BUFx12f_ASAP7_75t_L g1731 ( 
.A(n_1562),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1565),
.Y(n_1732)
);

AND2x2_ASAP7_75t_SL g1733 ( 
.A(n_1622),
.B(n_1323),
.Y(n_1733)
);

INVx2_ASAP7_75t_SL g1734 ( 
.A(n_1529),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1570),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1431),
.B(n_1365),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1585),
.Y(n_1737)
);

BUFx3_ASAP7_75t_L g1738 ( 
.A(n_1530),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1620),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1491),
.B(n_1584),
.Y(n_1740)
);

BUFx6f_ASAP7_75t_L g1741 ( 
.A(n_1507),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1594),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1609),
.A2(n_1365),
.B1(n_1427),
.B2(n_1327),
.Y(n_1743)
);

AND2x6_ASAP7_75t_SL g1744 ( 
.A(n_1577),
.B(n_1427),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1438),
.B(n_1323),
.Y(n_1745)
);

AOI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1623),
.A2(n_1427),
.B1(n_1421),
.B2(n_1327),
.Y(n_1746)
);

INVxp67_ASAP7_75t_L g1747 ( 
.A(n_1557),
.Y(n_1747)
);

NOR2xp67_ASAP7_75t_L g1748 ( 
.A(n_1613),
.B(n_1323),
.Y(n_1748)
);

BUFx3_ASAP7_75t_L g1749 ( 
.A(n_1530),
.Y(n_1749)
);

BUFx3_ASAP7_75t_L g1750 ( 
.A(n_1559),
.Y(n_1750)
);

BUFx3_ASAP7_75t_L g1751 ( 
.A(n_1559),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1596),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_SL g1753 ( 
.A(n_1434),
.B(n_1327),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1590),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1583),
.B(n_1344),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_SL g1756 ( 
.A(n_1532),
.B(n_1344),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1590),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_L g1758 ( 
.A1(n_1609),
.A2(n_1362),
.B1(n_1372),
.B2(n_1344),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1571),
.B(n_1362),
.Y(n_1759)
);

INVx5_ASAP7_75t_L g1760 ( 
.A(n_1507),
.Y(n_1760)
);

AOI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1456),
.A2(n_1372),
.B(n_1362),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1611),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1611),
.Y(n_1763)
);

BUFx8_ASAP7_75t_L g1764 ( 
.A(n_1592),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1447),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_1451),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1588),
.B(n_1372),
.Y(n_1767)
);

AOI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1549),
.A2(n_1421),
.B1(n_6),
.B2(n_4),
.Y(n_1768)
);

NAND2xp33_ASAP7_75t_L g1769 ( 
.A(n_1572),
.B(n_502),
.Y(n_1769)
);

BUFx6f_ASAP7_75t_L g1770 ( 
.A(n_1572),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1528),
.B(n_5),
.Y(n_1771)
);

OAI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1546),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1438),
.B(n_1454),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1447),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1533),
.Y(n_1775)
);

INVx2_ASAP7_75t_SL g1776 ( 
.A(n_1496),
.Y(n_1776)
);

OAI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1547),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1458),
.B(n_8),
.Y(n_1778)
);

CKINVDCx5p33_ASAP7_75t_R g1779 ( 
.A(n_1451),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1582),
.B(n_504),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1575),
.B(n_10),
.Y(n_1781)
);

INVx2_ASAP7_75t_SL g1782 ( 
.A(n_1562),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_R g1783 ( 
.A(n_1618),
.B(n_506),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1535),
.B(n_11),
.Y(n_1784)
);

INVx2_ASAP7_75t_SL g1785 ( 
.A(n_1587),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1536),
.Y(n_1786)
);

INVx5_ASAP7_75t_L g1787 ( 
.A(n_1473),
.Y(n_1787)
);

BUFx12f_ASAP7_75t_SL g1788 ( 
.A(n_1600),
.Y(n_1788)
);

BUFx3_ASAP7_75t_L g1789 ( 
.A(n_1504),
.Y(n_1789)
);

OR2x6_ASAP7_75t_L g1790 ( 
.A(n_1445),
.B(n_507),
.Y(n_1790)
);

NOR2xp67_ASAP7_75t_L g1791 ( 
.A(n_1550),
.B(n_508),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1537),
.Y(n_1792)
);

BUFx8_ASAP7_75t_L g1793 ( 
.A(n_1569),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1448),
.B(n_1473),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1482),
.B(n_1567),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1482),
.B(n_12),
.Y(n_1796)
);

AND2x4_ASAP7_75t_L g1797 ( 
.A(n_1593),
.B(n_511),
.Y(n_1797)
);

INVx3_ASAP7_75t_L g1798 ( 
.A(n_1504),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1591),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1602),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1522),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1468),
.B(n_13),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1440),
.B(n_14),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1488),
.B(n_14),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1602),
.Y(n_1805)
);

AOI22xp33_ASAP7_75t_L g1806 ( 
.A1(n_1623),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_1806)
);

O2A1O1Ixp5_ASAP7_75t_L g1807 ( 
.A1(n_1525),
.A2(n_18),
.B(n_16),
.C(n_17),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1519),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1489),
.B(n_18),
.Y(n_1809)
);

BUFx6f_ASAP7_75t_SL g1810 ( 
.A(n_1481),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1539),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1541),
.Y(n_1812)
);

NAND3xp33_ASAP7_75t_SL g1813 ( 
.A(n_1511),
.B(n_19),
.C(n_20),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1544),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_SL g1815 ( 
.A(n_1647),
.B(n_1432),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_SL g1816 ( 
.A(n_1715),
.B(n_1625),
.Y(n_1816)
);

NAND2xp33_ASAP7_75t_SL g1817 ( 
.A(n_1700),
.B(n_1474),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_SL g1818 ( 
.A(n_1688),
.B(n_1551),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1674),
.B(n_1509),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_SL g1820 ( 
.A(n_1634),
.B(n_1526),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1674),
.B(n_1492),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1650),
.B(n_1494),
.Y(n_1822)
);

NAND2xp33_ASAP7_75t_SL g1823 ( 
.A(n_1642),
.B(n_1540),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_SL g1824 ( 
.A(n_1740),
.B(n_1499),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_SL g1825 ( 
.A(n_1677),
.B(n_1500),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_SL g1826 ( 
.A(n_1676),
.B(n_1734),
.Y(n_1826)
);

NAND2xp33_ASAP7_75t_SL g1827 ( 
.A(n_1766),
.B(n_1779),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_SL g1828 ( 
.A(n_1643),
.B(n_1502),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1629),
.B(n_1490),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_SL g1830 ( 
.A(n_1643),
.B(n_1503),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_SL g1831 ( 
.A(n_1814),
.B(n_1578),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_SL g1832 ( 
.A(n_1801),
.B(n_1619),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_SL g1833 ( 
.A(n_1811),
.B(n_1619),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1730),
.B(n_1527),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1812),
.B(n_1621),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_SL g1836 ( 
.A(n_1723),
.B(n_1621),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_SL g1837 ( 
.A(n_1723),
.B(n_1545),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_SL g1838 ( 
.A(n_1716),
.B(n_1713),
.Y(n_1838)
);

NAND2xp33_ASAP7_75t_SL g1839 ( 
.A(n_1810),
.B(n_1699),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_SL g1840 ( 
.A(n_1667),
.B(n_1457),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_SL g1841 ( 
.A(n_1697),
.B(n_1606),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_SL g1842 ( 
.A(n_1708),
.B(n_1775),
.Y(n_1842)
);

NAND2xp33_ASAP7_75t_SL g1843 ( 
.A(n_1810),
.B(n_1471),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_SL g1844 ( 
.A(n_1786),
.B(n_1616),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_SL g1845 ( 
.A(n_1792),
.B(n_1616),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_SL g1846 ( 
.A(n_1747),
.B(n_1610),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_SL g1847 ( 
.A(n_1703),
.B(n_1597),
.Y(n_1847)
);

NAND2xp33_ASAP7_75t_SL g1848 ( 
.A(n_1638),
.B(n_1442),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1704),
.B(n_1505),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1666),
.B(n_1710),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1669),
.B(n_1472),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_SL g1852 ( 
.A(n_1703),
.B(n_1685),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_SL g1853 ( 
.A(n_1692),
.B(n_1597),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1639),
.B(n_1472),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_SL g1855 ( 
.A(n_1692),
.B(n_1601),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_SL g1856 ( 
.A(n_1785),
.B(n_1601),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_SL g1857 ( 
.A(n_1684),
.B(n_1598),
.Y(n_1857)
);

NAND2xp33_ASAP7_75t_SL g1858 ( 
.A(n_1644),
.B(n_1624),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_SL g1859 ( 
.A(n_1682),
.B(n_1443),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_SL g1860 ( 
.A(n_1780),
.B(n_1433),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_SL g1861 ( 
.A(n_1780),
.B(n_1604),
.Y(n_1861)
);

NAND2xp33_ASAP7_75t_SL g1862 ( 
.A(n_1741),
.B(n_19),
.Y(n_1862)
);

NAND2xp33_ASAP7_75t_SL g1863 ( 
.A(n_1741),
.B(n_20),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1759),
.B(n_21),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_SL g1865 ( 
.A(n_1797),
.B(n_21),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_SL g1866 ( 
.A(n_1797),
.B(n_22),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_SL g1867 ( 
.A(n_1678),
.B(n_22),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1641),
.B(n_23),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_SL g1869 ( 
.A(n_1678),
.B(n_23),
.Y(n_1869)
);

NAND2xp33_ASAP7_75t_SL g1870 ( 
.A(n_1741),
.B(n_24),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1706),
.B(n_1691),
.Y(n_1871)
);

NAND2xp33_ASAP7_75t_SL g1872 ( 
.A(n_1673),
.B(n_24),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_SL g1873 ( 
.A(n_1632),
.B(n_25),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_SL g1874 ( 
.A(n_1632),
.B(n_26),
.Y(n_1874)
);

NAND2xp33_ASAP7_75t_SL g1875 ( 
.A(n_1673),
.B(n_27),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_SL g1876 ( 
.A(n_1657),
.B(n_27),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_SL g1877 ( 
.A(n_1733),
.B(n_28),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_SL g1878 ( 
.A(n_1646),
.B(n_29),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_SL g1879 ( 
.A(n_1646),
.B(n_29),
.Y(n_1879)
);

NAND2xp33_ASAP7_75t_SL g1880 ( 
.A(n_1673),
.B(n_30),
.Y(n_1880)
);

NAND2xp33_ASAP7_75t_SL g1881 ( 
.A(n_1702),
.B(n_1776),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1691),
.B(n_30),
.Y(n_1882)
);

NAND2xp33_ASAP7_75t_SL g1883 ( 
.A(n_1702),
.B(n_31),
.Y(n_1883)
);

NAND2xp33_ASAP7_75t_SL g1884 ( 
.A(n_1702),
.B(n_32),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_SL g1885 ( 
.A(n_1671),
.B(n_32),
.Y(n_1885)
);

NAND2xp33_ASAP7_75t_SL g1886 ( 
.A(n_1783),
.B(n_33),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_SL g1887 ( 
.A(n_1651),
.B(n_33),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1709),
.B(n_1680),
.Y(n_1888)
);

NAND2xp33_ASAP7_75t_SL g1889 ( 
.A(n_1664),
.B(n_34),
.Y(n_1889)
);

NAND2xp33_ASAP7_75t_SL g1890 ( 
.A(n_1721),
.B(n_35),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_SL g1891 ( 
.A(n_1804),
.B(n_1809),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_SL g1892 ( 
.A(n_1804),
.B(n_35),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1722),
.B(n_36),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_SL g1894 ( 
.A(n_1809),
.B(n_36),
.Y(n_1894)
);

NAND2xp33_ASAP7_75t_SL g1895 ( 
.A(n_1729),
.B(n_37),
.Y(n_1895)
);

NAND2xp33_ASAP7_75t_SL g1896 ( 
.A(n_1803),
.B(n_1654),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_SL g1897 ( 
.A(n_1656),
.B(n_37),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_SL g1898 ( 
.A(n_1662),
.B(n_38),
.Y(n_1898)
);

NAND2xp33_ASAP7_75t_SL g1899 ( 
.A(n_1803),
.B(n_1768),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_SL g1900 ( 
.A(n_1755),
.B(n_39),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_SL g1901 ( 
.A(n_1767),
.B(n_39),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_L g1902 ( 
.A(n_1661),
.B(n_512),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_SL g1903 ( 
.A(n_1771),
.B(n_40),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1709),
.B(n_41),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_SL g1905 ( 
.A(n_1784),
.B(n_41),
.Y(n_1905)
);

AND2x2_ASAP7_75t_SL g1906 ( 
.A(n_1769),
.B(n_42),
.Y(n_1906)
);

NAND2xp33_ASAP7_75t_SL g1907 ( 
.A(n_1648),
.B(n_42),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_SL g1908 ( 
.A(n_1726),
.B(n_43),
.Y(n_1908)
);

NAND2xp33_ASAP7_75t_SL g1909 ( 
.A(n_1770),
.B(n_43),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1781),
.B(n_44),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_SL g1911 ( 
.A(n_1711),
.B(n_46),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_SL g1912 ( 
.A(n_1793),
.B(n_47),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_SL g1913 ( 
.A(n_1793),
.B(n_47),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1773),
.B(n_48),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_SL g1915 ( 
.A(n_1778),
.B(n_49),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_SL g1916 ( 
.A(n_1800),
.B(n_49),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_SL g1917 ( 
.A(n_1805),
.B(n_50),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1687),
.B(n_51),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_SL g1919 ( 
.A(n_1659),
.B(n_52),
.Y(n_1919)
);

AND2x4_ASAP7_75t_L g1920 ( 
.A(n_1652),
.B(n_515),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_SL g1921 ( 
.A(n_1640),
.B(n_53),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1773),
.B(n_54),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_SL g1923 ( 
.A(n_1640),
.B(n_55),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_SL g1924 ( 
.A(n_1787),
.B(n_56),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_SL g1925 ( 
.A(n_1787),
.B(n_57),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_SL g1926 ( 
.A(n_1787),
.B(n_1795),
.Y(n_1926)
);

NAND2xp33_ASAP7_75t_SL g1927 ( 
.A(n_1770),
.B(n_58),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_SL g1928 ( 
.A(n_1795),
.B(n_58),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1670),
.B(n_59),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_SL g1930 ( 
.A(n_1791),
.B(n_59),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_SL g1931 ( 
.A(n_1791),
.B(n_60),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_SL g1932 ( 
.A(n_1724),
.B(n_1770),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1652),
.B(n_516),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1754),
.B(n_63),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_SL g1935 ( 
.A(n_1724),
.B(n_65),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_SL g1936 ( 
.A(n_1714),
.B(n_65),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_SL g1937 ( 
.A(n_1719),
.B(n_66),
.Y(n_1937)
);

NAND2xp33_ASAP7_75t_SL g1938 ( 
.A(n_1806),
.B(n_66),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_SL g1939 ( 
.A(n_1727),
.B(n_67),
.Y(n_1939)
);

NAND2xp33_ASAP7_75t_SL g1940 ( 
.A(n_1782),
.B(n_67),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_SL g1941 ( 
.A(n_1732),
.B(n_1735),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_SL g1942 ( 
.A(n_1739),
.B(n_68),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_SL g1943 ( 
.A(n_1633),
.B(n_68),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_SL g1944 ( 
.A(n_1636),
.B(n_69),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_SL g1945 ( 
.A(n_1637),
.B(n_69),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_SL g1946 ( 
.A(n_1665),
.B(n_70),
.Y(n_1946)
);

AND2x4_ASAP7_75t_L g1947 ( 
.A(n_1652),
.B(n_518),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1757),
.B(n_72),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_SL g1949 ( 
.A(n_1737),
.B(n_72),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1762),
.B(n_73),
.Y(n_1950)
);

NAND2xp33_ASAP7_75t_SL g1951 ( 
.A(n_1758),
.B(n_74),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_SL g1952 ( 
.A(n_1660),
.B(n_76),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_SL g1953 ( 
.A(n_1660),
.B(n_76),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_SL g1954 ( 
.A(n_1698),
.B(n_77),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_SL g1955 ( 
.A(n_1701),
.B(n_77),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_SL g1956 ( 
.A(n_1796),
.B(n_78),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_SL g1957 ( 
.A(n_1796),
.B(n_79),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_SL g1958 ( 
.A(n_1763),
.B(n_79),
.Y(n_1958)
);

AND2x4_ASAP7_75t_L g1959 ( 
.A(n_1630),
.B(n_521),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1745),
.B(n_80),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_SL g1961 ( 
.A(n_1645),
.B(n_81),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_SL g1962 ( 
.A(n_1655),
.B(n_81),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1745),
.B(n_82),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1663),
.B(n_82),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_SL g1965 ( 
.A(n_1668),
.B(n_83),
.Y(n_1965)
);

NAND2xp33_ASAP7_75t_SL g1966 ( 
.A(n_1672),
.B(n_83),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_SL g1967 ( 
.A(n_1679),
.B(n_84),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1681),
.B(n_1686),
.Y(n_1968)
);

NAND2xp33_ASAP7_75t_SL g1969 ( 
.A(n_1672),
.B(n_1728),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_SL g1970 ( 
.A(n_1690),
.B(n_84),
.Y(n_1970)
);

NAND2xp33_ASAP7_75t_SL g1971 ( 
.A(n_1693),
.B(n_85),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_SL g1972 ( 
.A(n_1694),
.B(n_85),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_SL g1973 ( 
.A(n_1695),
.B(n_1705),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_SL g1974 ( 
.A(n_1712),
.B(n_86),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_SL g1975 ( 
.A(n_1748),
.B(n_86),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_SL g1976 ( 
.A(n_1748),
.B(n_87),
.Y(n_1976)
);

OR2x2_ASAP7_75t_L g1977 ( 
.A(n_1742),
.B(n_88),
.Y(n_1977)
);

NAND2xp33_ASAP7_75t_SL g1978 ( 
.A(n_1799),
.B(n_89),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1968),
.Y(n_1979)
);

INVxp67_ASAP7_75t_L g1980 ( 
.A(n_1826),
.Y(n_1980)
);

AND2x2_ASAP7_75t_SL g1981 ( 
.A(n_1906),
.B(n_1802),
.Y(n_1981)
);

NOR2x1_ASAP7_75t_L g1982 ( 
.A(n_1815),
.B(n_1756),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1973),
.Y(n_1983)
);

INVxp67_ASAP7_75t_L g1984 ( 
.A(n_1850),
.Y(n_1984)
);

AND2x4_ASAP7_75t_L g1985 ( 
.A(n_1920),
.B(n_1630),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1888),
.Y(n_1986)
);

CKINVDCx14_ASAP7_75t_R g1987 ( 
.A(n_1839),
.Y(n_1987)
);

BUFx12f_ASAP7_75t_L g1988 ( 
.A(n_1977),
.Y(n_1988)
);

HB1xp67_ASAP7_75t_L g1989 ( 
.A(n_1871),
.Y(n_1989)
);

AOI21xp5_ASAP7_75t_L g1990 ( 
.A1(n_1860),
.A2(n_1743),
.B(n_1794),
.Y(n_1990)
);

AND3x1_ASAP7_75t_SL g1991 ( 
.A(n_1889),
.B(n_1653),
.C(n_1788),
.Y(n_1991)
);

OR2x2_ASAP7_75t_L g1992 ( 
.A(n_1852),
.B(n_1736),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1868),
.B(n_1752),
.Y(n_1993)
);

AND2x4_ASAP7_75t_L g1994 ( 
.A(n_1920),
.B(n_1630),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1941),
.Y(n_1995)
);

AOI21xp5_ASAP7_75t_L g1996 ( 
.A1(n_1832),
.A2(n_1794),
.B(n_1761),
.Y(n_1996)
);

O2A1O1Ixp5_ASAP7_75t_L g1997 ( 
.A1(n_1876),
.A2(n_1777),
.B(n_1772),
.C(n_1802),
.Y(n_1997)
);

O2A1O1Ixp33_ASAP7_75t_L g1998 ( 
.A1(n_1915),
.A2(n_1813),
.B(n_1807),
.C(n_1753),
.Y(n_1998)
);

HB1xp67_ASAP7_75t_L g1999 ( 
.A(n_1926),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_SL g2000 ( 
.A(n_1824),
.B(n_1707),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1829),
.B(n_1834),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1891),
.B(n_1653),
.Y(n_2002)
);

HB1xp67_ASAP7_75t_L g2003 ( 
.A(n_1838),
.Y(n_2003)
);

NAND2x1p5_ASAP7_75t_L g2004 ( 
.A(n_1920),
.B(n_1635),
.Y(n_2004)
);

INVx5_ASAP7_75t_L g2005 ( 
.A(n_1933),
.Y(n_2005)
);

OAI22xp5_ASAP7_75t_SL g2006 ( 
.A1(n_1906),
.A2(n_1731),
.B1(n_1790),
.B2(n_1658),
.Y(n_2006)
);

OR2x2_ASAP7_75t_L g2007 ( 
.A(n_1960),
.B(n_1736),
.Y(n_2007)
);

A2O1A1Ixp33_ASAP7_75t_L g2008 ( 
.A1(n_1899),
.A2(n_1746),
.B(n_1808),
.C(n_1717),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1831),
.Y(n_2009)
);

NOR2xp33_ASAP7_75t_L g2010 ( 
.A(n_1842),
.B(n_1649),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1963),
.Y(n_2011)
);

INVx3_ASAP7_75t_L g2012 ( 
.A(n_1959),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1934),
.Y(n_2013)
);

BUFx2_ASAP7_75t_L g2014 ( 
.A(n_1969),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1821),
.B(n_1790),
.Y(n_2015)
);

AOI22xp33_ASAP7_75t_L g2016 ( 
.A1(n_1938),
.A2(n_1877),
.B1(n_1953),
.B2(n_1952),
.Y(n_2016)
);

INVx2_ASAP7_75t_SL g2017 ( 
.A(n_1932),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1948),
.Y(n_2018)
);

AOI21xp5_ASAP7_75t_L g2019 ( 
.A1(n_1833),
.A2(n_1720),
.B(n_1746),
.Y(n_2019)
);

XNOR2xp5_ASAP7_75t_L g2020 ( 
.A(n_1827),
.B(n_1718),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1950),
.Y(n_2021)
);

CKINVDCx5p33_ASAP7_75t_R g2022 ( 
.A(n_1822),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_SL g2023 ( 
.A(n_1825),
.B(n_1635),
.Y(n_2023)
);

A2O1A1Ixp33_ASAP7_75t_SL g2024 ( 
.A1(n_1902),
.A2(n_1798),
.B(n_1774),
.C(n_1765),
.Y(n_2024)
);

HB1xp67_ASAP7_75t_L g2025 ( 
.A(n_1841),
.Y(n_2025)
);

AOI21xp5_ASAP7_75t_L g2026 ( 
.A1(n_1835),
.A2(n_1845),
.B(n_1844),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1914),
.Y(n_2027)
);

INVx1_ASAP7_75t_SL g2028 ( 
.A(n_1893),
.Y(n_2028)
);

AOI21xp5_ASAP7_75t_L g2029 ( 
.A1(n_1836),
.A2(n_1683),
.B(n_1635),
.Y(n_2029)
);

BUFx6f_ASAP7_75t_L g2030 ( 
.A(n_1933),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1922),
.B(n_1744),
.Y(n_2031)
);

INVx4_ASAP7_75t_L g2032 ( 
.A(n_1933),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1964),
.Y(n_2033)
);

BUFx8_ASAP7_75t_SL g2034 ( 
.A(n_1864),
.Y(n_2034)
);

INVx4_ASAP7_75t_L g2035 ( 
.A(n_1947),
.Y(n_2035)
);

INVx8_ASAP7_75t_L g2036 ( 
.A(n_1947),
.Y(n_2036)
);

OR2x2_ASAP7_75t_L g2037 ( 
.A(n_1851),
.B(n_1675),
.Y(n_2037)
);

AOI22xp5_ASAP7_75t_L g2038 ( 
.A1(n_1823),
.A2(n_1764),
.B1(n_1749),
.B2(n_1750),
.Y(n_2038)
);

AOI22xp33_ASAP7_75t_L g2039 ( 
.A1(n_1886),
.A2(n_1789),
.B1(n_1764),
.B2(n_1751),
.Y(n_2039)
);

AND2x4_ASAP7_75t_L g2040 ( 
.A(n_1947),
.B(n_1760),
.Y(n_2040)
);

NOR2xp33_ASAP7_75t_L g2041 ( 
.A(n_1818),
.B(n_1738),
.Y(n_2041)
);

NOR2xp33_ASAP7_75t_L g2042 ( 
.A(n_1820),
.B(n_1744),
.Y(n_2042)
);

O2A1O1Ixp33_ASAP7_75t_L g2043 ( 
.A1(n_1840),
.A2(n_1696),
.B(n_1689),
.C(n_1683),
.Y(n_2043)
);

NAND2x1p5_ASAP7_75t_L g2044 ( 
.A(n_1959),
.B(n_1631),
.Y(n_2044)
);

BUFx6f_ASAP7_75t_L g2045 ( 
.A(n_1959),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1904),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1882),
.Y(n_2047)
);

INVx5_ASAP7_75t_L g2048 ( 
.A(n_1918),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1854),
.B(n_1689),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1849),
.Y(n_2050)
);

AOI221xp5_ASAP7_75t_L g2051 ( 
.A1(n_1890),
.A2(n_1696),
.B1(n_92),
.B2(n_90),
.C(n_91),
.Y(n_2051)
);

INVx3_ASAP7_75t_L g2052 ( 
.A(n_1910),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1853),
.Y(n_2053)
);

INVx5_ASAP7_75t_L g2054 ( 
.A(n_1858),
.Y(n_2054)
);

INVx3_ASAP7_75t_L g2055 ( 
.A(n_1881),
.Y(n_2055)
);

AOI21xp5_ASAP7_75t_L g2056 ( 
.A1(n_1855),
.A2(n_1725),
.B(n_523),
.Y(n_2056)
);

INVx6_ASAP7_75t_L g2057 ( 
.A(n_1817),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1856),
.Y(n_2058)
);

INVx1_ASAP7_75t_SL g2059 ( 
.A(n_1896),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_1885),
.B(n_1956),
.Y(n_2060)
);

O2A1O1Ixp33_ASAP7_75t_L g2061 ( 
.A1(n_1865),
.A2(n_1866),
.B(n_1905),
.C(n_1903),
.Y(n_2061)
);

NOR2xp33_ASAP7_75t_SL g2062 ( 
.A(n_1819),
.B(n_1725),
.Y(n_2062)
);

AOI222xp33_ASAP7_75t_SL g2063 ( 
.A1(n_1912),
.A2(n_96),
.B1(n_98),
.B2(n_90),
.C1(n_94),
.C2(n_97),
.Y(n_2063)
);

O2A1O1Ixp5_ASAP7_75t_SL g2064 ( 
.A1(n_1928),
.A2(n_97),
.B(n_94),
.C(n_96),
.Y(n_2064)
);

NOR2x1_ASAP7_75t_L g2065 ( 
.A(n_1828),
.B(n_1725),
.Y(n_2065)
);

INVx1_ASAP7_75t_SL g2066 ( 
.A(n_1816),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1892),
.B(n_522),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_1894),
.B(n_524),
.Y(n_2068)
);

BUFx6f_ASAP7_75t_L g2069 ( 
.A(n_1847),
.Y(n_2069)
);

BUFx3_ASAP7_75t_L g2070 ( 
.A(n_1848),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1957),
.Y(n_2071)
);

BUFx2_ASAP7_75t_L g2072 ( 
.A(n_1843),
.Y(n_2072)
);

AOI22xp5_ASAP7_75t_L g2073 ( 
.A1(n_1837),
.A2(n_1725),
.B1(n_101),
.B2(n_98),
.Y(n_2073)
);

AOI21xp5_ASAP7_75t_L g2074 ( 
.A1(n_1830),
.A2(n_526),
.B(n_525),
.Y(n_2074)
);

AOI21x1_ASAP7_75t_L g2075 ( 
.A1(n_1859),
.A2(n_529),
.B(n_527),
.Y(n_2075)
);

A2O1A1Ixp33_ASAP7_75t_L g2076 ( 
.A1(n_1951),
.A2(n_102),
.B(n_99),
.C(n_101),
.Y(n_2076)
);

INVx2_ASAP7_75t_SL g2077 ( 
.A(n_1924),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_1900),
.B(n_99),
.Y(n_2078)
);

AOI22xp5_ASAP7_75t_L g2079 ( 
.A1(n_1846),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_2079)
);

AND2x4_ASAP7_75t_L g2080 ( 
.A(n_1816),
.B(n_530),
.Y(n_2080)
);

AOI22xp33_ASAP7_75t_L g2081 ( 
.A1(n_1971),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.Y(n_2081)
);

OR2x6_ASAP7_75t_L g2082 ( 
.A(n_1975),
.B(n_531),
.Y(n_2082)
);

BUFx2_ASAP7_75t_L g2083 ( 
.A(n_1909),
.Y(n_2083)
);

OAI21xp5_ASAP7_75t_L g2084 ( 
.A1(n_1857),
.A2(n_1861),
.B(n_1930),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1921),
.Y(n_2085)
);

AOI21xp5_ASAP7_75t_L g2086 ( 
.A1(n_1976),
.A2(n_533),
.B(n_532),
.Y(n_2086)
);

INVx3_ASAP7_75t_L g2087 ( 
.A(n_1966),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_SL g2088 ( 
.A(n_1978),
.B(n_1927),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1923),
.Y(n_2089)
);

AND2x4_ASAP7_75t_L g2090 ( 
.A(n_1867),
.B(n_534),
.Y(n_2090)
);

O2A1O1Ixp33_ASAP7_75t_L g2091 ( 
.A1(n_1869),
.A2(n_108),
.B(n_105),
.C(n_106),
.Y(n_2091)
);

INVxp67_ASAP7_75t_SL g2092 ( 
.A(n_1919),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_1916),
.Y(n_2093)
);

BUFx6f_ASAP7_75t_L g2094 ( 
.A(n_1873),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1901),
.B(n_106),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_1989),
.B(n_1986),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1983),
.Y(n_2097)
);

NOR2xp33_ASAP7_75t_L g2098 ( 
.A(n_2001),
.B(n_1913),
.Y(n_2098)
);

NAND3xp33_ASAP7_75t_SL g2099 ( 
.A(n_2063),
.B(n_1907),
.C(n_1895),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1995),
.Y(n_2100)
);

A2O1A1Ixp33_ASAP7_75t_L g2101 ( 
.A1(n_2042),
.A2(n_1863),
.B(n_1870),
.C(n_1862),
.Y(n_2101)
);

INVx6_ASAP7_75t_L g2102 ( 
.A(n_2048),
.Y(n_2102)
);

AND2x4_ASAP7_75t_L g2103 ( 
.A(n_2005),
.B(n_1999),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2053),
.Y(n_2104)
);

INVxp67_ASAP7_75t_L g2105 ( 
.A(n_1993),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_2050),
.B(n_1929),
.Y(n_2106)
);

BUFx3_ASAP7_75t_L g2107 ( 
.A(n_1988),
.Y(n_2107)
);

AOI22xp33_ASAP7_75t_L g2108 ( 
.A1(n_1981),
.A2(n_1875),
.B1(n_1880),
.B2(n_1872),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1984),
.B(n_1908),
.Y(n_2109)
);

AO32x2_ASAP7_75t_L g2110 ( 
.A1(n_2006),
.A2(n_1879),
.A3(n_1878),
.B1(n_1955),
.B2(n_1954),
.Y(n_2110)
);

AND2x4_ASAP7_75t_L g2111 ( 
.A(n_2005),
.B(n_2053),
.Y(n_2111)
);

NAND2x1_ASAP7_75t_L g2112 ( 
.A(n_1982),
.B(n_1883),
.Y(n_2112)
);

INVx3_ASAP7_75t_L g2113 ( 
.A(n_1985),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2025),
.Y(n_2114)
);

AO31x2_ASAP7_75t_L g2115 ( 
.A1(n_1996),
.A2(n_2008),
.A3(n_2019),
.B(n_2026),
.Y(n_2115)
);

OAI21x1_ASAP7_75t_L g2116 ( 
.A1(n_1990),
.A2(n_1911),
.B(n_1931),
.Y(n_2116)
);

NOR2xp33_ASAP7_75t_L g2117 ( 
.A(n_2022),
.B(n_1935),
.Y(n_2117)
);

AOI21xp5_ASAP7_75t_L g2118 ( 
.A1(n_2005),
.A2(n_1917),
.B(n_1958),
.Y(n_2118)
);

AOI21xp5_ASAP7_75t_L g2119 ( 
.A1(n_2054),
.A2(n_1898),
.B(n_1897),
.Y(n_2119)
);

INVx3_ASAP7_75t_L g2120 ( 
.A(n_1985),
.Y(n_2120)
);

AOI21xp5_ASAP7_75t_L g2121 ( 
.A1(n_2054),
.A2(n_1884),
.B(n_1887),
.Y(n_2121)
);

OAI21x1_ASAP7_75t_L g2122 ( 
.A1(n_2075),
.A2(n_1937),
.B(n_1936),
.Y(n_2122)
);

A2O1A1Ixp33_ASAP7_75t_L g2123 ( 
.A1(n_1997),
.A2(n_1940),
.B(n_1874),
.C(n_1925),
.Y(n_2123)
);

AOI21xp5_ASAP7_75t_L g2124 ( 
.A1(n_2054),
.A2(n_1944),
.B(n_1943),
.Y(n_2124)
);

AOI21x1_ASAP7_75t_L g2125 ( 
.A1(n_2000),
.A2(n_1942),
.B(n_1939),
.Y(n_2125)
);

BUFx4_ASAP7_75t_R g2126 ( 
.A(n_1991),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_2015),
.B(n_1961),
.Y(n_2127)
);

NOR2xp33_ASAP7_75t_L g2128 ( 
.A(n_2010),
.B(n_1962),
.Y(n_2128)
);

OAI21x1_ASAP7_75t_L g2129 ( 
.A1(n_2029),
.A2(n_1946),
.B(n_1945),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1979),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2003),
.Y(n_2131)
);

AOI21xp5_ASAP7_75t_L g2132 ( 
.A1(n_1998),
.A2(n_1949),
.B(n_1965),
.Y(n_2132)
);

AO32x2_ASAP7_75t_L g2133 ( 
.A1(n_2077),
.A2(n_1972),
.A3(n_1974),
.B1(n_1970),
.B2(n_1967),
.Y(n_2133)
);

O2A1O1Ixp5_ASAP7_75t_L g2134 ( 
.A1(n_2088),
.A2(n_111),
.B(n_109),
.C(n_110),
.Y(n_2134)
);

BUFx6f_ASAP7_75t_L g2135 ( 
.A(n_1994),
.Y(n_2135)
);

AO31x2_ASAP7_75t_L g2136 ( 
.A1(n_2002),
.A2(n_112),
.A3(n_109),
.B(n_111),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_2052),
.B(n_112),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2009),
.Y(n_2138)
);

INVxp67_ASAP7_75t_SL g2139 ( 
.A(n_2058),
.Y(n_2139)
);

OR2x2_ASAP7_75t_L g2140 ( 
.A(n_2007),
.B(n_113),
.Y(n_2140)
);

BUFx6f_ASAP7_75t_L g2141 ( 
.A(n_1994),
.Y(n_2141)
);

O2A1O1Ixp33_ASAP7_75t_SL g2142 ( 
.A1(n_2076),
.A2(n_2051),
.B(n_2079),
.C(n_2024),
.Y(n_2142)
);

AOI22xp33_ASAP7_75t_L g2143 ( 
.A1(n_2084),
.A2(n_117),
.B1(n_113),
.B2(n_114),
.Y(n_2143)
);

O2A1O1Ixp33_ASAP7_75t_L g2144 ( 
.A1(n_2091),
.A2(n_118),
.B(n_114),
.C(n_117),
.Y(n_2144)
);

OAI21xp5_ASAP7_75t_L g2145 ( 
.A1(n_2086),
.A2(n_538),
.B(n_537),
.Y(n_2145)
);

OAI21x1_ASAP7_75t_L g2146 ( 
.A1(n_2056),
.A2(n_542),
.B(n_540),
.Y(n_2146)
);

OAI21xp5_ASAP7_75t_L g2147 ( 
.A1(n_2016),
.A2(n_544),
.B(n_543),
.Y(n_2147)
);

AOI21xp5_ASAP7_75t_L g2148 ( 
.A1(n_2036),
.A2(n_547),
.B(n_545),
.Y(n_2148)
);

AOI21xp5_ASAP7_75t_L g2149 ( 
.A1(n_2036),
.A2(n_549),
.B(n_548),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2018),
.Y(n_2150)
);

AO31x2_ASAP7_75t_L g2151 ( 
.A1(n_2085),
.A2(n_121),
.A3(n_118),
.B(n_119),
.Y(n_2151)
);

OAI21x1_ASAP7_75t_L g2152 ( 
.A1(n_2065),
.A2(n_551),
.B(n_550),
.Y(n_2152)
);

HB1xp67_ASAP7_75t_L g2153 ( 
.A(n_1992),
.Y(n_2153)
);

HB1xp67_ASAP7_75t_L g2154 ( 
.A(n_2066),
.Y(n_2154)
);

OAI21xp5_ASAP7_75t_L g2155 ( 
.A1(n_2074),
.A2(n_553),
.B(n_552),
.Y(n_2155)
);

OAI22x1_ASAP7_75t_L g2156 ( 
.A1(n_2072),
.A2(n_122),
.B1(n_119),
.B2(n_121),
.Y(n_2156)
);

AO32x2_ASAP7_75t_L g2157 ( 
.A1(n_2017),
.A2(n_124),
.A3(n_122),
.B1(n_123),
.B2(n_125),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2011),
.Y(n_2158)
);

AO31x2_ASAP7_75t_L g2159 ( 
.A1(n_2085),
.A2(n_127),
.A3(n_124),
.B(n_126),
.Y(n_2159)
);

INVxp67_ASAP7_75t_L g2160 ( 
.A(n_2028),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_2052),
.B(n_126),
.Y(n_2161)
);

OAI211xp5_ASAP7_75t_L g2162 ( 
.A1(n_2099),
.A2(n_2081),
.B(n_2073),
.C(n_2061),
.Y(n_2162)
);

OAI21x1_ASAP7_75t_L g2163 ( 
.A1(n_2116),
.A2(n_2023),
.B(n_2049),
.Y(n_2163)
);

OAI21x1_ASAP7_75t_L g2164 ( 
.A1(n_2129),
.A2(n_2043),
.B(n_2012),
.Y(n_2164)
);

OR2x2_ASAP7_75t_L g2165 ( 
.A(n_2153),
.B(n_2046),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2104),
.Y(n_2166)
);

AO21x2_ASAP7_75t_L g2167 ( 
.A1(n_2132),
.A2(n_2031),
.B(n_2089),
.Y(n_2167)
);

OA21x2_ASAP7_75t_L g2168 ( 
.A1(n_2122),
.A2(n_2071),
.B(n_2013),
.Y(n_2168)
);

HB1xp67_ASAP7_75t_L g2169 ( 
.A(n_2154),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2097),
.Y(n_2170)
);

OAI21x1_ASAP7_75t_L g2171 ( 
.A1(n_2152),
.A2(n_2146),
.B(n_2100),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2114),
.Y(n_2172)
);

INVx5_ASAP7_75t_L g2173 ( 
.A(n_2102),
.Y(n_2173)
);

AOI21xp5_ASAP7_75t_L g2174 ( 
.A1(n_2147),
.A2(n_2062),
.B(n_2082),
.Y(n_2174)
);

BUFx12f_ASAP7_75t_L g2175 ( 
.A(n_2140),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_2130),
.Y(n_2176)
);

BUFx3_ASAP7_75t_L g2177 ( 
.A(n_2102),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_2096),
.B(n_1980),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_2138),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_2158),
.Y(n_2180)
);

HB1xp67_ASAP7_75t_L g2181 ( 
.A(n_2131),
.Y(n_2181)
);

OAI21x1_ASAP7_75t_L g2182 ( 
.A1(n_2118),
.A2(n_2012),
.B(n_2087),
.Y(n_2182)
);

OAI22xp33_ASAP7_75t_L g2183 ( 
.A1(n_2112),
.A2(n_2082),
.B1(n_2048),
.B2(n_2087),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2139),
.Y(n_2184)
);

AOI21x1_ASAP7_75t_L g2185 ( 
.A1(n_2125),
.A2(n_2124),
.B(n_2119),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_2150),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_2115),
.Y(n_2187)
);

AOI21x1_ASAP7_75t_L g2188 ( 
.A1(n_2125),
.A2(n_2014),
.B(n_2060),
.Y(n_2188)
);

AOI22xp5_ASAP7_75t_L g2189 ( 
.A1(n_2143),
.A2(n_2090),
.B1(n_2080),
.B2(n_2092),
.Y(n_2189)
);

AND2x4_ASAP7_75t_L g2190 ( 
.A(n_2111),
.B(n_2032),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_2115),
.Y(n_2191)
);

OR2x6_ASAP7_75t_L g2192 ( 
.A(n_2111),
.B(n_2032),
.Y(n_2192)
);

OAI21x1_ASAP7_75t_L g2193 ( 
.A1(n_2121),
.A2(n_2064),
.B(n_2055),
.Y(n_2193)
);

NOR2xp67_ASAP7_75t_L g2194 ( 
.A(n_2113),
.B(n_2048),
.Y(n_2194)
);

AOI21x1_ASAP7_75t_L g2195 ( 
.A1(n_2106),
.A2(n_2083),
.B(n_2033),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2151),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_2105),
.B(n_2127),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_2103),
.Y(n_2198)
);

AND2x4_ASAP7_75t_L g2199 ( 
.A(n_2103),
.B(n_2035),
.Y(n_2199)
);

OAI21xp5_ASAP7_75t_L g2200 ( 
.A1(n_2123),
.A2(n_2059),
.B(n_2078),
.Y(n_2200)
);

AOI21xp33_ASAP7_75t_SL g2201 ( 
.A1(n_2156),
.A2(n_2041),
.B(n_2020),
.Y(n_2201)
);

AOI221xp5_ASAP7_75t_L g2202 ( 
.A1(n_2144),
.A2(n_2095),
.B1(n_2027),
.B2(n_2047),
.C(n_2021),
.Y(n_2202)
);

BUFx2_ASAP7_75t_L g2203 ( 
.A(n_2120),
.Y(n_2203)
);

AOI22xp33_ASAP7_75t_SL g2204 ( 
.A1(n_2128),
.A2(n_2080),
.B1(n_2090),
.B2(n_2057),
.Y(n_2204)
);

OAI21x1_ASAP7_75t_L g2205 ( 
.A1(n_2155),
.A2(n_2055),
.B(n_2004),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2109),
.B(n_2069),
.Y(n_2206)
);

AOI22xp33_ASAP7_75t_L g2207 ( 
.A1(n_2174),
.A2(n_2145),
.B1(n_2094),
.B2(n_2098),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2166),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_2169),
.B(n_2165),
.Y(n_2209)
);

NAND2xp33_ASAP7_75t_SL g2210 ( 
.A(n_2167),
.B(n_2035),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2165),
.B(n_2181),
.Y(n_2211)
);

AND2x2_ASAP7_75t_L g2212 ( 
.A(n_2198),
.B(n_2160),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2166),
.Y(n_2213)
);

NOR2xp67_ASAP7_75t_L g2214 ( 
.A(n_2173),
.B(n_2107),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_2178),
.B(n_2137),
.Y(n_2215)
);

AOI21xp5_ASAP7_75t_L g2216 ( 
.A1(n_2167),
.A2(n_2142),
.B(n_2148),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2170),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_2198),
.B(n_2157),
.Y(n_2218)
);

INVx2_ASAP7_75t_SL g2219 ( 
.A(n_2177),
.Y(n_2219)
);

AOI21xp5_ASAP7_75t_L g2220 ( 
.A1(n_2167),
.A2(n_2149),
.B(n_2101),
.Y(n_2220)
);

INVx6_ASAP7_75t_L g2221 ( 
.A(n_2173),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_2197),
.B(n_2157),
.Y(n_2222)
);

OAI22xp5_ASAP7_75t_L g2223 ( 
.A1(n_2189),
.A2(n_2108),
.B1(n_2070),
.B2(n_2057),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2184),
.B(n_2161),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2170),
.Y(n_2225)
);

AOI22xp33_ASAP7_75t_SL g2226 ( 
.A1(n_2162),
.A2(n_2094),
.B1(n_2069),
.B2(n_2030),
.Y(n_2226)
);

HB1xp67_ASAP7_75t_L g2227 ( 
.A(n_2184),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_2179),
.Y(n_2228)
);

CKINVDCx5p33_ASAP7_75t_R g2229 ( 
.A(n_2175),
.Y(n_2229)
);

OAI22xp5_ASAP7_75t_L g2230 ( 
.A1(n_2189),
.A2(n_2038),
.B1(n_1987),
.B2(n_2039),
.Y(n_2230)
);

AND2x2_ASAP7_75t_SL g2231 ( 
.A(n_2190),
.B(n_2030),
.Y(n_2231)
);

BUFx2_ASAP7_75t_SL g2232 ( 
.A(n_2194),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_2172),
.B(n_2136),
.Y(n_2233)
);

OAI22xp5_ASAP7_75t_L g2234 ( 
.A1(n_2207),
.A2(n_2204),
.B1(n_2183),
.B2(n_2201),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2208),
.Y(n_2235)
);

OAI22xp5_ASAP7_75t_SL g2236 ( 
.A1(n_2229),
.A2(n_2175),
.B1(n_2117),
.B2(n_2200),
.Y(n_2236)
);

OA21x2_ASAP7_75t_L g2237 ( 
.A1(n_2216),
.A2(n_2191),
.B(n_2187),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_2211),
.B(n_2172),
.Y(n_2238)
);

INVx4_ASAP7_75t_L g2239 ( 
.A(n_2229),
.Y(n_2239)
);

AO21x2_ASAP7_75t_L g2240 ( 
.A1(n_2220),
.A2(n_2188),
.B(n_2185),
.Y(n_2240)
);

INVx3_ASAP7_75t_L g2241 ( 
.A(n_2221),
.Y(n_2241)
);

OAI221xp5_ASAP7_75t_L g2242 ( 
.A1(n_2226),
.A2(n_2201),
.B1(n_2202),
.B2(n_2185),
.C(n_2206),
.Y(n_2242)
);

OAI221xp5_ASAP7_75t_L g2243 ( 
.A1(n_2230),
.A2(n_2194),
.B1(n_2134),
.B2(n_2196),
.C(n_2191),
.Y(n_2243)
);

BUFx2_ASAP7_75t_L g2244 ( 
.A(n_2221),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2235),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_2238),
.B(n_2212),
.Y(n_2246)
);

AND2x4_ASAP7_75t_L g2247 ( 
.A(n_2239),
.B(n_2214),
.Y(n_2247)
);

OR2x6_ASAP7_75t_L g2248 ( 
.A(n_2239),
.B(n_2236),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_2234),
.B(n_2212),
.Y(n_2249)
);

XNOR2xp5_ASAP7_75t_L g2250 ( 
.A(n_2242),
.B(n_2223),
.Y(n_2250)
);

AND2x4_ASAP7_75t_L g2251 ( 
.A(n_2239),
.B(n_2219),
.Y(n_2251)
);

AND2x4_ASAP7_75t_L g2252 ( 
.A(n_2247),
.B(n_2241),
.Y(n_2252)
);

AND2x4_ASAP7_75t_L g2253 ( 
.A(n_2251),
.B(n_2241),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_2248),
.B(n_2241),
.Y(n_2254)
);

OAI22xp5_ASAP7_75t_L g2255 ( 
.A1(n_2250),
.A2(n_2243),
.B1(n_2221),
.B2(n_2244),
.Y(n_2255)
);

AOI22xp33_ASAP7_75t_L g2256 ( 
.A1(n_2250),
.A2(n_2240),
.B1(n_2094),
.B2(n_2210),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_2249),
.B(n_2222),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_2248),
.B(n_2244),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2245),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2246),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2245),
.Y(n_2261)
);

NAND4xp25_ASAP7_75t_L g2262 ( 
.A(n_2255),
.B(n_2256),
.C(n_2258),
.D(n_2257),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2260),
.B(n_2222),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_2254),
.B(n_2219),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2253),
.B(n_2218),
.Y(n_2265)
);

NOR3xp33_ASAP7_75t_L g2266 ( 
.A(n_2252),
.B(n_2210),
.C(n_2193),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_2252),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2260),
.B(n_2235),
.Y(n_2268)
);

NAND3xp33_ASAP7_75t_L g2269 ( 
.A(n_2256),
.B(n_2233),
.C(n_2196),
.Y(n_2269)
);

AOI22xp33_ASAP7_75t_L g2270 ( 
.A1(n_2252),
.A2(n_2240),
.B1(n_2221),
.B2(n_2205),
.Y(n_2270)
);

OAI21xp5_ASAP7_75t_L g2271 ( 
.A1(n_2253),
.A2(n_2205),
.B(n_2193),
.Y(n_2271)
);

AOI22xp33_ASAP7_75t_L g2272 ( 
.A1(n_2259),
.A2(n_2240),
.B1(n_2187),
.B2(n_2231),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2268),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2267),
.B(n_2261),
.Y(n_2274)
);

NAND2x1_ASAP7_75t_L g2275 ( 
.A(n_2265),
.B(n_2261),
.Y(n_2275)
);

AND2x4_ASAP7_75t_L g2276 ( 
.A(n_2264),
.B(n_2177),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2263),
.B(n_2262),
.Y(n_2277)
);

HB1xp67_ASAP7_75t_L g2278 ( 
.A(n_2262),
.Y(n_2278)
);

AND2x2_ASAP7_75t_L g2279 ( 
.A(n_2270),
.B(n_2197),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_2269),
.B(n_2218),
.Y(n_2280)
);

BUFx3_ASAP7_75t_L g2281 ( 
.A(n_2272),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_2276),
.B(n_2271),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_2275),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_2276),
.B(n_2266),
.Y(n_2284)
);

OR2x2_ASAP7_75t_L g2285 ( 
.A(n_2277),
.B(n_2278),
.Y(n_2285)
);

AND2x2_ASAP7_75t_L g2286 ( 
.A(n_2283),
.B(n_2273),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_2285),
.B(n_2277),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2284),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2282),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_2286),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2289),
.B(n_2274),
.Y(n_2291)
);

AND2x4_ASAP7_75t_L g2292 ( 
.A(n_2286),
.B(n_2288),
.Y(n_2292)
);

OAI221xp5_ASAP7_75t_L g2293 ( 
.A1(n_2287),
.A2(n_2281),
.B1(n_2280),
.B2(n_2279),
.C(n_2232),
.Y(n_2293)
);

NOR2xp33_ASAP7_75t_L g2294 ( 
.A(n_2288),
.B(n_2034),
.Y(n_2294)
);

INVx3_ASAP7_75t_L g2295 ( 
.A(n_2286),
.Y(n_2295)
);

OR2x2_ASAP7_75t_L g2296 ( 
.A(n_2295),
.B(n_2290),
.Y(n_2296)
);

INVx2_ASAP7_75t_SL g2297 ( 
.A(n_2292),
.Y(n_2297)
);

INVx2_ASAP7_75t_SL g2298 ( 
.A(n_2292),
.Y(n_2298)
);

AND2x4_ASAP7_75t_L g2299 ( 
.A(n_2294),
.B(n_2209),
.Y(n_2299)
);

NOR2xp33_ASAP7_75t_L g2300 ( 
.A(n_2291),
.B(n_2126),
.Y(n_2300)
);

INVx1_ASAP7_75t_SL g2301 ( 
.A(n_2293),
.Y(n_2301)
);

INVxp67_ASAP7_75t_L g2302 ( 
.A(n_2294),
.Y(n_2302)
);

NOR2xp33_ASAP7_75t_L g2303 ( 
.A(n_2294),
.B(n_2215),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_2295),
.B(n_2227),
.Y(n_2304)
);

AOI22xp33_ASAP7_75t_L g2305 ( 
.A1(n_2293),
.A2(n_2232),
.B1(n_2177),
.B2(n_2173),
.Y(n_2305)
);

NOR2xp33_ASAP7_75t_SL g2306 ( 
.A(n_2297),
.B(n_2173),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2298),
.B(n_2217),
.Y(n_2307)
);

OAI221xp5_ASAP7_75t_SL g2308 ( 
.A1(n_2305),
.A2(n_2192),
.B1(n_2037),
.B2(n_2068),
.C(n_2067),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_2296),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2304),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2300),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2301),
.B(n_2299),
.Y(n_2312)
);

AOI32xp33_ASAP7_75t_L g2313 ( 
.A1(n_2303),
.A2(n_2040),
.A3(n_2157),
.B1(n_2182),
.B2(n_2203),
.Y(n_2313)
);

AND2x4_ASAP7_75t_L g2314 ( 
.A(n_2302),
.B(n_2224),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2297),
.B(n_2225),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2297),
.Y(n_2316)
);

NAND2x1p5_ASAP7_75t_L g2317 ( 
.A(n_2297),
.B(n_2040),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2297),
.B(n_2213),
.Y(n_2318)
);

OAI21xp33_ASAP7_75t_L g2319 ( 
.A1(n_2316),
.A2(n_2195),
.B(n_2231),
.Y(n_2319)
);

OAI21xp5_ASAP7_75t_L g2320 ( 
.A1(n_2312),
.A2(n_2182),
.B(n_2164),
.Y(n_2320)
);

OAI21xp33_ASAP7_75t_L g2321 ( 
.A1(n_2306),
.A2(n_2195),
.B(n_2188),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2309),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2311),
.B(n_2237),
.Y(n_2323)
);

OAI22xp5_ASAP7_75t_L g2324 ( 
.A1(n_2308),
.A2(n_2173),
.B1(n_2237),
.B2(n_2069),
.Y(n_2324)
);

OR2x2_ASAP7_75t_L g2325 ( 
.A(n_2307),
.B(n_2136),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2315),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2314),
.B(n_2317),
.Y(n_2327)
);

HB1xp67_ASAP7_75t_L g2328 ( 
.A(n_2318),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2310),
.Y(n_2329)
);

O2A1O1Ixp33_ASAP7_75t_L g2330 ( 
.A1(n_2313),
.A2(n_129),
.B(n_127),
.C(n_128),
.Y(n_2330)
);

OAI21xp33_ASAP7_75t_SL g2331 ( 
.A1(n_2316),
.A2(n_2164),
.B(n_2192),
.Y(n_2331)
);

AOI22xp33_ASAP7_75t_L g2332 ( 
.A1(n_2316),
.A2(n_2173),
.B1(n_2168),
.B2(n_2237),
.Y(n_2332)
);

INVxp33_ASAP7_75t_L g2333 ( 
.A(n_2316),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2322),
.Y(n_2334)
);

AOI222xp33_ASAP7_75t_L g2335 ( 
.A1(n_2333),
.A2(n_2093),
.B1(n_131),
.B2(n_133),
.C1(n_129),
.C2(n_130),
.Y(n_2335)
);

INVxp67_ASAP7_75t_L g2336 ( 
.A(n_2327),
.Y(n_2336)
);

OAI21xp5_ASAP7_75t_L g2337 ( 
.A1(n_2330),
.A2(n_2163),
.B(n_2171),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2328),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2329),
.B(n_2203),
.Y(n_2339)
);

INVx3_ASAP7_75t_L g2340 ( 
.A(n_2325),
.Y(n_2340)
);

AOI21xp5_ASAP7_75t_L g2341 ( 
.A1(n_2323),
.A2(n_2168),
.B(n_130),
.Y(n_2341)
);

O2A1O1Ixp33_ASAP7_75t_SL g2342 ( 
.A1(n_2326),
.A2(n_134),
.B(n_132),
.C(n_133),
.Y(n_2342)
);

AND2x2_ASAP7_75t_L g2343 ( 
.A(n_2319),
.B(n_2190),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2324),
.Y(n_2344)
);

INVxp33_ASAP7_75t_L g2345 ( 
.A(n_2321),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2331),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2320),
.Y(n_2347)
);

OAI21x1_ASAP7_75t_L g2348 ( 
.A1(n_2346),
.A2(n_2332),
.B(n_2171),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2342),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2339),
.B(n_2168),
.Y(n_2350)
);

AOI211x1_ASAP7_75t_L g2351 ( 
.A1(n_2341),
.A2(n_136),
.B(n_132),
.C(n_135),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2334),
.B(n_2168),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_2336),
.B(n_2151),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_2335),
.B(n_2159),
.Y(n_2354)
);

O2A1O1Ixp33_ASAP7_75t_L g2355 ( 
.A1(n_2338),
.A2(n_138),
.B(n_135),
.C(n_137),
.Y(n_2355)
);

OAI21xp33_ASAP7_75t_L g2356 ( 
.A1(n_2345),
.A2(n_2192),
.B(n_2190),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2340),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2340),
.Y(n_2358)
);

NOR2xp33_ASAP7_75t_R g2359 ( 
.A(n_2344),
.B(n_137),
.Y(n_2359)
);

NOR3xp33_ASAP7_75t_L g2360 ( 
.A(n_2347),
.B(n_139),
.C(n_140),
.Y(n_2360)
);

AOI221xp5_ASAP7_75t_L g2361 ( 
.A1(n_2343),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.C(n_142),
.Y(n_2361)
);

AOI22xp5_ASAP7_75t_L g2362 ( 
.A1(n_2337),
.A2(n_2190),
.B1(n_2199),
.B2(n_2192),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2339),
.Y(n_2363)
);

AOI22xp5_ASAP7_75t_L g2364 ( 
.A1(n_2336),
.A2(n_2199),
.B1(n_2192),
.B2(n_2228),
.Y(n_2364)
);

OAI22xp5_ASAP7_75t_L g2365 ( 
.A1(n_2336),
.A2(n_2044),
.B1(n_2228),
.B2(n_2030),
.Y(n_2365)
);

OR2x2_ASAP7_75t_L g2366 ( 
.A(n_2334),
.B(n_141),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2342),
.Y(n_2367)
);

O2A1O1Ixp33_ASAP7_75t_SL g2368 ( 
.A1(n_2346),
.A2(n_144),
.B(n_142),
.C(n_143),
.Y(n_2368)
);

O2A1O1Ixp5_ASAP7_75t_L g2369 ( 
.A1(n_2346),
.A2(n_146),
.B(n_144),
.C(n_145),
.Y(n_2369)
);

INVx5_ASAP7_75t_L g2370 ( 
.A(n_2363),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2366),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2349),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_2367),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2368),
.Y(n_2374)
);

BUFx2_ASAP7_75t_L g2375 ( 
.A(n_2359),
.Y(n_2375)
);

INVx2_ASAP7_75t_SL g2376 ( 
.A(n_2357),
.Y(n_2376)
);

INVxp33_ASAP7_75t_L g2377 ( 
.A(n_2360),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2369),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2358),
.Y(n_2379)
);

NOR2xp33_ASAP7_75t_L g2380 ( 
.A(n_2355),
.B(n_145),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2351),
.Y(n_2381)
);

INVxp33_ASAP7_75t_SL g2382 ( 
.A(n_2361),
.Y(n_2382)
);

INVxp67_ASAP7_75t_L g2383 ( 
.A(n_2353),
.Y(n_2383)
);

BUFx2_ASAP7_75t_L g2384 ( 
.A(n_2348),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2354),
.Y(n_2385)
);

NAND2x1_ASAP7_75t_SL g2386 ( 
.A(n_2364),
.B(n_146),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2352),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2356),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2350),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2365),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_2362),
.Y(n_2391)
);

INVx8_ASAP7_75t_L g2392 ( 
.A(n_2357),
.Y(n_2392)
);

INVx2_ASAP7_75t_SL g2393 ( 
.A(n_2349),
.Y(n_2393)
);

INVx5_ASAP7_75t_L g2394 ( 
.A(n_2363),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2366),
.Y(n_2395)
);

BUFx2_ASAP7_75t_L g2396 ( 
.A(n_2349),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2366),
.Y(n_2397)
);

INVx1_ASAP7_75t_SL g2398 ( 
.A(n_2349),
.Y(n_2398)
);

NOR2xp33_ASAP7_75t_L g2399 ( 
.A(n_2349),
.B(n_147),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2366),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2366),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2366),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2366),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2366),
.Y(n_2404)
);

NOR2xp33_ASAP7_75t_L g2405 ( 
.A(n_2349),
.B(n_148),
.Y(n_2405)
);

INVx1_ASAP7_75t_SL g2406 ( 
.A(n_2349),
.Y(n_2406)
);

NOR2xp33_ASAP7_75t_L g2407 ( 
.A(n_2398),
.B(n_149),
.Y(n_2407)
);

OAI22xp5_ASAP7_75t_L g2408 ( 
.A1(n_2406),
.A2(n_2045),
.B1(n_2179),
.B2(n_2176),
.Y(n_2408)
);

INVx2_ASAP7_75t_L g2409 ( 
.A(n_2392),
.Y(n_2409)
);

NOR2xp33_ASAP7_75t_L g2410 ( 
.A(n_2370),
.B(n_149),
.Y(n_2410)
);

NOR5xp2_ASAP7_75t_L g2411 ( 
.A(n_2383),
.B(n_152),
.C(n_150),
.D(n_151),
.E(n_153),
.Y(n_2411)
);

AOI211xp5_ASAP7_75t_L g2412 ( 
.A1(n_2399),
.A2(n_153),
.B(n_150),
.C(n_152),
.Y(n_2412)
);

OAI211xp5_ASAP7_75t_L g2413 ( 
.A1(n_2405),
.A2(n_156),
.B(n_154),
.C(n_155),
.Y(n_2413)
);

OAI31xp33_ASAP7_75t_L g2414 ( 
.A1(n_2374),
.A2(n_2396),
.A3(n_2378),
.B(n_2372),
.Y(n_2414)
);

CKINVDCx16_ASAP7_75t_R g2415 ( 
.A(n_2375),
.Y(n_2415)
);

OR2x2_ASAP7_75t_L g2416 ( 
.A(n_2393),
.B(n_154),
.Y(n_2416)
);

AOI221xp5_ASAP7_75t_L g2417 ( 
.A1(n_2379),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.C(n_158),
.Y(n_2417)
);

OAI22xp5_ASAP7_75t_L g2418 ( 
.A1(n_2376),
.A2(n_2045),
.B1(n_2176),
.B2(n_2199),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_2392),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2384),
.Y(n_2420)
);

OAI221xp5_ASAP7_75t_SL g2421 ( 
.A1(n_2373),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.C(n_160),
.Y(n_2421)
);

AOI221xp5_ASAP7_75t_L g2422 ( 
.A1(n_2380),
.A2(n_163),
.B1(n_161),
.B2(n_162),
.C(n_164),
.Y(n_2422)
);

AOI21xp33_ASAP7_75t_L g2423 ( 
.A1(n_2377),
.A2(n_161),
.B(n_162),
.Y(n_2423)
);

OAI221xp5_ASAP7_75t_L g2424 ( 
.A1(n_2388),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.C(n_169),
.Y(n_2424)
);

A2O1A1Ixp33_ASAP7_75t_SL g2425 ( 
.A1(n_2371),
.A2(n_169),
.B(n_165),
.C(n_166),
.Y(n_2425)
);

AOI22xp33_ASAP7_75t_SL g2426 ( 
.A1(n_2370),
.A2(n_2394),
.B1(n_2382),
.B2(n_2381),
.Y(n_2426)
);

AOI221xp5_ASAP7_75t_L g2427 ( 
.A1(n_2385),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.C(n_173),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2370),
.Y(n_2428)
);

OR2x2_ASAP7_75t_L g2429 ( 
.A(n_2395),
.B(n_170),
.Y(n_2429)
);

OAI21x1_ASAP7_75t_L g2430 ( 
.A1(n_2386),
.A2(n_2163),
.B(n_171),
.Y(n_2430)
);

XNOR2xp5_ASAP7_75t_L g2431 ( 
.A(n_2397),
.B(n_2400),
.Y(n_2431)
);

AOI322xp5_ASAP7_75t_L g2432 ( 
.A1(n_2391),
.A2(n_2159),
.A3(n_2110),
.B1(n_2199),
.B2(n_175),
.C1(n_176),
.C2(n_177),
.Y(n_2432)
);

AOI211xp5_ASAP7_75t_SL g2433 ( 
.A1(n_2401),
.A2(n_174),
.B(n_172),
.C(n_173),
.Y(n_2433)
);

BUFx4f_ASAP7_75t_SL g2434 ( 
.A(n_2402),
.Y(n_2434)
);

A2O1A1Ixp33_ASAP7_75t_L g2435 ( 
.A1(n_2390),
.A2(n_178),
.B(n_176),
.C(n_177),
.Y(n_2435)
);

AOI21xp5_ASAP7_75t_L g2436 ( 
.A1(n_2394),
.A2(n_178),
.B(n_179),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2394),
.Y(n_2437)
);

OAI22xp5_ASAP7_75t_L g2438 ( 
.A1(n_2403),
.A2(n_2045),
.B1(n_2186),
.B2(n_2180),
.Y(n_2438)
);

BUFx2_ASAP7_75t_L g2439 ( 
.A(n_2404),
.Y(n_2439)
);

NOR2xp67_ASAP7_75t_L g2440 ( 
.A(n_2389),
.B(n_179),
.Y(n_2440)
);

AOI21xp33_ASAP7_75t_SL g2441 ( 
.A1(n_2387),
.A2(n_180),
.B(n_181),
.Y(n_2441)
);

OAI22xp5_ASAP7_75t_L g2442 ( 
.A1(n_2398),
.A2(n_2186),
.B1(n_2180),
.B2(n_2135),
.Y(n_2442)
);

NOR2xp33_ASAP7_75t_L g2443 ( 
.A(n_2398),
.B(n_180),
.Y(n_2443)
);

OR2x2_ASAP7_75t_L g2444 ( 
.A(n_2374),
.B(n_181),
.Y(n_2444)
);

AOI211xp5_ASAP7_75t_L g2445 ( 
.A1(n_2407),
.A2(n_186),
.B(n_184),
.C(n_185),
.Y(n_2445)
);

AOI221xp5_ASAP7_75t_SL g2446 ( 
.A1(n_2420),
.A2(n_187),
.B1(n_184),
.B2(n_185),
.C(n_188),
.Y(n_2446)
);

AOI221xp5_ASAP7_75t_L g2447 ( 
.A1(n_2443),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.C(n_190),
.Y(n_2447)
);

AOI221xp5_ASAP7_75t_SL g2448 ( 
.A1(n_2428),
.A2(n_191),
.B1(n_189),
.B2(n_190),
.C(n_192),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2433),
.B(n_2440),
.Y(n_2449)
);

O2A1O1Ixp33_ASAP7_75t_L g2450 ( 
.A1(n_2425),
.A2(n_193),
.B(n_191),
.C(n_192),
.Y(n_2450)
);

OAI211xp5_ASAP7_75t_L g2451 ( 
.A1(n_2414),
.A2(n_195),
.B(n_193),
.C(n_194),
.Y(n_2451)
);

AOI221xp5_ASAP7_75t_L g2452 ( 
.A1(n_2410),
.A2(n_197),
.B1(n_194),
.B2(n_196),
.C(n_198),
.Y(n_2452)
);

NOR2x1_ASAP7_75t_L g2453 ( 
.A(n_2437),
.B(n_196),
.Y(n_2453)
);

AOI222xp33_ASAP7_75t_L g2454 ( 
.A1(n_2434),
.A2(n_199),
.B1(n_201),
.B2(n_197),
.C1(n_198),
.C2(n_200),
.Y(n_2454)
);

OAI211xp5_ASAP7_75t_L g2455 ( 
.A1(n_2426),
.A2(n_201),
.B(n_199),
.C(n_200),
.Y(n_2455)
);

NOR2xp33_ASAP7_75t_L g2456 ( 
.A(n_2415),
.B(n_2444),
.Y(n_2456)
);

NOR4xp25_ASAP7_75t_L g2457 ( 
.A(n_2409),
.B(n_204),
.C(n_202),
.D(n_203),
.Y(n_2457)
);

INVxp67_ASAP7_75t_L g2458 ( 
.A(n_2429),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2416),
.Y(n_2459)
);

OAI21xp5_ASAP7_75t_L g2460 ( 
.A1(n_2431),
.A2(n_202),
.B(n_203),
.Y(n_2460)
);

OAI211xp5_ASAP7_75t_SL g2461 ( 
.A1(n_2419),
.A2(n_207),
.B(n_204),
.C(n_206),
.Y(n_2461)
);

AOI211xp5_ASAP7_75t_L g2462 ( 
.A1(n_2441),
.A2(n_209),
.B(n_206),
.C(n_208),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2439),
.Y(n_2463)
);

AOI221xp5_ASAP7_75t_L g2464 ( 
.A1(n_2427),
.A2(n_210),
.B1(n_208),
.B2(n_209),
.C(n_212),
.Y(n_2464)
);

NOR2xp33_ASAP7_75t_R g2465 ( 
.A(n_2412),
.B(n_210),
.Y(n_2465)
);

O2A1O1Ixp33_ASAP7_75t_L g2466 ( 
.A1(n_2435),
.A2(n_214),
.B(n_212),
.C(n_213),
.Y(n_2466)
);

AOI221x1_ASAP7_75t_SL g2467 ( 
.A1(n_2423),
.A2(n_216),
.B1(n_214),
.B2(n_215),
.C(n_217),
.Y(n_2467)
);

AOI21xp5_ASAP7_75t_L g2468 ( 
.A1(n_2436),
.A2(n_216),
.B(n_218),
.Y(n_2468)
);

AOI221xp5_ASAP7_75t_L g2469 ( 
.A1(n_2408),
.A2(n_220),
.B1(n_218),
.B2(n_219),
.C(n_221),
.Y(n_2469)
);

NOR3xp33_ASAP7_75t_L g2470 ( 
.A(n_2422),
.B(n_2424),
.C(n_2413),
.Y(n_2470)
);

A2O1A1Ixp33_ASAP7_75t_L g2471 ( 
.A1(n_2411),
.A2(n_2430),
.B(n_2421),
.C(n_2417),
.Y(n_2471)
);

NAND4xp25_ASAP7_75t_SL g2472 ( 
.A(n_2432),
.B(n_2442),
.C(n_2418),
.D(n_2438),
.Y(n_2472)
);

AOI211xp5_ASAP7_75t_L g2473 ( 
.A1(n_2407),
.A2(n_221),
.B(n_219),
.C(n_220),
.Y(n_2473)
);

AOI321xp33_ASAP7_75t_L g2474 ( 
.A1(n_2409),
.A2(n_222),
.A3(n_223),
.B1(n_224),
.B2(n_225),
.C(n_226),
.Y(n_2474)
);

NOR3xp33_ASAP7_75t_L g2475 ( 
.A(n_2415),
.B(n_222),
.C(n_223),
.Y(n_2475)
);

AOI221x1_ASAP7_75t_L g2476 ( 
.A1(n_2420),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.C(n_227),
.Y(n_2476)
);

AOI22xp5_ASAP7_75t_L g2477 ( 
.A1(n_2415),
.A2(n_2141),
.B1(n_2135),
.B2(n_230),
.Y(n_2477)
);

AOI21xp33_ASAP7_75t_L g2478 ( 
.A1(n_2420),
.A2(n_228),
.B(n_229),
.Y(n_2478)
);

O2A1O1Ixp33_ASAP7_75t_L g2479 ( 
.A1(n_2425),
.A2(n_230),
.B(n_228),
.C(n_229),
.Y(n_2479)
);

AOI211xp5_ASAP7_75t_L g2480 ( 
.A1(n_2407),
.A2(n_234),
.B(n_232),
.C(n_233),
.Y(n_2480)
);

AOI211xp5_ASAP7_75t_L g2481 ( 
.A1(n_2407),
.A2(n_234),
.B(n_232),
.C(n_233),
.Y(n_2481)
);

OAI21xp5_ASAP7_75t_SL g2482 ( 
.A1(n_2414),
.A2(n_235),
.B(n_236),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2433),
.B(n_235),
.Y(n_2483)
);

AOI211xp5_ASAP7_75t_L g2484 ( 
.A1(n_2407),
.A2(n_239),
.B(n_237),
.C(n_238),
.Y(n_2484)
);

AOI211xp5_ASAP7_75t_L g2485 ( 
.A1(n_2407),
.A2(n_240),
.B(n_238),
.C(n_239),
.Y(n_2485)
);

AND3x1_ASAP7_75t_L g2486 ( 
.A(n_2414),
.B(n_240),
.C(n_241),
.Y(n_2486)
);

OAI221xp5_ASAP7_75t_SL g2487 ( 
.A1(n_2414),
.A2(n_244),
.B1(n_242),
.B2(n_243),
.C(n_245),
.Y(n_2487)
);

OAI21xp33_ASAP7_75t_SL g2488 ( 
.A1(n_2414),
.A2(n_242),
.B(n_244),
.Y(n_2488)
);

AOI21xp5_ASAP7_75t_L g2489 ( 
.A1(n_2428),
.A2(n_245),
.B(n_246),
.Y(n_2489)
);

NAND4xp25_ASAP7_75t_L g2490 ( 
.A(n_2414),
.B(n_248),
.C(n_246),
.D(n_247),
.Y(n_2490)
);

OAI211xp5_ASAP7_75t_L g2491 ( 
.A1(n_2414),
.A2(n_249),
.B(n_247),
.C(n_248),
.Y(n_2491)
);

OAI221xp5_ASAP7_75t_L g2492 ( 
.A1(n_2414),
.A2(n_251),
.B1(n_249),
.B2(n_250),
.C(n_252),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_2433),
.B(n_250),
.Y(n_2493)
);

AOI222xp33_ASAP7_75t_L g2494 ( 
.A1(n_2434),
.A2(n_251),
.B1(n_253),
.B2(n_254),
.C1(n_256),
.C2(n_257),
.Y(n_2494)
);

NAND3x1_ASAP7_75t_L g2495 ( 
.A(n_2414),
.B(n_253),
.C(n_256),
.Y(n_2495)
);

OAI21xp33_ASAP7_75t_L g2496 ( 
.A1(n_2431),
.A2(n_2141),
.B(n_258),
.Y(n_2496)
);

AOI211xp5_ASAP7_75t_L g2497 ( 
.A1(n_2407),
.A2(n_261),
.B(n_259),
.C(n_260),
.Y(n_2497)
);

O2A1O1Ixp33_ASAP7_75t_L g2498 ( 
.A1(n_2425),
.A2(n_261),
.B(n_259),
.C(n_260),
.Y(n_2498)
);

OR2x2_ASAP7_75t_L g2499 ( 
.A(n_2444),
.B(n_262),
.Y(n_2499)
);

AOI31xp33_ASAP7_75t_L g2500 ( 
.A1(n_2426),
.A2(n_264),
.A3(n_262),
.B(n_263),
.Y(n_2500)
);

AOI211xp5_ASAP7_75t_L g2501 ( 
.A1(n_2407),
.A2(n_265),
.B(n_263),
.C(n_264),
.Y(n_2501)
);

OAI221xp5_ASAP7_75t_L g2502 ( 
.A1(n_2414),
.A2(n_267),
.B1(n_265),
.B2(n_266),
.C(n_268),
.Y(n_2502)
);

AOI22xp5_ASAP7_75t_L g2503 ( 
.A1(n_2415),
.A2(n_269),
.B1(n_267),
.B2(n_268),
.Y(n_2503)
);

OAI31xp33_ASAP7_75t_L g2504 ( 
.A1(n_2425),
.A2(n_271),
.A3(n_269),
.B(n_270),
.Y(n_2504)
);

NAND3xp33_ASAP7_75t_L g2505 ( 
.A(n_2414),
.B(n_270),
.C(n_271),
.Y(n_2505)
);

OR2x2_ASAP7_75t_L g2506 ( 
.A(n_2444),
.B(n_272),
.Y(n_2506)
);

XNOR2x1_ASAP7_75t_L g2507 ( 
.A(n_2486),
.B(n_273),
.Y(n_2507)
);

AOI22xp33_ASAP7_75t_SL g2508 ( 
.A1(n_2463),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2453),
.Y(n_2509)
);

BUFx6f_ASAP7_75t_L g2510 ( 
.A(n_2456),
.Y(n_2510)
);

AOI22xp5_ASAP7_75t_L g2511 ( 
.A1(n_2496),
.A2(n_277),
.B1(n_274),
.B2(n_276),
.Y(n_2511)
);

OAI21xp5_ASAP7_75t_L g2512 ( 
.A1(n_2495),
.A2(n_276),
.B(n_277),
.Y(n_2512)
);

AOI211x1_ASAP7_75t_SL g2513 ( 
.A1(n_2505),
.A2(n_280),
.B(n_278),
.C(n_279),
.Y(n_2513)
);

AOI22xp5_ASAP7_75t_SL g2514 ( 
.A1(n_2449),
.A2(n_281),
.B1(n_279),
.B2(n_280),
.Y(n_2514)
);

OAI21xp5_ASAP7_75t_SL g2515 ( 
.A1(n_2482),
.A2(n_281),
.B(n_282),
.Y(n_2515)
);

XNOR2x1_ASAP7_75t_L g2516 ( 
.A(n_2499),
.B(n_282),
.Y(n_2516)
);

AOI22xp5_ASAP7_75t_L g2517 ( 
.A1(n_2470),
.A2(n_285),
.B1(n_283),
.B2(n_284),
.Y(n_2517)
);

NOR3xp33_ASAP7_75t_SL g2518 ( 
.A(n_2451),
.B(n_285),
.C(n_286),
.Y(n_2518)
);

OAI22xp5_ASAP7_75t_L g2519 ( 
.A1(n_2477),
.A2(n_288),
.B1(n_286),
.B2(n_287),
.Y(n_2519)
);

AOI22xp5_ASAP7_75t_L g2520 ( 
.A1(n_2490),
.A2(n_291),
.B1(n_287),
.B2(n_290),
.Y(n_2520)
);

AOI221xp5_ASAP7_75t_L g2521 ( 
.A1(n_2492),
.A2(n_290),
.B1(n_291),
.B2(n_292),
.C(n_293),
.Y(n_2521)
);

OAI222xp33_ASAP7_75t_L g2522 ( 
.A1(n_2487),
.A2(n_292),
.B1(n_294),
.B2(n_295),
.C1(n_296),
.C2(n_297),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_2457),
.B(n_294),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2448),
.B(n_295),
.Y(n_2524)
);

CKINVDCx20_ASAP7_75t_R g2525 ( 
.A(n_2465),
.Y(n_2525)
);

OAI211xp5_ASAP7_75t_L g2526 ( 
.A1(n_2488),
.A2(n_298),
.B(n_296),
.C(n_297),
.Y(n_2526)
);

AOI21xp5_ASAP7_75t_L g2527 ( 
.A1(n_2483),
.A2(n_299),
.B(n_300),
.Y(n_2527)
);

AOI222xp33_ASAP7_75t_L g2528 ( 
.A1(n_2491),
.A2(n_2502),
.B1(n_2458),
.B2(n_2459),
.C1(n_2471),
.C2(n_2493),
.Y(n_2528)
);

AOI221xp5_ASAP7_75t_L g2529 ( 
.A1(n_2450),
.A2(n_299),
.B1(n_301),
.B2(n_302),
.C(n_303),
.Y(n_2529)
);

NAND4xp25_ASAP7_75t_SL g2530 ( 
.A(n_2479),
.B(n_304),
.C(n_302),
.D(n_303),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2506),
.Y(n_2531)
);

NOR3x1_ASAP7_75t_L g2532 ( 
.A(n_2455),
.B(n_304),
.C(n_305),
.Y(n_2532)
);

O2A1O1Ixp33_ASAP7_75t_L g2533 ( 
.A1(n_2500),
.A2(n_307),
.B(n_305),
.C(n_306),
.Y(n_2533)
);

NOR4xp25_ASAP7_75t_SL g2534 ( 
.A(n_2464),
.B(n_308),
.C(n_306),
.D(n_307),
.Y(n_2534)
);

AOI221xp5_ASAP7_75t_L g2535 ( 
.A1(n_2498),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.C(n_311),
.Y(n_2535)
);

INVx1_ASAP7_75t_SL g2536 ( 
.A(n_2489),
.Y(n_2536)
);

OAI211xp5_ASAP7_75t_SL g2537 ( 
.A1(n_2504),
.A2(n_313),
.B(n_310),
.C(n_312),
.Y(n_2537)
);

AOI221xp5_ASAP7_75t_L g2538 ( 
.A1(n_2466),
.A2(n_312),
.B1(n_313),
.B2(n_314),
.C(n_315),
.Y(n_2538)
);

OAI222xp33_ASAP7_75t_L g2539 ( 
.A1(n_2468),
.A2(n_315),
.B1(n_316),
.B2(n_317),
.C1(n_318),
.C2(n_319),
.Y(n_2539)
);

OAI221xp5_ASAP7_75t_L g2540 ( 
.A1(n_2467),
.A2(n_2469),
.B1(n_2446),
.B2(n_2462),
.C(n_2460),
.Y(n_2540)
);

OAI211xp5_ASAP7_75t_SL g2541 ( 
.A1(n_2445),
.A2(n_318),
.B(n_316),
.C(n_317),
.Y(n_2541)
);

AOI21xp33_ASAP7_75t_L g2542 ( 
.A1(n_2461),
.A2(n_319),
.B(n_320),
.Y(n_2542)
);

NAND3xp33_ASAP7_75t_L g2543 ( 
.A(n_2473),
.B(n_321),
.C(n_322),
.Y(n_2543)
);

AOI211x1_ASAP7_75t_L g2544 ( 
.A1(n_2472),
.A2(n_324),
.B(n_322),
.C(n_323),
.Y(n_2544)
);

NAND4xp25_ASAP7_75t_L g2545 ( 
.A(n_2476),
.B(n_326),
.C(n_323),
.D(n_325),
.Y(n_2545)
);

AOI221xp5_ASAP7_75t_L g2546 ( 
.A1(n_2478),
.A2(n_326),
.B1(n_327),
.B2(n_328),
.C(n_329),
.Y(n_2546)
);

AOI211xp5_ASAP7_75t_L g2547 ( 
.A1(n_2475),
.A2(n_330),
.B(n_327),
.C(n_328),
.Y(n_2547)
);

OAI211xp5_ASAP7_75t_SL g2548 ( 
.A1(n_2480),
.A2(n_333),
.B(n_331),
.C(n_332),
.Y(n_2548)
);

AO22x2_ASAP7_75t_L g2549 ( 
.A1(n_2481),
.A2(n_334),
.B1(n_332),
.B2(n_333),
.Y(n_2549)
);

XNOR2xp5_ASAP7_75t_L g2550 ( 
.A(n_2484),
.B(n_2485),
.Y(n_2550)
);

AOI21xp33_ASAP7_75t_L g2551 ( 
.A1(n_2454),
.A2(n_335),
.B(n_336),
.Y(n_2551)
);

AOI221x1_ASAP7_75t_L g2552 ( 
.A1(n_2497),
.A2(n_335),
.B1(n_336),
.B2(n_337),
.C(n_338),
.Y(n_2552)
);

AOI221xp5_ASAP7_75t_L g2553 ( 
.A1(n_2447),
.A2(n_337),
.B1(n_340),
.B2(n_341),
.C(n_342),
.Y(n_2553)
);

A2O1A1Ixp33_ASAP7_75t_L g2554 ( 
.A1(n_2501),
.A2(n_344),
.B(n_341),
.C(n_343),
.Y(n_2554)
);

AND4x1_ASAP7_75t_L g2555 ( 
.A(n_2494),
.B(n_347),
.C(n_343),
.D(n_345),
.Y(n_2555)
);

AOI21xp33_ASAP7_75t_SL g2556 ( 
.A1(n_2503),
.A2(n_345),
.B(n_347),
.Y(n_2556)
);

OAI22xp33_ASAP7_75t_L g2557 ( 
.A1(n_2452),
.A2(n_350),
.B1(n_348),
.B2(n_349),
.Y(n_2557)
);

AOI21xp33_ASAP7_75t_SL g2558 ( 
.A1(n_2474),
.A2(n_348),
.B(n_349),
.Y(n_2558)
);

AOI211xp5_ASAP7_75t_L g2559 ( 
.A1(n_2487),
.A2(n_353),
.B(n_351),
.C(n_352),
.Y(n_2559)
);

OAI221xp5_ASAP7_75t_L g2560 ( 
.A1(n_2504),
.A2(n_351),
.B1(n_352),
.B2(n_353),
.C(n_354),
.Y(n_2560)
);

OAI211xp5_ASAP7_75t_L g2561 ( 
.A1(n_2488),
.A2(n_354),
.B(n_355),
.C(n_356),
.Y(n_2561)
);

AOI221xp5_ASAP7_75t_L g2562 ( 
.A1(n_2492),
.A2(n_355),
.B1(n_357),
.B2(n_358),
.C(n_359),
.Y(n_2562)
);

NOR2xp33_ASAP7_75t_L g2563 ( 
.A(n_2490),
.B(n_358),
.Y(n_2563)
);

HB1xp67_ASAP7_75t_L g2564 ( 
.A(n_2453),
.Y(n_2564)
);

O2A1O1Ixp33_ASAP7_75t_SL g2565 ( 
.A1(n_2471),
.A2(n_359),
.B(n_360),
.C(n_361),
.Y(n_2565)
);

AOI211xp5_ASAP7_75t_L g2566 ( 
.A1(n_2487),
.A2(n_360),
.B(n_361),
.C(n_362),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_2499),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2453),
.Y(n_2568)
);

AOI221xp5_ASAP7_75t_L g2569 ( 
.A1(n_2492),
.A2(n_362),
.B1(n_363),
.B2(n_364),
.C(n_365),
.Y(n_2569)
);

INVx2_ASAP7_75t_SL g2570 ( 
.A(n_2453),
.Y(n_2570)
);

AOI221xp5_ASAP7_75t_L g2571 ( 
.A1(n_2492),
.A2(n_363),
.B1(n_364),
.B2(n_365),
.C(n_366),
.Y(n_2571)
);

AOI221xp5_ASAP7_75t_L g2572 ( 
.A1(n_2492),
.A2(n_366),
.B1(n_367),
.B2(n_368),
.C(n_369),
.Y(n_2572)
);

CKINVDCx5p33_ASAP7_75t_R g2573 ( 
.A(n_2456),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2549),
.Y(n_2574)
);

AOI22xp5_ASAP7_75t_L g2575 ( 
.A1(n_2573),
.A2(n_2563),
.B1(n_2530),
.B2(n_2525),
.Y(n_2575)
);

OAI22xp33_ASAP7_75t_SL g2576 ( 
.A1(n_2523),
.A2(n_367),
.B1(n_369),
.B2(n_370),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2549),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2507),
.Y(n_2578)
);

AO22x1_ASAP7_75t_L g2579 ( 
.A1(n_2512),
.A2(n_370),
.B1(n_372),
.B2(n_373),
.Y(n_2579)
);

AOI22xp5_ASAP7_75t_L g2580 ( 
.A1(n_2510),
.A2(n_372),
.B1(n_373),
.B2(n_374),
.Y(n_2580)
);

NAND3xp33_ASAP7_75t_SL g2581 ( 
.A(n_2534),
.B(n_374),
.C(n_375),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_SL g2582 ( 
.A(n_2510),
.B(n_375),
.Y(n_2582)
);

INVxp67_ASAP7_75t_SL g2583 ( 
.A(n_2514),
.Y(n_2583)
);

HB1xp67_ASAP7_75t_L g2584 ( 
.A(n_2564),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2565),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2516),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2524),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2544),
.Y(n_2588)
);

NOR2x1_ASAP7_75t_L g2589 ( 
.A(n_2509),
.B(n_2568),
.Y(n_2589)
);

AOI22xp5_ASAP7_75t_SL g2590 ( 
.A1(n_2570),
.A2(n_377),
.B1(n_378),
.B2(n_379),
.Y(n_2590)
);

AOI22xp5_ASAP7_75t_L g2591 ( 
.A1(n_2510),
.A2(n_377),
.B1(n_378),
.B2(n_379),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2533),
.Y(n_2592)
);

INVx2_ASAP7_75t_L g2593 ( 
.A(n_2532),
.Y(n_2593)
);

OAI21xp5_ASAP7_75t_SL g2594 ( 
.A1(n_2515),
.A2(n_380),
.B(n_381),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2555),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2526),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2561),
.Y(n_2597)
);

AOI22xp5_ASAP7_75t_L g2598 ( 
.A1(n_2537),
.A2(n_380),
.B1(n_381),
.B2(n_382),
.Y(n_2598)
);

INVx1_ASAP7_75t_SL g2599 ( 
.A(n_2536),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2520),
.Y(n_2600)
);

INVx2_ASAP7_75t_L g2601 ( 
.A(n_2567),
.Y(n_2601)
);

AOI22xp5_ASAP7_75t_L g2602 ( 
.A1(n_2541),
.A2(n_383),
.B1(n_384),
.B2(n_385),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2545),
.Y(n_2603)
);

NOR2x1_ASAP7_75t_L g2604 ( 
.A(n_2539),
.B(n_383),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_L g2605 ( 
.A(n_2558),
.B(n_2529),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2518),
.Y(n_2606)
);

AOI22xp5_ASAP7_75t_L g2607 ( 
.A1(n_2548),
.A2(n_384),
.B1(n_385),
.B2(n_386),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2560),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2511),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_2535),
.B(n_386),
.Y(n_2610)
);

HB1xp67_ASAP7_75t_L g2611 ( 
.A(n_2513),
.Y(n_2611)
);

INVx2_ASAP7_75t_L g2612 ( 
.A(n_2531),
.Y(n_2612)
);

AOI22xp33_ASAP7_75t_L g2613 ( 
.A1(n_2543),
.A2(n_387),
.B1(n_388),
.B2(n_389),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2552),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2554),
.Y(n_2615)
);

NOR2xp67_ASAP7_75t_L g2616 ( 
.A(n_2517),
.B(n_387),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2550),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2547),
.Y(n_2618)
);

AOI22xp5_ASAP7_75t_L g2619 ( 
.A1(n_2519),
.A2(n_388),
.B1(n_389),
.B2(n_390),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2559),
.Y(n_2620)
);

AOI22xp5_ASAP7_75t_L g2621 ( 
.A1(n_2528),
.A2(n_390),
.B1(n_391),
.B2(n_392),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2566),
.Y(n_2622)
);

INVxp67_ASAP7_75t_SL g2623 ( 
.A(n_2508),
.Y(n_2623)
);

AND2x4_ASAP7_75t_L g2624 ( 
.A(n_2527),
.B(n_391),
.Y(n_2624)
);

AOI22xp5_ASAP7_75t_SL g2625 ( 
.A1(n_2522),
.A2(n_392),
.B1(n_393),
.B2(n_394),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_2540),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2556),
.Y(n_2627)
);

BUFx2_ASAP7_75t_L g2628 ( 
.A(n_2546),
.Y(n_2628)
);

HB1xp67_ASAP7_75t_L g2629 ( 
.A(n_2538),
.Y(n_2629)
);

AOI22xp5_ASAP7_75t_L g2630 ( 
.A1(n_2521),
.A2(n_393),
.B1(n_395),
.B2(n_396),
.Y(n_2630)
);

INVx2_ASAP7_75t_L g2631 ( 
.A(n_2542),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2557),
.Y(n_2632)
);

AND2x2_ASAP7_75t_L g2633 ( 
.A(n_2551),
.B(n_2110),
.Y(n_2633)
);

INVx2_ASAP7_75t_L g2634 ( 
.A(n_2572),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2562),
.Y(n_2635)
);

NOR2x1_ASAP7_75t_L g2636 ( 
.A(n_2581),
.B(n_2569),
.Y(n_2636)
);

NAND2x1_ASAP7_75t_L g2637 ( 
.A(n_2585),
.B(n_2571),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2625),
.Y(n_2638)
);

NOR2x1_ASAP7_75t_L g2639 ( 
.A(n_2614),
.B(n_2553),
.Y(n_2639)
);

BUFx6f_ASAP7_75t_L g2640 ( 
.A(n_2612),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2582),
.Y(n_2641)
);

OR2x2_ASAP7_75t_L g2642 ( 
.A(n_2588),
.B(n_395),
.Y(n_2642)
);

NAND4xp25_ASAP7_75t_L g2643 ( 
.A(n_2598),
.B(n_396),
.C(n_397),
.D(n_398),
.Y(n_2643)
);

NAND4xp25_ASAP7_75t_L g2644 ( 
.A(n_2575),
.B(n_397),
.C(n_398),
.D(n_399),
.Y(n_2644)
);

NOR2x1_ASAP7_75t_L g2645 ( 
.A(n_2589),
.B(n_399),
.Y(n_2645)
);

NAND4xp75_ASAP7_75t_L g2646 ( 
.A(n_2589),
.B(n_400),
.C(n_401),
.D(n_402),
.Y(n_2646)
);

INVx1_ASAP7_75t_SL g2647 ( 
.A(n_2590),
.Y(n_2647)
);

BUFx6f_ASAP7_75t_L g2648 ( 
.A(n_2601),
.Y(n_2648)
);

OAI22xp33_ASAP7_75t_SL g2649 ( 
.A1(n_2574),
.A2(n_400),
.B1(n_401),
.B2(n_402),
.Y(n_2649)
);

AND2x2_ASAP7_75t_L g2650 ( 
.A(n_2583),
.B(n_2110),
.Y(n_2650)
);

OR2x2_ASAP7_75t_L g2651 ( 
.A(n_2621),
.B(n_403),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2579),
.Y(n_2652)
);

NAND4xp75_ASAP7_75t_L g2653 ( 
.A(n_2596),
.B(n_403),
.C(n_404),
.D(n_405),
.Y(n_2653)
);

NOR4xp75_ASAP7_75t_SL g2654 ( 
.A(n_2605),
.B(n_405),
.C(n_406),
.D(n_407),
.Y(n_2654)
);

INVxp67_ASAP7_75t_L g2655 ( 
.A(n_2584),
.Y(n_2655)
);

NAND4xp75_ASAP7_75t_L g2656 ( 
.A(n_2597),
.B(n_406),
.C(n_407),
.D(n_409),
.Y(n_2656)
);

NOR2xp33_ASAP7_75t_R g2657 ( 
.A(n_2606),
.B(n_409),
.Y(n_2657)
);

XNOR2x1_ASAP7_75t_L g2658 ( 
.A(n_2604),
.B(n_410),
.Y(n_2658)
);

OR2x2_ASAP7_75t_L g2659 ( 
.A(n_2595),
.B(n_411),
.Y(n_2659)
);

BUFx2_ASAP7_75t_L g2660 ( 
.A(n_2577),
.Y(n_2660)
);

OR2x2_ASAP7_75t_L g2661 ( 
.A(n_2594),
.B(n_411),
.Y(n_2661)
);

NAND5xp2_ASAP7_75t_L g2662 ( 
.A(n_2617),
.B(n_412),
.C(n_413),
.D(n_414),
.E(n_415),
.Y(n_2662)
);

OR2x2_ASAP7_75t_L g2663 ( 
.A(n_2593),
.B(n_413),
.Y(n_2663)
);

OAI22xp5_ASAP7_75t_L g2664 ( 
.A1(n_2602),
.A2(n_414),
.B1(n_415),
.B2(n_416),
.Y(n_2664)
);

INVxp33_ASAP7_75t_SL g2665 ( 
.A(n_2629),
.Y(n_2665)
);

OR2x2_ASAP7_75t_L g2666 ( 
.A(n_2607),
.B(n_416),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_SL g2667 ( 
.A(n_2576),
.B(n_417),
.Y(n_2667)
);

INVx1_ASAP7_75t_SL g2668 ( 
.A(n_2624),
.Y(n_2668)
);

AOI21xp5_ASAP7_75t_L g2669 ( 
.A1(n_2610),
.A2(n_417),
.B(n_418),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_2613),
.B(n_419),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_L g2671 ( 
.A(n_2624),
.B(n_419),
.Y(n_2671)
);

OR5x1_ASAP7_75t_L g2672 ( 
.A(n_2623),
.B(n_421),
.C(n_422),
.D(n_423),
.E(n_424),
.Y(n_2672)
);

OAI211xp5_ASAP7_75t_SL g2673 ( 
.A1(n_2627),
.A2(n_421),
.B(n_423),
.C(n_424),
.Y(n_2673)
);

AND2x2_ASAP7_75t_L g2674 ( 
.A(n_2611),
.B(n_2133),
.Y(n_2674)
);

BUFx2_ASAP7_75t_L g2675 ( 
.A(n_2603),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2616),
.Y(n_2676)
);

NOR2xp33_ASAP7_75t_L g2677 ( 
.A(n_2592),
.B(n_425),
.Y(n_2677)
);

NAND4xp25_ASAP7_75t_L g2678 ( 
.A(n_2630),
.B(n_425),
.C(n_426),
.D(n_427),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_2619),
.B(n_427),
.Y(n_2679)
);

NOR3xp33_ASAP7_75t_SL g2680 ( 
.A(n_2667),
.B(n_2622),
.C(n_2620),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_SL g2681 ( 
.A(n_2654),
.B(n_2626),
.Y(n_2681)
);

NOR2xp33_ASAP7_75t_R g2682 ( 
.A(n_2638),
.B(n_2578),
.Y(n_2682)
);

NOR2xp33_ASAP7_75t_R g2683 ( 
.A(n_2648),
.B(n_2615),
.Y(n_2683)
);

NOR2xp33_ASAP7_75t_R g2684 ( 
.A(n_2648),
.B(n_2632),
.Y(n_2684)
);

NOR2xp33_ASAP7_75t_R g2685 ( 
.A(n_2640),
.B(n_2586),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_SL g2686 ( 
.A(n_2640),
.B(n_2599),
.Y(n_2686)
);

NOR2xp33_ASAP7_75t_R g2687 ( 
.A(n_2652),
.B(n_2600),
.Y(n_2687)
);

NOR2xp33_ASAP7_75t_R g2688 ( 
.A(n_2642),
.B(n_2587),
.Y(n_2688)
);

NAND3xp33_ASAP7_75t_L g2689 ( 
.A(n_2655),
.B(n_2645),
.C(n_2660),
.Y(n_2689)
);

NAND3xp33_ASAP7_75t_L g2690 ( 
.A(n_2658),
.B(n_2608),
.C(n_2635),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_SL g2691 ( 
.A(n_2665),
.B(n_2631),
.Y(n_2691)
);

NAND2xp33_ASAP7_75t_SL g2692 ( 
.A(n_2657),
.B(n_2609),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_SL g2693 ( 
.A(n_2649),
.B(n_2634),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_SL g2694 ( 
.A(n_2664),
.B(n_2618),
.Y(n_2694)
);

NOR2xp33_ASAP7_75t_R g2695 ( 
.A(n_2671),
.B(n_2628),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_SL g2696 ( 
.A(n_2647),
.B(n_2580),
.Y(n_2696)
);

NAND2xp33_ASAP7_75t_SL g2697 ( 
.A(n_2661),
.B(n_2633),
.Y(n_2697)
);

NOR2xp33_ASAP7_75t_R g2698 ( 
.A(n_2641),
.B(n_2591),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_L g2699 ( 
.A(n_2677),
.B(n_2646),
.Y(n_2699)
);

NAND3xp33_ASAP7_75t_L g2700 ( 
.A(n_2669),
.B(n_428),
.C(n_429),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_L g2701 ( 
.A(n_2663),
.B(n_428),
.Y(n_2701)
);

NAND3xp33_ASAP7_75t_SL g2702 ( 
.A(n_2668),
.B(n_429),
.C(n_430),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_SL g2703 ( 
.A(n_2675),
.B(n_430),
.Y(n_2703)
);

NAND3xp33_ASAP7_75t_SL g2704 ( 
.A(n_2637),
.B(n_431),
.C(n_432),
.Y(n_2704)
);

NOR2xp33_ASAP7_75t_R g2705 ( 
.A(n_2676),
.B(n_431),
.Y(n_2705)
);

NAND2xp33_ASAP7_75t_SL g2706 ( 
.A(n_2651),
.B(n_2666),
.Y(n_2706)
);

NOR2xp33_ASAP7_75t_R g2707 ( 
.A(n_2670),
.B(n_432),
.Y(n_2707)
);

NAND2xp33_ASAP7_75t_SL g2708 ( 
.A(n_2679),
.B(n_433),
.Y(n_2708)
);

NOR2xp33_ASAP7_75t_R g2709 ( 
.A(n_2659),
.B(n_433),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2653),
.B(n_434),
.Y(n_2710)
);

NOR2xp33_ASAP7_75t_R g2711 ( 
.A(n_2650),
.B(n_435),
.Y(n_2711)
);

NAND2xp33_ASAP7_75t_SL g2712 ( 
.A(n_2672),
.B(n_435),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_SL g2713 ( 
.A(n_2639),
.B(n_437),
.Y(n_2713)
);

NAND2xp33_ASAP7_75t_SL g2714 ( 
.A(n_2674),
.B(n_437),
.Y(n_2714)
);

NOR2xp33_ASAP7_75t_R g2715 ( 
.A(n_2662),
.B(n_438),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_SL g2716 ( 
.A(n_2636),
.B(n_438),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2656),
.B(n_440),
.Y(n_2717)
);

OR3x1_ASAP7_75t_L g2718 ( 
.A(n_2704),
.B(n_2643),
.C(n_2678),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2710),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2717),
.Y(n_2720)
);

OAI211xp5_ASAP7_75t_L g2721 ( 
.A1(n_2709),
.A2(n_2644),
.B(n_2673),
.C(n_444),
.Y(n_2721)
);

NAND4xp25_ASAP7_75t_SL g2722 ( 
.A(n_2689),
.B(n_442),
.C(n_443),
.D(n_444),
.Y(n_2722)
);

O2A1O1Ixp33_ASAP7_75t_L g2723 ( 
.A1(n_2713),
.A2(n_2716),
.B(n_2686),
.C(n_2681),
.Y(n_2723)
);

BUFx2_ASAP7_75t_L g2724 ( 
.A(n_2705),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2701),
.Y(n_2725)
);

AND2x2_ASAP7_75t_SL g2726 ( 
.A(n_2699),
.B(n_443),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2703),
.Y(n_2727)
);

NOR3xp33_ASAP7_75t_L g2728 ( 
.A(n_2691),
.B(n_445),
.C(n_446),
.Y(n_2728)
);

A2O1A1Ixp33_ASAP7_75t_L g2729 ( 
.A1(n_2714),
.A2(n_446),
.B(n_447),
.C(n_448),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_L g2730 ( 
.A(n_2711),
.B(n_447),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2700),
.Y(n_2731)
);

XNOR2xp5_ASAP7_75t_L g2732 ( 
.A(n_2690),
.B(n_449),
.Y(n_2732)
);

AOI22xp5_ASAP7_75t_L g2733 ( 
.A1(n_2692),
.A2(n_449),
.B1(n_450),
.B2(n_451),
.Y(n_2733)
);

INVx3_ASAP7_75t_L g2734 ( 
.A(n_2684),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2712),
.Y(n_2735)
);

INVx3_ASAP7_75t_L g2736 ( 
.A(n_2708),
.Y(n_2736)
);

NAND3xp33_ASAP7_75t_SL g2737 ( 
.A(n_2682),
.B(n_450),
.C(n_451),
.Y(n_2737)
);

OAI21xp5_ASAP7_75t_SL g2738 ( 
.A1(n_2702),
.A2(n_452),
.B(n_453),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_2693),
.Y(n_2739)
);

AOI221xp5_ASAP7_75t_L g2740 ( 
.A1(n_2735),
.A2(n_2697),
.B1(n_2706),
.B2(n_2696),
.C(n_2687),
.Y(n_2740)
);

AOI22xp33_ASAP7_75t_L g2741 ( 
.A1(n_2739),
.A2(n_2715),
.B1(n_2685),
.B2(n_2683),
.Y(n_2741)
);

OAI222xp33_ASAP7_75t_L g2742 ( 
.A1(n_2734),
.A2(n_2694),
.B1(n_2680),
.B2(n_2695),
.C1(n_2698),
.C2(n_2688),
.Y(n_2742)
);

INVx1_ASAP7_75t_SL g2743 ( 
.A(n_2726),
.Y(n_2743)
);

CKINVDCx20_ASAP7_75t_R g2744 ( 
.A(n_2724),
.Y(n_2744)
);

XOR2xp5_ASAP7_75t_L g2745 ( 
.A(n_2732),
.B(n_2707),
.Y(n_2745)
);

AND2x2_ASAP7_75t_L g2746 ( 
.A(n_2728),
.B(n_2133),
.Y(n_2746)
);

AOI221xp5_ASAP7_75t_L g2747 ( 
.A1(n_2738),
.A2(n_452),
.B1(n_453),
.B2(n_454),
.C(n_455),
.Y(n_2747)
);

CKINVDCx5p33_ASAP7_75t_R g2748 ( 
.A(n_2725),
.Y(n_2748)
);

NOR3xp33_ASAP7_75t_L g2749 ( 
.A(n_2723),
.B(n_454),
.C(n_456),
.Y(n_2749)
);

NOR3xp33_ASAP7_75t_L g2750 ( 
.A(n_2736),
.B(n_456),
.C(n_458),
.Y(n_2750)
);

CKINVDCx20_ASAP7_75t_R g2751 ( 
.A(n_2727),
.Y(n_2751)
);

OR2x2_ASAP7_75t_L g2752 ( 
.A(n_2737),
.B(n_458),
.Y(n_2752)
);

BUFx2_ASAP7_75t_L g2753 ( 
.A(n_2729),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2752),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_L g2755 ( 
.A(n_2749),
.B(n_2730),
.Y(n_2755)
);

NOR2xp33_ASAP7_75t_L g2756 ( 
.A(n_2742),
.B(n_2721),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2747),
.B(n_2733),
.Y(n_2757)
);

NOR2xp33_ASAP7_75t_L g2758 ( 
.A(n_2743),
.B(n_2731),
.Y(n_2758)
);

XNOR2xp5_ASAP7_75t_L g2759 ( 
.A(n_2745),
.B(n_2718),
.Y(n_2759)
);

OR2x2_ASAP7_75t_L g2760 ( 
.A(n_2753),
.B(n_2722),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2751),
.Y(n_2761)
);

INVx2_ASAP7_75t_L g2762 ( 
.A(n_2744),
.Y(n_2762)
);

OAI21x1_ASAP7_75t_L g2763 ( 
.A1(n_2762),
.A2(n_2741),
.B(n_2740),
.Y(n_2763)
);

NOR2xp33_ASAP7_75t_L g2764 ( 
.A(n_2761),
.B(n_2719),
.Y(n_2764)
);

NOR2x1_ASAP7_75t_L g2765 ( 
.A(n_2760),
.B(n_2720),
.Y(n_2765)
);

INVx2_ASAP7_75t_SL g2766 ( 
.A(n_2759),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2755),
.Y(n_2767)
);

AOI22xp5_ASAP7_75t_L g2768 ( 
.A1(n_2758),
.A2(n_2748),
.B1(n_2750),
.B2(n_2746),
.Y(n_2768)
);

AOI22xp5_ASAP7_75t_L g2769 ( 
.A1(n_2766),
.A2(n_2756),
.B1(n_2754),
.B2(n_2757),
.Y(n_2769)
);

CKINVDCx5p33_ASAP7_75t_R g2770 ( 
.A(n_2768),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2763),
.Y(n_2771)
);

INVx3_ASAP7_75t_L g2772 ( 
.A(n_2767),
.Y(n_2772)
);

AOI31xp33_ASAP7_75t_L g2773 ( 
.A1(n_2771),
.A2(n_2765),
.A3(n_2764),
.B(n_461),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2773),
.Y(n_2774)
);

XNOR2x1_ASAP7_75t_SL g2775 ( 
.A(n_2774),
.B(n_2772),
.Y(n_2775)
);

AOI222xp33_ASAP7_75t_L g2776 ( 
.A1(n_2775),
.A2(n_2770),
.B1(n_2769),
.B2(n_461),
.C1(n_462),
.C2(n_463),
.Y(n_2776)
);

NOR2x1_ASAP7_75t_SL g2777 ( 
.A(n_2776),
.B(n_459),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2777),
.Y(n_2778)
);

AOI221xp5_ASAP7_75t_L g2779 ( 
.A1(n_2778),
.A2(n_459),
.B1(n_460),
.B2(n_462),
.C(n_464),
.Y(n_2779)
);

AOI22xp5_ASAP7_75t_L g2780 ( 
.A1(n_2779),
.A2(n_460),
.B1(n_465),
.B2(n_466),
.Y(n_2780)
);

AOI22xp33_ASAP7_75t_L g2781 ( 
.A1(n_2780),
.A2(n_465),
.B1(n_466),
.B2(n_467),
.Y(n_2781)
);


endmodule