module fake_jpeg_25683_n_125 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_125);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_36),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx6f_ASAP7_75t_SL g46 ( 
.A(n_5),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_11),
.B(n_13),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_20),
.B(n_38),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_49),
.Y(n_70)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_52),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_59),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_0),
.Y(n_72)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_43),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_55),
.B(n_39),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_68),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_62),
.B(n_40),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_70),
.A2(n_19),
.B(n_37),
.Y(n_89)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_3),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_1),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_62),
.B(n_53),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_1),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_76),
.A2(n_48),
.B1(n_45),
.B2(n_42),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_84),
.B1(n_85),
.B2(n_91),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_82),
.Y(n_101)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_41),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_83),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_51),
.B1(n_49),
.B2(n_54),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_51),
.B1(n_24),
.B2(n_25),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_43),
.Y(n_86)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_90),
.C(n_3),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_75),
.B(n_2),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_79),
.A2(n_74),
.B1(n_66),
.B2(n_26),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_96),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_77),
.A2(n_17),
.B1(n_34),
.B2(n_32),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_4),
.Y(n_102)
);

A2O1A1O1Ixp25_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_12),
.B(n_31),
.C(n_30),
.D(n_7),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_100),
.B(n_21),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_102),
.A2(n_103),
.B(n_106),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_87),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_98),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_104),
.A2(n_107),
.B1(n_108),
.B2(n_6),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_4),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_95),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_92),
.C(n_94),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_111),
.Y(n_116)
);

HAxp5_ASAP7_75t_SL g111 ( 
.A(n_103),
.B(n_87),
.CON(n_111),
.SN(n_111)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_113),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_105),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_117),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_118),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_119),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_116),
.C(n_115),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_114),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_111),
.C(n_9),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_10),
.B(n_27),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_28),
.Y(n_125)
);


endmodule