module fake_jpeg_26084_n_291 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_291);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_291;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_40),
.B(n_46),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

HAxp5_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_45),
.CON(n_53),
.SN(n_53)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_9),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_25),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_23),
.A2(n_0),
.B(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_32),
.Y(n_52)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_33),
.B1(n_36),
.B2(n_32),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_51),
.A2(n_57),
.B1(n_58),
.B2(n_66),
.Y(n_84)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_52),
.A2(n_72),
.B(n_11),
.Y(n_109)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_56),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_33),
.B1(n_38),
.B2(n_29),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_33),
.B1(n_38),
.B2(n_29),
.Y(n_58)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_30),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_74),
.Y(n_94)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_22),
.B1(n_21),
.B2(n_26),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_47),
.Y(n_67)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_42),
.A2(n_22),
.B1(n_26),
.B2(n_20),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_68),
.A2(n_70),
.B1(n_78),
.B2(n_23),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_40),
.A2(n_28),
.B1(n_25),
.B2(n_20),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_27),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_73),
.B(n_76),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_30),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_46),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_SL g77 ( 
.A1(n_44),
.A2(n_27),
.B(n_20),
.Y(n_77)
);

NAND2xp33_ASAP7_75t_SL g96 ( 
.A(n_77),
.B(n_37),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_46),
.A2(n_28),
.B1(n_25),
.B2(n_31),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_35),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_23),
.Y(n_99)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_53),
.A2(n_23),
.B1(n_35),
.B2(n_34),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_82),
.B(n_98),
.Y(n_135)
);

HAxp5_ASAP7_75t_SL g85 ( 
.A(n_61),
.B(n_52),
.CON(n_85),
.SN(n_85)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_85),
.A2(n_113),
.B(n_94),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_53),
.A2(n_31),
.B1(n_28),
.B2(n_34),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_88),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_92),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_76),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_56),
.A2(n_31),
.B1(n_35),
.B2(n_12),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_95),
.A2(n_96),
.B1(n_101),
.B2(n_109),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_105),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_54),
.A2(n_11),
.B1(n_17),
.B2(n_16),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_62),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_104),
.Y(n_132)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_37),
.Y(n_105)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_74),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_110),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_49),
.A2(n_0),
.B(n_1),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_34),
.C(n_19),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_59),
.C(n_64),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_63),
.B(n_37),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_65),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_118),
.A2(n_128),
.B(n_4),
.Y(n_168)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_121),
.B(n_143),
.Y(n_178)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_125),
.B(n_127),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_140),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_108),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_105),
.A2(n_0),
.B(n_2),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_129),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_90),
.A2(n_49),
.B1(n_80),
.B2(n_71),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_133),
.B(n_136),
.Y(n_158)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_141),
.Y(n_177)
);

AND2x6_ASAP7_75t_L g136 ( 
.A(n_85),
.B(n_13),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_59),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_147),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_99),
.A2(n_60),
.B1(n_50),
.B2(n_67),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_140),
.A2(n_144),
.B1(n_114),
.B2(n_86),
.Y(n_148)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_84),
.A2(n_67),
.B1(n_75),
.B2(n_19),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_145),
.B(n_2),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_83),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_146),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_88),
.B(n_113),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_148),
.A2(n_149),
.B1(n_152),
.B2(n_153),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_82),
.B1(n_114),
.B2(n_106),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_156),
.C(n_169),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_147),
.A2(n_82),
.B1(n_116),
.B2(n_106),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_82),
.B1(n_104),
.B2(n_97),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_132),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_155),
.B(n_166),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_112),
.C(n_89),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_100),
.B1(n_97),
.B2(n_103),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_157),
.A2(n_159),
.B1(n_160),
.B2(n_162),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_103),
.B1(n_93),
.B2(n_115),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_144),
.A2(n_139),
.B1(n_125),
.B2(n_130),
.Y(n_160)
);

AO21x1_ASAP7_75t_L g161 ( 
.A1(n_130),
.A2(n_19),
.B(n_115),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_161),
.A2(n_123),
.B(n_121),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_118),
.A2(n_93),
.B1(n_115),
.B2(n_107),
.Y(n_162)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_2),
.B(n_17),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_164),
.A2(n_170),
.B(n_175),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_133),
.A2(n_131),
.B1(n_126),
.B2(n_137),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_168),
.A2(n_8),
.B(n_10),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_4),
.C(n_5),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_141),
.A2(n_4),
.B(n_6),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_128),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_174)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_136),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_146),
.A2(n_124),
.B1(n_142),
.B2(n_127),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_176),
.B(n_142),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_124),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_179),
.B(n_183),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_145),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_185),
.A2(n_188),
.B(n_189),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_168),
.A2(n_134),
.B(n_123),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_L g191 ( 
.A1(n_173),
.A2(n_12),
.B(n_13),
.Y(n_191)
);

NOR4xp25_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_163),
.C(n_187),
.D(n_184),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_143),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_201),
.C(n_180),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_167),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_194),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_177),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_198),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_121),
.Y(n_196)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_196),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_120),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_204),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_120),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_202),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_167),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_200),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_127),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_161),
.Y(n_202)
);

BUFx24_ASAP7_75t_SL g203 ( 
.A(n_158),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_164),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_158),
.A2(n_129),
.B(n_15),
.Y(n_204)
);

BUFx24_ASAP7_75t_SL g241 ( 
.A(n_206),
.Y(n_241)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_197),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_211),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_190),
.A2(n_153),
.B1(n_149),
.B2(n_148),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_209),
.A2(n_224),
.B1(n_225),
.B2(n_186),
.Y(n_226)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_193),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_181),
.A2(n_152),
.B1(n_151),
.B2(n_157),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_215),
.A2(n_223),
.B1(n_189),
.B2(n_198),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_221),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_176),
.C(n_172),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_222),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_170),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_180),
.B(n_172),
.C(n_160),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_181),
.A2(n_154),
.B1(n_159),
.B2(n_177),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_192),
.A2(n_175),
.B1(n_174),
.B2(n_154),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_190),
.A2(n_161),
.B1(n_178),
.B2(n_169),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_226),
.A2(n_227),
.B1(n_231),
.B2(n_239),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_209),
.A2(n_186),
.B1(n_196),
.B2(n_201),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_217),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_228),
.B(n_229),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_212),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_230),
.B(n_235),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_225),
.A2(n_196),
.B1(n_202),
.B2(n_179),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_234),
.C(n_208),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_208),
.B(n_204),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_212),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_240),
.B1(n_242),
.B2(n_205),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_224),
.A2(n_187),
.B1(n_182),
.B2(n_200),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_205),
.A2(n_182),
.B1(n_178),
.B2(n_188),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_223),
.A2(n_119),
.B1(n_167),
.B2(n_16),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_232),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_249),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_231),
.A2(n_214),
.B(n_210),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_244),
.A2(n_251),
.B(n_253),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_234),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_219),
.Y(n_247)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_247),
.Y(n_258)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_242),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_219),
.Y(n_250)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_250),
.Y(n_264)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_227),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_222),
.C(n_213),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_237),
.C(n_233),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_238),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_236),
.A2(n_216),
.B1(n_214),
.B2(n_207),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_255),
.A2(n_254),
.B1(n_251),
.B2(n_243),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_256),
.B(n_215),
.Y(n_259)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_259),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_262),
.C(n_263),
.Y(n_273)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_261),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_220),
.C(n_226),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_216),
.C(n_211),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_248),
.Y(n_272)
);

AO21x1_ASAP7_75t_L g267 ( 
.A1(n_265),
.A2(n_244),
.B(n_256),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_267),
.B(n_254),
.Y(n_274)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_257),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_270),
.B(n_271),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_264),
.A2(n_241),
.B1(n_249),
.B2(n_206),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_119),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_276),
.Y(n_281)
);

OAI321xp33_ASAP7_75t_L g276 ( 
.A1(n_267),
.A2(n_246),
.A3(n_258),
.B1(n_259),
.B2(n_266),
.C(n_263),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_260),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_277),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_268),
.A2(n_262),
.B1(n_119),
.B2(n_15),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_278),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_279),
.B(n_269),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_282),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_281),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_274),
.Y(n_285)
);

A2O1A1Ixp33_ASAP7_75t_L g287 ( 
.A1(n_286),
.A2(n_275),
.B(n_283),
.C(n_273),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_287),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_288),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_13),
.Y(n_291)
);


endmodule