module real_jpeg_5380_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_286;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

OAI22xp33_ASAP7_75t_L g157 ( 
.A1(n_0),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_0),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_0),
.A2(n_158),
.B1(n_296),
.B2(n_299),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g391 ( 
.A1(n_0),
.A2(n_158),
.B1(n_392),
.B2(n_394),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_0),
.A2(n_72),
.B1(n_158),
.B2(n_426),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_1),
.A2(n_85),
.B1(n_89),
.B2(n_92),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_1),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_1),
.A2(n_92),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g403 ( 
.A1(n_1),
.A2(n_92),
.B1(n_206),
.B2(n_404),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_1),
.A2(n_92),
.B1(n_440),
.B2(n_442),
.Y(n_439)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_2),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_2),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_2),
.Y(n_258)
);

INVx8_ASAP7_75t_L g268 ( 
.A(n_2),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g300 ( 
.A(n_2),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_2),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_2),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_3),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_4),
.A2(n_95),
.B1(n_98),
.B2(n_102),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_4),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_4),
.A2(n_102),
.B1(n_131),
.B2(n_134),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_4),
.A2(n_102),
.B1(n_333),
.B2(n_371),
.Y(n_410)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_5),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_5),
.Y(n_159)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_5),
.Y(n_162)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_5),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_5),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_5),
.Y(n_461)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_6),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_6),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_6),
.B(n_127),
.C(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_6),
.B(n_73),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_6),
.B(n_222),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_6),
.B(n_129),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_6),
.B(n_97),
.Y(n_288)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_7),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_7),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_7),
.A2(n_207),
.B1(n_280),
.B2(n_282),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g387 ( 
.A1(n_7),
.A2(n_207),
.B1(n_323),
.B2(n_388),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_7),
.A2(n_159),
.B1(n_207),
.B2(n_435),
.Y(n_434)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g354 ( 
.A(n_8),
.Y(n_354)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_9),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_10),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_10),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_10),
.A2(n_194),
.B1(n_224),
.B2(n_227),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_10),
.A2(n_173),
.B1(n_194),
.B2(n_291),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_10),
.A2(n_194),
.B1(n_382),
.B2(n_383),
.Y(n_381)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_11),
.Y(n_113)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_11),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_11),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_11),
.Y(n_127)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_12),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_13),
.Y(n_122)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_13),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_13),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_14),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_14),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_14),
.A2(n_57),
.B1(n_169),
.B2(n_172),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g369 ( 
.A1(n_14),
.A2(n_57),
.B1(n_332),
.B2(n_370),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_14),
.A2(n_57),
.B1(n_417),
.B2(n_419),
.Y(n_416)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_16),
.A2(n_32),
.B1(n_48),
.B2(n_50),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_16),
.A2(n_50),
.B1(n_332),
.B2(n_334),
.Y(n_331)
);

OAI22xp33_ASAP7_75t_SL g412 ( 
.A1(n_16),
.A2(n_50),
.B1(n_232),
.B2(n_413),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_SL g430 ( 
.A1(n_16),
.A2(n_50),
.B1(n_291),
.B2(n_431),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_17),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_17),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_17),
.A2(n_233),
.B1(n_251),
.B2(n_254),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_17),
.A2(n_233),
.B1(n_321),
.B2(n_323),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_17),
.A2(n_48),
.B1(n_233),
.B2(n_460),
.Y(n_459)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_538),
.B(n_541),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_176),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_174),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_149),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_23),
.B(n_149),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_138),
.B2(n_139),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_58),
.C(n_103),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_26),
.B(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_47),
.B1(n_51),
.B2(n_53),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_27),
.A2(n_51),
.B1(n_53),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_27),
.A2(n_47),
.B1(n_51),
.B2(n_156),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_27),
.A2(n_380),
.B(n_434),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_27),
.A2(n_51),
.B1(n_434),
.B2(n_459),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_28),
.A2(n_378),
.B(n_379),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_28),
.B(n_381),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_38),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_34),
.Y(n_145)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_39),
.B1(n_42),
.B2(n_45),
.Y(n_38)
);

INVx6_ASAP7_75t_L g356 ( 
.A(n_36),
.Y(n_356)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_44),
.Y(n_173)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_44),
.Y(n_291)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp33_ASAP7_75t_SL g378 ( 
.A1(n_48),
.A2(n_189),
.B(n_359),
.Y(n_378)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_51),
.B(n_189),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_51),
.A2(n_459),
.B(n_483),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_52),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_52),
.B(n_157),
.Y(n_482)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_58),
.A2(n_103),
.B1(n_104),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_58),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_84),
.B1(n_93),
.B2(n_94),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g141 ( 
.A(n_59),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_59),
.A2(n_84),
.B1(n_93),
.B2(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_59),
.A2(n_93),
.B1(n_320),
.B2(n_387),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_59),
.A2(n_93),
.B1(n_425),
.B2(n_430),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_73),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_65),
.B1(n_69),
.B2(n_71),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_68),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g302 ( 
.A(n_68),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_68),
.Y(n_429)
);

NAND2xp33_ASAP7_75t_SL g309 ( 
.A(n_69),
.B(n_133),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_73),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_73),
.A2(n_141),
.B(n_142),
.Y(n_140)
);

AOI22x1_ASAP7_75t_L g462 ( 
.A1(n_73),
.A2(n_141),
.B1(n_327),
.B2(n_463),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_73),
.A2(n_141),
.B1(n_168),
.B2(n_471),
.Y(n_470)
);

AO22x2_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_78),
.B2(n_81),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g234 ( 
.A(n_75),
.Y(n_234)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g199 ( 
.A(n_77),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_77),
.Y(n_418)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_79),
.Y(n_393)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_83),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g325 ( 
.A(n_88),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_88),
.Y(n_432)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_93),
.B(n_290),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_93),
.A2(n_320),
.B(n_326),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

INVx6_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_101),
.Y(n_286)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_101),
.Y(n_348)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_101),
.Y(n_358)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_101),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_103),
.B(n_155),
.C(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_103),
.A2(n_104),
.B1(n_165),
.B2(n_166),
.Y(n_527)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_128),
.B(n_130),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_105),
.A2(n_186),
.B(n_190),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_105),
.A2(n_128),
.B1(n_231),
.B2(n_279),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_105),
.A2(n_190),
.B(n_279),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_105),
.A2(n_128),
.B1(n_391),
.B2(n_452),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_106),
.B(n_191),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_106),
.A2(n_129),
.B1(n_412),
.B2(n_416),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_106),
.A2(n_129),
.B1(n_416),
.B2(n_439),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_106),
.A2(n_129),
.B1(n_439),
.B2(n_474),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_117),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_111),
.B1(n_114),
.B2(n_116),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_110),
.Y(n_415)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx5_ASAP7_75t_SL g232 ( 
.A(n_116),
.Y(n_232)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_117),
.A2(n_231),
.B(n_235),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_120),
.B1(n_123),
.B2(n_126),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_120),
.Y(n_227)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g206 ( 
.A(n_122),
.Y(n_206)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_122),
.Y(n_226)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx8_ASAP7_75t_L g255 ( 
.A(n_124),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_125),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_125),
.Y(n_212)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_128),
.A2(n_235),
.B(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_129),
.B(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_130),
.Y(n_474)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_133),
.Y(n_441)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_134),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_136),
.Y(n_305)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_137),
.Y(n_188)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_137),
.Y(n_193)
);

INVx6_ASAP7_75t_L g422 ( 
.A(n_137),
.Y(n_422)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_141),
.A2(n_285),
.B(n_289),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_141),
.B(n_327),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_141),
.A2(n_289),
.B(n_496),
.Y(n_495)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_154),
.C(n_163),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_150),
.A2(n_151),
.B1(n_154),
.B2(n_155),
.Y(n_533)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_154),
.A2(n_155),
.B1(n_527),
.B2(n_528),
.Y(n_526)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx8_ASAP7_75t_L g361 ( 
.A(n_159),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_161),
.Y(n_160)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_163),
.A2(n_164),
.B1(n_532),
.B2(n_533),
.Y(n_531)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g322 ( 
.A(n_171),
.Y(n_322)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_522),
.B(n_535),
.Y(n_177)
);

OAI311xp33_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_397),
.A3(n_498),
.B1(n_516),
.C1(n_521),
.Y(n_178)
);

AOI21x1_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_339),
.B(n_396),
.Y(n_179)
);

AO21x1_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_311),
.B(n_338),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_273),
.B(n_310),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_238),
.B(n_272),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_203),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_184),
.B(n_203),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_196),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_185),
.A2(n_196),
.B1(n_197),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_185),
.Y(n_270)
);

INVx11_ASAP7_75t_L g195 ( 
.A(n_188),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_189),
.A2(n_213),
.B(n_220),
.Y(n_247)
);

OAI21xp33_ASAP7_75t_SL g285 ( 
.A1(n_189),
.A2(n_286),
.B(n_287),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_189),
.B(n_360),
.Y(n_359)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_193),
.Y(n_281)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_195),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

INVx3_ASAP7_75t_SL g198 ( 
.A(n_199),
.Y(n_198)
);

INVx5_ASAP7_75t_L g443 ( 
.A(n_199),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_201),
.Y(n_334)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_202),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_228),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_204),
.B(n_229),
.C(n_237),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_213),
.B(n_220),
.Y(n_204)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_205),
.Y(n_265)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx4_ASAP7_75t_SL g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_210),
.Y(n_299)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_212),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_212),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_213),
.A2(n_364),
.B1(n_365),
.B2(n_368),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_213),
.A2(n_403),
.B1(n_407),
.B2(n_410),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_213),
.A2(n_410),
.B(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_214),
.B(n_223),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_214),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_214),
.A2(n_295),
.B1(n_331),
.B2(n_335),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_214),
.A2(n_369),
.B1(n_454),
.B2(n_455),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_217),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_226),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_236),
.B2(n_237),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_232),
.Y(n_282)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_262),
.B(n_271),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_248),
.B(n_261),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_247),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_246),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx5_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

BUFx8_ASAP7_75t_L g298 ( 
.A(n_245),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_260),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_260),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_256),
.B(n_259),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_250),
.Y(n_264)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx3_ASAP7_75t_SL g256 ( 
.A(n_257),
.Y(n_256)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_258),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_259),
.A2(n_294),
.B(n_300),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_269),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_269),
.Y(n_271)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_268),
.Y(n_367)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_268),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_274),
.B(n_275),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_292),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_283),
.B2(n_284),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_278),
.B(n_283),
.C(n_292),
.Y(n_312)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVxp33_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

AOI32xp33_ASAP7_75t_L g301 ( 
.A1(n_288),
.A2(n_302),
.A3(n_303),
.B1(n_306),
.B2(n_309),
.Y(n_301)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_290),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_301),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_301),
.Y(n_317)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx8_ASAP7_75t_L g371 ( 
.A(n_298),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx8_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_312),
.B(n_313),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_318),
.B2(n_337),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_316),
.B(n_317),
.C(n_337),
.Y(n_340)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_318),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_328),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_319),
.B(n_329),
.C(n_330),
.Y(n_372)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_331),
.Y(n_364)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_340),
.B(n_341),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_375),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_343),
.A2(n_372),
.B1(n_373),
.B2(n_374),
.Y(n_342)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_343),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_344),
.A2(n_345),
.B1(n_362),
.B2(n_363),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_345),
.B(n_362),
.Y(n_494)
);

OAI32xp33_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_349),
.A3(n_352),
.B1(n_355),
.B2(n_359),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_372),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_372),
.B(n_373),
.C(n_375),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_376),
.A2(n_377),
.B1(n_385),
.B2(n_395),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_376),
.B(n_386),
.C(n_390),
.Y(n_507)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_382),
.Y(n_384)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_382),
.Y(n_435)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_385),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_386),
.B(n_390),
.Y(n_385)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_387),
.Y(n_496)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

NAND2xp33_ASAP7_75t_SL g397 ( 
.A(n_398),
.B(n_484),
.Y(n_397)
);

A2O1A1Ixp33_ASAP7_75t_SL g516 ( 
.A1(n_398),
.A2(n_484),
.B(n_517),
.C(n_520),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_464),
.Y(n_398)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_399),
.B(n_464),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_436),
.C(n_449),
.Y(n_399)
);

FAx1_ASAP7_75t_SL g497 ( 
.A(n_400),
.B(n_436),
.CI(n_449),
.CON(n_497),
.SN(n_497)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_423),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_401),
.B(n_424),
.C(n_433),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_411),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_402),
.B(n_411),
.Y(n_490)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_403),
.Y(n_454)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx6_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_412),
.Y(n_452)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx5_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx8_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_433),
.Y(n_423)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_425),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_427),
.Y(n_426)
);

INVx5_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_430),
.Y(n_471)
);

INVx4_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_437),
.A2(n_438),
.B1(n_444),
.B2(n_448),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_438),
.B(n_444),
.Y(n_478)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_444),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_444),
.A2(n_448),
.B1(n_480),
.B2(n_481),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_444),
.A2(n_478),
.B(n_481),
.Y(n_525)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx4_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_457),
.C(n_462),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_450),
.B(n_488),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_451),
.B(n_453),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_451),
.B(n_453),
.Y(n_506)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_457),
.A2(n_458),
.B1(n_462),
.B2(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_462),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_466),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_465),
.B(n_468),
.C(n_476),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_467),
.A2(n_468),
.B1(n_476),
.B2(n_477),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_469),
.A2(n_472),
.B(n_475),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_470),
.B(n_473),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

FAx1_ASAP7_75t_SL g524 ( 
.A(n_475),
.B(n_525),
.CI(n_526),
.CON(n_524),
.SN(n_524)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_475),
.B(n_525),
.C(n_526),
.Y(n_534)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_479),
.Y(n_477)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_483),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_497),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_485),
.B(n_497),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_490),
.C(n_491),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_486),
.A2(n_487),
.B1(n_490),
.B2(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_490),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_491),
.B(n_509),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_494),
.C(n_495),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_492),
.A2(n_493),
.B1(n_495),
.B2(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_494),
.B(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_495),
.Y(n_504)
);

BUFx24_ASAP7_75t_SL g544 ( 
.A(n_497),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_499),
.B(n_511),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_500),
.A2(n_518),
.B(n_519),
.Y(n_517)
);

NOR2x1_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_508),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_501),
.B(n_508),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_505),
.C(n_507),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_502),
.B(n_514),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_505),
.A2(n_506),
.B1(n_507),
.B2(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_507),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_513),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_512),
.B(n_513),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_530),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_524),
.B(n_529),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_524),
.B(n_529),
.Y(n_536)
);

BUFx24_ASAP7_75t_SL g546 ( 
.A(n_524),
.Y(n_546)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_527),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_530),
.A2(n_536),
.B(n_537),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_531),
.B(n_534),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_531),
.B(n_534),
.Y(n_537)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVx5_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx6_ASAP7_75t_L g542 ( 
.A(n_540),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_542),
.B(n_543),
.Y(n_541)
);


endmodule