module fake_jpeg_9191_n_342 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_5),
.B(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_40),
.Y(n_51)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_46),
.Y(n_59)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_26),
.Y(n_67)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_49),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_53),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_56),
.Y(n_74)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_62),
.Y(n_77)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_66),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_19),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_48),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_26),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_84),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_37),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_29),
.Y(n_119)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_33),
.B1(n_39),
.B2(n_48),
.Y(n_80)
);

NOR2x1p5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_97),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_26),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_25),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_85),
.B(n_87),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_63),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_25),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_22),
.C(n_21),
.Y(n_108)
);

CKINVDCx12_ASAP7_75t_R g91 ( 
.A(n_60),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_91),
.B(n_94),
.Y(n_131)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_52),
.A2(n_42),
.B(n_28),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_92),
.Y(n_111)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_93),
.Y(n_105)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_101),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_52),
.A2(n_17),
.B1(n_33),
.B2(n_44),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_96),
.A2(n_17),
.B1(n_22),
.B2(n_29),
.Y(n_109)
);

OAI32xp33_ASAP7_75t_L g97 ( 
.A1(n_56),
.A2(n_45),
.A3(n_21),
.B1(n_29),
.B2(n_22),
.Y(n_97)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_102),
.B(n_106),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_17),
.B1(n_33),
.B2(n_21),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_104),
.A2(n_99),
.B1(n_100),
.B2(n_34),
.Y(n_157)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_108),
.B(n_118),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_109),
.A2(n_99),
.B1(n_100),
.B2(n_93),
.Y(n_154)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_117),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_82),
.B(n_19),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_121),
.Y(n_143)
);

NAND2xp33_ASAP7_75t_SL g120 ( 
.A(n_78),
.B(n_18),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_120),
.A2(n_18),
.B1(n_30),
.B2(n_34),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_50),
.C(n_44),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_78),
.A2(n_20),
.B1(n_28),
.B2(n_27),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_122),
.A2(n_90),
.B1(n_25),
.B2(n_27),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_58),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_123),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_84),
.B(n_50),
.C(n_62),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_125),
.Y(n_134)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_75),
.B(n_20),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_127),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_73),
.C(n_64),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_129),
.Y(n_140)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_112),
.A2(n_85),
.B(n_80),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_142),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_136),
.B(n_145),
.Y(n_175)
);

MAJx2_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_80),
.C(n_83),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_144),
.C(n_128),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_114),
.A2(n_87),
.B1(n_53),
.B2(n_55),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_141),
.A2(n_129),
.B1(n_122),
.B2(n_126),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_112),
.A2(n_27),
.B(n_18),
.Y(n_142)
);

MAJx2_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_18),
.C(n_30),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_107),
.B(n_101),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_110),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_150),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_130),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_118),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_153),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_131),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_154),
.A2(n_157),
.B1(n_117),
.B2(n_105),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_109),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_156),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_158),
.A2(n_176),
.B(n_18),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_159),
.A2(n_169),
.B1(n_173),
.B2(n_136),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_156),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_160),
.B(n_161),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_152),
.B(n_125),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_164),
.Y(n_185)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_154),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_174),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_166),
.A2(n_113),
.B1(n_150),
.B2(n_135),
.Y(n_197)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_167),
.B(n_179),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_146),
.A2(n_121),
.B1(n_107),
.B2(n_124),
.Y(n_169)
);

A2O1A1O1Ixp25_ASAP7_75t_L g170 ( 
.A1(n_138),
.A2(n_142),
.B(n_133),
.C(n_144),
.D(n_146),
.Y(n_170)
);

A2O1A1O1Ixp25_ASAP7_75t_L g192 ( 
.A1(n_170),
.A2(n_132),
.B(n_148),
.C(n_153),
.D(n_137),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_148),
.A2(n_140),
.B1(n_147),
.B2(n_139),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_172),
.A2(n_182),
.B1(n_175),
.B2(n_178),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_140),
.A2(n_115),
.B1(n_103),
.B2(n_106),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_119),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_103),
.C(n_108),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_180),
.C(n_183),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_119),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_184),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_182),
.B(n_54),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_88),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_156),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_188),
.Y(n_225)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

INVx13_ASAP7_75t_L g189 ( 
.A(n_181),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_189),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_190),
.B(n_213),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_192),
.A2(n_196),
.B(n_198),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_132),
.Y(n_193)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_197),
.A2(n_81),
.B1(n_24),
.B2(n_34),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_137),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_199),
.B(n_202),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_169),
.A2(n_135),
.B1(n_113),
.B2(n_130),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_200),
.A2(n_210),
.B1(n_98),
.B2(n_151),
.Y(n_237)
);

NOR2x1_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_105),
.Y(n_201)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_201),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_75),
.Y(n_202)
);

INVx13_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_203),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_36),
.Y(n_204)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_0),
.Y(n_240)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_168),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_208),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_158),
.A2(n_70),
.B1(n_65),
.B2(n_72),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_207),
.A2(n_81),
.B1(n_24),
.B2(n_23),
.Y(n_221)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_168),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_75),
.C(n_81),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_0),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_170),
.A2(n_98),
.B1(n_151),
.B2(n_36),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_36),
.Y(n_211)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_179),
.Y(n_213)
);

AOI32xp33_ASAP7_75t_L g216 ( 
.A1(n_201),
.A2(n_176),
.A3(n_81),
.B1(n_23),
.B2(n_34),
.Y(n_216)
);

OAI21x1_ASAP7_75t_SL g252 ( 
.A1(n_216),
.A2(n_218),
.B(n_211),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_219),
.B(n_224),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_186),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_12),
.B(n_16),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_222),
.A2(n_228),
.B(n_236),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_185),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_187),
.B(n_11),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_226),
.B(n_10),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_194),
.A2(n_13),
.B(n_15),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_203),
.A2(n_151),
.B1(n_116),
.B2(n_98),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_230),
.A2(n_232),
.B1(n_197),
.B2(n_198),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_206),
.A2(n_23),
.B1(n_24),
.B2(n_3),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_36),
.Y(n_234)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_234),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_194),
.B(n_24),
.Y(n_235)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_235),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_212),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_237),
.A2(n_196),
.B1(n_207),
.B2(n_204),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_209),
.C(n_205),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_228),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_241),
.A2(n_227),
.B1(n_214),
.B2(n_220),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_231),
.A2(n_200),
.B1(n_210),
.B2(n_188),
.Y(n_242)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_242),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_246),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_217),
.A2(n_213),
.B1(n_208),
.B2(n_190),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_245),
.A2(n_217),
.B1(n_231),
.B2(n_237),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_191),
.Y(n_246)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_247),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_191),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_256),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_189),
.Y(n_249)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_249),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_225),
.Y(n_250)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_250),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_251),
.B(n_263),
.C(n_240),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_252),
.A2(n_259),
.B1(n_230),
.B2(n_232),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_225),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_255),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_192),
.Y(n_256)
);

NAND3xp33_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_8),
.C(n_14),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_261),
.Y(n_275)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_223),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_234),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_262),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_220),
.B(n_0),
.C(n_1),
.Y(n_263)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_264),
.Y(n_289)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_265),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_241),
.A2(n_227),
.B1(n_214),
.B2(n_219),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_269),
.A2(n_258),
.B1(n_244),
.B2(n_263),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_256),
.B(n_233),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_281),
.Y(n_287)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_272),
.Y(n_295)
);

FAx1_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_222),
.CI(n_233),
.CON(n_277),
.SN(n_277)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_277),
.A2(n_270),
.B(n_274),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_235),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_279),
.C(n_251),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_245),
.B(n_238),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_266),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_284),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g283 ( 
.A(n_277),
.Y(n_283)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_283),
.Y(n_310)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_264),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_292),
.C(n_268),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_286),
.B(n_291),
.Y(n_301)
);

BUFx12f_ASAP7_75t_L g288 ( 
.A(n_280),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_290),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_275),
.B(n_254),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_248),
.C(n_244),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_243),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_215),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_297),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_215),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_257),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_299),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_295),
.B(n_257),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_305),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_304),
.C(n_306),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_285),
.C(n_267),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_271),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_288),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_284),
.A2(n_268),
.B(n_267),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_294),
.A2(n_279),
.B1(n_281),
.B2(n_221),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_287),
.C(n_288),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_309),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_289),
.A2(n_8),
.B1(n_4),
.B2(n_6),
.Y(n_309)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_313),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_315),
.A2(n_316),
.B1(n_300),
.B2(n_304),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_287),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_317),
.A2(n_8),
.B(n_10),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_301),
.A2(n_9),
.B(n_4),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_320),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_310),
.A2(n_9),
.B1(n_4),
.B2(n_7),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_299),
.B(n_7),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_321),
.B(n_313),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_326),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_324),
.B(n_325),
.C(n_327),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_303),
.C(n_308),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_298),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_7),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_329),
.B(n_13),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_325),
.A2(n_318),
.B(n_10),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_330),
.B(n_331),
.Y(n_336)
);

A2O1A1Ixp33_ASAP7_75t_L g334 ( 
.A1(n_323),
.A2(n_13),
.B(n_15),
.C(n_1),
.Y(n_334)
);

O2A1O1Ixp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_328),
.B(n_329),
.C(n_1),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_335),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_332),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_338),
.B(n_333),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_339),
.A2(n_336),
.B(n_327),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_334),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_1),
.Y(n_342)
);


endmodule