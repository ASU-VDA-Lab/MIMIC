module fake_jpeg_14168_n_130 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_130);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx2_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_12),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_31),
.A2(n_38),
.B1(n_23),
.B2(n_22),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_43),
.Y(n_49)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_8),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_9),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_22),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_40),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_4),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_20),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_45),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_9),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_47),
.Y(n_54)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_13),
.B1(n_18),
.B2(n_23),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_69),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_56),
.B(n_57),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_20),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_16),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_60),
.B(n_61),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_46),
.B(n_16),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_21),
.Y(n_62)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_21),
.Y(n_65)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

NAND2x1p5_ASAP7_75t_L g66 ( 
.A(n_29),
.B(n_28),
.Y(n_66)
);

A2O1A1O1Ixp25_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_71),
.B(n_18),
.C(n_11),
.D(n_10),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_53),
.Y(n_82)
);

NOR2x1_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_24),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_33),
.B(n_10),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_59),
.A2(n_30),
.B1(n_41),
.B2(n_24),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_75),
.B1(n_81),
.B2(n_82),
.Y(n_95)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_61),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_68),
.A2(n_13),
.B1(n_63),
.B2(n_57),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_49),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_87),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_48),
.A2(n_53),
.B1(n_66),
.B2(n_69),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_54),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_85),
.C(n_81),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_53),
.A2(n_66),
.B1(n_69),
.B2(n_71),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_85),
.A2(n_64),
.B1(n_50),
.B2(n_58),
.Y(n_91)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_52),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_92),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_80),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_91),
.A2(n_88),
.B1(n_73),
.B2(n_86),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_52),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_55),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_100),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_55),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_99),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_64),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_67),
.B1(n_70),
.B2(n_82),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_101),
.A2(n_72),
.B1(n_87),
.B2(n_74),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_84),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_106),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_82),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_105),
.B(n_110),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_107),
.A2(n_94),
.B(n_98),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_83),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_98),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_109),
.A2(n_104),
.B1(n_97),
.B2(n_90),
.Y(n_114)
);

MAJx2_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_92),
.C(n_93),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_113),
.C(n_109),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_114),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_117),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_119),
.Y(n_125)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_120),
.A2(n_102),
.B(n_103),
.Y(n_123)
);

NOR3xp33_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_124),
.C(n_96),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_121),
.A2(n_112),
.B(n_111),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_118),
.B1(n_122),
.B2(n_96),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_126),
.A2(n_127),
.B(n_79),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_128),
.B(n_67),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_67),
.Y(n_130)
);


endmodule