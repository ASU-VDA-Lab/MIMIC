module fake_jpeg_32027_n_167 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_167);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

INVx11_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_24),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_6),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_29),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

BUFx4f_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_27),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_2),
.B(n_7),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_4),
.Y(n_72)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_0),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_77),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_20),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_82),
.Y(n_85)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_1),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_72),
.Y(n_89)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_17),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_77),
.A2(n_56),
.B1(n_51),
.B2(n_62),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_94),
.B1(n_97),
.B2(n_75),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_64),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_93),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_59),
.B1(n_69),
.B2(n_65),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_88),
.A2(n_56),
.B1(n_51),
.B2(n_50),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_89),
.B(n_95),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_57),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_69),
.B1(n_58),
.B2(n_52),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_79),
.B(n_70),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_73),
.A2(n_52),
.B1(n_58),
.B2(n_62),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_125)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_63),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_106),
.Y(n_120)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_111),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_1),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_3),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_115),
.Y(n_129)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

AO22x1_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_77),
.B1(n_68),
.B2(n_61),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_110),
.A2(n_53),
.B1(n_6),
.B2(n_7),
.Y(n_123)
);

OR2x2_ASAP7_75t_SL g111 ( 
.A(n_86),
.B(n_3),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_113),
.Y(n_122)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_94),
.B(n_54),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_114),
.B(n_116),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_4),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_5),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_117),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_123),
.A2(n_125),
.B1(n_11),
.B2(n_12),
.Y(n_141)
);

AND2x6_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_26),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_23),
.B(n_25),
.C(n_28),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_116),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_130),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_107),
.B(n_8),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_9),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_132),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_10),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_134),
.A2(n_33),
.B1(n_39),
.B2(n_40),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_34),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_99),
.B(n_31),
.C(n_45),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_13),
.Y(n_144)
);

XOR2x2_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_30),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_151),
.Y(n_152)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_141),
.A2(n_147),
.B1(n_149),
.B2(n_134),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_121),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_142),
.A2(n_150),
.B1(n_123),
.B2(n_144),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_143),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_145),
.Y(n_153)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_136),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_42),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_154),
.A2(n_148),
.B(n_129),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_155),
.Y(n_159)
);

AOI322xp5_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_138),
.A3(n_124),
.B1(n_126),
.B2(n_151),
.C1(n_146),
.C2(n_147),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_158),
.A2(n_152),
.B(n_153),
.Y(n_162)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

AOI322xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_159),
.A3(n_157),
.B1(n_154),
.B2(n_156),
.C1(n_120),
.C2(n_128),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_161),
.B(n_137),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_164),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_43),
.C(n_47),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_135),
.C(n_133),
.Y(n_167)
);


endmodule