module fake_jpeg_10405_n_112 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_112);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_112;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx11_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

BUFx10_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_2),
.B(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_0),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_32),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_30),
.A2(n_31),
.B1(n_22),
.B2(n_24),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_20),
.A2(n_1),
.B1(n_6),
.B2(n_7),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_34),
.A2(n_22),
.B1(n_18),
.B2(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_22),
.B1(n_21),
.B2(n_19),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_25),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_21),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_24),
.C(n_25),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_15),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_16),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_42),
.B(n_25),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_26),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_53),
.B1(n_62),
.B2(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

AOI222xp33_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_41),
.B1(n_38),
.B2(n_14),
.C1(n_15),
.C2(n_16),
.Y(n_55)
);

MAJx2_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_23),
.C(n_17),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_46),
.B(n_45),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_61),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_19),
.Y(n_58)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_63),
.A2(n_13),
.B(n_48),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_71),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_46),
.B(n_47),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_72),
.B(n_52),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_60),
.A2(n_29),
.B1(n_44),
.B2(n_48),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_74),
.B1(n_59),
.B2(n_61),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_62),
.A2(n_18),
.B1(n_23),
.B2(n_9),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_72),
.A2(n_55),
.B(n_54),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_82),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_SL g78 ( 
.A(n_69),
.B(n_56),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_85),
.C(n_74),
.Y(n_88)
);

CKINVDCx5p33_ASAP7_75t_R g82 ( 
.A(n_75),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_51),
.B(n_59),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_77),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_6),
.B(n_7),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_71),
.C(n_73),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_88),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_81),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_93),
.A2(n_68),
.B(n_70),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_98),
.Y(n_99)
);

NOR3xp33_ASAP7_75t_SL g98 ( 
.A(n_92),
.B(n_70),
.C(n_51),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_95),
.A2(n_93),
.B1(n_87),
.B2(n_86),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_101),
.Y(n_104)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

AOI31xp67_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_95),
.A3(n_10),
.B(n_75),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_103),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_100),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_99),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_108),
.A2(n_109),
.B(n_104),
.Y(n_110)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_107),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_57),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_10),
.Y(n_112)
);


endmodule