module fake_jpeg_16809_n_201 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_201);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_40),
.Y(n_58)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_33),
.C(n_24),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_43),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_0),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_17),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_28),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_41),
.A2(n_32),
.B1(n_27),
.B2(n_18),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_49),
.B1(n_55),
.B2(n_37),
.Y(n_70)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_48),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_41),
.A2(n_32),
.B1(n_27),
.B2(n_18),
.Y(n_49)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_57),
.Y(n_84)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_28),
.B1(n_30),
.B2(n_20),
.Y(n_55)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_20),
.B1(n_29),
.B2(n_26),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_60),
.A2(n_44),
.B1(n_40),
.B2(n_19),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_67),
.Y(n_94)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_63),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_29),
.B1(n_20),
.B2(n_30),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_68),
.A2(n_69),
.B(n_31),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_38),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_70),
.A2(n_75),
.B1(n_77),
.B2(n_81),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_60),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_73),
.Y(n_95)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_47),
.A2(n_39),
.B1(n_30),
.B2(n_28),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_63),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_76),
.B(n_89),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_52),
.A2(n_39),
.B1(n_29),
.B2(n_22),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_43),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_35),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_51),
.A2(n_45),
.B1(n_54),
.B2(n_57),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_79),
.A2(n_87),
.B1(n_16),
.B2(n_33),
.Y(n_110)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_50),
.A2(n_39),
.B1(n_22),
.B2(n_19),
.Y(n_81)
);

HAxp5_ASAP7_75t_SL g85 ( 
.A(n_62),
.B(n_43),
.CON(n_85),
.SN(n_85)
);

MAJIxp5_ASAP7_75t_SL g112 ( 
.A(n_85),
.B(n_23),
.C(n_33),
.Y(n_112)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_88),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_36),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_93),
.B(n_110),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_106),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_71),
.A2(n_26),
.B1(n_34),
.B2(n_31),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_104),
.B(n_64),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_56),
.C(n_24),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_111),
.C(n_103),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_56),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_113),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_21),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_21),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_108),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_16),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_69),
.A2(n_34),
.B1(n_56),
.B2(n_3),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_109),
.A2(n_82),
.B1(n_64),
.B2(n_90),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_23),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_112),
.A2(n_95),
.B(n_101),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_83),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_85),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_97),
.B1(n_113),
.B2(n_110),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_96),
.A2(n_65),
.B1(n_80),
.B2(n_83),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

OAI22x1_ASAP7_75t_SL g120 ( 
.A1(n_112),
.A2(n_72),
.B1(n_86),
.B2(n_66),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_120),
.A2(n_123),
.B1(n_105),
.B2(n_92),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_131),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_124),
.Y(n_149)
);

OAI22x1_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_67),
.B1(n_90),
.B2(n_88),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_98),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_125),
.B(n_129),
.Y(n_139)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

AO221x1_ASAP7_75t_L g146 ( 
.A1(n_126),
.A2(n_123),
.B1(n_120),
.B2(n_124),
.C(n_91),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_128),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_82),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_76),
.Y(n_130)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_130),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

FAx1_ASAP7_75t_SL g134 ( 
.A(n_127),
.B(n_104),
.CI(n_100),
.CON(n_134),
.SN(n_134)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_136),
.Y(n_161)
);

AOI221xp5_ASAP7_75t_L g165 ( 
.A1(n_135),
.A2(n_116),
.B1(n_117),
.B2(n_126),
.C(n_5),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_123),
.Y(n_155)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_105),
.C(n_91),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_151),
.Y(n_160)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_147),
.A2(n_122),
.B1(n_114),
.B2(n_117),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_125),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_13),
.C(n_11),
.Y(n_151)
);

MAJx2_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_128),
.C(n_118),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_161),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_151),
.B(n_115),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_154),
.B(n_159),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_155),
.A2(n_165),
.B1(n_148),
.B2(n_147),
.Y(n_169)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_164),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_114),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_136),
.C(n_142),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_163),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_115),
.Y(n_164)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_171),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_169),
.A2(n_156),
.B1(n_155),
.B2(n_159),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_137),
.C(n_138),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_139),
.C(n_116),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_175),
.Y(n_184)
);

NOR2xp67_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_144),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_176),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_143),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_1),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_2),
.C(n_5),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_167),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_179),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_126),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_2),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_174),
.A2(n_160),
.B(n_152),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_182),
.A2(n_174),
.B(n_4),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_13),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_185),
.A2(n_6),
.B(n_7),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_188),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_8),
.C(n_5),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_190),
.Y(n_193)
);

OAI321xp33_ASAP7_75t_L g196 ( 
.A1(n_191),
.A2(n_194),
.A3(n_6),
.B1(n_7),
.B2(n_181),
.C(n_184),
.Y(n_196)
);

A2O1A1Ixp33_ASAP7_75t_SL g194 ( 
.A1(n_186),
.A2(n_183),
.B(n_178),
.C(n_179),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_193),
.B(n_186),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_195),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_196),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_184),
.C(n_194),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_197),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_198),
.Y(n_201)
);


endmodule