module fake_jpeg_23388_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_145;
wire n_18;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_16),
.B1(n_28),
.B2(n_30),
.Y(n_48)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_48),
.A2(n_43),
.B1(n_32),
.B2(n_27),
.Y(n_90)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_58),
.Y(n_82)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_59),
.B(n_43),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_17),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_61),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_8),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_30),
.B1(n_34),
.B2(n_32),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_63),
.A2(n_72),
.B1(n_74),
.B2(n_85),
.Y(n_105)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_66),
.Y(n_100)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_68),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_50),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_50),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_69),
.A2(n_41),
.B1(n_49),
.B2(n_56),
.Y(n_98)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_71),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_53),
.A2(n_30),
.B1(n_19),
.B2(n_21),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_51),
.A2(n_23),
.B1(n_19),
.B2(n_21),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_60),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_76),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_60),
.Y(n_79)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_61),
.A2(n_32),
.B1(n_34),
.B2(n_19),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_87),
.Y(n_117)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_22),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_90),
.A2(n_92),
.B1(n_23),
.B2(n_22),
.Y(n_121)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_59),
.A2(n_42),
.B1(n_41),
.B2(n_37),
.Y(n_92)
);

AND2x4_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_38),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_94),
.A2(n_97),
.B(n_99),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_103),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_91),
.A2(n_36),
.B(n_56),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_98),
.A2(n_109),
.B1(n_121),
.B2(n_49),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_1),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_76),
.A2(n_81),
.B1(n_83),
.B2(n_21),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_90),
.A2(n_42),
.B1(n_54),
.B2(n_38),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_119),
.B1(n_67),
.B2(n_44),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_112),
.B(n_118),
.Y(n_123)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_116),
.Y(n_148)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_42),
.B1(n_54),
.B2(n_38),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_47),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_64),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_115),
.A2(n_71),
.B1(n_87),
.B2(n_84),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_124),
.A2(n_138),
.B1(n_108),
.B2(n_103),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_100),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_125),
.B(n_135),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_102),
.B1(n_107),
.B2(n_36),
.Y(n_156)
);

MAJx2_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_80),
.C(n_35),
.Y(n_129)
);

XNOR2x1_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_130),
.Y(n_155)
);

AOI32xp33_ASAP7_75t_L g130 ( 
.A1(n_94),
.A2(n_49),
.A3(n_44),
.B1(n_65),
.B2(n_70),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_131),
.B(n_139),
.Y(n_164)
);

AND2x4_ASAP7_75t_SL g132 ( 
.A(n_94),
.B(n_44),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_132),
.A2(n_133),
.B(n_137),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_75),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_134),
.B(n_150),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_97),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_95),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_136),
.B(n_140),
.Y(n_182)
);

O2A1O1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_44),
.B(n_27),
.C(n_66),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_96),
.B(n_86),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_94),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_142),
.Y(n_170)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_143),
.A2(n_108),
.B1(n_117),
.B2(n_113),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g144 ( 
.A(n_95),
.B(n_55),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_27),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_1),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_146),
.A2(n_147),
.B(n_31),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_2),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_86),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_149),
.B(n_12),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_99),
.B(n_78),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_135),
.A2(n_115),
.B1(n_102),
.B2(n_105),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_151),
.A2(n_156),
.B1(n_157),
.B2(n_159),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_121),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_123),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_141),
.A2(n_99),
.B1(n_122),
.B2(n_78),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_158),
.A2(n_140),
.B1(n_125),
.B2(n_126),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_93),
.B1(n_110),
.B2(n_113),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_138),
.A2(n_110),
.B1(n_93),
.B2(n_118),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_132),
.A2(n_57),
.B1(n_52),
.B2(n_46),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_132),
.A2(n_116),
.B1(n_101),
.B2(n_39),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_133),
.A2(n_101),
.B1(n_39),
.B2(n_35),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_165),
.A2(n_171),
.B1(n_172),
.B2(n_180),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_129),
.A2(n_18),
.B(n_16),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_166),
.A2(n_179),
.B(n_31),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_144),
.A2(n_39),
.B(n_35),
.C(n_29),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_167),
.A2(n_177),
.B(n_178),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_39),
.C(n_35),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_31),
.C(n_26),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_175),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_134),
.A2(n_16),
.B1(n_28),
.B2(n_22),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_137),
.A2(n_23),
.B1(n_28),
.B2(n_18),
.Y(n_172)
);

OA21x2_ASAP7_75t_R g175 ( 
.A1(n_147),
.A2(n_146),
.B(n_130),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_2),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_127),
.A2(n_31),
.B(n_25),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_146),
.A2(n_29),
.B1(n_25),
.B2(n_26),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_183),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_184),
.Y(n_223)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_182),
.Y(n_185)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_185),
.Y(n_232)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_186),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_187),
.B(n_189),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_176),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_188),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_147),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_165),
.Y(n_191)
);

INVxp67_ASAP7_75t_SL g238 ( 
.A(n_191),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_126),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_192),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_177),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_193),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_195),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_131),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_197),
.B(n_209),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_199),
.A2(n_204),
.B(n_211),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_151),
.A2(n_143),
.B1(n_142),
.B2(n_29),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_173),
.A2(n_142),
.B1(n_29),
.B2(n_25),
.Y(n_201)
);

AO22x2_ASAP7_75t_L g202 ( 
.A1(n_175),
.A2(n_25),
.B1(n_26),
.B2(n_24),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_203),
.A2(n_207),
.B1(n_214),
.B2(n_167),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_2),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_181),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_205),
.Y(n_239)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_163),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_173),
.A2(n_26),
.B1(n_24),
.B2(n_20),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_208),
.A2(n_156),
.B1(n_172),
.B2(n_167),
.Y(n_233)
);

XNOR2x1_ASAP7_75t_L g209 ( 
.A(n_152),
.B(n_166),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_213),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_178),
.A2(n_170),
.B(n_160),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_168),
.B(n_31),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_157),
.B(n_31),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_162),
.B(n_24),
.C(n_20),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_215),
.A2(n_180),
.B(n_179),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_167),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_216),
.A2(n_234),
.B(n_240),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_202),
.Y(n_219)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_219),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_221),
.B(n_230),
.Y(n_262)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_190),
.Y(n_225)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_225),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_206),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_228),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_204),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_194),
.Y(n_229)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_229),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_233),
.A2(n_200),
.B1(n_208),
.B2(n_198),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_211),
.A2(n_167),
.B(n_177),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_202),
.A2(n_169),
.B1(n_171),
.B2(n_24),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_235),
.A2(n_212),
.B1(n_213),
.B2(n_20),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_189),
.B(n_3),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_196),
.A2(n_10),
.B(n_15),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_241),
.A2(n_212),
.B(n_215),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_242),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_197),
.C(n_187),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_246),
.C(n_249),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_209),
.C(n_214),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_204),
.Y(n_247)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_198),
.Y(n_248)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_248),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_210),
.C(n_199),
.Y(n_249)
);

XNOR2x1_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_202),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_251),
.B(n_260),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_252),
.A2(n_258),
.B(n_234),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_20),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_230),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_225),
.A2(n_229),
.B1(n_221),
.B2(n_220),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_255),
.A2(n_218),
.B1(n_233),
.B2(n_216),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_256),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_3),
.C(n_4),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_241),
.C(n_239),
.Y(n_271)
);

A2O1A1Ixp33_ASAP7_75t_SL g258 ( 
.A1(n_216),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_258)
);

XOR2x2_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_10),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_245),
.B(n_237),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_265),
.B(n_277),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_266),
.A2(n_260),
.B1(n_259),
.B2(n_252),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_224),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_275),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_269),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_274),
.C(n_257),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_250),
.A2(n_235),
.B1(n_218),
.B2(n_222),
.Y(n_272)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_273),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_223),
.C(n_240),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_240),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_244),
.B(n_10),
.Y(n_277)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_278),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_246),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_258),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_281),
.A2(n_286),
.B(n_285),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_263),
.A2(n_255),
.B(n_261),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_282),
.A2(n_286),
.B(n_5),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_242),
.Y(n_283)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_283),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_259),
.C(n_254),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_253),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_294),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_291),
.A2(n_276),
.B1(n_273),
.B2(n_280),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g293 ( 
.A(n_266),
.Y(n_293)
);

AND2x2_ASAP7_75t_SL g303 ( 
.A(n_293),
.B(n_264),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_271),
.B(n_258),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_6),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_267),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_302),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_289),
.A2(n_270),
.B1(n_274),
.B2(n_276),
.Y(n_298)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_298),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_275),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_300),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_258),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_301),
.A2(n_305),
.B(n_308),
.Y(n_315)
);

AO21x1_ASAP7_75t_L g316 ( 
.A1(n_303),
.A2(n_304),
.B(n_295),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_290),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_281),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_292),
.A2(n_8),
.B(n_11),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_287),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_317),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_11),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_306),
.B(n_290),
.Y(n_314)
);

OAI21x1_ASAP7_75t_SL g323 ( 
.A1(n_314),
.A2(n_316),
.B(n_304),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_296),
.B(n_284),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_313),
.Y(n_318)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_318),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_312),
.A2(n_303),
.B(n_302),
.Y(n_319)
);

AOI21xp33_ASAP7_75t_L g327 ( 
.A1(n_319),
.A2(n_324),
.B(n_310),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_314),
.A2(n_303),
.B1(n_300),
.B2(n_307),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_320),
.A2(n_322),
.B(n_323),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_315),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_327),
.B(n_322),
.Y(n_328)
);

OAI321xp33_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_325),
.A3(n_321),
.B1(n_326),
.B2(n_12),
.C(n_11),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_13),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_13),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_13),
.Y(n_332)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_332),
.Y(n_333)
);


endmodule