module fake_netlist_1_4018_n_467 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_467);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_467;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_266;
wire n_84;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_444;
wire n_176;
wire n_123;
wire n_457;
wire n_223;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g71 ( .A(n_5), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_34), .Y(n_72) );
CKINVDCx16_ASAP7_75t_R g73 ( .A(n_7), .Y(n_73) );
INVx2_ASAP7_75t_L g74 ( .A(n_54), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_7), .Y(n_75) );
CKINVDCx5p33_ASAP7_75t_R g76 ( .A(n_29), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_19), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_53), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_26), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_47), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_59), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_15), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_14), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_30), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_61), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_69), .Y(n_86) );
HB1xp67_ASAP7_75t_L g87 ( .A(n_40), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_63), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_44), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_42), .Y(n_90) );
INVxp67_ASAP7_75t_SL g91 ( .A(n_70), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_33), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_24), .Y(n_93) );
INVxp33_ASAP7_75t_L g94 ( .A(n_0), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_20), .Y(n_95) );
INVxp33_ASAP7_75t_SL g96 ( .A(n_66), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_52), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_62), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_65), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_11), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_3), .Y(n_101) );
INVx1_ASAP7_75t_SL g102 ( .A(n_12), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_43), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_73), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_98), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_87), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_71), .Y(n_107) );
AND2x4_ASAP7_75t_L g108 ( .A(n_71), .B(n_0), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_102), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_72), .Y(n_110) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_74), .Y(n_111) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_94), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_96), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_74), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_72), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_77), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_75), .Y(n_117) );
AND2x6_ASAP7_75t_L g118 ( .A(n_77), .B(n_31), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_75), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_78), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_82), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_82), .Y(n_122) );
AND2x4_ASAP7_75t_L g123 ( .A(n_83), .B(n_1), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_76), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_78), .Y(n_125) );
BUFx3_ASAP7_75t_L g126 ( .A(n_118), .Y(n_126) );
INVx1_ASAP7_75t_SL g127 ( .A(n_112), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_120), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_120), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_120), .Y(n_130) );
AND2x6_ASAP7_75t_L g131 ( .A(n_108), .B(n_80), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_111), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_110), .B(n_89), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_118), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_120), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_120), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_118), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_110), .B(n_90), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_111), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_111), .Y(n_140) );
INVxp33_ASAP7_75t_L g141 ( .A(n_119), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_118), .Y(n_142) );
INVxp67_ASAP7_75t_SL g143 ( .A(n_116), .Y(n_143) );
BUFx3_ASAP7_75t_L g144 ( .A(n_118), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_111), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_108), .B(n_83), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_111), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_107), .B(n_101), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_134), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_143), .B(n_124), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_143), .B(n_124), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_141), .B(n_116), .Y(n_152) );
BUFx3_ASAP7_75t_L g153 ( .A(n_126), .Y(n_153) );
BUFx4f_ASAP7_75t_L g154 ( .A(n_131), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_128), .Y(n_155) );
INVx1_ASAP7_75t_SL g156 ( .A(n_127), .Y(n_156) );
OR2x2_ASAP7_75t_L g157 ( .A(n_127), .B(n_105), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_141), .B(n_125), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_128), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_146), .B(n_125), .Y(n_160) );
BUFx2_ASAP7_75t_L g161 ( .A(n_131), .Y(n_161) );
BUFx2_ASAP7_75t_L g162 ( .A(n_131), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_146), .B(n_113), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_129), .Y(n_164) );
AOI221xp5_ASAP7_75t_L g165 ( .A1(n_148), .A2(n_104), .B1(n_122), .B2(n_121), .C(n_117), .Y(n_165) );
AOI22xp5_ASAP7_75t_SL g166 ( .A1(n_131), .A2(n_106), .B1(n_109), .B2(n_104), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_146), .B(n_113), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_146), .Y(n_168) );
OR2x6_ASAP7_75t_L g169 ( .A(n_146), .B(n_108), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_148), .B(n_108), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_134), .Y(n_171) );
BUFx4f_ASAP7_75t_L g172 ( .A(n_131), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_148), .B(n_123), .Y(n_173) );
OR2x2_ASAP7_75t_L g174 ( .A(n_133), .B(n_123), .Y(n_174) );
AND3x1_ASAP7_75t_SL g175 ( .A(n_129), .B(n_101), .C(n_81), .Y(n_175) );
NAND2xp33_ASAP7_75t_SL g176 ( .A(n_134), .B(n_123), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_133), .B(n_123), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_131), .Y(n_178) );
OR2x2_ASAP7_75t_SL g179 ( .A(n_157), .B(n_134), .Y(n_179) );
INVx3_ASAP7_75t_SL g180 ( .A(n_156), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_149), .Y(n_181) );
INVx4_ASAP7_75t_L g182 ( .A(n_154), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_156), .B(n_131), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_176), .A2(n_126), .B(n_144), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_177), .B(n_131), .Y(n_185) );
OR2x6_ASAP7_75t_L g186 ( .A(n_161), .B(n_134), .Y(n_186) );
BUFx2_ASAP7_75t_L g187 ( .A(n_157), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_166), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_149), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_160), .A2(n_134), .B(n_142), .Y(n_190) );
AND2x4_ASAP7_75t_L g191 ( .A(n_161), .B(n_131), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_149), .Y(n_192) );
INVx2_ASAP7_75t_SL g193 ( .A(n_154), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g194 ( .A1(n_152), .A2(n_138), .B(n_115), .C(n_100), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_177), .B(n_131), .Y(n_195) );
INVx2_ASAP7_75t_SL g196 ( .A(n_154), .Y(n_196) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_149), .Y(n_197) );
BUFx3_ASAP7_75t_L g198 ( .A(n_172), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_168), .A2(n_118), .B1(n_126), .B2(n_144), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_168), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_169), .A2(n_118), .B1(n_126), .B2(n_144), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_149), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_171), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_169), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_169), .Y(n_205) );
OR2x2_ASAP7_75t_L g206 ( .A(n_158), .B(n_138), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_169), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_206), .B(n_170), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_200), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_206), .B(n_150), .Y(n_210) );
AOI221xp5_ASAP7_75t_L g211 ( .A1(n_187), .A2(n_165), .B1(n_163), .B2(n_194), .C(n_167), .Y(n_211) );
OAI22xp33_ASAP7_75t_L g212 ( .A1(n_180), .A2(n_151), .B1(n_169), .B2(n_172), .Y(n_212) );
NAND2xp33_ASAP7_75t_SL g213 ( .A(n_180), .B(n_162), .Y(n_213) );
NAND2xp33_ASAP7_75t_L g214 ( .A(n_180), .B(n_134), .Y(n_214) );
NAND3xp33_ASAP7_75t_L g215 ( .A(n_190), .B(n_166), .C(n_140), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_197), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_187), .B(n_174), .Y(n_217) );
OAI22xp33_ASAP7_75t_L g218 ( .A1(n_188), .A2(n_172), .B1(n_174), .B2(n_173), .Y(n_218) );
BUFx12f_ASAP7_75t_L g219 ( .A(n_183), .Y(n_219) );
BUFx2_ASAP7_75t_L g220 ( .A(n_183), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_197), .Y(n_221) );
AOI22xp33_ASAP7_75t_L g222 ( .A1(n_204), .A2(n_162), .B1(n_178), .B2(n_137), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_200), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_204), .Y(n_224) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_205), .A2(n_178), .B1(n_137), .B2(n_142), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_205), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_197), .Y(n_227) );
NAND2xp33_ASAP7_75t_R g228 ( .A(n_183), .B(n_175), .Y(n_228) );
AOI21x1_ASAP7_75t_L g229 ( .A1(n_190), .A2(n_140), .B(n_139), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_207), .B(n_153), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_197), .Y(n_231) );
NAND2xp33_ASAP7_75t_R g232 ( .A(n_210), .B(n_183), .Y(n_232) );
OAI22xp33_ASAP7_75t_L g233 ( .A1(n_228), .A2(n_185), .B1(n_195), .B2(n_207), .Y(n_233) );
OR2x2_ASAP7_75t_L g234 ( .A(n_208), .B(n_179), .Y(n_234) );
OA21x2_ASAP7_75t_L g235 ( .A1(n_229), .A2(n_203), .B(n_202), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_211), .A2(n_217), .B1(n_218), .B2(n_215), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_209), .Y(n_237) );
INVx3_ASAP7_75t_L g238 ( .A(n_230), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_209), .Y(n_239) );
BUFx2_ASAP7_75t_L g240 ( .A(n_219), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_217), .A2(n_115), .B1(n_114), .B2(n_185), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_208), .B(n_195), .Y(n_242) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_212), .A2(n_179), .B1(n_201), .B2(n_191), .Y(n_243) );
OAI21x1_ASAP7_75t_L g244 ( .A1(n_229), .A2(n_203), .B(n_202), .Y(n_244) );
OAI221xp5_ASAP7_75t_L g245 ( .A1(n_215), .A2(n_114), .B1(n_199), .B2(n_80), .C(n_95), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_220), .A2(n_88), .B1(n_81), .B2(n_97), .Y(n_246) );
NOR3xp33_ASAP7_75t_L g247 ( .A(n_213), .B(n_91), .C(n_103), .Y(n_247) );
OAI221xp5_ASAP7_75t_L g248 ( .A1(n_223), .A2(n_95), .B1(n_85), .B2(n_103), .C(n_86), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_223), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_220), .B(n_191), .Y(n_250) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_244), .Y(n_251) );
INVxp67_ASAP7_75t_L g252 ( .A(n_232), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_240), .B(n_219), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_237), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_237), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_237), .Y(n_256) );
BUFx3_ASAP7_75t_L g257 ( .A(n_240), .Y(n_257) );
AOI22xp33_ASAP7_75t_SL g258 ( .A1(n_243), .A2(n_219), .B1(n_214), .B2(n_226), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_249), .Y(n_259) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_239), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_239), .Y(n_261) );
NAND4xp25_ASAP7_75t_SL g262 ( .A(n_247), .B(n_85), .C(n_86), .D(n_88), .Y(n_262) );
INVx4_ASAP7_75t_L g263 ( .A(n_238), .Y(n_263) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_233), .A2(n_226), .B1(n_224), .B2(n_230), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_239), .Y(n_265) );
NAND3xp33_ASAP7_75t_L g266 ( .A(n_246), .B(n_97), .C(n_99), .Y(n_266) );
OAI221xp5_ASAP7_75t_L g267 ( .A1(n_236), .A2(n_224), .B1(n_222), .B2(n_99), .C(n_92), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_249), .Y(n_268) );
AO21x2_ASAP7_75t_L g269 ( .A1(n_244), .A2(n_231), .B(n_216), .Y(n_269) );
NOR2xp33_ASAP7_75t_R g270 ( .A(n_238), .B(n_191), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_269), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_269), .Y(n_272) );
AND2x4_ASAP7_75t_L g273 ( .A(n_265), .B(n_244), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_254), .B(n_238), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_254), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_255), .B(n_238), .Y(n_276) );
AOI211xp5_ASAP7_75t_SL g277 ( .A1(n_252), .A2(n_233), .B(n_243), .C(n_248), .Y(n_277) );
OAI22xp5_ASAP7_75t_L g278 ( .A1(n_258), .A2(n_236), .B1(n_234), .B2(n_248), .Y(n_278) );
INVx1_ASAP7_75t_SL g279 ( .A(n_257), .Y(n_279) );
BUFx2_ASAP7_75t_L g280 ( .A(n_260), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_255), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_256), .B(n_234), .Y(n_282) );
OAI31xp33_ASAP7_75t_SL g283 ( .A1(n_262), .A2(n_245), .A3(n_242), .B(n_250), .Y(n_283) );
AOI21xp5_ASAP7_75t_SL g284 ( .A1(n_264), .A2(n_245), .B(n_234), .Y(n_284) );
OAI221xp5_ASAP7_75t_L g285 ( .A1(n_266), .A2(n_241), .B1(n_246), .B2(n_247), .C(n_242), .Y(n_285) );
AOI221xp5_ASAP7_75t_L g286 ( .A1(n_267), .A2(n_242), .B1(n_241), .B2(n_92), .C(n_250), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_256), .B(n_235), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_261), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_261), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_259), .B(n_235), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_268), .B(n_235), .Y(n_291) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_265), .Y(n_292) );
OAI21xp5_ASAP7_75t_L g293 ( .A1(n_253), .A2(n_235), .B(n_225), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_263), .B(n_235), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_263), .B(n_250), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_263), .B(n_216), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_269), .B(n_230), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_251), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_257), .B(n_216), .Y(n_299) );
BUFx2_ASAP7_75t_L g300 ( .A(n_279), .Y(n_300) );
OAI211xp5_ASAP7_75t_SL g301 ( .A1(n_283), .A2(n_130), .B(n_135), .C(n_132), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_278), .B(n_1), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_287), .B(n_294), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_282), .B(n_251), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_280), .B(n_251), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_280), .B(n_251), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_287), .B(n_251), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_292), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_294), .B(n_2), .Y(n_309) );
NOR4xp25_ASAP7_75t_SL g310 ( .A(n_285), .B(n_79), .C(n_84), .D(n_93), .Y(n_310) );
INVxp67_ASAP7_75t_L g311 ( .A(n_279), .Y(n_311) );
INVxp67_ASAP7_75t_SL g312 ( .A(n_292), .Y(n_312) );
NAND2xp33_ASAP7_75t_SL g313 ( .A(n_278), .B(n_270), .Y(n_313) );
A2O1A1Ixp33_ASAP7_75t_L g314 ( .A1(n_283), .A2(n_230), .B(n_191), .C(n_227), .Y(n_314) );
INVx2_ASAP7_75t_SL g315 ( .A(n_299), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_285), .B(n_2), .Y(n_316) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_299), .Y(n_317) );
NAND3xp33_ASAP7_75t_L g318 ( .A(n_277), .B(n_132), .C(n_139), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_282), .B(n_3), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_297), .B(n_4), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_275), .Y(n_321) );
AND2x4_ASAP7_75t_L g322 ( .A(n_281), .B(n_221), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_281), .B(n_4), .Y(n_323) );
AOI221xp5_ASAP7_75t_L g324 ( .A1(n_284), .A2(n_130), .B1(n_135), .B2(n_136), .C(n_132), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_288), .B(n_5), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_288), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_289), .B(n_6), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_289), .B(n_6), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_274), .Y(n_329) );
NOR3xp33_ASAP7_75t_L g330 ( .A(n_286), .B(n_139), .C(n_145), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_274), .Y(n_331) );
NAND5xp2_ASAP7_75t_SL g332 ( .A(n_286), .B(n_8), .C(n_9), .D(n_10), .E(n_11), .Y(n_332) );
AOI21xp5_ASAP7_75t_L g333 ( .A1(n_284), .A2(n_231), .B(n_227), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_273), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_276), .Y(n_335) );
INVx2_ASAP7_75t_SL g336 ( .A(n_296), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_273), .B(n_8), .Y(n_337) );
NOR2xp33_ASAP7_75t_SL g338 ( .A(n_296), .B(n_182), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_290), .Y(n_339) );
OR2x6_ASAP7_75t_L g340 ( .A(n_297), .B(n_227), .Y(n_340) );
OAI222xp33_ASAP7_75t_L g341 ( .A1(n_309), .A2(n_295), .B1(n_291), .B2(n_290), .C1(n_271), .C2(n_272), .Y(n_341) );
NAND4xp25_ASAP7_75t_L g342 ( .A(n_313), .B(n_277), .C(n_293), .D(n_295), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_321), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_313), .A2(n_293), .B1(n_273), .B2(n_271), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_303), .B(n_271), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_326), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_309), .Y(n_347) );
AOI211xp5_ASAP7_75t_L g348 ( .A1(n_302), .A2(n_291), .B(n_272), .C(n_298), .Y(n_348) );
AOI221x1_ASAP7_75t_L g349 ( .A1(n_316), .A2(n_272), .B1(n_298), .B2(n_147), .C(n_145), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_317), .B(n_9), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_329), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_307), .B(n_10), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_336), .B(n_12), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_331), .Y(n_354) );
AOI322xp5_ASAP7_75t_L g355 ( .A1(n_319), .A2(n_13), .A3(n_14), .B1(n_15), .B2(n_16), .C1(n_17), .C2(n_18), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_307), .B(n_13), .Y(n_356) );
OAI322xp33_ASAP7_75t_L g357 ( .A1(n_320), .A2(n_335), .A3(n_339), .B1(n_319), .B2(n_311), .C1(n_336), .C2(n_327), .Y(n_357) );
OAI21xp5_ASAP7_75t_L g358 ( .A1(n_337), .A2(n_147), .B(n_145), .Y(n_358) );
INVxp67_ASAP7_75t_SL g359 ( .A(n_312), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_334), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_337), .Y(n_361) );
AND2x2_ASAP7_75t_SL g362 ( .A(n_300), .B(n_182), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_334), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_314), .A2(n_231), .B1(n_221), .B2(n_182), .Y(n_364) );
INVxp67_ASAP7_75t_L g365 ( .A(n_315), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_320), .B(n_16), .Y(n_366) );
AOI222xp33_ASAP7_75t_L g367 ( .A1(n_323), .A2(n_17), .B1(n_18), .B2(n_147), .C1(n_136), .C2(n_221), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_315), .B(n_136), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_308), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_304), .B(n_21), .Y(n_370) );
AOI322xp5_ASAP7_75t_L g371 ( .A1(n_323), .A2(n_136), .A3(n_193), .B1(n_196), .B2(n_198), .C1(n_202), .C2(n_192), .Y(n_371) );
AOI211xp5_ASAP7_75t_L g372 ( .A1(n_314), .A2(n_196), .B(n_193), .C(n_136), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_305), .Y(n_373) );
INVxp67_ASAP7_75t_L g374 ( .A(n_338), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_325), .B(n_22), .Y(n_375) );
AOI22xp5_ASAP7_75t_L g376 ( .A1(n_325), .A2(n_182), .B1(n_186), .B2(n_198), .Y(n_376) );
AOI22xp5_ASAP7_75t_L g377 ( .A1(n_327), .A2(n_186), .B1(n_198), .B2(n_192), .Y(n_377) );
OAI21xp5_ASAP7_75t_SL g378 ( .A1(n_328), .A2(n_184), .B(n_197), .Y(n_378) );
NAND3xp33_ASAP7_75t_L g379 ( .A(n_324), .B(n_203), .C(n_192), .Y(n_379) );
AOI221xp5_ASAP7_75t_L g380 ( .A1(n_332), .A2(n_164), .B1(n_159), .B2(n_155), .C(n_137), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_305), .Y(n_381) );
AOI211xp5_ASAP7_75t_L g382 ( .A1(n_328), .A2(n_142), .B(n_137), .C(n_189), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_306), .B(n_23), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_322), .Y(n_384) );
NOR2xp33_ASAP7_75t_SL g385 ( .A(n_322), .B(n_186), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_340), .B(n_25), .Y(n_386) );
NOR3xp33_ASAP7_75t_L g387 ( .A(n_366), .B(n_301), .C(n_318), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_346), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_362), .B(n_306), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_347), .B(n_322), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_351), .B(n_340), .Y(n_391) );
NAND3xp33_ASAP7_75t_SL g392 ( .A(n_372), .B(n_310), .C(n_330), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_343), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_342), .A2(n_340), .B1(n_333), .B2(n_186), .Y(n_394) );
NOR3xp33_ASAP7_75t_SL g395 ( .A(n_357), .B(n_340), .C(n_28), .Y(n_395) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_362), .B(n_197), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_343), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_354), .Y(n_398) );
NAND3xp33_ASAP7_75t_L g399 ( .A(n_348), .B(n_189), .C(n_181), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_345), .B(n_27), .Y(n_400) );
NAND3xp33_ASAP7_75t_L g401 ( .A(n_344), .B(n_189), .C(n_181), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_359), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_369), .Y(n_403) );
NOR2xp33_ASAP7_75t_R g404 ( .A(n_385), .B(n_32), .Y(n_404) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_344), .A2(n_186), .B(n_181), .Y(n_405) );
CKINVDCx20_ASAP7_75t_R g406 ( .A(n_365), .Y(n_406) );
XOR2xp5_ASAP7_75t_L g407 ( .A(n_361), .B(n_35), .Y(n_407) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_374), .A2(n_142), .B1(n_137), .B2(n_164), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_373), .B(n_36), .Y(n_409) );
INVxp67_ASAP7_75t_SL g410 ( .A(n_353), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_352), .B(n_37), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_381), .Y(n_412) );
OAI21xp5_ASAP7_75t_L g413 ( .A1(n_355), .A2(n_38), .B(n_39), .Y(n_413) );
NOR3xp33_ASAP7_75t_SL g414 ( .A(n_341), .B(n_41), .C(n_45), .Y(n_414) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_378), .A2(n_164), .B(n_159), .Y(n_415) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_352), .A2(n_159), .B1(n_142), .B2(n_137), .C(n_155), .Y(n_416) );
OAI322xp33_ASAP7_75t_L g417 ( .A1(n_350), .A2(n_46), .A3(n_48), .B1(n_49), .B2(n_50), .C1(n_51), .C2(n_55), .Y(n_417) );
INVx1_ASAP7_75t_SL g418 ( .A(n_353), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_403), .B(n_360), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g420 ( .A1(n_394), .A2(n_356), .B1(n_384), .B2(n_367), .Y(n_420) );
OAI211xp5_ASAP7_75t_L g421 ( .A1(n_395), .A2(n_350), .B(n_356), .C(n_358), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g422 ( .A1(n_410), .A2(n_363), .B1(n_364), .B2(n_375), .C(n_368), .Y(n_422) );
XNOR2xp5_ASAP7_75t_L g423 ( .A(n_406), .B(n_377), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_402), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_388), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_398), .Y(n_426) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_418), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_393), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_397), .B(n_349), .Y(n_429) );
NAND4xp25_ASAP7_75t_L g430 ( .A(n_413), .B(n_386), .C(n_376), .D(n_382), .Y(n_430) );
AOI321xp33_ASAP7_75t_L g431 ( .A1(n_410), .A2(n_370), .A3(n_383), .B1(n_371), .B2(n_380), .C(n_379), .Y(n_431) );
AO22x2_ASAP7_75t_L g432 ( .A1(n_389), .A2(n_370), .B1(n_57), .B2(n_58), .Y(n_432) );
NOR3xp33_ASAP7_75t_L g433 ( .A(n_392), .B(n_56), .C(n_60), .Y(n_433) );
INVxp67_ASAP7_75t_L g434 ( .A(n_391), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_412), .B(n_64), .Y(n_435) );
CKINVDCx16_ASAP7_75t_R g436 ( .A(n_404), .Y(n_436) );
OAI21xp33_ASAP7_75t_SL g437 ( .A1(n_389), .A2(n_67), .B(n_68), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_390), .Y(n_438) );
NOR2xp33_ASAP7_75t_R g439 ( .A(n_436), .B(n_411), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_424), .Y(n_440) );
O2A1O1Ixp33_ASAP7_75t_L g441 ( .A1(n_437), .A2(n_395), .B(n_387), .C(n_414), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_427), .Y(n_442) );
AOI222xp33_ASAP7_75t_L g443 ( .A1(n_421), .A2(n_423), .B1(n_432), .B2(n_422), .C1(n_425), .C2(n_426), .Y(n_443) );
AOI221xp5_ASAP7_75t_L g444 ( .A1(n_434), .A2(n_387), .B1(n_417), .B2(n_399), .C(n_401), .Y(n_444) );
NAND3xp33_ASAP7_75t_SL g445 ( .A(n_433), .B(n_404), .C(n_414), .Y(n_445) );
NOR2xp67_ASAP7_75t_L g446 ( .A(n_430), .B(n_396), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_419), .Y(n_447) );
NOR2xp67_ASAP7_75t_L g448 ( .A(n_429), .B(n_405), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_420), .A2(n_407), .B1(n_400), .B2(n_409), .Y(n_449) );
AND2x2_ASAP7_75t_SL g450 ( .A(n_429), .B(n_416), .Y(n_450) );
OAI221xp5_ASAP7_75t_L g451 ( .A1(n_431), .A2(n_408), .B1(n_415), .B2(n_137), .C(n_142), .Y(n_451) );
OAI221xp5_ASAP7_75t_L g452 ( .A1(n_438), .A2(n_153), .B1(n_171), .B2(n_419), .C(n_428), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g453 ( .A1(n_435), .A2(n_436), .B1(n_406), .B2(n_427), .Y(n_453) );
OAI211xp5_ASAP7_75t_SL g454 ( .A1(n_420), .A2(n_395), .B(n_421), .C(n_431), .Y(n_454) );
OAI211xp5_ASAP7_75t_L g455 ( .A1(n_437), .A2(n_421), .B(n_395), .C(n_420), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_447), .Y(n_456) );
NAND3xp33_ASAP7_75t_L g457 ( .A(n_443), .B(n_454), .C(n_455), .Y(n_457) );
CKINVDCx12_ASAP7_75t_R g458 ( .A(n_442), .Y(n_458) );
XNOR2xp5_ASAP7_75t_L g459 ( .A(n_453), .B(n_449), .Y(n_459) );
NOR2x1_ASAP7_75t_L g460 ( .A(n_457), .B(n_445), .Y(n_460) );
NAND3xp33_ASAP7_75t_L g461 ( .A(n_459), .B(n_443), .C(n_446), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_456), .B(n_450), .Y(n_462) );
INVx3_ASAP7_75t_L g463 ( .A(n_462), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_460), .Y(n_464) );
AO22x2_ASAP7_75t_L g465 ( .A1(n_464), .A2(n_461), .B1(n_458), .B2(n_440), .Y(n_465) );
AOI222xp33_ASAP7_75t_L g466 ( .A1(n_465), .A2(n_464), .B1(n_463), .B2(n_448), .C1(n_444), .C2(n_451), .Y(n_466) );
AOI221xp5_ASAP7_75t_L g467 ( .A1(n_466), .A2(n_463), .B1(n_439), .B2(n_441), .C(n_452), .Y(n_467) );
endmodule