module fake_jpeg_21369_n_103 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_103);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_103;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_20),
.B(n_6),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_28),
.Y(n_32)
);

BUFx2_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

AND2x4_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_27),
.B(n_30),
.Y(n_34)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_37),
.Y(n_59)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_42),
.Y(n_47)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_12),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_23),
.Y(n_42)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_40),
.B1(n_37),
.B2(n_41),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_46),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_19),
.B1(n_18),
.B2(n_16),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_48),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_39),
.B(n_23),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_51),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_19),
.B1(n_18),
.B2(n_16),
.Y(n_50)
);

NOR3xp33_ASAP7_75t_SL g65 ( 
.A(n_50),
.B(n_0),
.C(n_1),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_21),
.B1(n_12),
.B2(n_13),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_12),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_54),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_34),
.B(n_15),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_58),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_61),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_33),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_13),
.B(n_15),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_0),
.Y(n_62)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_SL g79 ( 
.A(n_62),
.B(n_60),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_51),
.B1(n_59),
.B2(n_48),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_3),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_4),
.Y(n_67)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_44),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_75),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_43),
.C(n_58),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_79),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_43),
.C(n_54),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_80),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_76),
.A2(n_73),
.B1(n_61),
.B2(n_65),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_68),
.B1(n_73),
.B2(n_70),
.Y(n_90)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_81),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_89),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_80),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_90),
.A2(n_91),
.B(n_92),
.Y(n_93)
);

NAND4xp25_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_69),
.C(n_62),
.D(n_79),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_86),
.C(n_84),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_95),
.C(n_57),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_86),
.C(n_43),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_7),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_99),
.C(n_8),
.Y(n_101)
);

AOI21xp33_ASAP7_75t_SL g99 ( 
.A1(n_93),
.A2(n_11),
.B(n_7),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_101),
.B(n_8),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);


endmodule