module fake_jpeg_30059_n_104 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_104);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_2),
.B(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

INVx2_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_22),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_26),
.B(n_2),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_0),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_48),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_49),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_38),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_1),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_52),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_51),
.A2(n_36),
.B(n_5),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_3),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_38),
.C(n_36),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_54),
.A2(n_56),
.B(n_57),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_51),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_58),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_45),
.B(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_49),
.B(n_44),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

AO21x2_ASAP7_75t_L g60 ( 
.A1(n_48),
.A2(n_40),
.B(n_35),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_61),
.B1(n_17),
.B2(n_18),
.Y(n_78)
);

OA21x2_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_37),
.B(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_50),
.B(n_4),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_63),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_SL g66 ( 
.A(n_64),
.B(n_6),
.C(n_8),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_66),
.B(n_68),
.Y(n_88)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_60),
.A2(n_37),
.B1(n_8),
.B2(n_6),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_69),
.A2(n_70),
.B1(n_76),
.B2(n_78),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_73),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_13),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_74),
.B(n_25),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_34),
.B1(n_15),
.B2(n_16),
.Y(n_76)
);

HAxp5_ASAP7_75t_SL g77 ( 
.A(n_57),
.B(n_14),
.CON(n_77),
.SN(n_77)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_65),
.A2(n_19),
.B(n_24),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_86),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_84),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_75),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_76),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_27),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_87),
.B(n_28),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_72),
.C(n_69),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_95),
.Y(n_98)
);

NAND2x1p5_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_79),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_86),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_94),
.A2(n_89),
.B1(n_81),
.B2(n_80),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_32),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_96),
.A2(n_92),
.B1(n_83),
.B2(n_91),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_97),
.A2(n_81),
.B(n_88),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_100),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_98),
.C(n_92),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_98),
.Y(n_104)
);


endmodule