module fake_aes_1214_n_605 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_605);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_605;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_73;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_593;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_243;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_89;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_446;
wire n_420;
wire n_423;
wire n_342;
wire n_165;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_493;
wire n_418;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g73 ( .A(n_32), .Y(n_73) );
CKINVDCx20_ASAP7_75t_R g74 ( .A(n_20), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_56), .Y(n_75) );
NOR2xp33_ASAP7_75t_L g76 ( .A(n_51), .B(n_21), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_40), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_68), .Y(n_78) );
INVxp67_ASAP7_75t_SL g79 ( .A(n_29), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_69), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_61), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_43), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_36), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_6), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_34), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_38), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_5), .Y(n_87) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_5), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_26), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_39), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_58), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_50), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_2), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_3), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_17), .Y(n_95) );
CKINVDCx16_ASAP7_75t_R g96 ( .A(n_49), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_27), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_7), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_19), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_67), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_16), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_11), .Y(n_102) );
INVxp67_ASAP7_75t_SL g103 ( .A(n_12), .Y(n_103) );
INVxp67_ASAP7_75t_L g104 ( .A(n_31), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_0), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_57), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_53), .Y(n_107) );
INVx3_ASAP7_75t_L g108 ( .A(n_70), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_12), .Y(n_109) );
CKINVDCx14_ASAP7_75t_R g110 ( .A(n_71), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_66), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_15), .Y(n_112) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_4), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_6), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_42), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_47), .Y(n_116) );
CKINVDCx16_ASAP7_75t_R g117 ( .A(n_8), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_24), .Y(n_118) );
NOR2xp67_ASAP7_75t_L g119 ( .A(n_63), .B(n_46), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_108), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_73), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_108), .Y(n_122) );
BUFx2_ASAP7_75t_L g123 ( .A(n_96), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g124 ( .A(n_108), .B(n_0), .Y(n_124) );
BUFx10_ASAP7_75t_L g125 ( .A(n_106), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_107), .Y(n_126) );
BUFx2_ASAP7_75t_L g127 ( .A(n_110), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_78), .Y(n_128) );
BUFx2_ASAP7_75t_L g129 ( .A(n_113), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_117), .Y(n_130) );
AND2x2_ASAP7_75t_SL g131 ( .A(n_73), .B(n_30), .Y(n_131) );
AND3x1_ASAP7_75t_L g132 ( .A(n_112), .B(n_1), .C(n_2), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_75), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_107), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_75), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_84), .B(n_1), .Y(n_136) );
INVxp67_ASAP7_75t_L g137 ( .A(n_84), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_116), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_105), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_116), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_77), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g142 ( .A(n_74), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_93), .B(n_3), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_77), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_80), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_104), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_93), .B(n_4), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_94), .B(n_7), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_80), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_81), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_94), .B(n_8), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_95), .B(n_9), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_81), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_95), .B(n_9), .Y(n_154) );
OAI21x1_ASAP7_75t_L g155 ( .A1(n_82), .A2(n_37), .B(n_72), .Y(n_155) );
INVxp67_ASAP7_75t_L g156 ( .A(n_123), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_127), .B(n_82), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_155), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_129), .B(n_112), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_150), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_128), .Y(n_161) );
NOR2x1p5_ASAP7_75t_L g162 ( .A(n_130), .B(n_103), .Y(n_162) );
NAND3x1_ASAP7_75t_L g163 ( .A(n_136), .B(n_154), .C(n_148), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_127), .B(n_97), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_150), .Y(n_165) );
AND2x4_ASAP7_75t_L g166 ( .A(n_129), .B(n_101), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_150), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_129), .B(n_101), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_127), .B(n_92), .Y(n_169) );
NAND2x1p5_ASAP7_75t_L g170 ( .A(n_131), .B(n_92), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_150), .Y(n_171) );
AND2x2_ASAP7_75t_SL g172 ( .A(n_131), .B(n_100), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_150), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_150), .Y(n_174) );
NAND2x1p5_ASAP7_75t_L g175 ( .A(n_131), .B(n_136), .Y(n_175) );
BUFx2_ASAP7_75t_L g176 ( .A(n_123), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_150), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_150), .Y(n_178) );
HB1xp67_ASAP7_75t_L g179 ( .A(n_123), .Y(n_179) );
INVx3_ASAP7_75t_L g180 ( .A(n_120), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_155), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_120), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_120), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_146), .B(n_97), .Y(n_184) );
AND2x4_ASAP7_75t_L g185 ( .A(n_122), .B(n_102), .Y(n_185) );
NOR2xp33_ASAP7_75t_SL g186 ( .A(n_131), .B(n_86), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_122), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_122), .Y(n_188) );
BUFx3_ASAP7_75t_L g189 ( .A(n_126), .Y(n_189) );
INVx4_ASAP7_75t_L g190 ( .A(n_141), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_141), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_141), .Y(n_192) );
INVx4_ASAP7_75t_SL g193 ( .A(n_121), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_126), .Y(n_194) );
BUFx3_ASAP7_75t_L g195 ( .A(n_126), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_146), .B(n_83), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_142), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_137), .B(n_102), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_137), .B(n_114), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_141), .Y(n_200) );
AND2x2_ASAP7_75t_SL g201 ( .A(n_132), .B(n_100), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_134), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_155), .Y(n_203) );
INVx6_ASAP7_75t_L g204 ( .A(n_125), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_141), .Y(n_205) );
BUFx2_ASAP7_75t_L g206 ( .A(n_139), .Y(n_206) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_136), .Y(n_207) );
INVx3_ASAP7_75t_L g208 ( .A(n_149), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g209 ( .A1(n_132), .A2(n_87), .B1(n_88), .B2(n_98), .Y(n_209) );
BUFx3_ASAP7_75t_L g210 ( .A(n_134), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_149), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_149), .Y(n_212) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_154), .A2(n_109), .B1(n_114), .B2(n_99), .Y(n_213) );
BUFx2_ASAP7_75t_L g214 ( .A(n_176), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_208), .Y(n_215) );
OAI21xp5_ASAP7_75t_L g216 ( .A1(n_191), .A2(n_133), .B(n_153), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_208), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_198), .B(n_125), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_208), .Y(n_219) );
AND2x4_ASAP7_75t_L g220 ( .A(n_166), .B(n_154), .Y(n_220) );
NAND3xp33_ASAP7_75t_SL g221 ( .A(n_161), .B(n_142), .C(n_152), .Y(n_221) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_176), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_166), .B(n_124), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_172), .A2(n_153), .B1(n_133), .B2(n_135), .Y(n_224) );
INVx4_ASAP7_75t_L g225 ( .A(n_193), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_169), .B(n_125), .Y(n_226) );
NOR3xp33_ASAP7_75t_SL g227 ( .A(n_197), .B(n_152), .C(n_151), .Y(n_227) );
NOR3xp33_ASAP7_75t_SL g228 ( .A(n_184), .B(n_151), .C(n_148), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_158), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_188), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_190), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_188), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_L g233 ( .A1(n_172), .A2(n_149), .B(n_121), .C(n_144), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_190), .Y(n_234) );
NOR3xp33_ASAP7_75t_SL g235 ( .A(n_196), .B(n_143), .C(n_147), .Y(n_235) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_158), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_190), .Y(n_237) );
BUFx3_ASAP7_75t_L g238 ( .A(n_204), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_198), .B(n_125), .Y(n_239) );
NOR2xp33_ASAP7_75t_R g240 ( .A(n_206), .B(n_125), .Y(n_240) );
BUFx3_ASAP7_75t_L g241 ( .A(n_204), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_190), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_182), .Y(n_243) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_179), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_191), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_182), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g247 ( .A1(n_186), .A2(n_144), .B1(n_135), .B2(n_124), .Y(n_247) );
NOR3xp33_ASAP7_75t_SL g248 ( .A(n_164), .B(n_143), .C(n_147), .Y(n_248) );
BUFx3_ASAP7_75t_L g249 ( .A(n_204), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_183), .Y(n_250) );
INVxp67_ASAP7_75t_L g251 ( .A(n_206), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_199), .B(n_149), .Y(n_252) );
BUFx3_ASAP7_75t_L g253 ( .A(n_204), .Y(n_253) );
BUFx2_ASAP7_75t_L g254 ( .A(n_156), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_172), .A2(n_145), .B1(n_109), .B2(n_138), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_L g256 ( .A1(n_207), .A2(n_145), .B(n_140), .C(n_138), .Y(n_256) );
INVx1_ASAP7_75t_SL g257 ( .A(n_166), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_192), .Y(n_258) );
BUFx2_ASAP7_75t_L g259 ( .A(n_166), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_192), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_200), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_199), .B(n_145), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_168), .Y(n_263) );
NOR3xp33_ASAP7_75t_SL g264 ( .A(n_157), .B(n_76), .C(n_79), .Y(n_264) );
OAI21xp5_ASAP7_75t_L g265 ( .A1(n_200), .A2(n_111), .B(n_85), .Y(n_265) );
NOR2x1p5_ASAP7_75t_L g266 ( .A(n_168), .B(n_111), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_168), .B(n_140), .Y(n_267) );
NAND2x1_ASAP7_75t_L g268 ( .A(n_205), .B(n_211), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_205), .Y(n_269) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_168), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_175), .B(n_138), .Y(n_271) );
NOR2xp67_ASAP7_75t_L g272 ( .A(n_180), .B(n_140), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_211), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_162), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_183), .Y(n_275) );
CKINVDCx14_ASAP7_75t_R g276 ( .A(n_240), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_270), .Y(n_277) );
INVx3_ASAP7_75t_L g278 ( .A(n_225), .Y(n_278) );
OR2x6_ASAP7_75t_L g279 ( .A(n_214), .B(n_175), .Y(n_279) );
CKINVDCx12_ASAP7_75t_R g280 ( .A(n_271), .Y(n_280) );
INVx1_ASAP7_75t_SL g281 ( .A(n_214), .Y(n_281) );
INVx3_ASAP7_75t_L g282 ( .A(n_225), .Y(n_282) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_218), .A2(n_158), .B(n_203), .Y(n_283) );
O2A1O1Ixp33_ASAP7_75t_L g284 ( .A1(n_233), .A2(n_175), .B(n_170), .C(n_159), .Y(n_284) );
INVx3_ASAP7_75t_L g285 ( .A(n_225), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_251), .B(n_159), .Y(n_286) );
NAND3xp33_ASAP7_75t_L g287 ( .A(n_248), .B(n_209), .C(n_213), .Y(n_287) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_229), .Y(n_288) );
AOI22xp33_ASAP7_75t_SL g289 ( .A1(n_263), .A2(n_170), .B1(n_201), .B2(n_220), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_220), .B(n_163), .Y(n_290) );
OR2x2_ASAP7_75t_L g291 ( .A(n_244), .B(n_222), .Y(n_291) );
NAND3xp33_ASAP7_75t_L g292 ( .A(n_228), .B(n_209), .C(n_201), .Y(n_292) );
NOR2xp67_ASAP7_75t_SL g293 ( .A(n_225), .B(n_193), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_259), .Y(n_294) );
BUFx12f_ASAP7_75t_L g295 ( .A(n_274), .Y(n_295) );
A2O1A1Ixp33_ASAP7_75t_L g296 ( .A1(n_256), .A2(n_185), .B(n_194), .C(n_187), .Y(n_296) );
BUFx4f_ASAP7_75t_L g297 ( .A(n_220), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_220), .B(n_163), .Y(n_298) );
NAND2xp5_ASAP7_75t_SL g299 ( .A(n_231), .B(n_193), .Y(n_299) );
AOI21xp33_ASAP7_75t_L g300 ( .A1(n_263), .A2(n_170), .B(n_201), .Y(n_300) );
OR2x6_ASAP7_75t_L g301 ( .A(n_259), .B(n_162), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_254), .Y(n_302) );
AND2x4_ASAP7_75t_L g303 ( .A(n_266), .B(n_159), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_262), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_223), .B(n_159), .Y(n_305) );
AOI22xp33_ASAP7_75t_SL g306 ( .A1(n_257), .A2(n_185), .B1(n_181), .B2(n_203), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_223), .B(n_212), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_254), .Y(n_308) );
NAND2x1p5_ASAP7_75t_L g309 ( .A(n_271), .B(n_185), .Y(n_309) );
NAND2xp5_ASAP7_75t_SL g310 ( .A(n_231), .B(n_193), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g311 ( .A(n_274), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_267), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_229), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_245), .Y(n_314) );
BUFx2_ASAP7_75t_L g315 ( .A(n_223), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_245), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_230), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_223), .A2(n_185), .B1(n_210), .B2(n_189), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_230), .Y(n_319) );
AND2x4_ASAP7_75t_L g320 ( .A(n_227), .B(n_193), .Y(n_320) );
CKINVDCx11_ASAP7_75t_R g321 ( .A(n_238), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_317), .Y(n_322) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_288), .Y(n_323) );
AOI221xp5_ASAP7_75t_L g324 ( .A1(n_287), .A2(n_235), .B1(n_264), .B2(n_221), .C(n_252), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_302), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_281), .B(n_239), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_319), .Y(n_327) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_308), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_288), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_289), .A2(n_224), .B1(n_255), .B2(n_247), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_304), .B(n_232), .Y(n_331) );
AOI22xp33_ASAP7_75t_SL g332 ( .A1(n_276), .A2(n_265), .B1(n_232), .B2(n_203), .Y(n_332) );
AO31x2_ASAP7_75t_L g333 ( .A1(n_296), .A2(n_134), .A3(n_187), .B(n_194), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_309), .B(n_216), .Y(n_334) );
OR2x4_ASAP7_75t_L g335 ( .A(n_291), .B(n_226), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_308), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_288), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_305), .B(n_258), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_288), .Y(n_339) );
CKINVDCx6p67_ASAP7_75t_R g340 ( .A(n_280), .Y(n_340) );
BUFx2_ASAP7_75t_L g341 ( .A(n_309), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g342 ( .A1(n_292), .A2(n_247), .B1(n_272), .B2(n_273), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_314), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_289), .A2(n_234), .B1(n_242), .B2(n_237), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_303), .A2(n_237), .B1(n_242), .B2(n_273), .Y(n_345) );
A2O1A1Ixp33_ASAP7_75t_L g346 ( .A1(n_284), .A2(n_305), .B(n_316), .C(n_296), .Y(n_346) );
INVx4_ASAP7_75t_L g347 ( .A(n_297), .Y(n_347) );
INVx3_ASAP7_75t_L g348 ( .A(n_278), .Y(n_348) );
A2O1A1Ixp33_ASAP7_75t_L g349 ( .A1(n_283), .A2(n_272), .B(n_260), .C(n_269), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_297), .B(n_189), .Y(n_350) );
OAI21x1_ASAP7_75t_L g351 ( .A1(n_329), .A2(n_299), .B(n_310), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_331), .B(n_312), .Y(n_352) );
AOI21x1_ASAP7_75t_L g353 ( .A1(n_329), .A2(n_119), .B(n_310), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_323), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_324), .A2(n_303), .B1(n_301), .B2(n_279), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_330), .A2(n_301), .B1(n_279), .B2(n_300), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_330), .A2(n_301), .B1(n_279), .B2(n_315), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_323), .Y(n_358) );
AOI221xp5_ASAP7_75t_L g359 ( .A1(n_338), .A2(n_286), .B1(n_298), .B2(n_290), .C(n_277), .Y(n_359) );
AOI22xp33_ASAP7_75t_SL g360 ( .A1(n_336), .A2(n_311), .B1(n_295), .B2(n_320), .Y(n_360) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_323), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_334), .A2(n_321), .B1(n_320), .B2(n_294), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_323), .Y(n_363) );
AOI22xp5_ASAP7_75t_L g364 ( .A1(n_334), .A2(n_318), .B1(n_306), .B2(n_307), .Y(n_364) );
INVxp67_ASAP7_75t_L g365 ( .A(n_328), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_331), .B(n_318), .Y(n_366) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_336), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_332), .A2(n_306), .B1(n_195), .B2(n_189), .Y(n_368) );
OA21x2_ASAP7_75t_L g369 ( .A1(n_349), .A2(n_115), .B(n_83), .Y(n_369) );
AOI21xp5_ASAP7_75t_L g370 ( .A1(n_346), .A2(n_313), .B(n_229), .Y(n_370) );
OAI21x1_ASAP7_75t_L g371 ( .A1(n_329), .A2(n_299), .B(n_278), .Y(n_371) );
OAI22x1_ASAP7_75t_L g372 ( .A1(n_325), .A2(n_115), .B1(n_118), .B2(n_91), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_338), .A2(n_258), .B1(n_269), .B2(n_261), .Y(n_373) );
AOI21xp5_ASAP7_75t_L g374 ( .A1(n_337), .A2(n_313), .B(n_229), .Y(n_374) );
OAI21x1_ASAP7_75t_L g375 ( .A1(n_337), .A2(n_282), .B(n_285), .Y(n_375) );
AOI322xp5_ASAP7_75t_L g376 ( .A1(n_355), .A2(n_322), .A3(n_327), .B1(n_332), .B2(n_341), .C1(n_343), .C2(n_118), .Y(n_376) );
NAND2xp5_ASAP7_75t_SL g377 ( .A(n_360), .B(n_343), .Y(n_377) );
OAI221xp5_ASAP7_75t_L g378 ( .A1(n_356), .A2(n_326), .B1(n_344), .B2(n_345), .C(n_342), .Y(n_378) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_367), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_352), .Y(n_380) );
AOI21xp33_ASAP7_75t_L g381 ( .A1(n_352), .A2(n_342), .B(n_326), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_357), .A2(n_347), .B1(n_322), .B2(n_327), .Y(n_382) );
INVx2_ASAP7_75t_SL g383 ( .A(n_366), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_354), .Y(n_384) );
AOI21xp5_ASAP7_75t_L g385 ( .A1(n_370), .A2(n_313), .B(n_323), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_354), .Y(n_386) );
AO21x2_ASAP7_75t_L g387 ( .A1(n_370), .A2(n_337), .B(n_339), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_365), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_373), .A2(n_335), .B1(n_340), .B2(n_347), .Y(n_389) );
INVx3_ASAP7_75t_L g390 ( .A(n_361), .Y(n_390) );
NOR2xp33_ASAP7_75t_R g391 ( .A(n_362), .B(n_340), .Y(n_391) );
A2O1A1Ixp33_ASAP7_75t_L g392 ( .A1(n_373), .A2(n_350), .B(n_253), .C(n_348), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_353), .Y(n_393) );
OAI21xp5_ASAP7_75t_L g394 ( .A1(n_368), .A2(n_260), .B(n_261), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_354), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_375), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_364), .A2(n_335), .B1(n_347), .B2(n_348), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_366), .A2(n_335), .B1(n_347), .B2(n_348), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_375), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_359), .B(n_195), .Y(n_400) );
NAND3xp33_ASAP7_75t_L g401 ( .A(n_369), .B(n_91), .C(n_90), .Y(n_401) );
INVx2_ASAP7_75t_SL g402 ( .A(n_361), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_359), .A2(n_348), .B1(n_202), .B2(n_210), .Y(n_403) );
AOI22xp33_ASAP7_75t_SL g404 ( .A1(n_368), .A2(n_339), .B1(n_323), .B2(n_90), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_372), .A2(n_195), .B1(n_202), .B2(n_210), .Y(n_405) );
AO21x2_ASAP7_75t_L g406 ( .A1(n_358), .A2(n_339), .B(n_85), .Y(n_406) );
BUFx3_ASAP7_75t_L g407 ( .A(n_361), .Y(n_407) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_372), .A2(n_180), .B1(n_89), .B2(n_202), .C(n_212), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_396), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_396), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_383), .B(n_333), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_383), .B(n_333), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g413 ( .A1(n_389), .A2(n_180), .B1(n_158), .B2(n_181), .C(n_203), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_399), .Y(n_414) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_379), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_380), .B(n_333), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_380), .B(n_333), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_399), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_384), .Y(n_419) );
AND2x4_ASAP7_75t_L g420 ( .A(n_407), .B(n_358), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_384), .Y(n_421) );
BUFx3_ASAP7_75t_L g422 ( .A(n_407), .Y(n_422) );
NOR2x1_ASAP7_75t_L g423 ( .A(n_389), .B(n_369), .Y(n_423) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_388), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_386), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_386), .B(n_333), .Y(n_426) );
HB1xp67_ASAP7_75t_SL g427 ( .A(n_398), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_398), .B(n_333), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_395), .Y(n_429) );
BUFx2_ASAP7_75t_L g430 ( .A(n_407), .Y(n_430) );
XNOR2xp5_ASAP7_75t_L g431 ( .A(n_377), .B(n_10), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_395), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_404), .A2(n_369), .B1(n_358), .B2(n_363), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_387), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_394), .B(n_369), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_387), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_381), .B(n_363), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_387), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_376), .B(n_363), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_393), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_394), .B(n_371), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_393), .Y(n_442) );
NAND2x1p5_ASAP7_75t_L g443 ( .A(n_390), .B(n_361), .Y(n_443) );
OAI33xp33_ASAP7_75t_L g444 ( .A1(n_397), .A2(n_13), .A3(n_14), .B1(n_15), .B2(n_16), .B3(n_17), .Y(n_444) );
AOI211x1_ASAP7_75t_L g445 ( .A1(n_378), .A2(n_13), .B(n_14), .C(n_18), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_390), .Y(n_446) );
INVx1_ASAP7_75t_SL g447 ( .A(n_391), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_390), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_402), .B(n_371), .Y(n_449) );
BUFx2_ASAP7_75t_L g450 ( .A(n_402), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_382), .B(n_351), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_406), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_406), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_406), .Y(n_454) );
OR2x2_ASAP7_75t_SL g455 ( .A(n_401), .B(n_361), .Y(n_455) );
AOI322xp5_ASAP7_75t_L g456 ( .A1(n_405), .A2(n_18), .A3(n_19), .B1(n_20), .B2(n_21), .C1(n_158), .C2(n_203), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_411), .B(n_401), .Y(n_457) );
NOR3xp33_ASAP7_75t_L g458 ( .A(n_444), .B(n_408), .C(n_400), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_431), .B(n_392), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_415), .B(n_403), .Y(n_460) );
NAND4xp25_ASAP7_75t_L g461 ( .A(n_445), .B(n_385), .C(n_167), .D(n_171), .Y(n_461) );
BUFx4f_ASAP7_75t_L g462 ( .A(n_443), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_431), .B(n_181), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_424), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_412), .B(n_181), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_426), .B(n_22), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_419), .B(n_275), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_423), .B(n_374), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_419), .B(n_275), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_442), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_421), .B(n_250), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_442), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_421), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_441), .B(n_23), .Y(n_474) );
OR2x6_ASAP7_75t_L g475 ( .A(n_423), .B(n_313), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_441), .B(n_25), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_416), .B(n_28), .Y(n_477) );
BUFx8_ASAP7_75t_SL g478 ( .A(n_430), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_417), .B(n_33), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_439), .B(n_246), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_417), .B(n_35), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_429), .B(n_246), .Y(n_482) );
BUFx2_ASAP7_75t_L g483 ( .A(n_450), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_425), .B(n_41), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_432), .B(n_243), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_432), .B(n_243), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_409), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_425), .B(n_44), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_414), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_447), .A2(n_229), .B1(n_236), .B2(n_217), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_435), .A2(n_236), .B1(n_217), .B2(n_215), .Y(n_491) );
AOI21xp33_ASAP7_75t_L g492 ( .A1(n_437), .A2(n_236), .B(n_177), .Y(n_492) );
NOR2xp33_ASAP7_75t_R g493 ( .A(n_427), .B(n_45), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_428), .B(n_48), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_445), .B(n_236), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_450), .B(n_52), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_440), .Y(n_497) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_430), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_456), .B(n_215), .Y(n_499) );
INVx1_ASAP7_75t_SL g500 ( .A(n_422), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_422), .B(n_54), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_456), .B(n_219), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_409), .Y(n_503) );
NAND2x1_ASAP7_75t_L g504 ( .A(n_453), .B(n_293), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_464), .Y(n_505) );
NOR4xp25_ASAP7_75t_L g506 ( .A(n_459), .B(n_433), .C(n_413), .D(n_451), .Y(n_506) );
OAI21xp33_ASAP7_75t_SL g507 ( .A1(n_494), .A2(n_452), .B(n_428), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_463), .A2(n_458), .B1(n_460), .B2(n_457), .Y(n_508) );
AOI31xp33_ASAP7_75t_L g509 ( .A1(n_493), .A2(n_452), .A3(n_454), .B(n_453), .Y(n_509) );
OAI322xp33_ASAP7_75t_L g510 ( .A1(n_463), .A2(n_434), .A3(n_436), .B1(n_438), .B2(n_410), .C1(n_418), .C2(n_448), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_483), .B(n_410), .Y(n_511) );
NAND3xp33_ASAP7_75t_SL g512 ( .A(n_493), .B(n_453), .C(n_454), .Y(n_512) );
NOR2xp33_ASAP7_75t_SL g513 ( .A(n_478), .B(n_422), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_470), .Y(n_514) );
NAND3xp33_ASAP7_75t_SL g515 ( .A(n_496), .B(n_454), .C(n_438), .Y(n_515) );
OAI21xp5_ASAP7_75t_L g516 ( .A1(n_461), .A2(n_448), .B(n_446), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_494), .A2(n_455), .B1(n_410), .B2(n_418), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_472), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_498), .B(n_420), .Y(n_519) );
NOR3xp33_ASAP7_75t_L g520 ( .A(n_480), .B(n_438), .C(n_436), .Y(n_520) );
NOR2xp33_ASAP7_75t_R g521 ( .A(n_500), .B(n_55), .Y(n_521) );
OAI21xp33_ASAP7_75t_L g522 ( .A1(n_474), .A2(n_436), .B(n_434), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_489), .Y(n_523) );
AOI32xp33_ASAP7_75t_L g524 ( .A1(n_474), .A2(n_449), .A3(n_434), .B1(n_420), .B2(n_253), .Y(n_524) );
AOI32xp33_ASAP7_75t_L g525 ( .A1(n_476), .A2(n_449), .A3(n_420), .B1(n_253), .B2(n_282), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_462), .B(n_443), .Y(n_526) );
INVxp67_ASAP7_75t_L g527 ( .A(n_478), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_473), .Y(n_528) );
INVx1_ASAP7_75t_SL g529 ( .A(n_501), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_487), .Y(n_530) );
NAND3xp33_ASAP7_75t_L g531 ( .A(n_468), .B(n_178), .C(n_177), .Y(n_531) );
NOR2x1_ASAP7_75t_L g532 ( .A(n_504), .B(n_249), .Y(n_532) );
OAI221xp5_ASAP7_75t_L g533 ( .A1(n_491), .A2(n_249), .B1(n_241), .B2(n_238), .C(n_178), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_497), .B(n_173), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_503), .B(n_173), .Y(n_535) );
OAI21xp5_ASAP7_75t_L g536 ( .A1(n_477), .A2(n_479), .B(n_481), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_487), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_465), .B(n_59), .Y(n_538) );
OAI221xp5_ASAP7_75t_L g539 ( .A1(n_491), .A2(n_268), .B1(n_174), .B2(n_165), .C(n_160), .Y(n_539) );
OAI221xp5_ASAP7_75t_L g540 ( .A1(n_499), .A2(n_174), .B1(n_165), .B2(n_160), .C(n_65), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_467), .Y(n_541) );
NAND3xp33_ASAP7_75t_SL g542 ( .A(n_490), .B(n_60), .C(n_62), .Y(n_542) );
OAI221xp5_ASAP7_75t_L g543 ( .A1(n_508), .A2(n_502), .B1(n_490), .B2(n_468), .C(n_475), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_509), .A2(n_462), .B1(n_475), .B2(n_479), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_530), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_505), .Y(n_546) );
AOI21xp33_ASAP7_75t_SL g547 ( .A1(n_527), .A2(n_475), .B(n_481), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_512), .A2(n_462), .B(n_495), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_541), .B(n_477), .Y(n_549) );
INVx2_ASAP7_75t_SL g550 ( .A(n_521), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_514), .B(n_466), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_518), .Y(n_552) );
OAI21xp5_ASAP7_75t_SL g553 ( .A1(n_525), .A2(n_488), .B(n_484), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_523), .Y(n_554) );
CKINVDCx16_ASAP7_75t_R g555 ( .A(n_513), .Y(n_555) );
NOR2x1_ASAP7_75t_L g556 ( .A(n_542), .B(n_482), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_528), .Y(n_557) );
XNOR2x2_ASAP7_75t_L g558 ( .A(n_536), .B(n_488), .Y(n_558) );
INVxp67_ASAP7_75t_L g559 ( .A(n_511), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_537), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_520), .B(n_471), .Y(n_561) );
BUFx2_ASAP7_75t_L g562 ( .A(n_519), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_506), .B(n_469), .Y(n_563) );
NOR2x1_ASAP7_75t_L g564 ( .A(n_542), .B(n_486), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_529), .B(n_492), .Y(n_565) );
NOR3xp33_ASAP7_75t_SL g566 ( .A(n_507), .B(n_540), .C(n_515), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_510), .B(n_484), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_516), .B(n_485), .Y(n_568) );
INVx2_ASAP7_75t_SL g569 ( .A(n_555), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_566), .A2(n_517), .B1(n_524), .B2(n_522), .Y(n_570) );
INVxp67_ASAP7_75t_L g571 ( .A(n_563), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_550), .B(n_526), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_545), .Y(n_573) );
INVx8_ASAP7_75t_L g574 ( .A(n_556), .Y(n_574) );
NAND3xp33_ASAP7_75t_L g575 ( .A(n_566), .B(n_517), .C(n_540), .Y(n_575) );
INVxp67_ASAP7_75t_L g576 ( .A(n_564), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_562), .B(n_532), .Y(n_577) );
AND2x4_ASAP7_75t_L g578 ( .A(n_559), .B(n_538), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_560), .B(n_534), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_558), .A2(n_531), .B1(n_539), .B2(n_533), .Y(n_580) );
INVxp67_ASAP7_75t_L g581 ( .A(n_543), .Y(n_581) );
OAI22x1_ASAP7_75t_L g582 ( .A1(n_569), .A2(n_567), .B1(n_559), .B2(n_546), .Y(n_582) );
AO22x2_ASAP7_75t_L g583 ( .A1(n_571), .A2(n_544), .B1(n_548), .B2(n_552), .Y(n_583) );
CKINVDCx16_ASAP7_75t_R g584 ( .A(n_572), .Y(n_584) );
NOR4xp25_ASAP7_75t_L g585 ( .A(n_571), .B(n_557), .C(n_554), .D(n_553), .Y(n_585) );
INVx1_ASAP7_75t_SL g586 ( .A(n_578), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_576), .B(n_561), .Y(n_587) );
AOI21xp33_ASAP7_75t_SL g588 ( .A1(n_574), .A2(n_568), .B(n_565), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_581), .A2(n_565), .B1(n_549), .B2(n_551), .Y(n_589) );
INVx2_ASAP7_75t_SL g590 ( .A(n_574), .Y(n_590) );
AOI32xp33_ASAP7_75t_L g591 ( .A1(n_570), .A2(n_64), .A3(n_535), .B1(n_577), .B2(n_580), .Y(n_591) );
NAND4xp75_ASAP7_75t_L g592 ( .A(n_579), .B(n_569), .C(n_550), .D(n_566), .Y(n_592) );
NAND4xp25_ASAP7_75t_SL g593 ( .A(n_573), .B(n_575), .C(n_447), .D(n_547), .Y(n_593) );
XNOR2x2_ASAP7_75t_L g594 ( .A(n_575), .B(n_558), .Y(n_594) );
INVx1_ASAP7_75t_SL g595 ( .A(n_590), .Y(n_595) );
AND2x2_ASAP7_75t_SL g596 ( .A(n_585), .B(n_584), .Y(n_596) );
XOR2xp5_ASAP7_75t_L g597 ( .A(n_592), .B(n_594), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_595), .B(n_587), .Y(n_598) );
XNOR2xp5_ASAP7_75t_L g599 ( .A(n_597), .B(n_589), .Y(n_599) );
NOR3xp33_ASAP7_75t_L g600 ( .A(n_598), .B(n_595), .C(n_593), .Y(n_600) );
NOR3xp33_ASAP7_75t_SL g601 ( .A(n_599), .B(n_596), .C(n_591), .Y(n_601) );
BUFx2_ASAP7_75t_L g602 ( .A(n_601), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_600), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_602), .A2(n_582), .B1(n_583), .B2(n_586), .Y(n_604) );
AOI221xp5_ASAP7_75t_L g605 ( .A1(n_604), .A2(n_602), .B1(n_603), .B2(n_583), .C(n_588), .Y(n_605) );
endmodule