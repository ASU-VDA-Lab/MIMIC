module fake_ariane_53_n_234 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_38, n_2, n_18, n_32, n_28, n_37, n_9, n_11, n_34, n_26, n_3, n_14, n_0, n_36, n_33, n_19, n_30, n_39, n_31, n_16, n_5, n_12, n_15, n_21, n_23, n_35, n_10, n_25, n_234);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_38;
input n_2;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_11;
input n_34;
input n_26;
input n_3;
input n_14;
input n_0;
input n_36;
input n_33;
input n_19;
input n_30;
input n_39;
input n_31;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_35;
input n_10;
input n_25;

output n_234;

wire n_83;
wire n_233;
wire n_56;
wire n_60;
wire n_170;
wire n_190;
wire n_160;
wire n_64;
wire n_179;
wire n_180;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_195;
wire n_213;
wire n_47;
wire n_110;
wire n_153;
wire n_197;
wire n_221;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_203;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_40;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_205;
wire n_71;
wire n_109;
wire n_208;
wire n_96;
wire n_156;
wire n_209;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_187;
wire n_132;
wire n_62;
wire n_210;
wire n_147;
wire n_204;
wire n_225;
wire n_200;
wire n_51;
wire n_166;
wire n_76;
wire n_218;
wire n_103;
wire n_79;
wire n_226;
wire n_46;
wire n_220;
wire n_84;
wire n_199;
wire n_91;
wire n_159;
wire n_107;
wire n_189;
wire n_72;
wire n_105;
wire n_128;
wire n_217;
wire n_44;
wire n_224;
wire n_82;
wire n_178;
wire n_42;
wire n_131;
wire n_57;
wire n_201;
wire n_229;
wire n_70;
wire n_222;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_144;
wire n_130;
wire n_214;
wire n_227;
wire n_48;
wire n_94;
wire n_101;
wire n_134;
wire n_188;
wire n_185;
wire n_58;
wire n_65;
wire n_123;
wire n_212;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_198;
wire n_148;
wire n_232;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_228;
wire n_118;
wire n_93;
wire n_121;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_196;
wire n_125;
wire n_168;
wire n_43;
wire n_81;
wire n_87;
wire n_206;
wire n_207;
wire n_41;
wire n_219;
wire n_140;
wire n_55;
wire n_191;
wire n_151;
wire n_136;
wire n_231;
wire n_192;
wire n_80;
wire n_146;
wire n_230;
wire n_211;
wire n_194;
wire n_97;
wire n_154;
wire n_215;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_202;
wire n_145;
wire n_78;
wire n_193;
wire n_59;
wire n_63;
wire n_99;
wire n_216;
wire n_155;
wire n_127;
wire n_223;
wire n_54;

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVxp33_ASAP7_75t_SL g44 ( 
.A(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVxp67_ASAP7_75t_SL g57 ( 
.A(n_11),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_8),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_12),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_13),
.Y(n_70)
);

INVxp67_ASAP7_75t_SL g71 ( 
.A(n_29),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_0),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_46),
.Y(n_73)
);

AND2x6_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_17),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_0),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_1),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_2),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_4),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

OA21x2_ASAP7_75t_L g83 ( 
.A1(n_45),
.A2(n_4),
.B(n_5),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_44),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

AND2x4_ASAP7_75t_L g96 ( 
.A(n_47),
.B(n_9),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_63),
.Y(n_100)
);

NAND2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_58),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_96),
.B(n_44),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_49),
.B1(n_58),
.B2(n_69),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_60),
.B(n_70),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g105 ( 
.A(n_88),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_68),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_67),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_66),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_R g111 ( 
.A(n_89),
.B(n_65),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_65),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

INVx4_ASAP7_75t_SL g117 ( 
.A(n_74),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_102),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_96),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_79),
.B1(n_90),
.B2(n_76),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_79),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_95),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_111),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_94),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_82),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_93),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_105),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

INVxp67_ASAP7_75t_SL g137 ( 
.A(n_128),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_101),
.B(n_80),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_72),
.Y(n_140)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_122),
.A2(n_105),
.B1(n_85),
.B2(n_78),
.Y(n_142)
);

CKINVDCx11_ASAP7_75t_R g143 ( 
.A(n_134),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_72),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_134),
.B(n_123),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_119),
.A2(n_75),
.B1(n_77),
.B2(n_71),
.Y(n_146)
);

AND2x4_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_117),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_77),
.Y(n_148)
);

AO21x2_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_101),
.B(n_112),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_122),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_98),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_153),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_144),
.A2(n_130),
.B1(n_57),
.B2(n_121),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_153),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_155),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_126),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

CKINVDCx6p67_ASAP7_75t_R g171 ( 
.A(n_143),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_163),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_161),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_148),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_137),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_142),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

AOI222xp33_ASAP7_75t_L g190 ( 
.A1(n_181),
.A2(n_142),
.B1(n_152),
.B2(n_143),
.C1(n_145),
.C2(n_146),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_184),
.A2(n_139),
.B(n_157),
.Y(n_191)
);

NAND3xp33_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_154),
.C(n_167),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_171),
.Y(n_193)
);

OAI33xp33_ASAP7_75t_L g194 ( 
.A1(n_175),
.A2(n_168),
.A3(n_170),
.B1(n_126),
.B2(n_172),
.B3(n_52),
.Y(n_194)
);

INVx4_ASAP7_75t_SL g195 ( 
.A(n_179),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_180),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_162),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_196),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_197),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_192),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_182),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_177),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_185),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_198),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_204),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_83),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_199),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_177),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_203),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_186),
.Y(n_213)
);

OAI33xp33_ASAP7_75t_L g214 ( 
.A1(n_205),
.A2(n_52),
.A3(n_186),
.B1(n_176),
.B2(n_173),
.B3(n_194),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_195),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_198),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_210),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_206),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_208),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_216),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_211),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_217),
.A2(n_194),
.B1(n_176),
.B2(n_173),
.Y(n_224)
);

AOI211xp5_ASAP7_75t_L g225 ( 
.A1(n_223),
.A2(n_82),
.B(n_97),
.C(n_209),
.Y(n_225)
);

NOR3xp33_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_221),
.C(n_219),
.Y(n_226)
);

NAND3xp33_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_222),
.C(n_220),
.Y(n_227)
);

NAND3xp33_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_225),
.C(n_224),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_228),
.Y(n_229)
);

OAI221xp5_ASAP7_75t_L g230 ( 
.A1(n_229),
.A2(n_129),
.B1(n_150),
.B2(n_141),
.C(n_74),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_230),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_231),
.A2(n_149),
.B(n_20),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_232),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_233),
.A2(n_149),
.B(n_39),
.Y(n_234)
);


endmodule