module fake_jpeg_15031_n_123 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_123);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_123;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_58),
.Y(n_66)
);

BUFx4f_ASAP7_75t_SL g58 ( 
.A(n_44),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_56),
.B(n_42),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_67),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_53),
.A2(n_41),
.B1(n_44),
.B2(n_51),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_43),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_71),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_45),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_1),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_40),
.B1(n_37),
.B2(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_73),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_49),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_46),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_69),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_80),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_78),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_91)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_83),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_67),
.Y(n_83)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_85),
.A2(n_73),
.B1(n_47),
.B2(n_7),
.Y(n_98)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_87),
.Y(n_95)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_4),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_91),
.A2(n_98),
.B1(n_75),
.B2(n_85),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_76),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_92),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_63),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_94),
.C(n_75),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_40),
.C(n_37),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_84),
.C(n_47),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_99),
.A2(n_103),
.B(n_97),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_102),
.Y(n_106)
);

BUFx4f_ASAP7_75t_SL g102 ( 
.A(n_89),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_87),
.B1(n_79),
.B2(n_96),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_104),
.A2(n_107),
.B1(n_108),
.B2(n_5),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_25),
.C(n_36),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_99),
.A2(n_98),
.B1(n_90),
.B2(n_95),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_106),
.B(n_94),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_104),
.A2(n_23),
.B(n_32),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_113),
.A2(n_111),
.B1(n_112),
.B2(n_6),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_114),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_13),
.B1(n_15),
.B2(n_17),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_18),
.C(n_20),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_22),
.B(n_26),
.C(n_28),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_120),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_29),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_30),
.Y(n_123)
);


endmodule