module fake_jpeg_23165_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_43),
.B1(n_17),
.B2(n_26),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_40),
.Y(n_45)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_42),
.Y(n_49)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_17),
.B1(n_30),
.B2(n_23),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_28),
.B1(n_43),
.B2(n_26),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_18),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

NAND2xp33_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_23),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_59),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_18),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_16),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_28),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_27),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_58),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_27),
.Y(n_59)
);

HAxp5_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_17),
.CON(n_60),
.SN(n_60)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_33),
.B1(n_34),
.B2(n_28),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_47),
.B(n_32),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_71),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_63),
.A2(n_73),
.B1(n_75),
.B2(n_88),
.Y(n_117)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_64),
.B(n_69),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_16),
.Y(n_66)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

AO22x1_ASAP7_75t_L g68 ( 
.A1(n_60),
.A2(n_33),
.B1(n_44),
.B2(n_38),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_68),
.A2(n_84),
.B1(n_57),
.B2(n_61),
.Y(n_92)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_70),
.A2(n_49),
.B1(n_45),
.B2(n_59),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_47),
.B(n_32),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_56),
.A2(n_26),
.B1(n_41),
.B2(n_33),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_58),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_50),
.A2(n_41),
.B1(n_31),
.B2(n_32),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_45),
.B1(n_59),
.B2(n_61),
.Y(n_98)
);

CKINVDCx5p33_ASAP7_75t_R g82 ( 
.A(n_61),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_82),
.Y(n_120)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_46),
.A2(n_20),
.B1(n_29),
.B2(n_25),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_22),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_45),
.B(n_20),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_90),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_69),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_96),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_92),
.A2(n_98),
.B1(n_105),
.B2(n_63),
.Y(n_126)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_77),
.B1(n_76),
.B2(n_85),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_111),
.Y(n_140)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_80),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_103),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_77),
.A2(n_56),
.B1(n_52),
.B2(n_51),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_68),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_108),
.B(n_110),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_58),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_80),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_113),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_35),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_114),
.B(n_89),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_75),
.Y(n_118)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_118),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_121),
.A2(n_146),
.B1(n_148),
.B2(n_109),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_67),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_122),
.A2(n_124),
.B(n_132),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_123),
.Y(n_152)
);

AND2x4_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_67),
.Y(n_124)
);

BUFx8_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_127),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_126),
.A2(n_133),
.B1(n_142),
.B2(n_144),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_131),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_67),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_98),
.A2(n_81),
.B1(n_84),
.B2(n_70),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_72),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_138),
.C(n_145),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_72),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_95),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_110),
.A2(n_70),
.B1(n_88),
.B2(n_52),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_108),
.A2(n_70),
.B1(n_51),
.B2(n_52),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_97),
.B(n_101),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_105),
.A2(n_51),
.B1(n_52),
.B2(n_87),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_112),
.A2(n_71),
.B(n_62),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_147),
.A2(n_114),
.B(n_115),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_100),
.A2(n_51),
.B1(n_83),
.B2(n_90),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_149),
.B(n_150),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_124),
.A2(n_112),
.B(n_109),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_151),
.A2(n_155),
.B1(n_157),
.B2(n_172),
.Y(n_185)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_153),
.B(n_162),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_135),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_154),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_148),
.A2(n_117),
.B1(n_115),
.B2(n_113),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_156),
.B(n_161),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_124),
.A2(n_119),
.B1(n_95),
.B2(n_103),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_143),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_160),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_123),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_163),
.B(n_167),
.Y(n_211)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_140),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_169),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_124),
.B(n_134),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_129),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_178),
.Y(n_191)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_125),
.Y(n_171)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_126),
.A2(n_94),
.B1(n_93),
.B2(n_99),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_116),
.C(n_93),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_147),
.C(n_132),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_141),
.A2(n_120),
.B(n_29),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_179),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_142),
.Y(n_177)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_122),
.A2(n_99),
.B(n_116),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_128),
.B(n_94),
.Y(n_180)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_128),
.B(n_118),
.Y(n_181)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_184),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_163),
.A2(n_133),
.B1(n_132),
.B2(n_122),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_187),
.A2(n_193),
.B1(n_173),
.B2(n_179),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_188),
.B(n_152),
.C(n_171),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_168),
.A2(n_127),
.B1(n_145),
.B2(n_107),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_118),
.B1(n_137),
.B2(n_130),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_195),
.A2(n_196),
.B1(n_198),
.B2(n_199),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_175),
.A2(n_49),
.B1(n_102),
.B2(n_24),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_177),
.A2(n_49),
.B1(n_24),
.B2(n_19),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_178),
.A2(n_49),
.B1(n_24),
.B2(n_19),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_164),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_161),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_27),
.Y(n_204)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_204),
.Y(n_214)
);

XNOR2x1_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_44),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_166),
.Y(n_216)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_207),
.B(n_209),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_149),
.B(n_27),
.Y(n_208)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_208),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_154),
.B(n_25),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_162),
.A2(n_38),
.B1(n_36),
.B2(n_35),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_210),
.A2(n_212),
.B1(n_213),
.B2(n_159),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_151),
.A2(n_36),
.B1(n_34),
.B2(n_16),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_155),
.A2(n_34),
.B1(n_16),
.B2(n_2),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_190),
.A2(n_176),
.B1(n_157),
.B2(n_150),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_215),
.A2(n_225),
.B1(n_198),
.B2(n_200),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_220),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_183),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_217),
.Y(n_247)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_218),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_202),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_219),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_158),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_221),
.A2(n_195),
.B1(n_212),
.B2(n_213),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_158),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_224),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_191),
.A2(n_208),
.B(n_205),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_190),
.A2(n_160),
.B1(n_156),
.B2(n_166),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_189),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_236),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_191),
.B(n_169),
.Y(n_229)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_204),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_234),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_194),
.C(n_210),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_182),
.B(n_152),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_233),
.B(n_238),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_184),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_193),
.B(n_200),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_34),
.Y(n_260)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_197),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_237),
.A2(n_231),
.B1(n_226),
.B2(n_185),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_182),
.B(n_206),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_187),
.B(n_167),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_188),
.Y(n_248)
);

AND2x4_ASAP7_75t_L g240 ( 
.A(n_239),
.B(n_229),
.Y(n_240)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_240),
.Y(n_266)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_241),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_251),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_215),
.B(n_203),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_250),
.B(n_236),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_192),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_252),
.A2(n_254),
.B1(n_231),
.B2(n_228),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_226),
.A2(n_201),
.B1(n_192),
.B2(n_196),
.Y(n_253)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_253),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_257),
.C(n_258),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_223),
.B(n_232),
.C(n_221),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_199),
.C(n_153),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_234),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_249),
.B(n_225),
.Y(n_262)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_262),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_263),
.A2(n_275),
.B1(n_240),
.B2(n_258),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_218),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_268),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_224),
.C(n_216),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_273),
.C(n_274),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_230),
.Y(n_268)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_269),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_227),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_271),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_214),
.C(n_222),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_214),
.C(n_1),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_240),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_8),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_8),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_251),
.C(n_240),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_260),
.C(n_253),
.Y(n_289)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_279),
.Y(n_299)
);

BUFx24_ASAP7_75t_SL g281 ( 
.A(n_269),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_281),
.B(n_284),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_272),
.A2(n_255),
.B1(n_254),
.B2(n_256),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_283),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_273),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_242),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_285),
.B(n_291),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_266),
.A2(n_246),
.B(n_243),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_286),
.A2(n_292),
.B(n_9),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_261),
.Y(n_294)
);

MAJx2_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_246),
.C(n_241),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_290),
.B(n_0),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_8),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_304),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_261),
.C(n_264),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_295),
.A2(n_297),
.B(n_301),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_280),
.A2(n_264),
.B(n_1),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_298),
.B(n_300),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_293),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_289),
.C(n_285),
.Y(n_301)
);

XOR2x2_ASAP7_75t_SL g309 ( 
.A(n_302),
.B(n_10),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_290),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_282),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_284),
.A2(n_0),
.B(n_4),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_305),
.A2(n_10),
.B1(n_15),
.B2(n_11),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_312),
.Y(n_317)
);

AOI21x1_ASAP7_75t_L g319 ( 
.A1(n_309),
.A2(n_302),
.B(n_304),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_313),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_287),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_10),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_11),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_306),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_299),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_321),
.Y(n_325)
);

NOR2x1_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_309),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_320),
.A2(n_322),
.B(n_311),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_296),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_308),
.A2(n_295),
.B(n_297),
.Y(n_322)
);

NAND4xp25_ASAP7_75t_SL g326 ( 
.A(n_323),
.B(n_324),
.C(n_311),
.D(n_317),
.Y(n_326)
);

OAI21xp33_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_316),
.B(n_325),
.Y(n_327)
);

OAI321xp33_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_15),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C(n_4),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_328),
.A2(n_4),
.B(n_5),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_15),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_7),
.Y(n_331)
);


endmodule