module real_jpeg_7868_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_17;
wire n_57;
wire n_43;
wire n_37;
wire n_21;
wire n_54;
wire n_65;
wire n_35;
wire n_38;
wire n_33;
wire n_50;
wire n_29;
wire n_55;
wire n_69;
wire n_49;
wire n_52;
wire n_31;
wire n_58;
wire n_67;
wire n_63;
wire n_12;
wire n_68;
wire n_24;
wire n_66;
wire n_34;
wire n_72;
wire n_28;
wire n_44;
wire n_60;
wire n_46;
wire n_62;
wire n_59;
wire n_64;
wire n_23;
wire n_47;
wire n_11;
wire n_14;
wire n_51;
wire n_45;
wire n_25;
wire n_71;
wire n_61;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_39;
wire n_40;
wire n_36;
wire n_70;
wire n_41;
wire n_26;
wire n_56;
wire n_20;
wire n_48;
wire n_19;
wire n_32;
wire n_30;
wire n_27;
wire n_16;
wire n_15;
wire n_13;

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_0),
.A2(n_16),
.B1(n_17),
.B2(n_23),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_1),
.A2(n_28),
.B(n_30),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_1),
.B(n_28),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_SL g63 ( 
.A(n_5),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_7),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_7),
.A2(n_18),
.B1(n_28),
.B2(n_29),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_8),
.A2(n_16),
.B1(n_17),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_8),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_9),
.A2(n_16),
.B1(n_17),
.B2(n_37),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_57),
.Y(n_10)
);

AOI21xp5_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_43),
.B(n_56),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_24),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_13),
.B(n_24),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_15),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_20),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_16),
.A2(n_17),
.B1(n_32),
.B2(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_16),
.B(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_16),
.B(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_17),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_19),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_20),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_22),
.A2(n_47),
.B1(n_48),
.B2(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_38),
.B2(n_42),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_25),
.B(n_42),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_31),
.B1(n_34),
.B2(n_36),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_SL g31 ( 
.A1(n_28),
.A2(n_32),
.B(n_33),
.C(n_34),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_32),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_28),
.A2(n_29),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_31),
.A2(n_34),
.B1(n_36),
.B2(n_66),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_32),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_34),
.B(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_38),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_51),
.B(n_55),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_49),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_50),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_71),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_70),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_70),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx24_ASAP7_75t_SL g73 ( 
.A(n_60),
.Y(n_73)
);

FAx1_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_65),
.CI(n_67),
.CON(n_60),
.SN(n_60)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_63),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);


endmodule