module real_jpeg_31877_n_17 (n_8, n_0, n_141, n_2, n_139, n_142, n_143, n_10, n_137, n_9, n_12, n_135, n_134, n_6, n_136, n_133, n_11, n_14, n_138, n_7, n_3, n_5, n_4, n_1, n_140, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_141;
input n_2;
input n_139;
input n_142;
input n_143;
input n_10;
input n_137;
input n_9;
input n_12;
input n_135;
input n_134;
input n_6;
input n_136;
input n_133;
input n_11;
input n_14;
input n_138;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_140;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

AOI221xp5_ASAP7_75t_L g49 ( 
.A1(n_0),
.A2(n_14),
.B1(n_50),
.B2(n_55),
.C(n_58),
.Y(n_49)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_1),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_2),
.B(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_3),
.A2(n_19),
.B1(n_20),
.B2(n_25),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_5),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_5),
.B(n_124),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_6),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_21),
.Y(n_20)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_9),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_9),
.B(n_108),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_10),
.B(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_10),
.Y(n_120)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_11),
.Y(n_100)
);

AOI322xp5_ASAP7_75t_L g116 ( 
.A1(n_11),
.A2(n_95),
.A3(n_97),
.B1(n_102),
.B2(n_117),
.C1(n_119),
.C2(n_143),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_12),
.B(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_13),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_13),
.B(n_83),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_14),
.B(n_50),
.C(n_55),
.Y(n_61)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_15),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_15),
.B(n_104),
.Y(n_115)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_26),
.Y(n_17)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_35),
.B(n_130),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_34),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_29),
.B(n_34),
.Y(n_131)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp67_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_122),
.B(n_129),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_79),
.B(n_112),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_73),
.C(n_74),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_62),
.B(n_72),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_49),
.B1(n_60),
.B2(n_61),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_51),
.B(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_135),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_71),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_71),
.Y(n_72)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NOR4xp25_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_88),
.C(n_101),
.D(n_107),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_87),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_105),
.Y(n_104)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_88),
.A2(n_113),
.B(n_116),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_95),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NOR3xp33_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_107),
.C(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_100),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_140),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OA21x2_ASAP7_75t_SL g113 ( 
.A1(n_101),
.A2(n_114),
.B(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_106),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2x1_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_128),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_133),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_134),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_136),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_137),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_138),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_139),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_141),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_142),
.Y(n_109)
);


endmodule