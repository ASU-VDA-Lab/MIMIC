module fake_jpeg_31300_n_408 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_408);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_408;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx8_ASAP7_75t_SL g42 ( 
.A(n_17),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_19),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_57),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

BUFx4f_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVxp67_ASAP7_75t_SL g105 ( 
.A(n_63),
.Y(n_105)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_22),
.B(n_50),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_79),
.Y(n_98)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_31),
.B(n_10),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_78),
.Y(n_91)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_74),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_36),
.B(n_0),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_38),
.C(n_43),
.Y(n_93)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

HAxp5_ASAP7_75t_SL g78 ( 
.A(n_27),
.B(n_0),
.CON(n_78),
.SN(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_22),
.B(n_10),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_48),
.Y(n_117)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_93),
.B(n_121),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_59),
.A2(n_24),
.B1(n_48),
.B2(n_47),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_95),
.A2(n_102),
.B1(n_104),
.B2(n_111),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_50),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_100),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_78),
.A2(n_38),
.B1(n_49),
.B2(n_46),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_84),
.A2(n_49),
.B1(n_46),
.B2(n_44),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_34),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_107),
.B(n_42),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_23),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_109),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_58),
.A2(n_49),
.B1(n_44),
.B2(n_45),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_66),
.A2(n_34),
.B1(n_33),
.B2(n_43),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_116),
.A2(n_23),
.B1(n_41),
.B2(n_47),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_73),
.B(n_33),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_67),
.A2(n_48),
.B1(n_47),
.B2(n_24),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_117),
.B1(n_95),
.B2(n_87),
.Y(n_146)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_131),
.Y(n_187)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_123),
.A2(n_55),
.B1(n_60),
.B2(n_62),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_135),
.A2(n_141),
.B1(n_146),
.B2(n_147),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

INVx11_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_99),
.A2(n_80),
.B1(n_42),
.B2(n_86),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_127),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_149),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_140),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_87),
.A2(n_24),
.B1(n_26),
.B2(n_28),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_142),
.Y(n_183)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_143),
.Y(n_167)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

INVxp67_ASAP7_75t_SL g149 ( 
.A(n_96),
.Y(n_149)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_97),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_153),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_99),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_115),
.A2(n_26),
.B1(n_28),
.B2(n_61),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_155),
.Y(n_178)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_90),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_157),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_92),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_106),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_161),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_115),
.A2(n_26),
.B1(n_28),
.B2(n_63),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_160),
.B(n_72),
.Y(n_174)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_91),
.A2(n_63),
.B(n_25),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g181 ( 
.A1(n_162),
.A2(n_163),
.B(n_164),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_118),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_91),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_172),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_119),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_174),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_98),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_180),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_148),
.B(n_122),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_132),
.B(n_128),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_163),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_102),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_148),
.C(n_147),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_173),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_198),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_168),
.A2(n_132),
.B1(n_145),
.B2(n_146),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_191),
.A2(n_195),
.B1(n_206),
.B2(n_182),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_194),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_185),
.A2(n_104),
.B1(n_111),
.B2(n_130),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_171),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_182),
.A2(n_164),
.B1(n_129),
.B2(n_89),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_200),
.A2(n_139),
.B(n_157),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_173),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_201),
.Y(n_225)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_172),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_207),
.Y(n_216)
);

OA21x2_ASAP7_75t_L g204 ( 
.A1(n_178),
.A2(n_159),
.B(n_153),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_204),
.A2(n_186),
.B(n_184),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_202),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_174),
.A2(n_128),
.B1(n_156),
.B2(n_155),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_209),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_175),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_189),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_226),
.C(n_208),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_202),
.B(n_189),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_211),
.B(n_223),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_192),
.A2(n_167),
.B1(n_188),
.B2(n_181),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_212),
.A2(n_219),
.B1(n_203),
.B2(n_191),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_195),
.A2(n_188),
.B1(n_180),
.B2(n_178),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_214),
.A2(n_221),
.B1(n_229),
.B2(n_207),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_208),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_217),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_218),
.A2(n_216),
.B(n_222),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_205),
.A2(n_165),
.B1(n_177),
.B2(n_167),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_192),
.A2(n_150),
.B1(n_179),
.B2(n_134),
.Y(n_221)
);

A2O1A1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_197),
.A2(n_158),
.B(n_134),
.C(n_173),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_205),
.A2(n_157),
.B(n_183),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_224),
.B(n_206),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_197),
.Y(n_228)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_228),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_231),
.B(n_249),
.Y(n_273)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_213),
.Y(n_233)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_213),
.Y(n_234)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_234),
.Y(n_268)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_227),
.Y(n_235)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_235),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_242),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_238),
.A2(n_212),
.B1(n_219),
.B2(n_206),
.Y(n_266)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_227),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_244),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_240),
.A2(n_237),
.B(n_234),
.Y(n_262)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_196),
.C(n_198),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_224),
.Y(n_256)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_246),
.Y(n_261)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_216),
.Y(n_247)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_247),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_214),
.A2(n_204),
.B1(n_198),
.B2(n_196),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_248),
.A2(n_254),
.B1(n_204),
.B2(n_225),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_170),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_222),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_250),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_218),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_251),
.A2(n_223),
.B(n_215),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_220),
.B(n_204),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_252),
.B(n_253),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_170),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_228),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_256),
.B(n_278),
.C(n_235),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_251),
.A2(n_231),
.B1(n_229),
.B2(n_254),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_259),
.A2(n_265),
.B1(n_269),
.B2(n_140),
.Y(n_304)
);

NAND2x1p5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_218),
.Y(n_260)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_262),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_232),
.A2(n_229),
.B1(n_221),
.B2(n_211),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_266),
.A2(n_272),
.B1(n_190),
.B2(n_176),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_243),
.A2(n_226),
.B1(n_210),
.B2(n_225),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_267),
.A2(n_247),
.B1(n_233),
.B2(n_232),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_270),
.A2(n_246),
.B(n_244),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_243),
.A2(n_223),
.B(n_210),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_271),
.A2(n_113),
.B(n_137),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_250),
.A2(n_204),
.B1(n_200),
.B2(n_201),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_236),
.B(n_183),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_277),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_245),
.B(n_144),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_240),
.B(n_190),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_258),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_279),
.A2(n_295),
.B1(n_299),
.B2(n_302),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_282),
.B(n_288),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_257),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_283),
.A2(n_286),
.B(n_287),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_241),
.Y(n_284)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_284),
.Y(n_307)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_276),
.Y(n_285)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_285),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_270),
.A2(n_241),
.B(n_239),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_170),
.Y(n_289)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_289),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_290),
.A2(n_297),
.B1(n_265),
.B2(n_260),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_261),
.Y(n_291)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_291),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_255),
.B(n_176),
.Y(n_292)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_292),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_271),
.A2(n_166),
.B(n_179),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_293),
.B(n_298),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_268),
.B(n_176),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_294),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_262),
.B(n_16),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_261),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_263),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_273),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_278),
.C(n_259),
.Y(n_305)
);

NAND3xp33_ASAP7_75t_L g301 ( 
.A(n_274),
.B(n_131),
.C(n_11),
.Y(n_301)
);

AOI21xp33_ASAP7_75t_L g326 ( 
.A1(n_301),
.A2(n_16),
.B(n_20),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_274),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_260),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_303),
.A2(n_281),
.B1(n_287),
.B2(n_296),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_304),
.A2(n_166),
.B1(n_140),
.B2(n_136),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_305),
.B(n_284),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_263),
.C(n_256),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_306),
.B(n_308),
.C(n_313),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_277),
.C(n_266),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_310),
.B(n_314),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_311),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_312),
.A2(n_320),
.B1(n_283),
.B2(n_286),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_280),
.B(n_110),
.C(n_114),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_280),
.B(n_187),
.C(n_136),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_296),
.A2(n_166),
.B1(n_187),
.B2(n_120),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_315),
.B(n_323),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_304),
.A2(n_187),
.B1(n_126),
.B2(n_101),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_303),
.A2(n_101),
.B1(n_124),
.B2(n_83),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_326),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_281),
.A2(n_71),
.B1(n_77),
.B2(n_56),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_327),
.B(n_118),
.Y(n_341)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_307),
.Y(n_328)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_328),
.Y(n_347)
);

FAx1_ASAP7_75t_SL g329 ( 
.A(n_322),
.B(n_282),
.CI(n_293),
.CON(n_329),
.SN(n_329)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_329),
.B(n_334),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_330),
.A2(n_338),
.B1(n_344),
.B2(n_327),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_331),
.B(n_343),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_316),
.A2(n_297),
.B(n_291),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_333),
.B(n_345),
.Y(n_348)
);

FAx1_ASAP7_75t_SL g334 ( 
.A(n_322),
.B(n_300),
.CI(n_294),
.CON(n_334),
.SN(n_334)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_309),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_336),
.B(n_337),
.Y(n_350)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_317),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_318),
.A2(n_285),
.B1(n_292),
.B2(n_15),
.Y(n_338)
);

XNOR2x1_ASAP7_75t_L g351 ( 
.A(n_341),
.B(n_305),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_324),
.B(n_105),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_312),
.A2(n_12),
.B1(n_20),
.B2(n_19),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_308),
.B(n_105),
.Y(n_345)
);

XOR2x1_ASAP7_75t_L g349 ( 
.A(n_335),
.B(n_311),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_349),
.B(n_351),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_340),
.B(n_315),
.Y(n_352)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_352),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_335),
.A2(n_325),
.B1(n_323),
.B2(n_321),
.Y(n_354)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_354),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_332),
.A2(n_319),
.B(n_306),
.Y(n_355)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_355),
.Y(n_362)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_356),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_332),
.B(n_313),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_339),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_331),
.Y(n_358)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_358),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_330),
.A2(n_320),
.B1(n_314),
.B2(n_324),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_359),
.B(n_329),
.C(n_334),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_358),
.B(n_342),
.C(n_345),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_363),
.B(n_370),
.C(n_69),
.Y(n_383)
);

FAx1_ASAP7_75t_SL g364 ( 
.A(n_353),
.B(n_346),
.CI(n_348),
.CON(n_364),
.SN(n_364)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_364),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_365),
.B(n_368),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_351),
.B(n_343),
.C(n_339),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_369),
.B(n_350),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_346),
.B(n_341),
.C(n_76),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_364),
.B(n_362),
.Y(n_374)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_374),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_375),
.B(n_376),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_363),
.B(n_347),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_371),
.B(n_349),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_377),
.B(n_378),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_360),
.B(n_11),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_367),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_379),
.B(n_383),
.Y(n_389)
);

AOI21x1_ASAP7_75t_L g380 ( 
.A1(n_366),
.A2(n_11),
.B(n_19),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_380),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_366),
.B(n_9),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_381),
.B(n_8),
.Y(n_388)
);

NOR3xp33_ASAP7_75t_SL g382 ( 
.A(n_361),
.B(n_9),
.C(n_13),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_SL g391 ( 
.A(n_382),
.B(n_8),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_388),
.B(n_390),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_372),
.B(n_370),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_391),
.B(n_392),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_373),
.B(n_6),
.Y(n_392)
);

O2A1O1Ixp33_ASAP7_75t_SL g393 ( 
.A1(n_385),
.A2(n_382),
.B(n_381),
.C(n_383),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_393),
.A2(n_394),
.B(n_398),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_387),
.A2(n_389),
.B(n_386),
.Y(n_394)
);

OAI211xp5_ASAP7_75t_L g396 ( 
.A1(n_384),
.A2(n_6),
.B(n_12),
.C(n_17),
.Y(n_396)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_396),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_387),
.A2(n_5),
.B(n_17),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_395),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_400),
.B(n_397),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_402),
.B(n_403),
.C(n_52),
.Y(n_404)
);

AO221x1_ASAP7_75t_L g403 ( 
.A1(n_399),
.A2(n_401),
.B1(n_5),
.B2(n_9),
.C(n_3),
.Y(n_403)
);

AOI321xp33_ASAP7_75t_SL g405 ( 
.A1(n_404),
.A2(n_25),
.A3(n_4),
.B1(n_3),
.B2(n_5),
.C(n_16),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_405),
.A2(n_0),
.B(n_1),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_406),
.B(n_0),
.C(n_1),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_407),
.A2(n_2),
.B(n_394),
.Y(n_408)
);


endmodule