module fake_jpeg_1285_n_653 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_653);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_653;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_58),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_24),
.B(n_8),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_59),
.B(n_62),
.Y(n_133)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_61),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_63),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_64),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_24),
.B(n_8),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_65),
.B(n_77),
.Y(n_137)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_66),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_67),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_68),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_28),
.B(n_0),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_69),
.B(n_74),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_70),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_37),
.Y(n_71)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_71),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_72),
.Y(n_196)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_73),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_0),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_75),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_39),
.B(n_1),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_76),
.B(n_123),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_32),
.B(n_10),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_78),
.Y(n_165)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_79),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_80),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_81),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_22),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_82),
.B(n_84),
.Y(n_140)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_83),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_38),
.B(n_10),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_85),
.Y(n_223)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_86),
.Y(n_199)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_88),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_22),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_89),
.B(n_91),
.Y(n_152)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_90),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_25),
.Y(n_91)
);

INVx4_ASAP7_75t_SL g92 ( 
.A(n_53),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_92),
.B(n_45),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_93),
.Y(n_216)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_94),
.Y(n_183)
);

BUFx4f_ASAP7_75t_SL g95 ( 
.A(n_39),
.Y(n_95)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_95),
.Y(n_225)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_96),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_97),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_48),
.B(n_1),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_98),
.B(n_2),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_99),
.Y(n_160)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_100),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_47),
.B(n_10),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_101),
.B(n_106),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_102),
.Y(n_180)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_103),
.Y(n_192)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_104),
.Y(n_209)
);

BUFx12_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

BUFx2_ASAP7_75t_R g153 ( 
.A(n_105),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_41),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_25),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_107),
.B(n_109),
.Y(n_162)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_108),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_25),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_41),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_110),
.B(n_113),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_111),
.Y(n_174)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_112),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_57),
.Y(n_113)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_114),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_48),
.Y(n_115)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_115),
.Y(n_215)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_116),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_34),
.Y(n_117)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_117),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_34),
.Y(n_118)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_118),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_35),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_119),
.B(n_125),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_34),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_120),
.Y(n_186)
);

CKINVDCx9p33_ASAP7_75t_R g121 ( 
.A(n_35),
.Y(n_121)
);

INVx11_ASAP7_75t_L g207 ( 
.A(n_121),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_46),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_122),
.Y(n_213)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_36),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_54),
.Y(n_124)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_41),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_54),
.B(n_11),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_126),
.B(n_12),
.Y(n_175)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_43),
.Y(n_128)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_128),
.Y(n_226)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_43),
.Y(n_129)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_46),
.Y(n_130)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_130),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_74),
.A2(n_56),
.B1(n_52),
.B2(n_42),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_132),
.A2(n_212),
.B1(n_117),
.B2(n_120),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_76),
.A2(n_41),
.B(n_56),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_136),
.A2(n_180),
.B(n_217),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_69),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_139),
.B(n_175),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_121),
.A2(n_46),
.B1(n_53),
.B2(n_43),
.Y(n_142)
);

OAI21xp33_ASAP7_75t_SL g308 ( 
.A1(n_142),
.A2(n_150),
.B(n_155),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_144),
.B(n_122),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_92),
.A2(n_53),
.B1(n_43),
.B2(n_55),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_98),
.B(n_21),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_154),
.B(n_177),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_96),
.A2(n_42),
.B1(n_52),
.B2(n_40),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_76),
.A2(n_40),
.B1(n_21),
.B2(n_44),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_158),
.A2(n_172),
.B1(n_189),
.B2(n_136),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_114),
.A2(n_99),
.B1(n_81),
.B2(n_72),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_166),
.A2(n_194),
.B1(n_201),
.B2(n_218),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_61),
.A2(n_53),
.B1(n_43),
.B2(n_44),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_170),
.A2(n_171),
.B1(n_173),
.B2(n_208),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_90),
.A2(n_33),
.B1(n_29),
.B2(n_49),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_115),
.A2(n_49),
.B1(n_27),
.B2(n_29),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_112),
.A2(n_33),
.B1(n_20),
.B2(n_45),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_60),
.B(n_2),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_178),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_108),
.B(n_2),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_179),
.B(n_187),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_127),
.B(n_11),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_184),
.B(n_188),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_73),
.B(n_2),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_71),
.B(n_11),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_58),
.A2(n_20),
.B1(n_13),
.B2(n_14),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_68),
.B(n_13),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_190),
.B(n_197),
.Y(n_238)
);

OA22x2_ASAP7_75t_L g191 ( 
.A1(n_104),
.A2(n_20),
.B1(n_4),
.B2(n_5),
.Y(n_191)
);

O2A1O1Ixp33_ASAP7_75t_SL g264 ( 
.A1(n_191),
.A2(n_105),
.B(n_78),
.C(n_100),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_63),
.A2(n_20),
.B1(n_13),
.B2(n_14),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_68),
.B(n_18),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_64),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_102),
.B(n_95),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_203),
.B(n_204),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_128),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_102),
.B(n_17),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_206),
.B(n_211),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_94),
.A2(n_116),
.B1(n_88),
.B2(n_86),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_95),
.B(n_17),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_70),
.A2(n_7),
.B1(n_13),
.B2(n_5),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_79),
.Y(n_214)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_214),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_85),
.A2(n_7),
.B1(n_4),
.B2(n_5),
.Y(n_218)
);

A2O1A1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_83),
.A2(n_7),
.B(n_4),
.C(n_6),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_219),
.B(n_3),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_93),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_221),
.A2(n_224),
.B1(n_207),
.B2(n_192),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_111),
.A2(n_3),
.B1(n_6),
.B2(n_130),
.Y(n_224)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_228),
.Y(n_229)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_229),
.Y(n_317)
);

BUFx12f_ASAP7_75t_L g230 ( 
.A(n_151),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_230),
.Y(n_313)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_228),
.Y(n_231)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_231),
.Y(n_324)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_141),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_233),
.B(n_248),
.Y(n_321)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_234),
.Y(n_330)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_205),
.Y(n_235)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_235),
.Y(n_328)
);

INVx13_ASAP7_75t_L g236 ( 
.A(n_153),
.Y(n_236)
);

BUFx2_ASAP7_75t_SL g327 ( 
.A(n_236),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_240),
.B(n_263),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_241),
.A2(n_312),
.B(n_255),
.Y(n_369)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_243),
.Y(n_329)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_148),
.Y(n_244)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_244),
.Y(n_339)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_149),
.Y(n_245)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_245),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_135),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_246),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_247),
.B(n_250),
.Y(n_315)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_143),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_L g249 ( 
.A1(n_172),
.A2(n_129),
.B1(n_97),
.B2(n_118),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_249),
.A2(n_264),
.B1(n_272),
.B2(n_274),
.Y(n_323)
);

OAI32xp33_ASAP7_75t_L g250 ( 
.A1(n_138),
.A2(n_105),
.A3(n_103),
.B1(n_123),
.B2(n_75),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_149),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_251),
.Y(n_319)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_220),
.Y(n_252)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_252),
.Y(n_331)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_147),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_253),
.B(n_265),
.Y(n_325)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_182),
.Y(n_256)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_256),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_225),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_257),
.Y(n_322)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_148),
.Y(n_258)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_258),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_259),
.A2(n_267),
.B1(n_292),
.B2(n_293),
.Y(n_326)
);

INVx11_ASAP7_75t_L g261 ( 
.A(n_207),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_261),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_138),
.B(n_3),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_162),
.Y(n_265)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_165),
.Y(n_266)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_266),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_131),
.A2(n_225),
.B1(n_156),
.B2(n_192),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_152),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_268),
.B(n_269),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_178),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_164),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_270),
.B(n_279),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_167),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_271),
.B(n_275),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_133),
.B(n_3),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_273),
.Y(n_344)
);

OAI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_158),
.A2(n_67),
.B1(n_80),
.B2(n_6),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_179),
.Y(n_275)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_165),
.Y(n_276)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_276),
.Y(n_346)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_135),
.Y(n_277)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_277),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_145),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_278),
.Y(n_349)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_227),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_131),
.B(n_177),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_280),
.B(n_285),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_154),
.B(n_6),
.C(n_144),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_281),
.B(n_294),
.C(n_311),
.Y(n_358)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_182),
.Y(n_282)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_282),
.Y(n_350)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_185),
.Y(n_283)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_283),
.Y(n_352)
);

INVx6_ASAP7_75t_L g284 ( 
.A(n_145),
.Y(n_284)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_284),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_131),
.B(n_187),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_209),
.Y(n_286)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_286),
.Y(n_362)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_169),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_287),
.B(n_290),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_146),
.Y(n_288)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_288),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_186),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_185),
.Y(n_291)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_291),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_159),
.A2(n_137),
.B1(n_198),
.B2(n_140),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_198),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_134),
.B(n_161),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_161),
.A2(n_193),
.B1(n_195),
.B2(n_222),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_295),
.A2(n_301),
.B1(n_303),
.B2(n_309),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_153),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_296),
.B(n_297),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_134),
.B(n_183),
.Y(n_297)
);

INVx5_ASAP7_75t_SL g298 ( 
.A(n_146),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_298),
.B(n_305),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_219),
.B(n_191),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_300),
.B(n_302),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_195),
.A2(n_168),
.B1(n_222),
.B2(n_183),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_191),
.B(n_200),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_168),
.A2(n_216),
.B1(n_213),
.B2(n_199),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_157),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_304),
.Y(n_336)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_200),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_191),
.B(n_209),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_306),
.B(n_223),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_226),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_307),
.Y(n_342)
);

O2A1O1Ixp33_ASAP7_75t_SL g309 ( 
.A1(n_189),
.A2(n_216),
.B(n_163),
.C(n_217),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_163),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_310),
.A2(n_151),
.B1(n_176),
.B2(n_296),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_202),
.B(n_180),
.C(n_199),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_306),
.A2(n_174),
.B1(n_160),
.B2(n_215),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_314),
.A2(n_333),
.B1(n_249),
.B2(n_293),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_239),
.B(n_280),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_318),
.B(n_359),
.C(n_358),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_302),
.A2(n_174),
.B1(n_160),
.B2(n_215),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_272),
.A2(n_196),
.B1(n_157),
.B2(n_210),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_337),
.A2(n_354),
.B1(n_360),
.B2(n_336),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_340),
.B(n_284),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_242),
.B(n_202),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_343),
.B(n_348),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_242),
.B(n_181),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_300),
.A2(n_181),
.B1(n_196),
.B2(n_210),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_239),
.B(n_223),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_357),
.B(n_366),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_280),
.B(n_176),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_363),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_264),
.A2(n_254),
.B1(n_260),
.B2(n_231),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_364),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_240),
.B(n_263),
.Y(n_366)
);

OAI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_299),
.A2(n_312),
.B1(n_250),
.B2(n_289),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_367),
.A2(n_294),
.B1(n_298),
.B2(n_236),
.Y(n_388)
);

AO21x1_ASAP7_75t_L g416 ( 
.A1(n_369),
.A2(n_261),
.B(n_230),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_344),
.B(n_237),
.Y(n_373)
);

CKINVDCx14_ASAP7_75t_R g428 ( 
.A(n_373),
.Y(n_428)
);

INVx5_ASAP7_75t_L g374 ( 
.A(n_313),
.Y(n_374)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_374),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_325),
.B(n_338),
.Y(n_376)
);

CKINVDCx14_ASAP7_75t_R g433 ( 
.A(n_376),
.Y(n_433)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_377),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_315),
.A2(n_308),
.B1(n_285),
.B2(n_238),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_378),
.A2(n_380),
.B1(n_383),
.B2(n_402),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_318),
.B(n_285),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_379),
.B(n_396),
.C(n_332),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_315),
.A2(n_229),
.B1(n_309),
.B2(n_281),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_325),
.B(n_262),
.Y(n_381)
);

CKINVDCx14_ASAP7_75t_R g447 ( 
.A(n_381),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_338),
.B(n_251),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_382),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_315),
.A2(n_294),
.B1(n_311),
.B2(n_234),
.Y(n_383)
);

BUFx5_ASAP7_75t_L g385 ( 
.A(n_327),
.Y(n_385)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_385),
.Y(n_457)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_317),
.Y(n_386)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_386),
.Y(n_431)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_317),
.Y(n_387)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_387),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_388),
.A2(n_416),
.B(n_346),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_359),
.B(n_293),
.Y(n_390)
);

CKINVDCx14_ASAP7_75t_R g430 ( 
.A(n_390),
.Y(n_430)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_324),
.Y(n_391)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_391),
.Y(n_440)
);

FAx1_ASAP7_75t_SL g392 ( 
.A(n_320),
.B(n_232),
.CI(n_286),
.CON(n_392),
.SN(n_392)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_392),
.B(n_398),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_340),
.B(n_252),
.Y(n_393)
);

AND2x2_ASAP7_75t_SL g444 ( 
.A(n_393),
.B(n_394),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_320),
.B(n_243),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_395),
.B(n_405),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_335),
.B(n_305),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_369),
.A2(n_310),
.B(n_257),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_397),
.A2(n_360),
.B(n_334),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_366),
.B(n_282),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_368),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_400),
.B(n_401),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_321),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_323),
.A2(n_235),
.B1(n_291),
.B2(n_283),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_365),
.B(n_245),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_403),
.B(n_322),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_321),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_404),
.B(n_406),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_335),
.B(n_256),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_345),
.B(n_288),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_323),
.A2(n_304),
.B1(n_278),
.B2(n_246),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_407),
.A2(n_408),
.B1(n_417),
.B2(n_419),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_337),
.A2(n_244),
.B1(n_258),
.B2(n_266),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_348),
.B(n_276),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_409),
.B(n_410),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_343),
.B(n_277),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_324),
.Y(n_411)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_411),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_316),
.Y(n_412)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_412),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_413),
.B(n_372),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_357),
.B(n_230),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_414),
.B(n_415),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_355),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_314),
.A2(n_333),
.B1(n_354),
.B2(n_358),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_418),
.A2(n_362),
.B1(n_336),
.B2(n_342),
.Y(n_425)
);

AOI22x1_ASAP7_75t_L g419 ( 
.A1(n_372),
.A2(n_326),
.B1(n_351),
.B2(n_361),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_372),
.A2(n_361),
.B1(n_355),
.B2(n_368),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_420),
.A2(n_342),
.B1(n_362),
.B2(n_334),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_SL g424 ( 
.A1(n_384),
.A2(n_389),
.B1(n_418),
.B2(n_400),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_424),
.A2(n_449),
.B1(n_450),
.B2(n_456),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_425),
.A2(n_441),
.B1(n_446),
.B2(n_386),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_426),
.B(n_460),
.C(n_405),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_413),
.B(n_345),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g464 ( 
.A(n_429),
.B(n_443),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_434),
.B(n_404),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_437),
.A2(n_452),
.B(n_416),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_379),
.B(n_371),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_380),
.A2(n_356),
.B1(n_347),
.B2(n_341),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_383),
.A2(n_356),
.B1(n_347),
.B2(n_341),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_407),
.A2(n_417),
.B1(n_402),
.B2(n_378),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_375),
.B(n_332),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_451),
.B(n_458),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_403),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_455),
.B(n_401),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_394),
.A2(n_346),
.B1(n_349),
.B2(n_339),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_375),
.B(n_371),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_459),
.B(n_420),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_396),
.B(n_352),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_462),
.B(n_465),
.Y(n_509)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_431),
.Y(n_463)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_463),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_436),
.B(n_415),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_L g517 ( 
.A1(n_466),
.A2(n_477),
.B1(n_480),
.B2(n_482),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_467),
.B(n_489),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_432),
.B(n_399),
.Y(n_468)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_468),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_432),
.B(n_399),
.Y(n_469)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_469),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_451),
.B(n_409),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_470),
.B(n_471),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_458),
.B(n_410),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_455),
.B(n_394),
.Y(n_473)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_473),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_474),
.B(n_444),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_436),
.B(n_414),
.Y(n_475)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_475),
.Y(n_524)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_431),
.Y(n_476)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_476),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_428),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_438),
.Y(n_478)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_478),
.Y(n_528)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_438),
.Y(n_479)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_479),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_445),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_439),
.A2(n_397),
.B1(n_389),
.B2(n_419),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_481),
.A2(n_490),
.B1(n_498),
.B2(n_430),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_442),
.B(n_387),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_426),
.B(n_460),
.C(n_459),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_483),
.B(n_487),
.C(n_493),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_421),
.A2(n_419),
.B1(n_388),
.B2(n_377),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_484),
.A2(n_485),
.B1(n_430),
.B2(n_435),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_421),
.A2(n_395),
.B1(n_390),
.B2(n_393),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_447),
.B(n_411),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_486),
.B(n_488),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_445),
.B(n_398),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_427),
.B(n_392),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_439),
.A2(n_390),
.B1(n_392),
.B2(n_393),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_491),
.A2(n_497),
.B(n_452),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_453),
.B(n_391),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_492),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_429),
.B(n_370),
.C(n_352),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_440),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_494),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_427),
.B(n_416),
.Y(n_495)
);

CKINVDCx16_ASAP7_75t_R g505 ( 
.A(n_495),
.Y(n_505)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_440),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_496),
.A2(n_448),
.B1(n_434),
.B2(n_422),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_433),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_435),
.A2(n_384),
.B1(n_408),
.B2(n_374),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_483),
.B(n_443),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_499),
.B(n_502),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_500),
.A2(n_485),
.B1(n_466),
.B2(n_465),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_483),
.B(n_423),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_503),
.A2(n_508),
.B1(n_518),
.B2(n_522),
.Y(n_536)
);

XNOR2x1_ASAP7_75t_L g504 ( 
.A(n_474),
.B(n_423),
.Y(n_504)
);

XNOR2x1_ASAP7_75t_L g553 ( 
.A(n_504),
.B(n_525),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_L g548 ( 
.A1(n_506),
.A2(n_526),
.B(n_462),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_472),
.A2(n_450),
.B1(n_446),
.B2(n_441),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_512),
.B(n_515),
.C(n_519),
.Y(n_535)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_513),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_487),
.B(n_444),
.C(n_449),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_472),
.A2(n_437),
.B1(n_425),
.B2(n_453),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_464),
.B(n_444),
.C(n_448),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_484),
.A2(n_444),
.B1(n_456),
.B2(n_422),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_464),
.B(n_493),
.C(n_480),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_523),
.B(n_533),
.C(n_479),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_SL g525 ( 
.A(n_464),
.B(n_350),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_491),
.A2(n_495),
.B(n_481),
.Y(n_526)
);

OA21x2_ASAP7_75t_L g531 ( 
.A1(n_491),
.A2(n_454),
.B(n_457),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_531),
.B(n_494),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_468),
.B(n_370),
.C(n_339),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_510),
.B(n_477),
.Y(n_534)
);

CKINVDCx16_ASAP7_75t_R g585 ( 
.A(n_534),
.Y(n_585)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_517),
.Y(n_537)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_537),
.Y(n_569)
);

CKINVDCx16_ASAP7_75t_R g538 ( 
.A(n_513),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_538),
.B(n_543),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_539),
.B(n_559),
.Y(n_577)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_511),
.Y(n_540)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_540),
.Y(n_580)
);

FAx1_ASAP7_75t_L g541 ( 
.A(n_526),
.B(n_490),
.CI(n_467),
.CON(n_541),
.SN(n_541)
);

OAI21xp5_ASAP7_75t_SL g574 ( 
.A1(n_541),
.A2(n_544),
.B(n_548),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_508),
.A2(n_469),
.B1(n_489),
.B2(n_461),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_542),
.A2(n_546),
.B1(n_547),
.B2(n_551),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_510),
.B(n_497),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_507),
.B(n_475),
.C(n_473),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_545),
.B(n_557),
.C(n_512),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_500),
.A2(n_470),
.B1(n_461),
.B2(n_498),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_503),
.A2(n_471),
.B1(n_488),
.B2(n_482),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_514),
.A2(n_492),
.B1(n_486),
.B2(n_478),
.Y(n_551)
);

CKINVDCx16_ASAP7_75t_R g552 ( 
.A(n_509),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_552),
.A2(n_556),
.B1(n_561),
.B2(n_530),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_554),
.B(n_531),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_514),
.A2(n_496),
.B1(n_476),
.B2(n_463),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_555),
.A2(n_521),
.B1(n_454),
.B2(n_412),
.Y(n_584)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_527),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_507),
.B(n_499),
.C(n_515),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_524),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_558),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_502),
.B(n_350),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_529),
.B(n_457),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_560),
.Y(n_563)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_528),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_533),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_562),
.B(n_523),
.Y(n_567)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_548),
.A2(n_506),
.B(n_518),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_565),
.A2(n_549),
.B(n_554),
.Y(n_587)
);

OAI21x1_ASAP7_75t_L g602 ( 
.A1(n_567),
.A2(n_331),
.B(n_328),
.Y(n_602)
);

A2O1A1O1Ixp25_ASAP7_75t_L g568 ( 
.A1(n_541),
.A2(n_519),
.B(n_514),
.C(n_516),
.D(n_501),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_L g596 ( 
.A1(n_568),
.A2(n_559),
.B(n_558),
.Y(n_596)
);

OA22x2_ASAP7_75t_L g570 ( 
.A1(n_541),
.A2(n_522),
.B1(n_531),
.B2(n_501),
.Y(n_570)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_570),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_571),
.B(n_573),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_572),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_550),
.B(n_504),
.C(n_525),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_550),
.B(n_532),
.C(n_505),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_575),
.B(n_583),
.C(n_539),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_555),
.B(n_532),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_576),
.B(n_579),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_535),
.B(n_520),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_SL g594 ( 
.A(n_578),
.B(n_535),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_542),
.B(n_520),
.Y(n_579)
);

INVxp33_ASAP7_75t_SL g590 ( 
.A(n_581),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_557),
.B(n_521),
.C(n_313),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_SL g597 ( 
.A1(n_584),
.A2(n_561),
.B1(n_412),
.B2(n_316),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_SL g614 ( 
.A1(n_587),
.A2(n_591),
.B(n_592),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_SL g588 ( 
.A1(n_564),
.A2(n_536),
.B1(n_549),
.B2(n_547),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_SL g617 ( 
.A1(n_588),
.A2(n_572),
.B1(n_566),
.B2(n_570),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_589),
.B(n_595),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_574),
.A2(n_536),
.B(n_551),
.Y(n_591)
);

AOI21xp5_ASAP7_75t_L g592 ( 
.A1(n_574),
.A2(n_546),
.B(n_544),
.Y(n_592)
);

XOR2xp5_ASAP7_75t_L g610 ( 
.A(n_594),
.B(n_573),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_585),
.B(n_545),
.Y(n_595)
);

AOI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_596),
.A2(n_598),
.B(n_572),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g618 ( 
.A(n_597),
.Y(n_618)
);

OAI21xp5_ASAP7_75t_L g598 ( 
.A1(n_565),
.A2(n_553),
.B(n_313),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_583),
.B(n_316),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_599),
.B(n_601),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_571),
.B(n_553),
.C(n_328),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_602),
.B(n_580),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_578),
.B(n_329),
.C(n_331),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_603),
.B(n_600),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_L g605 ( 
.A1(n_590),
.A2(n_566),
.B1(n_569),
.B2(n_579),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_605),
.A2(n_617),
.B1(n_592),
.B2(n_604),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_606),
.B(n_607),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_589),
.B(n_567),
.Y(n_607)
);

XOR2xp5_ASAP7_75t_L g631 ( 
.A(n_608),
.B(n_610),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_609),
.B(n_616),
.Y(n_627)
);

XOR2xp5_ASAP7_75t_L g612 ( 
.A(n_596),
.B(n_575),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_612),
.B(n_613),
.C(n_604),
.Y(n_629)
);

XOR2xp5_ASAP7_75t_L g613 ( 
.A(n_591),
.B(n_577),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_594),
.B(n_577),
.C(n_576),
.Y(n_616)
);

CKINVDCx16_ASAP7_75t_R g619 ( 
.A(n_586),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_619),
.B(n_620),
.Y(n_622)
);

OAI21xp5_ASAP7_75t_SL g620 ( 
.A1(n_587),
.A2(n_568),
.B(n_570),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_611),
.B(n_603),
.C(n_601),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_621),
.B(n_623),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_615),
.B(n_563),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g634 ( 
.A(n_625),
.B(n_629),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_616),
.B(n_563),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_626),
.B(n_628),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_612),
.B(n_588),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_613),
.B(n_593),
.C(n_586),
.Y(n_630)
);

OAI21xp5_ASAP7_75t_L g636 ( 
.A1(n_630),
.A2(n_632),
.B(n_620),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_614),
.B(n_582),
.Y(n_632)
);

OAI21x1_ASAP7_75t_SL g635 ( 
.A1(n_622),
.A2(n_609),
.B(n_608),
.Y(n_635)
);

AO21x1_ASAP7_75t_L g645 ( 
.A1(n_635),
.A2(n_584),
.B(n_582),
.Y(n_645)
);

AOI31xp33_ASAP7_75t_L g641 ( 
.A1(n_636),
.A2(n_621),
.A3(n_630),
.B(n_631),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_SL g637 ( 
.A1(n_624),
.A2(n_614),
.B(n_593),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_SL g642 ( 
.A1(n_637),
.A2(n_638),
.B(n_618),
.Y(n_642)
);

OAI21xp5_ASAP7_75t_SL g638 ( 
.A1(n_627),
.A2(n_618),
.B(n_598),
.Y(n_638)
);

XOR2xp5_ASAP7_75t_L g639 ( 
.A(n_631),
.B(n_617),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_639),
.B(n_570),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_L g648 ( 
.A1(n_641),
.A2(n_642),
.B(n_643),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_640),
.B(n_610),
.C(n_597),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_SL g646 ( 
.A1(n_644),
.A2(n_645),
.B(n_633),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g649 ( 
.A(n_646),
.B(n_634),
.C(n_353),
.Y(n_649)
);

OAI311xp33_ASAP7_75t_L g647 ( 
.A1(n_644),
.A2(n_639),
.A3(n_634),
.B1(n_385),
.C1(n_322),
.Y(n_647)
);

AOI221xp5_ASAP7_75t_L g650 ( 
.A1(n_647),
.A2(n_319),
.B1(n_329),
.B2(n_330),
.C(n_353),
.Y(n_650)
);

INVxp33_ASAP7_75t_L g651 ( 
.A(n_649),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_651),
.B(n_648),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_652),
.B(n_650),
.Y(n_653)
);


endmodule