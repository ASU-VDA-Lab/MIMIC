module fake_jpeg_8299_n_269 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_269);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_269;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx5_ASAP7_75t_SL g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_17),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_25),
.C(n_24),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_26),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_42),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_22),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_41),
.B(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_46),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_50),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_41),
.B(n_33),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_17),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_20),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_54),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_19),
.B1(n_28),
.B2(n_31),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_23),
.B1(n_31),
.B2(n_32),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_27),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_64),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_18),
.C(n_29),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_37),
.A2(n_28),
.B1(n_19),
.B2(n_23),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_61),
.A2(n_63),
.B1(n_23),
.B2(n_31),
.Y(n_83)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

OAI21xp33_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_20),
.B(n_28),
.Y(n_63)
);

INVx5_ASAP7_75t_SL g64 ( 
.A(n_37),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_65),
.B(n_68),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_52),
.B(n_38),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_78),
.Y(n_97)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_25),
.Y(n_101)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_79),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_83),
.B1(n_32),
.B2(n_30),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_59),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_30),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_80),
.B(n_82),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_18),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_86),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_29),
.Y(n_85)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_55),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_58),
.Y(n_98)
);

OAI32xp33_ASAP7_75t_L g89 ( 
.A1(n_87),
.A2(n_78),
.A3(n_68),
.B1(n_65),
.B2(n_80),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_89),
.B(n_72),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_56),
.B1(n_36),
.B2(n_42),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_90),
.A2(n_79),
.B1(n_64),
.B2(n_47),
.Y(n_131)
);

INVx6_ASAP7_75t_SL g92 ( 
.A(n_66),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_109),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_75),
.B1(n_82),
.B2(n_58),
.Y(n_118)
);

AND2x4_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_88),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_96),
.B(n_106),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_102),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_84),
.A2(n_32),
.B1(n_30),
.B2(n_64),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_101),
.B(n_111),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_55),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_38),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_69),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_34),
.Y(n_106)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_70),
.Y(n_132)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_75),
.A2(n_36),
.B(n_42),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_74),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_114),
.B(n_115),
.Y(n_144)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_116),
.B(n_117),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_107),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_131),
.B1(n_135),
.B2(n_108),
.Y(n_141)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_119),
.B(n_122),
.Y(n_156)
);

NOR3xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_113),
.C(n_96),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_124),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_110),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_128),
.Y(n_155)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_92),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_129),
.A2(n_133),
.B1(n_109),
.B2(n_66),
.Y(n_164)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_74),
.B1(n_36),
.B2(n_42),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_96),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_73),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_137),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_139),
.B(n_34),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_106),
.C(n_97),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_142),
.C(n_165),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_141),
.A2(n_151),
.B1(n_164),
.B2(n_47),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_97),
.C(n_96),
.Y(n_142)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_128),
.B(n_93),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_147),
.B(n_155),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_94),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_149),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_94),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_150),
.B(n_157),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_126),
.A2(n_100),
.B1(n_89),
.B2(n_49),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_101),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_160),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_125),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_158),
.B(n_159),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_100),
.B(n_101),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_162),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_116),
.B(n_38),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_138),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_138),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_130),
.Y(n_166)
);

INVx13_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_158),
.A2(n_121),
.B1(n_130),
.B2(n_114),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_167),
.A2(n_182),
.B1(n_188),
.B2(n_152),
.Y(n_197)
);

NAND5xp2_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_139),
.C(n_118),
.D(n_121),
.E(n_35),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_169),
.B(n_38),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_162),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_181),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_160),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_172),
.A2(n_146),
.B(n_148),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_173),
.B(n_147),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_176),
.A2(n_152),
.B1(n_143),
.B2(n_157),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_62),
.C(n_48),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_184),
.C(n_35),
.Y(n_209)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_166),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_180),
.Y(n_201)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_144),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_151),
.A2(n_47),
.B1(n_70),
.B2(n_43),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_62),
.C(n_48),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_143),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_86),
.Y(n_202)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_187),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_141),
.A2(n_27),
.B1(n_24),
.B2(n_20),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_190),
.B(n_197),
.Y(n_211)
);

A2O1A1Ixp33_ASAP7_75t_SL g223 ( 
.A1(n_191),
.A2(n_189),
.B(n_35),
.C(n_86),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_149),
.Y(n_192)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_156),
.Y(n_193)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_140),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_206),
.C(n_209),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_153),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_179),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_196),
.A2(n_199),
.B1(n_203),
.B2(n_205),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_175),
.A2(n_183),
.B1(n_169),
.B2(n_172),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_167),
.A2(n_154),
.B1(n_142),
.B2(n_16),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_200),
.B(n_202),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_175),
.A2(n_59),
.B1(n_69),
.B2(n_103),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_181),
.B(n_15),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_204),
.B(n_0),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_168),
.A2(n_16),
.B1(n_69),
.B2(n_3),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_38),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_177),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_217),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_198),
.A2(n_184),
.B(n_186),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_216),
.A2(n_192),
.B(n_201),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_186),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_178),
.C(n_187),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_220),
.Y(n_237)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_219),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_178),
.Y(n_220)
);

FAx1_ASAP7_75t_SL g221 ( 
.A(n_193),
.B(n_172),
.CI(n_180),
.CON(n_221),
.SN(n_221)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_221),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_222),
.Y(n_235)
);

A2O1A1Ixp33_ASAP7_75t_SL g229 ( 
.A1(n_223),
.A2(n_207),
.B(n_191),
.C(n_203),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_189),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_208),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_211),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_225),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_229),
.A2(n_223),
.B1(n_210),
.B2(n_224),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_230),
.A2(n_233),
.B(n_226),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_223),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_218),
.A2(n_196),
.B(n_195),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_223),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_213),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_236),
.B(n_214),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_212),
.C(n_227),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_242),
.C(n_243),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_239),
.A2(n_240),
.B1(n_247),
.B2(n_3),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_241),
.A2(n_244),
.B(n_246),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_212),
.C(n_215),
.Y(n_242)
);

INVxp33_ASAP7_75t_L g252 ( 
.A(n_245),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_231),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_230),
.B(n_229),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_243),
.A2(n_229),
.B1(n_35),
.B2(n_4),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_255),
.C(n_8),
.Y(n_259)
);

NOR2x1_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_2),
.Y(n_251)
);

OAI21x1_ASAP7_75t_L g257 ( 
.A1(n_251),
.A2(n_8),
.B(n_9),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_7),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_238),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_254),
.A2(n_8),
.B(n_10),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_247),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_255)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

AOI31xp67_ASAP7_75t_SL g262 ( 
.A1(n_257),
.A2(n_251),
.A3(n_248),
.B(n_252),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_12),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_259),
.B(n_260),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_252),
.B(n_10),
.Y(n_260)
);

AOI322xp5_ASAP7_75t_L g265 ( 
.A1(n_262),
.A2(n_263),
.A3(n_264),
.B1(n_261),
.B2(n_13),
.C1(n_12),
.C2(n_250),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_265),
.B(n_266),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_249),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_267),
.B(n_249),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_13),
.Y(n_269)
);


endmodule