module fake_jpeg_18587_n_253 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_253);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_253;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVxp33_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_34),
.Y(n_56)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_8),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_38),
.Y(n_45)
);

AOI21xp33_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_8),
.B(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_21),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

HAxp5_ASAP7_75t_SL g43 ( 
.A(n_37),
.B(n_32),
.CON(n_43),
.SN(n_43)
);

OR2x4_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_33),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_35),
.A2(n_20),
.B1(n_29),
.B2(n_26),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_49),
.B1(n_59),
.B2(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_53),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_20),
.B1(n_29),
.B2(n_26),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_20),
.B1(n_29),
.B2(n_28),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_17),
.B1(n_18),
.B2(n_27),
.Y(n_75)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_30),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_40),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_60),
.Y(n_70)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_20),
.B1(n_27),
.B2(n_18),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_26),
.Y(n_60)
);

NOR2x1_ASAP7_75t_R g96 ( 
.A(n_62),
.B(n_73),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_65),
.A2(n_49),
.B1(n_48),
.B2(n_52),
.Y(n_89)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_41),
.C(n_42),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_83),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_39),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_74),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_84),
.Y(n_94)
);

FAx1_ASAP7_75t_SL g73 ( 
.A(n_45),
.B(n_39),
.CI(n_41),
.CON(n_73),
.SN(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_75),
.A2(n_79),
.B1(n_17),
.B2(n_18),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_45),
.A2(n_24),
.B(n_33),
.C(n_22),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_78),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_23),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_44),
.A2(n_24),
.B1(n_22),
.B2(n_33),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_36),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_81),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_47),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_22),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_50),
.A2(n_24),
.B1(n_19),
.B2(n_23),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_78),
.B1(n_72),
.B2(n_71),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_59),
.B(n_41),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_41),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_59),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_40),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_98),
.B1(n_100),
.B2(n_106),
.Y(n_113)
);

BUFx8_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVxp67_ASAP7_75t_SL g114 ( 
.A(n_91),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_93),
.B(n_104),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_81),
.A2(n_59),
.B(n_17),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_103),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_19),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_74),
.A2(n_57),
.B1(n_48),
.B2(n_46),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_41),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_68),
.C(n_80),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_23),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_109),
.B(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_42),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_78),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_25),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_87),
.A2(n_57),
.B1(n_52),
.B2(n_51),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_112),
.A2(n_75),
.B1(n_57),
.B2(n_69),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_115),
.A2(n_128),
.B1(n_42),
.B2(n_36),
.Y(n_160)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_96),
.A2(n_73),
.B(n_62),
.C(n_77),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_127),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_SL g119 ( 
.A(n_96),
.B(n_73),
.C(n_79),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_119),
.A2(n_28),
.B(n_25),
.Y(n_152)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_123),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_110),
.Y(n_122)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_86),
.C(n_41),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_89),
.A2(n_69),
.B1(n_76),
.B2(n_63),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_41),
.C(n_36),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_131),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_105),
.A2(n_64),
.B1(n_52),
.B2(n_63),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_130),
.A2(n_58),
.B1(n_91),
.B2(n_61),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_67),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_95),
.B(n_76),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_138),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_67),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_112),
.Y(n_149)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_66),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_128),
.B(n_101),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_145),
.A2(n_150),
.B(n_152),
.Y(n_177)
);

OAI32xp33_ASAP7_75t_L g146 ( 
.A1(n_131),
.A2(n_90),
.A3(n_103),
.B1(n_108),
.B2(n_100),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_149),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_90),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_147),
.B(n_155),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_125),
.A2(n_93),
.B1(n_97),
.B2(n_27),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_91),
.B(n_97),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_153),
.A2(n_156),
.B(n_1),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_25),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_119),
.A2(n_91),
.B(n_2),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_42),
.Y(n_157)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_113),
.A2(n_58),
.B1(n_42),
.B2(n_36),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_158),
.A2(n_161),
.B1(n_124),
.B2(n_123),
.Y(n_165)
);

INVxp33_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_160),
.A2(n_163),
.B1(n_137),
.B2(n_114),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_113),
.A2(n_8),
.B1(n_15),
.B2(n_3),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_115),
.A2(n_16),
.B1(n_61),
.B2(n_1),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_165),
.A2(n_167),
.B1(n_162),
.B2(n_148),
.Y(n_187)
);

OAI21x1_ASAP7_75t_L g166 ( 
.A1(n_145),
.A2(n_152),
.B(n_118),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_166),
.A2(n_182),
.B(n_184),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_149),
.A2(n_124),
.B1(n_121),
.B2(n_129),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_136),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_142),
.Y(n_188)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_171),
.Y(n_201)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

NOR3xp33_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_120),
.C(n_116),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_173),
.A2(n_179),
.B1(n_180),
.B2(n_185),
.Y(n_204)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_141),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_178),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_160),
.A2(n_133),
.B1(n_132),
.B2(n_3),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_154),
.A2(n_133),
.B1(n_10),
.B2(n_4),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_153),
.A2(n_1),
.B(n_2),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_16),
.Y(n_183)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_143),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_139),
.B(n_16),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_186),
.A2(n_150),
.B1(n_142),
.B2(n_161),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_188),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_192),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_181),
.B1(n_163),
.B2(n_167),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_190),
.A2(n_195),
.B1(n_173),
.B2(n_179),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_181),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_148),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_198),
.C(n_203),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_194),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_146),
.B1(n_157),
.B2(n_158),
.Y(n_195)
);

OAI21xp33_ASAP7_75t_L g197 ( 
.A1(n_176),
.A2(n_143),
.B(n_1),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_16),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_164),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_186),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_201),
.Y(n_206)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_206),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_196),
.B(n_168),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_208),
.B(n_210),
.Y(n_218)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_200),
.Y(n_211)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_211),
.Y(n_228)
);

FAx1_ASAP7_75t_SL g212 ( 
.A(n_193),
.B(n_180),
.CI(n_176),
.CON(n_212),
.SN(n_212)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_215),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_204),
.A2(n_164),
.B1(n_5),
.B2(n_6),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_214),
.A2(n_191),
.B1(n_195),
.B2(n_202),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_191),
.A2(n_4),
.B(n_5),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_189),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_4),
.C(n_6),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_207),
.C(n_209),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_222),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_217),
.B(n_203),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_213),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_225),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_205),
.A2(n_199),
.B(n_212),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_224),
.A2(n_212),
.B(n_215),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_213),
.A2(n_198),
.B1(n_197),
.B2(n_188),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_226),
.A2(n_214),
.B1(n_215),
.B2(n_10),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_11),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_229),
.A2(n_218),
.B(n_219),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_209),
.C(n_207),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_233),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_236),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_220),
.A2(n_6),
.B1(n_7),
.B2(n_11),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_220),
.A2(n_7),
.B(n_11),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_225),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_240),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_231),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_234),
.A2(n_228),
.B(n_224),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_233),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_242),
.A2(n_232),
.B(n_229),
.Y(n_243)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_12),
.C(n_13),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_245),
.B(n_246),
.Y(n_249)
);

FAx1_ASAP7_75t_SL g246 ( 
.A(n_237),
.B(n_230),
.CI(n_226),
.CON(n_246),
.SN(n_246)
);

OAI31xp33_ASAP7_75t_SL g247 ( 
.A1(n_244),
.A2(n_241),
.A3(n_235),
.B(n_239),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_248),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_249),
.B(n_246),
.C(n_12),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_250),
.C(n_12),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_13),
.Y(n_253)
);


endmodule