module real_aes_7076_n_207 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_174, n_156, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_183, n_205, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_3, n_41, n_140, n_153, n_75, n_178, n_19, n_71, n_180, n_40, n_49, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_81, n_133, n_48, n_204, n_37, n_117, n_97, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_207);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_97;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_207;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_364;
wire n_421;
wire n_555;
wire n_319;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_216;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_236;
wire n_278;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_533;
wire n_366;
wire n_346;
wire n_649;
wire n_397;
wire n_293;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_498;
wire n_691;
wire n_481;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_456;
wire n_359;
wire n_312;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_371;
wire n_541;
wire n_224;
wire n_639;
wire n_546;
wire n_587;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_208;
wire n_215;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g627 ( .A(n_0), .Y(n_627) );
AOI22xp5_ASAP7_75t_SL g335 ( .A1(n_1), .A2(n_175), .B1(n_336), .B2(n_337), .Y(n_335) );
AOI22xp33_ASAP7_75t_SL g673 ( .A1(n_2), .A2(n_12), .B1(n_349), .B2(n_455), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_3), .A2(n_92), .B1(n_344), .B2(n_671), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_4), .A2(n_13), .B1(n_412), .B2(n_433), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g382 ( .A(n_5), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_6), .A2(n_46), .B1(n_350), .B2(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g612 ( .A(n_7), .Y(n_612) );
INVx1_ASAP7_75t_L g394 ( .A(n_8), .Y(n_394) );
CKINVDCx20_ASAP7_75t_R g386 ( .A(n_9), .Y(n_386) );
CKINVDCx20_ASAP7_75t_R g422 ( .A(n_10), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_11), .A2(n_117), .B1(n_447), .B2(n_553), .Y(n_582) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_14), .A2(n_89), .B1(n_276), .B2(n_412), .C(n_413), .Y(n_411) );
CKINVDCx20_ASAP7_75t_R g341 ( .A(n_15), .Y(n_341) );
CKINVDCx20_ASAP7_75t_R g248 ( .A(n_16), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g378 ( .A(n_17), .Y(n_378) );
AOI222xp33_ASAP7_75t_L g453 ( .A1(n_18), .A2(n_66), .B1(n_114), .B2(n_454), .C1(n_455), .C2(n_456), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_19), .A2(n_57), .B1(n_519), .B2(n_520), .Y(n_518) );
AOI22xp33_ASAP7_75t_SL g554 ( .A1(n_20), .A2(n_130), .B1(n_486), .B2(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_21), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g620 ( .A(n_22), .Y(n_620) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_23), .Y(n_369) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_24), .B(n_548), .Y(n_547) );
AO22x2_ASAP7_75t_L g229 ( .A1(n_25), .A2(n_70), .B1(n_230), .B2(n_231), .Y(n_229) );
INVx1_ASAP7_75t_L g660 ( .A(n_25), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_26), .A2(n_127), .B1(n_506), .B2(n_508), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_27), .Y(n_504) );
AOI22xp33_ASAP7_75t_SL g347 ( .A1(n_28), .A2(n_157), .B1(n_348), .B2(n_349), .Y(n_347) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_29), .A2(n_126), .B1(n_277), .B2(n_333), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_30), .A2(n_206), .B1(n_534), .B2(n_553), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_31), .A2(n_190), .B1(n_330), .B2(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g617 ( .A(n_32), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g220 ( .A1(n_33), .A2(n_221), .B1(n_321), .B2(n_322), .Y(n_220) );
INVx1_ASAP7_75t_L g321 ( .A(n_33), .Y(n_321) );
INVx1_ASAP7_75t_L g572 ( .A(n_34), .Y(n_572) );
AOI22xp33_ASAP7_75t_SL g549 ( .A1(n_35), .A2(n_135), .B1(n_350), .B2(n_550), .Y(n_549) );
AO22x2_ASAP7_75t_L g233 ( .A1(n_36), .A2(n_75), .B1(n_230), .B2(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g661 ( .A(n_36), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g365 ( .A1(n_37), .A2(n_107), .B1(n_306), .B2(n_345), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_38), .A2(n_128), .B1(n_336), .B2(n_446), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_39), .A2(n_195), .B1(n_353), .B2(n_420), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_40), .A2(n_129), .B1(n_268), .B2(n_277), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_41), .A2(n_67), .B1(n_441), .B2(n_442), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_42), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_43), .A2(n_74), .B1(n_250), .B2(n_257), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_44), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g302 ( .A(n_45), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_47), .A2(n_58), .B1(n_446), .B2(n_579), .Y(n_604) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_48), .Y(n_240) );
AOI22xp5_ASAP7_75t_SL g331 ( .A1(n_49), .A2(n_123), .B1(n_332), .B2(n_333), .Y(n_331) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_50), .Y(n_468) );
AOI221xp5_ASAP7_75t_L g418 ( .A1(n_51), .A2(n_82), .B1(n_419), .B2(n_420), .C(n_421), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_52), .A2(n_402), .B1(n_403), .B2(n_426), .Y(n_401) );
INVx1_ASAP7_75t_L g426 ( .A(n_52), .Y(n_426) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_53), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_54), .A2(n_200), .B1(n_488), .B2(n_489), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_55), .Y(n_514) );
AOI22xp33_ASAP7_75t_SL g552 ( .A1(n_56), .A2(n_149), .B1(n_489), .B2(n_553), .Y(n_552) );
AOI22xp5_ASAP7_75t_SL g328 ( .A1(n_59), .A2(n_113), .B1(n_329), .B2(n_330), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_60), .A2(n_166), .B1(n_353), .B2(n_356), .Y(n_352) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_61), .Y(n_472) );
AO22x2_ASAP7_75t_L g464 ( .A1(n_62), .A2(n_465), .B1(n_493), .B2(n_494), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_62), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_63), .A2(n_174), .B1(n_251), .B2(n_486), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g281 ( .A(n_64), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_65), .A2(n_168), .B1(n_419), .B2(n_450), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_68), .A2(n_118), .B1(n_534), .B2(n_558), .Y(n_677) );
INVx1_ASAP7_75t_L g583 ( .A(n_69), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g373 ( .A(n_71), .Y(n_373) );
AOI222xp33_ASAP7_75t_L g424 ( .A1(n_72), .A2(n_91), .B1(n_111), .B2(n_299), .C1(n_304), .C2(n_425), .Y(n_424) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_73), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_76), .A2(n_153), .B1(n_258), .B2(n_269), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g297 ( .A(n_77), .Y(n_297) );
INVx1_ASAP7_75t_L g215 ( .A(n_78), .Y(n_215) );
INVx1_ASAP7_75t_L g605 ( .A(n_79), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_80), .A2(n_112), .B1(n_444), .B2(n_447), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_81), .A2(n_108), .B1(n_273), .B2(n_276), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_83), .B(n_636), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_84), .A2(n_152), .B1(n_553), .B2(n_581), .Y(n_678) );
INVx1_ASAP7_75t_L g211 ( .A(n_85), .Y(n_211) );
AOI22xp33_ASAP7_75t_SL g544 ( .A1(n_86), .A2(n_116), .B1(n_306), .B2(n_348), .Y(n_544) );
AOI22xp33_ASAP7_75t_SL g680 ( .A1(n_87), .A2(n_131), .B1(n_273), .B2(n_523), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_88), .B(n_420), .Y(n_568) );
INVx1_ASAP7_75t_L g367 ( .A(n_90), .Y(n_367) );
CKINVDCx20_ASAP7_75t_R g357 ( .A(n_93), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_94), .A2(n_164), .B1(n_348), .B2(n_349), .Y(n_593) );
CKINVDCx20_ASAP7_75t_R g314 ( .A(n_95), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_96), .B(n_567), .Y(n_592) );
INVx1_ASAP7_75t_L g629 ( .A(n_97), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_98), .A2(n_188), .B1(n_530), .B2(n_533), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_99), .A2(n_136), .B1(n_491), .B2(n_558), .Y(n_599) );
INVx1_ASAP7_75t_L g640 ( .A(n_100), .Y(n_640) );
CKINVDCx20_ASAP7_75t_R g286 ( .A(n_101), .Y(n_286) );
INVx1_ASAP7_75t_L g416 ( .A(n_102), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_103), .A2(n_608), .B1(n_641), .B2(n_642), .Y(n_607) );
CKINVDCx16_ASAP7_75t_R g641 ( .A(n_103), .Y(n_641) );
INVx1_ASAP7_75t_L g595 ( .A(n_104), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_105), .A2(n_180), .B1(n_526), .B2(n_528), .Y(n_525) );
INVx1_ASAP7_75t_L g396 ( .A(n_106), .Y(n_396) );
AOI221xp5_ASAP7_75t_L g405 ( .A1(n_109), .A2(n_148), .B1(n_329), .B2(n_406), .C(n_407), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g343 ( .A1(n_110), .A2(n_139), .B1(n_344), .B2(n_345), .Y(n_343) );
AND2x2_ASAP7_75t_L g214 ( .A(n_115), .B(n_215), .Y(n_214) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_119), .A2(n_172), .B1(n_345), .B2(n_452), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g265 ( .A(n_120), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_121), .A2(n_155), .B1(n_257), .B2(n_522), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_122), .A2(n_181), .B1(n_622), .B2(n_624), .Y(n_621) );
AND2x6_ASAP7_75t_L g210 ( .A(n_124), .B(n_211), .Y(n_210) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_124), .Y(n_654) );
AO22x2_ASAP7_75t_L g237 ( .A1(n_125), .A2(n_171), .B1(n_230), .B2(n_234), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g371 ( .A(n_132), .Y(n_371) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_133), .Y(n_383) );
AOI22xp33_ASAP7_75t_SL g580 ( .A1(n_134), .A2(n_192), .B1(n_277), .B2(n_581), .Y(n_580) );
AOI22xp33_ASAP7_75t_SL g602 ( .A1(n_137), .A2(n_151), .B1(n_523), .B2(n_603), .Y(n_602) );
CKINVDCx20_ASAP7_75t_R g692 ( .A(n_138), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_140), .A2(n_191), .B1(n_491), .B2(n_492), .Y(n_490) );
AO22x1_ASAP7_75t_L g407 ( .A1(n_141), .A2(n_169), .B1(n_408), .B2(n_410), .Y(n_407) );
AOI22xp33_ASAP7_75t_SL g557 ( .A1(n_142), .A2(n_184), .B1(n_534), .B2(n_558), .Y(n_557) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_143), .A2(n_664), .B1(n_665), .B2(n_682), .Y(n_663) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_143), .Y(n_682) );
CKINVDCx20_ASAP7_75t_R g560 ( .A(n_144), .Y(n_560) );
AO22x2_ASAP7_75t_L g239 ( .A1(n_145), .A2(n_183), .B1(n_230), .B2(n_231), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_146), .A2(n_196), .B1(n_344), .B2(n_550), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_147), .A2(n_185), .B1(n_475), .B2(n_476), .Y(n_474) );
INVx1_ASAP7_75t_L g364 ( .A(n_150), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_154), .A2(n_202), .B1(n_305), .B2(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g391 ( .A(n_156), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_158), .B(n_567), .Y(n_566) );
AOI22xp33_ASAP7_75t_SL g559 ( .A1(n_159), .A2(n_186), .B1(n_329), .B2(n_333), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_160), .A2(n_205), .B1(n_436), .B2(n_438), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g379 ( .A(n_161), .B(n_337), .Y(n_379) );
AOI211xp5_ASAP7_75t_L g207 ( .A1(n_162), .A2(n_208), .B(n_216), .C(n_662), .Y(n_207) );
INVx1_ASAP7_75t_L g634 ( .A(n_163), .Y(n_634) );
CKINVDCx20_ASAP7_75t_R g271 ( .A(n_165), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_167), .Y(n_482) );
AOI22xp33_ASAP7_75t_SL g578 ( .A1(n_170), .A2(n_176), .B1(n_409), .B2(n_579), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_171), .B(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_173), .B(n_420), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_177), .Y(n_388) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_178), .Y(n_470) );
INVx1_ASAP7_75t_L g639 ( .A(n_179), .Y(n_639) );
INVx1_ASAP7_75t_L g414 ( .A(n_182), .Y(n_414) );
INVx1_ASAP7_75t_L g657 ( .A(n_183), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_187), .Y(n_515) );
INVx1_ASAP7_75t_L g614 ( .A(n_189), .Y(n_614) );
CKINVDCx20_ASAP7_75t_R g423 ( .A(n_193), .Y(n_423) );
INVx1_ASAP7_75t_L g230 ( .A(n_194), .Y(n_230) );
INVx1_ASAP7_75t_L g232 ( .A(n_194), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g310 ( .A(n_197), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g308 ( .A(n_198), .Y(n_308) );
INVx1_ASAP7_75t_L g632 ( .A(n_199), .Y(n_632) );
OA22x2_ASAP7_75t_L g428 ( .A1(n_201), .A2(n_429), .B1(n_430), .B2(n_457), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_201), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g669 ( .A(n_203), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_204), .A2(n_498), .B1(n_535), .B2(n_536), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_204), .Y(n_535) );
INVx1_ASAP7_75t_SL g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_210), .B(n_212), .Y(n_209) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_211), .Y(n_653) );
OAI21xp5_ASAP7_75t_L g690 ( .A1(n_212), .A2(n_652), .B(n_691), .Y(n_690) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_213), .Y(n_212) );
INVxp67_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AOI221xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_459), .B1(n_647), .B2(n_648), .C(n_649), .Y(n_216) );
INVx1_ASAP7_75t_L g648 ( .A(n_217), .Y(n_648) );
AOI22xp5_ASAP7_75t_SL g217 ( .A1(n_218), .A2(n_398), .B1(n_399), .B2(n_458), .Y(n_217) );
INVx1_ASAP7_75t_L g458 ( .A(n_218), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_323), .B1(n_324), .B2(n_397), .Y(n_218) );
INVx3_ASAP7_75t_L g397 ( .A(n_219), .Y(n_397) );
BUFx3_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g322 ( .A(n_221), .Y(n_322) );
AND2x2_ASAP7_75t_SL g221 ( .A(n_222), .B(n_279), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_223), .B(n_261), .Y(n_222) );
OAI221xp5_ASAP7_75t_SL g223 ( .A1(n_224), .A2(n_240), .B1(n_241), .B2(n_248), .C(n_249), .Y(n_223) );
INVx3_ASAP7_75t_L g329 ( .A(n_224), .Y(n_329) );
INVx2_ASAP7_75t_SL g442 ( .A(n_224), .Y(n_442) );
INVx11_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx11_ASAP7_75t_L g395 ( .A(n_225), .Y(n_395) );
AND2x6_ASAP7_75t_L g225 ( .A(n_226), .B(n_235), .Y(n_225) );
AND2x4_ASAP7_75t_L g355 ( .A(n_226), .B(n_270), .Y(n_355) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
OR2x2_ASAP7_75t_L g284 ( .A(n_227), .B(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_233), .Y(n_227) );
AND2x2_ASAP7_75t_L g246 ( .A(n_228), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g256 ( .A(n_228), .B(n_233), .Y(n_256) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g296 ( .A(n_229), .B(n_237), .Y(n_296) );
AND2x2_ASAP7_75t_L g301 ( .A(n_229), .B(n_233), .Y(n_301) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g234 ( .A(n_232), .Y(n_234) );
INVx2_ASAP7_75t_L g247 ( .A(n_233), .Y(n_247) );
INVx1_ASAP7_75t_L g260 ( .A(n_233), .Y(n_260) );
AND2x2_ASAP7_75t_L g264 ( .A(n_235), .B(n_246), .Y(n_264) );
AND2x4_ASAP7_75t_L g275 ( .A(n_235), .B(n_256), .Y(n_275) );
AND2x6_ASAP7_75t_L g300 ( .A(n_235), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_238), .Y(n_235) );
AND2x2_ASAP7_75t_L g270 ( .A(n_236), .B(n_239), .Y(n_270) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_237), .B(n_239), .Y(n_245) );
AND2x2_ASAP7_75t_L g254 ( .A(n_237), .B(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g255 ( .A(n_239), .Y(n_255) );
INVx1_ASAP7_75t_L g295 ( .A(n_239), .Y(n_295) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_242), .Y(n_410) );
BUFx3_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
BUFx3_ASAP7_75t_L g336 ( .A(n_243), .Y(n_336) );
INVx1_ASAP7_75t_L g387 ( .A(n_243), .Y(n_387) );
BUFx2_ASAP7_75t_L g447 ( .A(n_243), .Y(n_447) );
BUFx3_ASAP7_75t_L g492 ( .A(n_243), .Y(n_492) );
BUFx3_ASAP7_75t_L g534 ( .A(n_243), .Y(n_534) );
AND2x4_ASAP7_75t_L g243 ( .A(n_244), .B(n_246), .Y(n_243) );
AND2x2_ASAP7_75t_L g337 ( .A(n_244), .B(n_313), .Y(n_337) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
OR2x6_ASAP7_75t_L g259 ( .A(n_245), .B(n_260), .Y(n_259) );
AND2x4_ASAP7_75t_L g269 ( .A(n_246), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g278 ( .A(n_246), .B(n_254), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_246), .B(n_254), .Y(n_392) );
AND2x2_ASAP7_75t_L g294 ( .A(n_247), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g313 ( .A(n_247), .Y(n_313) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx3_ASAP7_75t_L g330 ( .A(n_252), .Y(n_330) );
INVx4_ASAP7_75t_L g437 ( .A(n_252), .Y(n_437) );
INVx5_ASAP7_75t_L g523 ( .A(n_252), .Y(n_523) );
INVx1_ASAP7_75t_L g555 ( .A(n_252), .Y(n_555) );
BUFx3_ASAP7_75t_L g623 ( .A(n_252), .Y(n_623) );
INVx8_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_256), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_254), .B(n_256), .Y(n_389) );
INVx1_ASAP7_75t_L g320 ( .A(n_255), .Y(n_320) );
NAND2x1p5_ASAP7_75t_L g289 ( .A(n_256), .B(n_270), .Y(n_289) );
AND2x6_ASAP7_75t_L g356 ( .A(n_256), .B(n_270), .Y(n_356) );
CKINVDCx20_ASAP7_75t_R g417 ( .A(n_257), .Y(n_417) );
BUFx4f_ASAP7_75t_SL g257 ( .A(n_258), .Y(n_257) );
BUFx2_ASAP7_75t_L g438 ( .A(n_258), .Y(n_438) );
BUFx2_ASAP7_75t_L g486 ( .A(n_258), .Y(n_486) );
INVx6_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
INVx1_ASAP7_75t_SL g579 ( .A(n_259), .Y(n_579) );
INVx1_ASAP7_75t_SL g624 ( .A(n_259), .Y(n_624) );
INVx1_ASAP7_75t_L g351 ( .A(n_260), .Y(n_351) );
OAI221xp5_ASAP7_75t_SL g261 ( .A1(n_262), .A2(n_265), .B1(n_266), .B2(n_271), .C(n_272), .Y(n_261) );
INVx3_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_263), .Y(n_406) );
BUFx3_ASAP7_75t_L g441 ( .A(n_263), .Y(n_441) );
BUFx3_ASAP7_75t_L g519 ( .A(n_263), .Y(n_519) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
BUFx2_ASAP7_75t_SL g332 ( .A(n_264), .Y(n_332) );
INVx2_ASAP7_75t_L g381 ( .A(n_264), .Y(n_381) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
BUFx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g377 ( .A(n_269), .Y(n_377) );
BUFx3_ASAP7_75t_L g409 ( .A(n_269), .Y(n_409) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_269), .Y(n_446) );
BUFx3_ASAP7_75t_L g489 ( .A(n_269), .Y(n_489) );
INVx1_ASAP7_75t_L g285 ( .A(n_270), .Y(n_285) );
INVx3_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OAI22xp5_ASAP7_75t_SL g380 ( .A1(n_274), .A2(n_381), .B1(n_382), .B2(n_383), .Y(n_380) );
INVx2_ASAP7_75t_L g412 ( .A(n_274), .Y(n_412) );
INVx2_ASAP7_75t_L g528 ( .A(n_274), .Y(n_528) );
INVx2_ASAP7_75t_L g577 ( .A(n_274), .Y(n_577) );
OAI221xp5_ASAP7_75t_SL g616 ( .A1(n_274), .A2(n_617), .B1(n_618), .B2(n_620), .C(n_621), .Y(n_616) );
INVx6_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
BUFx3_ASAP7_75t_L g333 ( .A(n_275), .Y(n_333) );
BUFx3_ASAP7_75t_L g603 ( .A(n_275), .Y(n_603) );
BUFx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g434 ( .A(n_277), .Y(n_434) );
BUFx3_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
BUFx3_ASAP7_75t_L g532 ( .A(n_278), .Y(n_532) );
BUFx3_ASAP7_75t_L g558 ( .A(n_278), .Y(n_558) );
NOR3xp33_ASAP7_75t_L g279 ( .A(n_280), .B(n_290), .C(n_309), .Y(n_279) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .B1(n_286), .B2(n_287), .Y(n_280) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g469 ( .A(n_283), .Y(n_469) );
INVx1_ASAP7_75t_SL g628 ( .A(n_283), .Y(n_628) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OAI21xp5_ASAP7_75t_L g363 ( .A1(n_284), .A2(n_364), .B(n_365), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_287), .A2(n_468), .B1(n_469), .B2(n_470), .Y(n_467) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx3_ASAP7_75t_L g368 ( .A(n_289), .Y(n_368) );
OAI222xp33_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_297), .B1(n_298), .B2(n_302), .C1(n_303), .C2(n_308), .Y(n_290) );
OAI222xp33_ASAP7_75t_L g511 ( .A1(n_291), .A2(n_303), .B1(n_512), .B2(n_513), .C1(n_514), .C2(n_515), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_292), .Y(n_291) );
BUFx6f_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_293), .Y(n_348) );
BUFx4f_ASAP7_75t_SL g455 ( .A(n_293), .Y(n_455) );
BUFx2_ASAP7_75t_L g475 ( .A(n_293), .Y(n_475) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_293), .Y(n_570) );
AND2x4_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
INVx1_ASAP7_75t_L g307 ( .A(n_295), .Y(n_307) );
AND2x4_ASAP7_75t_L g306 ( .A(n_296), .B(n_307), .Y(n_306) );
NAND2x1p5_ASAP7_75t_L g312 ( .A(n_296), .B(n_313), .Y(n_312) );
AND2x4_ASAP7_75t_L g350 ( .A(n_296), .B(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_SL g631 ( .A(n_299), .Y(n_631) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g342 ( .A(n_300), .Y(n_342) );
INVx2_ASAP7_75t_SL g372 ( .A(n_300), .Y(n_372) );
BUFx3_ASAP7_75t_L g454 ( .A(n_300), .Y(n_454) );
INVx2_ASAP7_75t_L g513 ( .A(n_300), .Y(n_513) );
INVx1_ASAP7_75t_L g318 ( .A(n_301), .Y(n_318) );
AND2x4_ASAP7_75t_L g345 ( .A(n_301), .B(n_320), .Y(n_345) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx3_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx12f_ASAP7_75t_L g344 ( .A(n_306), .Y(n_344) );
BUFx6f_ASAP7_75t_L g637 ( .A(n_306), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_311), .B1(n_314), .B2(n_315), .Y(n_309) );
BUFx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_312), .A2(n_367), .B1(n_368), .B2(n_369), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_312), .A2(n_315), .B1(n_422), .B2(n_423), .Y(n_421) );
INVx4_ASAP7_75t_L g481 ( .A(n_312), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_315), .A2(n_480), .B1(n_639), .B2(n_640), .Y(n_638) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
CKINVDCx16_ASAP7_75t_R g316 ( .A(n_317), .Y(n_316) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_317), .A2(n_479), .B1(n_480), .B2(n_482), .Y(n_478) );
OR2x6_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI22xp5_ASAP7_75t_SL g324 ( .A1(n_325), .A2(n_326), .B1(n_358), .B2(n_359), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
XOR2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_357), .Y(n_326) );
NAND4xp75_ASAP7_75t_SL g327 ( .A(n_328), .B(n_331), .C(n_334), .D(n_339), .Y(n_327) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_338), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_340), .B(n_346), .Y(n_339) );
OAI21xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_342), .B(n_343), .Y(n_340) );
BUFx4f_ASAP7_75t_SL g456 ( .A(n_344), .Y(n_456) );
INVx2_ASAP7_75t_L g477 ( .A(n_344), .Y(n_477) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_345), .Y(n_510) );
BUFx3_ASAP7_75t_L g550 ( .A(n_345), .Y(n_550) );
BUFx2_ASAP7_75t_SL g574 ( .A(n_345), .Y(n_574) );
BUFx2_ASAP7_75t_SL g671 ( .A(n_345), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_352), .Y(n_346) );
INVx4_ASAP7_75t_L g374 ( .A(n_348), .Y(n_374) );
BUFx3_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx2_ASAP7_75t_L g452 ( .A(n_350), .Y(n_452) );
INVx1_ASAP7_75t_L g507 ( .A(n_350), .Y(n_507) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_353), .Y(n_419) );
INVx5_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g548 ( .A(n_354), .Y(n_548) );
INVx2_ASAP7_75t_L g567 ( .A(n_354), .Y(n_567) );
INVx4_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx4f_ASAP7_75t_L g420 ( .A(n_356), .Y(n_420) );
BUFx2_ASAP7_75t_L g450 ( .A(n_356), .Y(n_450) );
BUFx2_ASAP7_75t_L g591 ( .A(n_356), .Y(n_591) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
BUFx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
XNOR2x1_ASAP7_75t_L g360 ( .A(n_361), .B(n_396), .Y(n_360) );
AND3x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_375), .C(n_384), .Y(n_361) );
NOR3xp33_ASAP7_75t_L g362 ( .A(n_363), .B(n_366), .C(n_370), .Y(n_362) );
INVx2_ASAP7_75t_L g503 ( .A(n_368), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_368), .A2(n_627), .B1(n_628), .B2(n_629), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_372), .B1(n_373), .B2(n_374), .Y(n_370) );
INVx3_ASAP7_75t_L g425 ( .A(n_374), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_376), .B(n_380), .Y(n_375) );
OAI21xp5_ASAP7_75t_SL g376 ( .A1(n_377), .A2(n_378), .B(n_379), .Y(n_376) );
INVx1_ASAP7_75t_L g520 ( .A(n_377), .Y(n_520) );
INVx3_ASAP7_75t_L g488 ( .A(n_381), .Y(n_488) );
INVx3_ASAP7_75t_L g553 ( .A(n_381), .Y(n_553) );
NOR3xp33_ASAP7_75t_L g384 ( .A(n_385), .B(n_390), .C(n_393), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B1(n_388), .B2(n_389), .Y(n_385) );
BUFx2_ASAP7_75t_R g415 ( .A(n_389), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVx1_ASAP7_75t_L g619 ( .A(n_392), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx2_ASAP7_75t_SL g491 ( .A(n_395), .Y(n_491) );
INVx5_ASAP7_75t_SL g581 ( .A(n_395), .Y(n_581) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
OAI22xp5_ASAP7_75t_SL g399 ( .A1(n_400), .A2(n_401), .B1(n_427), .B2(n_428), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AND4x1_ASAP7_75t_L g404 ( .A(n_405), .B(n_411), .C(n_418), .D(n_424), .Y(n_404) );
INVx1_ASAP7_75t_SL g611 ( .A(n_406), .Y(n_611) );
BUFx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_415), .B1(n_416), .B2(n_417), .Y(n_413) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_SL g457 ( .A(n_430), .Y(n_457) );
NAND4xp75_ASAP7_75t_L g430 ( .A(n_431), .B(n_439), .C(n_448), .D(n_453), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_435), .Y(n_431) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_443), .Y(n_439) );
INVx1_ASAP7_75t_L g613 ( .A(n_442), .Y(n_613) );
INVx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx4_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_SL g448 ( .A(n_449), .B(n_451), .Y(n_448) );
INVx3_ASAP7_75t_L g473 ( .A(n_454), .Y(n_473) );
INVx1_ASAP7_75t_L g647 ( .A(n_459), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B1(n_537), .B2(n_646), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
XOR2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_495), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_SL g493 ( .A(n_465), .Y(n_493) );
AND2x2_ASAP7_75t_SL g465 ( .A(n_466), .B(n_483), .Y(n_465) );
NOR3xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_471), .C(n_478), .Y(n_466) );
OAI221xp5_ASAP7_75t_L g500 ( .A1(n_469), .A2(n_501), .B1(n_502), .B2(n_504), .C(n_505), .Y(n_500) );
OAI21xp33_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B(n_474), .Y(n_471) );
INVx1_ASAP7_75t_L g633 ( .A(n_475), .Y(n_633) );
INVx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AND4x1_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .C(n_487), .D(n_490), .Y(n_483) );
INVx1_ASAP7_75t_L g527 ( .A(n_491), .Y(n_527) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_SL g536 ( .A(n_498), .Y(n_536) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_516), .Y(n_498) );
NOR2xp33_ASAP7_75t_SL g499 ( .A(n_500), .B(n_511), .Y(n_499) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_SL g509 ( .A(n_510), .Y(n_509) );
OAI21xp5_ASAP7_75t_SL g542 ( .A1(n_513), .A2(n_543), .B(n_544), .Y(n_542) );
OAI21xp5_ASAP7_75t_L g571 ( .A1(n_513), .A2(n_572), .B(n_573), .Y(n_571) );
OAI21xp5_ASAP7_75t_SL g594 ( .A1(n_513), .A2(n_595), .B(n_596), .Y(n_594) );
OAI21xp5_ASAP7_75t_L g668 ( .A1(n_513), .A2(n_669), .B(n_670), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_517), .B(n_524), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_521), .Y(n_517) );
BUFx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_525), .B(n_529), .Y(n_524) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
BUFx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g646 ( .A(n_537), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_539), .B1(n_561), .B2(n_645), .Y(n_537) );
INVx4_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
XOR2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_560), .Y(n_539) );
NAND3x1_ASAP7_75t_L g540 ( .A(n_541), .B(n_551), .C(n_556), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_545), .Y(n_541) );
NAND3xp33_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .C(n_549), .Y(n_545) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_554), .Y(n_551) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_559), .Y(n_556) );
INVx1_ASAP7_75t_L g645 ( .A(n_561), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_584), .B1(n_643), .B2(n_644), .Y(n_561) );
INVx1_ASAP7_75t_L g643 ( .A(n_562), .Y(n_643) );
XOR2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_583), .Y(n_562) );
NAND4xp75_ASAP7_75t_SL g563 ( .A(n_564), .B(n_575), .C(n_580), .D(n_582), .Y(n_563) );
NOR2xp67_ASAP7_75t_SL g564 ( .A(n_565), .B(n_571), .Y(n_564) );
NAND3xp33_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .C(n_569), .Y(n_565) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_578), .Y(n_575) );
INVx1_ASAP7_75t_SL g644 ( .A(n_584), .Y(n_644) );
XOR2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_606), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
XOR2x2_ASAP7_75t_SL g586 ( .A(n_587), .B(n_605), .Y(n_586) );
NAND2x1p5_ASAP7_75t_L g587 ( .A(n_588), .B(n_597), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_589), .B(n_594), .Y(n_588) );
NAND3xp33_ASAP7_75t_L g589 ( .A(n_590), .B(n_592), .C(n_593), .Y(n_589) );
NOR2x1_ASAP7_75t_L g597 ( .A(n_598), .B(n_601), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g642 ( .A(n_608), .Y(n_642) );
AND2x2_ASAP7_75t_SL g608 ( .A(n_609), .B(n_625), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_610), .B(n_616), .Y(n_609) );
OAI221xp5_ASAP7_75t_SL g610 ( .A1(n_611), .A2(n_612), .B1(n_613), .B2(n_614), .C(n_615), .Y(n_610) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx3_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NOR3xp33_ASAP7_75t_L g625 ( .A(n_626), .B(n_630), .C(n_638), .Y(n_625) );
OAI221xp5_ASAP7_75t_SL g630 ( .A1(n_631), .A2(n_632), .B1(n_633), .B2(n_634), .C(n_635), .Y(n_630) );
BUFx4f_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
NOR2x1_ASAP7_75t_L g650 ( .A(n_651), .B(n_655), .Y(n_650) );
OR2x2_ASAP7_75t_SL g696 ( .A(n_651), .B(n_656), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .Y(n_651) );
CKINVDCx20_ASAP7_75t_R g684 ( .A(n_652), .Y(n_684) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_653), .B(n_688), .Y(n_691) );
CKINVDCx16_ASAP7_75t_R g688 ( .A(n_654), .Y(n_688) );
CKINVDCx20_ASAP7_75t_R g655 ( .A(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
OAI322xp33_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_683), .A3(n_685), .B1(n_689), .B2(n_692), .C1(n_693), .C2(n_694), .Y(n_662) );
CKINVDCx20_ASAP7_75t_R g664 ( .A(n_665), .Y(n_664) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
XOR2x2_ASAP7_75t_L g693 ( .A(n_666), .B(n_692), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g666 ( .A(n_667), .B(n_675), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_668), .B(n_672), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_679), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
BUFx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_690), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g694 ( .A(n_695), .Y(n_694) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_696), .Y(n_695) );
endmodule