module fake_jpeg_31116_n_545 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_545);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_545;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_15),
.B(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_52),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_53),
.Y(n_148)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_57),
.Y(n_165)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_59),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_63),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_18),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_64),
.B(n_72),
.Y(n_119)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_69),
.Y(n_150)
);

BUFx4f_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_19),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_73),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_38),
.B(n_18),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_74),
.B(n_88),
.Y(n_129)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_77),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_80),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_82),
.B(n_103),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_85),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_86),
.Y(n_138)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_87),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_46),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_19),
.B(n_18),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_89),
.B(n_92),
.Y(n_155)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_94),
.Y(n_140)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_96),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_97),
.Y(n_164)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_20),
.Y(n_101)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_20),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_72),
.A2(n_51),
.B1(n_27),
.B2(n_30),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_107),
.B(n_118),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_64),
.A2(n_51),
.B1(n_27),
.B2(n_30),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_108),
.A2(n_109),
.B1(n_133),
.B2(n_154),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_21),
.B1(n_26),
.B2(n_39),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_46),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_111),
.B(n_139),
.Y(n_200)
);

OR2x4_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_45),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_96),
.A2(n_40),
.B1(n_47),
.B2(n_43),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_63),
.A2(n_95),
.B1(n_91),
.B2(n_84),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_137),
.A2(n_50),
.B1(n_47),
.B2(n_36),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_67),
.A2(n_21),
.B1(n_26),
.B2(n_39),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_52),
.B(n_45),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_163),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_53),
.B(n_44),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_156),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_57),
.A2(n_102),
.B1(n_60),
.B2(n_97),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_100),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_66),
.B(n_44),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_162),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_83),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_78),
.B(n_46),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_117),
.A2(n_40),
.B1(n_47),
.B2(n_43),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_167),
.A2(n_184),
.B1(n_204),
.B2(n_215),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_137),
.A2(n_94),
.B1(n_86),
.B2(n_81),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_168),
.A2(n_214),
.B1(n_165),
.B2(n_128),
.Y(n_274)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_170),
.Y(n_264)
);

AND2x2_ASAP7_75t_SL g172 ( 
.A(n_104),
.B(n_79),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_172),
.B(n_177),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_166),
.A2(n_33),
.B(n_25),
.Y(n_173)
);

O2A1O1Ixp33_ASAP7_75t_L g270 ( 
.A1(n_173),
.A2(n_34),
.B(n_128),
.C(n_164),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_174),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_122),
.Y(n_175)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_175),
.Y(n_276)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_106),
.Y(n_176)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_176),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_124),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_178),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_130),
.A2(n_50),
.B1(n_47),
.B2(n_48),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_179),
.A2(n_138),
.B1(n_164),
.B2(n_140),
.Y(n_254)
);

INVx5_ASAP7_75t_SL g180 ( 
.A(n_161),
.Y(n_180)
);

CKINVDCx6p67_ASAP7_75t_R g252 ( 
.A(n_180),
.Y(n_252)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_110),
.Y(n_182)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_182),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_125),
.A2(n_40),
.B1(n_50),
.B2(n_25),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_185),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_112),
.Y(n_186)
);

INVx13_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_166),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_187),
.B(n_192),
.Y(n_234)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_121),
.Y(n_188)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_188),
.Y(n_247)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_189),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_119),
.A2(n_50),
.B1(n_48),
.B2(n_25),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_191),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_111),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_157),
.Y(n_193)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_193),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_129),
.B(n_46),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_194),
.B(n_207),
.Y(n_243)
);

INVx11_ASAP7_75t_L g195 ( 
.A(n_110),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_195),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_105),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_196),
.B(n_198),
.Y(n_273)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_146),
.Y(n_197)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_197),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_105),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_148),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g233 ( 
.A(n_199),
.Y(n_233)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_116),
.Y(n_201)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_201),
.Y(n_242)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_123),
.Y(n_202)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_202),
.Y(n_265)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_152),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_203),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_113),
.A2(n_40),
.B1(n_48),
.B2(n_33),
.Y(n_204)
);

A2O1A1Ixp33_ASAP7_75t_L g205 ( 
.A1(n_119),
.A2(n_33),
.B(n_17),
.C(n_16),
.Y(n_205)
);

OR2x2_ASAP7_75t_SL g240 ( 
.A(n_205),
.B(n_32),
.Y(n_240)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_126),
.Y(n_206)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_206),
.Y(n_269)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_132),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_131),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_208),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_155),
.B(n_17),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_217),
.Y(n_232)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_115),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_210),
.B(n_212),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g239 ( 
.A(n_211),
.Y(n_239)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_135),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_134),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_213),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_133),
.A2(n_40),
.B1(n_36),
.B2(n_34),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_147),
.A2(n_34),
.B1(n_32),
.B2(n_36),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_136),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_216),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_155),
.B(n_34),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_150),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_218),
.B(n_222),
.Y(n_250)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_159),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_223),
.Y(n_251)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_149),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_220),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_129),
.B(n_34),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_32),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_137),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_160),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_120),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_225),
.Y(n_258)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_161),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_120),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_226),
.Y(n_238)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_138),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_226),
.Y(n_262)
);

NAND2xp33_ASAP7_75t_SL g311 ( 
.A(n_236),
.B(n_240),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_222),
.A2(n_141),
.B1(n_135),
.B2(n_140),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_245),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_254),
.A2(n_250),
.B1(n_252),
.B2(n_264),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_183),
.B(n_144),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_266),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_200),
.B(n_32),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_261),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_200),
.B(n_32),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_263),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_171),
.B(n_190),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_173),
.B(n_114),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_181),
.B(n_114),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_169),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_270),
.A2(n_218),
.B(n_186),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_208),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_277),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_274),
.A2(n_177),
.B1(n_172),
.B2(n_185),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_275),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_181),
.B(n_0),
.Y(n_277)
);

CKINVDCx12_ASAP7_75t_R g278 ( 
.A(n_188),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_188),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_192),
.C(n_200),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_281),
.B(n_287),
.C(n_302),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_282),
.B(n_303),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_284),
.B(n_297),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_232),
.B(n_172),
.C(n_214),
.Y(n_287)
);

OAI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_270),
.A2(n_205),
.B1(n_180),
.B2(n_212),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_288),
.A2(n_305),
.B1(n_325),
.B2(n_247),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_289),
.B(n_327),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_290),
.A2(n_294),
.B1(n_319),
.B2(n_272),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_232),
.B(n_225),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_291),
.B(n_299),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_276),
.Y(n_292)
);

BUFx12f_ASAP7_75t_L g358 ( 
.A(n_292),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_243),
.B(n_223),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_293),
.B(n_300),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_230),
.A2(n_201),
.B1(n_206),
.B2(n_189),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_242),
.Y(n_295)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_295),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_250),
.A2(n_178),
.B(n_203),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_296),
.A2(n_301),
.B(n_307),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_266),
.B(n_216),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_236),
.B(n_268),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_298),
.B(n_304),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_234),
.B(n_197),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_273),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_250),
.A2(n_219),
.B(n_210),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_260),
.B(n_213),
.C(n_220),
.Y(n_302)
);

NAND2x1_ASAP7_75t_SL g303 ( 
.A(n_252),
.B(n_195),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_230),
.B(n_182),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_240),
.A2(n_211),
.B1(n_199),
.B2(n_175),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_242),
.Y(n_306)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_306),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_237),
.A2(n_0),
.B(n_1),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_256),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_308),
.B(n_316),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_230),
.B(n_261),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_309),
.B(n_314),
.Y(n_357)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_269),
.Y(n_310)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_310),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_260),
.B(n_174),
.C(n_2),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_312),
.B(n_326),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_313),
.A2(n_324),
.B1(n_231),
.B2(n_271),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_261),
.B(n_0),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_279),
.B(n_2),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_315),
.B(n_318),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_279),
.B(n_3),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_269),
.Y(n_317)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_317),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_264),
.B(n_3),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_274),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_276),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_320),
.Y(n_337)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_252),
.Y(n_321)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_321),
.Y(n_356)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_252),
.Y(n_322)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_322),
.Y(n_360)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_235),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_323),
.B(n_246),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_254),
.B(n_8),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_233),
.Y(n_327)
);

AO22x1_ASAP7_75t_L g331 ( 
.A1(n_283),
.A2(n_248),
.B1(n_246),
.B2(n_251),
.Y(n_331)
);

OA21x2_ASAP7_75t_L g391 ( 
.A1(n_331),
.A2(n_301),
.B(n_318),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_332),
.A2(n_354),
.B1(n_321),
.B2(n_322),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_283),
.A2(n_309),
.B(n_282),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_335),
.A2(n_340),
.B(n_364),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_280),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_338),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_SL g339 ( 
.A(n_311),
.B(n_241),
.C(n_247),
.Y(n_339)
);

OAI21x1_ASAP7_75t_SL g402 ( 
.A1(n_339),
.A2(n_320),
.B(n_233),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_304),
.A2(n_258),
.B(n_241),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_298),
.B(n_253),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_343),
.B(n_285),
.C(n_314),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_344),
.B(n_367),
.Y(n_378)
);

OAI21xp33_ASAP7_75t_L g346 ( 
.A1(n_291),
.A2(n_259),
.B(n_228),
.Y(n_346)
);

OA21x2_ASAP7_75t_SL g400 ( 
.A1(n_346),
.A2(n_331),
.B(n_341),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_303),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_347),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_300),
.B(n_231),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_350),
.B(n_353),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_286),
.B(n_256),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_284),
.A2(n_228),
.B1(n_267),
.B2(n_255),
.Y(n_354)
);

BUFx24_ASAP7_75t_SL g359 ( 
.A(n_299),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_359),
.B(n_316),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_281),
.B(n_259),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_361),
.B(n_312),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_363),
.A2(n_365),
.B1(n_290),
.B2(n_294),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_297),
.A2(n_238),
.B(n_244),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_326),
.A2(n_249),
.B1(n_238),
.B2(n_272),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_307),
.A2(n_244),
.B(n_265),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_366),
.A2(n_369),
.B(n_233),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_287),
.B(n_235),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_368),
.B(n_302),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_296),
.A2(n_265),
.B(n_229),
.Y(n_369)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_329),
.Y(n_371)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_371),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_345),
.B(n_315),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_373),
.B(n_390),
.Y(n_417)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_329),
.Y(n_374)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_374),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_330),
.B(n_285),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_375),
.B(n_330),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_376),
.A2(n_395),
.B1(n_343),
.B2(n_348),
.Y(n_411)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_334),
.Y(n_377)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_377),
.Y(n_433)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_356),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_379),
.B(n_380),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_382),
.A2(n_363),
.B1(n_364),
.B2(n_365),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_345),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_384),
.Y(n_414)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_334),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_385),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_386),
.B(n_375),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_387),
.B(n_333),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_367),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_388),
.Y(n_430)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_349),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_389),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_391),
.B(n_392),
.Y(n_425)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_349),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_351),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_393),
.B(n_398),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_332),
.A2(n_326),
.B1(n_285),
.B2(n_325),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_394),
.A2(n_401),
.B1(n_347),
.B2(n_344),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_342),
.A2(n_319),
.B1(n_306),
.B2(n_295),
.Y(n_395)
);

NAND2x1_ASAP7_75t_L g396 ( 
.A(n_339),
.B(n_331),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_396),
.A2(n_400),
.B(n_402),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_338),
.B(n_308),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_397),
.B(n_399),
.Y(n_434)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_351),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_348),
.B(n_327),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_354),
.A2(n_317),
.B1(n_310),
.B2(n_303),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_403),
.A2(n_328),
.B(n_366),
.Y(n_420)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_356),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_SL g422 ( 
.A1(n_404),
.A2(n_360),
.B1(n_358),
.B2(n_337),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_405),
.B(n_416),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_406),
.B(n_428),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_407),
.A2(n_408),
.B1(n_424),
.B2(n_391),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_411),
.A2(n_415),
.B1(n_429),
.B2(n_432),
.Y(n_458)
);

OA21x2_ASAP7_75t_L g413 ( 
.A1(n_400),
.A2(n_352),
.B(n_342),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_413),
.B(n_431),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_376),
.A2(n_328),
.B1(n_368),
.B2(n_362),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_380),
.B(n_335),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_418),
.B(n_426),
.C(n_427),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_420),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_422),
.A2(n_398),
.B(n_393),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_394),
.A2(n_378),
.B1(n_382),
.B2(n_383),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_386),
.B(n_352),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_381),
.B(n_362),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_370),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_395),
.A2(n_328),
.B1(n_355),
.B2(n_360),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_402),
.A2(n_341),
.B1(n_340),
.B2(n_369),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_384),
.A2(n_355),
.B1(n_357),
.B2(n_336),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_435),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_436),
.B(n_441),
.Y(n_472)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_435),
.Y(n_439)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_439),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_414),
.B(n_372),
.Y(n_440)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_440),
.Y(n_477)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_419),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_430),
.B(n_388),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_442),
.B(n_443),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_430),
.B(n_434),
.Y(n_443)
);

NOR3xp33_ASAP7_75t_SL g444 ( 
.A(n_417),
.B(n_372),
.C(n_378),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g480 ( 
.A(n_444),
.Y(n_480)
);

NOR3xp33_ASAP7_75t_L g445 ( 
.A(n_414),
.B(n_383),
.C(n_396),
.Y(n_445)
);

AOI21x1_ASAP7_75t_L g482 ( 
.A1(n_445),
.A2(n_455),
.B(n_462),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_405),
.B(n_416),
.C(n_427),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_446),
.B(n_459),
.C(n_418),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_426),
.B(n_373),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_448),
.B(n_453),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_449),
.A2(n_452),
.B1(n_431),
.B2(n_429),
.Y(n_463)
);

NAND5xp2_ASAP7_75t_L g450 ( 
.A(n_425),
.B(n_396),
.C(n_381),
.D(n_391),
.E(n_401),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_450),
.A2(n_461),
.B(n_433),
.Y(n_469)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_419),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_451),
.A2(n_456),
.B1(n_457),
.B2(n_433),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_424),
.A2(n_391),
.B1(n_403),
.B2(n_404),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_413),
.B(n_377),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_409),
.B(n_379),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_423),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_423),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_415),
.B(n_357),
.C(n_336),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_425),
.A2(n_392),
.B(n_389),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_463),
.B(n_469),
.Y(n_497)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_464),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_449),
.A2(n_411),
.B1(n_409),
.B2(n_413),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_465),
.B(n_466),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_452),
.A2(n_408),
.B1(n_410),
.B2(n_420),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_467),
.B(n_454),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_460),
.B(n_410),
.C(n_421),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_468),
.B(n_476),
.C(n_479),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_469),
.A2(n_470),
.B(n_455),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_438),
.A2(n_385),
.B(n_374),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_458),
.A2(n_412),
.B1(n_371),
.B2(n_337),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_473),
.A2(n_443),
.B1(n_450),
.B2(n_451),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_462),
.A2(n_358),
.B1(n_292),
.B2(n_320),
.Y(n_474)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_474),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_439),
.A2(n_358),
.B1(n_249),
.B2(n_323),
.Y(n_475)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_475),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_460),
.B(n_229),
.C(n_358),
.Y(n_476)
);

FAx1_ASAP7_75t_SL g478 ( 
.A(n_454),
.B(n_8),
.CI(n_9),
.CON(n_478),
.SN(n_478)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_478),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_446),
.B(n_233),
.C(n_239),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_437),
.B(n_239),
.C(n_9),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_484),
.B(n_442),
.C(n_438),
.Y(n_490)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_477),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_485),
.B(n_495),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_468),
.B(n_437),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_489),
.B(n_493),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_490),
.B(n_494),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_467),
.B(n_461),
.C(n_459),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_491),
.B(n_500),
.C(n_479),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_480),
.A2(n_447),
.B1(n_444),
.B2(n_454),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_497),
.B(n_466),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_498),
.B(n_482),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_481),
.B(n_457),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_499),
.B(n_478),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_476),
.B(n_456),
.C(n_441),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_503),
.B(n_505),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_492),
.A2(n_483),
.B1(n_473),
.B2(n_471),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_504),
.A2(n_496),
.B1(n_488),
.B2(n_501),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_493),
.A2(n_463),
.B1(n_465),
.B2(n_482),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_506),
.A2(n_486),
.B1(n_497),
.B2(n_490),
.Y(n_517)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_507),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_494),
.B(n_481),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_508),
.B(n_512),
.C(n_515),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_491),
.A2(n_470),
.B(n_472),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_511),
.A2(n_513),
.B(n_498),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_487),
.B(n_483),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_486),
.A2(n_472),
.B(n_484),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_514),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_487),
.B(n_474),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_516),
.B(n_517),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_509),
.A2(n_500),
.B(n_485),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_520),
.A2(n_524),
.B(n_525),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_522),
.B(n_525),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_506),
.A2(n_464),
.B(n_478),
.Y(n_524)
);

OAI22x1_ASAP7_75t_L g525 ( 
.A1(n_507),
.A2(n_475),
.B1(n_489),
.B2(n_239),
.Y(n_525)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_527),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_518),
.B(n_512),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_529),
.B(n_531),
.Y(n_532)
);

XNOR2x1_ASAP7_75t_L g530 ( 
.A(n_521),
.B(n_502),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_530),
.B(n_521),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_518),
.B(n_523),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_528),
.A2(n_519),
.B(n_510),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_533),
.A2(n_526),
.B(n_503),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_535),
.B(n_502),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_536),
.B(n_537),
.C(n_535),
.Y(n_539)
);

OAI321xp33_ASAP7_75t_L g538 ( 
.A1(n_536),
.A2(n_534),
.A3(n_532),
.B1(n_524),
.B2(n_515),
.C(n_505),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_SL g540 ( 
.A1(n_538),
.A2(n_539),
.B(n_508),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_540),
.B(n_239),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_541),
.A2(n_8),
.B(n_10),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g543 ( 
.A1(n_542),
.A2(n_10),
.B(n_11),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_543),
.B(n_11),
.C(n_13),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_544),
.B(n_11),
.C(n_13),
.Y(n_545)
);


endmodule