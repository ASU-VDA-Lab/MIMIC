module fake_aes_1979_n_42 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_42);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_42;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_30;
wire n_13;
wire n_33;
wire n_26;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
AND2x4_ASAP7_75t_L g11 ( .A(n_3), .B(n_4), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_0), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_4), .B(n_8), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_0), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_6), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_7), .B(n_5), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_6), .Y(n_17) );
INVx3_ASAP7_75t_L g18 ( .A(n_11), .Y(n_18) );
CKINVDCx16_ASAP7_75t_R g19 ( .A(n_11), .Y(n_19) );
CKINVDCx20_ASAP7_75t_R g20 ( .A(n_14), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_11), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_11), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_12), .Y(n_23) );
AOI22xp33_ASAP7_75t_L g24 ( .A1(n_21), .A2(n_15), .B1(n_17), .B2(n_12), .Y(n_24) );
AOI22xp33_ASAP7_75t_L g25 ( .A1(n_21), .A2(n_15), .B1(n_14), .B2(n_16), .Y(n_25) );
BUFx3_ASAP7_75t_L g26 ( .A(n_18), .Y(n_26) );
AND2x2_ASAP7_75t_L g27 ( .A(n_19), .B(n_13), .Y(n_27) );
AOI22xp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_18), .B1(n_22), .B2(n_20), .Y(n_28) );
OR2x6_ASAP7_75t_L g29 ( .A(n_27), .B(n_22), .Y(n_29) );
NAND3xp33_ASAP7_75t_L g30 ( .A(n_25), .B(n_20), .C(n_23), .Y(n_30) );
INVx2_ASAP7_75t_SL g31 ( .A(n_29), .Y(n_31) );
NAND2x1_ASAP7_75t_L g32 ( .A(n_28), .B(n_24), .Y(n_32) );
NOR2xp33_ASAP7_75t_L g33 ( .A(n_31), .B(n_30), .Y(n_33) );
INVxp67_ASAP7_75t_SL g34 ( .A(n_31), .Y(n_34) );
INVx1_ASAP7_75t_SL g35 ( .A(n_33), .Y(n_35) );
AOI221xp5_ASAP7_75t_L g36 ( .A1(n_34), .A2(n_32), .B1(n_26), .B2(n_3), .C(n_5), .Y(n_36) );
AOI221x1_ASAP7_75t_L g37 ( .A1(n_33), .A2(n_1), .B1(n_2), .B2(n_9), .C(n_10), .Y(n_37) );
CKINVDCx5p33_ASAP7_75t_R g38 ( .A(n_35), .Y(n_38) );
NAND2xp5_ASAP7_75t_L g39 ( .A(n_36), .B(n_26), .Y(n_39) );
NOR2x1_ASAP7_75t_L g40 ( .A(n_39), .B(n_37), .Y(n_40) );
HB1xp67_ASAP7_75t_L g41 ( .A(n_38), .Y(n_41) );
NAND3xp33_ASAP7_75t_L g42 ( .A(n_40), .B(n_41), .C(n_1), .Y(n_42) );
endmodule