module fake_jpeg_21022_n_88 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_88);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_88;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_82;

INVx6_ASAP7_75t_SL g33 ( 
.A(n_15),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_8),
.B(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_46),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_1),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_49),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_1),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_50),
.A2(n_35),
.B1(n_33),
.B2(n_5),
.Y(n_56)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_48),
.B(n_40),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_55),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_56),
.A2(n_38),
.B1(n_4),
.B2(n_5),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_6),
.Y(n_64)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_59),
.B(n_3),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_62),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_64),
.B(n_66),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_65),
.Y(n_74)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_11),
.B(n_13),
.C(n_16),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_22),
.B(n_24),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_18),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_68),
.B(n_69),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_21),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_76),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_78),
.A2(n_71),
.B(n_61),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_74),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_80),
.A2(n_77),
.B(n_75),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_81),
.C(n_75),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_83),
.B(n_73),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_84),
.B(n_67),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_25),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_86),
.A2(n_26),
.B(n_29),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_30),
.B(n_31),
.Y(n_88)
);


endmodule