module real_jpeg_25245_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g112 ( 
.A(n_0),
.Y(n_112)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_0),
.Y(n_113)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_0),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_0),
.B(n_2),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_2),
.A2(n_22),
.B1(n_26),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_2),
.A2(n_34),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_2),
.A2(n_34),
.B1(n_53),
.B2(n_56),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_34),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_2),
.A2(n_60),
.B(n_204),
.C(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_2),
.B(n_58),
.Y(n_220)
);

O2A1O1Ixp33_ASAP7_75t_L g230 ( 
.A1(n_2),
.A2(n_38),
.B(n_44),
.C(n_231),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_2),
.B(n_24),
.C(n_28),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_2),
.B(n_98),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_2),
.B(n_27),
.Y(n_275)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_5),
.A2(n_50),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_5),
.A2(n_22),
.B1(n_26),
.B2(n_50),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_50),
.Y(n_136)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_7),
.A2(n_53),
.B1(n_54),
.B2(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_7),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_7),
.A2(n_43),
.B1(n_44),
.B2(n_146),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_7),
.A2(n_22),
.B1(n_26),
.B2(n_146),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_146),
.Y(n_260)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_11),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_11),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_11),
.A2(n_43),
.B1(n_44),
.B2(n_55),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_11),
.A2(n_22),
.B1(n_26),
.B2(n_55),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_55),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_92),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_90),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_77),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_15),
.B(n_77),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_17),
.B1(n_68),
.B2(n_76),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_35),
.C(n_51),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_18),
.A2(n_35),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_18),
.A2(n_81),
.B1(n_86),
.B2(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_18),
.A2(n_81),
.B1(n_188),
.B2(n_216),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_31),
.B(n_32),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_19),
.A2(n_117),
.B(n_118),
.Y(n_116)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_20),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_20),
.B(n_33),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_20),
.B(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_27),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_21)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_22),
.A2(n_26),
.B1(n_38),
.B2(n_40),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_22),
.B(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_23),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp33_ASAP7_75t_L g231 ( 
.A1(n_26),
.A2(n_34),
.B(n_40),
.Y(n_231)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_27),
.B(n_103),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_27),
.B(n_235),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_28),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_28),
.B(n_271),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_31),
.B(n_32),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_31),
.A2(n_102),
.B(n_117),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

OAI21xp33_ASAP7_75t_L g204 ( 
.A1(n_34),
.A2(n_44),
.B(n_59),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_35),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_46),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_36),
.B(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_41),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_48),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_37),
.A2(n_41),
.B(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_37),
.B(n_49),
.Y(n_89)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_42),
.B(n_87),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_44),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx6p67_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_46),
.A2(n_88),
.B(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_46),
.B(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_49),
.Y(n_46)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_47),
.B(n_198),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_58),
.B(n_61),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_52),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_53),
.A2(n_54),
.B1(n_59),
.B2(n_60),
.Y(n_64)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_53),
.Y(n_205)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_65),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_58),
.B(n_84),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_58),
.B(n_145),
.Y(n_174)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_62),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_63),
.B(n_145),
.Y(n_144)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_74),
.B2(n_75),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_69),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_69),
.B(n_164),
.C(n_173),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_69),
.A2(n_74),
.B1(n_173),
.B2(n_304),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_70),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_72),
.B(n_73),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_71),
.A2(n_121),
.B(n_122),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_73),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_73),
.B(n_144),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_82),
.C(n_85),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_78),
.A2(n_82),
.B1(n_107),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_78),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_82),
.C(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_81),
.B(n_186),
.C(n_188),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_105),
.B1(n_107),
.B2(n_108),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_83),
.B(n_174),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_85),
.B(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B(n_89),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_89),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_89),
.B(n_197),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI211xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_147),
.B(n_153),
.C(n_315),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_123),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_94),
.B(n_123),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_109),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_104),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_96),
.A2(n_97),
.B(n_99),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_96),
.B(n_104),
.C(n_109),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_98),
.B(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_100),
.B(n_233),
.Y(n_232)
);

INVxp33_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_102),
.B(n_245),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_105),
.Y(n_108)
);

AOI21xp33_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_115),
.B(n_119),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_110),
.A2(n_119),
.B1(n_120),
.B2(n_127),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_110),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_110),
.A2(n_116),
.B1(n_127),
.B2(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_110),
.B(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_110),
.A2(n_127),
.B1(n_230),
.B2(n_287),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_113),
.B(n_114),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_111),
.A2(n_167),
.B(n_168),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_111),
.B(n_114),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_111),
.B(n_259),
.Y(n_258)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_116),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_118),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_118),
.B(n_234),
.Y(n_253)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.C(n_129),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_124),
.A2(n_125),
.B1(n_128),
.B2(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_128),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_138),
.C(n_141),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_137),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_131),
.B(n_137),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_132),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_133),
.B(n_260),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_135),
.A2(n_167),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_135),
.B(n_265),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_138),
.A2(n_141),
.B1(n_142),
.B2(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_140),
.B(n_190),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NAND3xp33_ASAP7_75t_SL g153 ( 
.A(n_148),
.B(n_154),
.C(n_155),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_149),
.B(n_150),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_178),
.B(n_314),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_175),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_157),
.B(n_175),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.C(n_163),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_158),
.B(n_161),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_163),
.B(n_312),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_164),
.A2(n_165),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_171),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_171),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_169),
.B(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_169),
.B(n_258),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_172),
.B(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_173),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_309),
.B(n_313),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_223),
.B(n_296),
.C(n_308),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_211),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_181),
.B(n_211),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_194),
.B2(n_210),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_192),
.B2(n_193),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_184),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_184),
.B(n_193),
.C(n_210),
.Y(n_297)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_185),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_187),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_188),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

INVxp67_ASAP7_75t_SL g198 ( 
.A(n_191),
.Y(n_198)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_202),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_195)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_196),
.B(n_201),
.C(n_202),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_199),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_206),
.Y(n_217)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_217),
.C(n_218),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_212),
.A2(n_213),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_218),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.C(n_221),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_228),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_221),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_222),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_295),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_239),
.B(n_294),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_236),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_226),
.B(n_236),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.C(n_232),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_227),
.B(n_292),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_229),
.B(n_232),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_230),
.Y(n_287)
);

INVxp33_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_289),
.B(n_293),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_280),
.B(n_288),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_262),
.B(n_279),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_249),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_243),
.B(n_249),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_244),
.A2(n_246),
.B1(n_247),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_244),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_256),
.B2(n_261),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_252),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_255),
.C(n_261),
.Y(n_281)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_253),
.Y(n_255)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_256),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_268),
.B(n_278),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_264),
.B(n_266),
.Y(n_278)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_265),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_274),
.B(n_277),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_272),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_275),
.B(n_276),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_281),
.B(n_282),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_286),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_285),
.C(n_286),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_290),
.B(n_291),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_297),
.B(n_298),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_307),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_305),
.B2(n_306),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_306),
.C(n_307),
.Y(n_310)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_310),
.B(n_311),
.Y(n_313)
);


endmodule