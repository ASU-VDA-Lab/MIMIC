module fake_jpeg_814_n_218 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_218);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_218;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_5),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_41),
.B(n_5),
.Y(n_67)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_29),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_27),
.Y(n_71)
);

INVx11_ASAP7_75t_SL g72 ( 
.A(n_15),
.Y(n_72)
);

INVx8_ASAP7_75t_SL g73 ( 
.A(n_37),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_52),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_1),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_42),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_4),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_1),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_44),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_58),
.B(n_2),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_81),
.B(n_77),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_61),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_76),
.B1(n_63),
.B2(n_68),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_77),
.B1(n_75),
.B2(n_80),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g107 ( 
.A(n_91),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_67),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_99),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_88),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_94),
.B(n_96),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_67),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_85),
.A2(n_68),
.B1(n_76),
.B2(n_79),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_101),
.A2(n_82),
.B1(n_61),
.B2(n_74),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_91),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_110),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_59),
.Y(n_108)
);

NOR3xp33_ASAP7_75t_SL g124 ( 
.A(n_108),
.B(n_117),
.C(n_119),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_60),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_71),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_113),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_70),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_116),
.A2(n_120),
.B1(n_101),
.B2(n_75),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_62),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

AOI21xp33_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_73),
.B(n_69),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_66),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_128),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_106),
.A2(n_112),
.B(n_108),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_115),
.A2(n_69),
.B(n_86),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_107),
.A2(n_88),
.B1(n_78),
.B2(n_61),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_134),
.B1(n_141),
.B2(n_23),
.Y(n_150)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_78),
.B1(n_64),
.B2(n_82),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_114),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_138),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_103),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_109),
.A2(n_64),
.B1(n_82),
.B2(n_97),
.Y(n_141)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_142),
.Y(n_157)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_133),
.A2(n_132),
.B1(n_124),
.B2(n_130),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_150),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_124),
.B(n_56),
.Y(n_149)
);

MAJx2_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_31),
.C(n_50),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_140),
.B(n_129),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_158),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_133),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_154),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_127),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_154)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_25),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_11),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_139),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_162),
.Y(n_182)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_8),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_164),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_9),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_125),
.B(n_10),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_165),
.A2(n_12),
.B(n_13),
.Y(n_175)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_166),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_169),
.B(n_175),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_144),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_172),
.A2(n_180),
.B1(n_163),
.B2(n_157),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

MAJx2_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_30),
.C(n_49),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_14),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_161),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_176),
.B(n_178),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_147),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_155),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_183),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_184),
.A2(n_177),
.B1(n_172),
.B2(n_16),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_168),
.A2(n_144),
.B1(n_145),
.B2(n_151),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_185),
.A2(n_189),
.B1(n_191),
.B2(n_192),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_168),
.A2(n_145),
.B1(n_151),
.B2(n_33),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_170),
.A2(n_26),
.B(n_48),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_24),
.B(n_47),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_194),
.B(n_169),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_181),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_196),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_167),
.C(n_173),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_198),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_190),
.Y(n_199)
);

NOR2xp67_ASAP7_75t_SL g206 ( 
.A(n_199),
.B(n_200),
.Y(n_206)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_174),
.C(n_171),
.Y(n_201)
);

MAJx2_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_186),
.C(n_194),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_202),
.B(n_177),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_201),
.C(n_195),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_207),
.B(n_189),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_197),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_208),
.B(n_209),
.Y(n_211)
);

AOI21x1_ASAP7_75t_L g212 ( 
.A1(n_211),
.A2(n_206),
.B(n_203),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_212),
.A2(n_210),
.B(n_32),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_22),
.C(n_46),
.Y(n_214)
);

OA22x2_ASAP7_75t_L g215 ( 
.A1(n_214),
.A2(n_21),
.B1(n_45),
.B2(n_35),
.Y(n_215)
);

AOI21x1_ASAP7_75t_L g216 ( 
.A1(n_215),
.A2(n_19),
.B(n_20),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_34),
.C(n_54),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_16),
.Y(n_218)
);


endmodule