module real_jpeg_2944_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_244;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

INVx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_1),
.B(n_55),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_1),
.B(n_30),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_1),
.B(n_53),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_1),
.B(n_28),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_1),
.B(n_48),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_2),
.B(n_30),
.Y(n_68)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_2),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_2),
.B(n_63),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_4),
.B(n_34),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_4),
.B(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_4),
.B(n_55),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_4),
.B(n_38),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_4),
.B(n_53),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_4),
.B(n_30),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_4),
.B(n_28),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_4),
.B(n_48),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_5),
.B(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_5),
.B(n_34),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_5),
.B(n_63),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_5),
.B(n_55),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_8),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_8),
.B(n_38),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_8),
.B(n_63),
.Y(n_91)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_8),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_8),
.B(n_55),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_8),
.B(n_53),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_9),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_9),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_9),
.B(n_55),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_9),
.B(n_28),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_9),
.B(n_63),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_9),
.B(n_34),
.Y(n_277)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_11),
.B(n_28),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_11),
.B(n_30),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_11),
.B(n_53),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_11),
.B(n_55),
.Y(n_265)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_14),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_14),
.B(n_53),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_14),
.B(n_63),
.Y(n_111)
);

AND2x2_ASAP7_75t_SL g153 ( 
.A(n_14),
.B(n_30),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_14),
.B(n_34),
.Y(n_240)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_14),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_248),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_245),
.Y(n_17)
);

INVxp33_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_208),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_130),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_94),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_22),
.B(n_94),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_58),
.C(n_83),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_23),
.B(n_205),
.Y(n_204)
);

BUFx24_ASAP7_75t_SL g285 ( 
.A(n_23),
.Y(n_285)
);

FAx1_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_40),
.CI(n_44),
.CON(n_23),
.SN(n_23)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_24),
.B(n_40),
.C(n_44),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_33),
.C(n_37),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_25),
.A2(n_26),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_26),
.A2(n_76),
.B(n_148),
.C(n_227),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_27),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_27),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_27),
.A2(n_29),
.B1(n_76),
.B2(n_148),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_27),
.A2(n_148),
.B1(n_152),
.B2(n_153),
.Y(n_256)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_29),
.A2(n_73),
.B1(n_76),
.B2(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_31),
.B(n_129),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_33),
.B(n_37),
.Y(n_201)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_34),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_SL g221 ( 
.A(n_38),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B(n_43),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_42),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_43),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_43),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_50),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_45),
.B(n_52),
.C(n_54),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_46),
.B(n_74),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_46),
.B(n_105),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_47),
.B(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_57),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_51),
.A2(n_52),
.B1(n_264),
.B2(n_267),
.Y(n_263)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_55),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_58),
.B(n_83),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_70),
.B2(n_82),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_71),
.C(n_78),
.Y(n_96)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_65),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_61),
.B(n_67),
.C(n_69),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_64),
.B(n_221),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_66),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_77),
.B2(n_78),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_75),
.B(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.C(n_81),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_79),
.A2(n_81),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_79),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_88),
.C(n_92),
.Y(n_83)
);

FAx1_ASAP7_75t_SL g195 ( 
.A(n_84),
.B(n_88),
.CI(n_92),
.CON(n_195),
.SN(n_195)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.C(n_91),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_89),
.B(n_91),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_90),
.B(n_141),
.Y(n_140)
);

BUFx24_ASAP7_75t_SL g288 ( 
.A(n_94),
.Y(n_288)
);

FAx1_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_116),
.CI(n_117),
.CON(n_94),
.SN(n_94)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_95),
.B(n_116),
.C(n_117),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_96),
.B(n_99),
.C(n_106),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_106),
.B2(n_107),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_100),
.B(n_102),
.C(n_104),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_114),
.B2(n_115),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_111),
.B(n_112),
.C(n_114),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_112),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_114),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.Y(n_117)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_119),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_119),
.B(n_120),
.C(n_122),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_128),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_124),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_127),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_124),
.B(n_126),
.C(n_128),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_203),
.B(n_207),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_191),
.B(n_202),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_163),
.B(n_190),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_154),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_134),
.B(n_154),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_144),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_140),
.B1(n_142),
.B2(n_143),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_136),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.C(n_139),
.Y(n_136)
);

FAx1_ASAP7_75t_SL g155 ( 
.A(n_137),
.B(n_138),
.CI(n_139),
.CON(n_155),
.SN(n_155)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_140),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_140),
.B(n_142),
.C(n_144),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_149),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_145),
.B(n_150),
.C(n_151),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.C(n_162),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_187),
.Y(n_186)
);

BUFx24_ASAP7_75t_SL g289 ( 
.A(n_155),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_156),
.A2(n_157),
.B1(n_162),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_184),
.B(n_189),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_175),
.B(n_183),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_171),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_171),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_169),
.C(n_170),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_172),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_178),
.B(n_182),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_180),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_186),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_192),
.B(n_193),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_198),
.C(n_199),
.Y(n_206)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx24_ASAP7_75t_SL g290 ( 
.A(n_195),
.Y(n_290)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_204),
.B(n_206),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_209),
.A2(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_244),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_244),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_211),
.B(n_213),
.C(n_229),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_228),
.B2(n_229),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx24_ASAP7_75t_SL g287 ( 
.A(n_214),
.Y(n_287)
);

FAx1_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_224),
.CI(n_225),
.CON(n_214),
.SN(n_214)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_215),
.B(n_224),
.C(n_225),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_216),
.B(n_220),
.C(n_222),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_222),
.B2(n_223),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_221),
.B(n_258),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_222),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_234),
.C(n_235),
.Y(n_251)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_242),
.B2(n_243),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_240),
.C(n_242),
.Y(n_272)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_240),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_283),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_282),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_250),
.B(n_282),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_268),
.B2(n_281),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_261),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_259),
.B2(n_260),
.Y(n_255)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_256),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_257),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_264),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_268),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_280),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_271),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_279),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_276),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_277),
.Y(n_279)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);


endmodule