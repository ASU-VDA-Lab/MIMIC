module fake_jpeg_5743_n_10 (n_3, n_2, n_1, n_0, n_4, n_10);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_10;

wire n_8;
wire n_9;
wire n_6;
wire n_5;
wire n_7;

INVx5_ASAP7_75t_L g5 ( 
.A(n_3),
.Y(n_5)
);

INVx1_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

AOI21xp5_ASAP7_75t_SL g7 ( 
.A1(n_5),
.A2(n_0),
.B(n_1),
.Y(n_7)
);

CKINVDCx14_ASAP7_75t_R g8 ( 
.A(n_7),
.Y(n_8)
);

AOI21x1_ASAP7_75t_L g9 ( 
.A1(n_8),
.A2(n_5),
.B(n_6),
.Y(n_9)
);

A2O1A1O1Ixp25_ASAP7_75t_L g10 ( 
.A1(n_9),
.A2(n_0),
.B(n_1),
.C(n_2),
.D(n_8),
.Y(n_10)
);


endmodule