module fake_jpeg_15519_n_109 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_109);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_109;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_21),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_24),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_23),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_37),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_29),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_14),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_48),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_44),
.Y(n_69)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_63),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_63),
.A2(n_45),
.B1(n_46),
.B2(n_52),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_65),
.A2(n_67),
.B(n_1),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_58),
.A2(n_46),
.B1(n_53),
.B2(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_41),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_0),
.Y(n_70)
);

AO22x1_ASAP7_75t_L g86 ( 
.A1(n_70),
.A2(n_43),
.B1(n_50),
.B2(n_8),
.Y(n_86)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_74),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_77),
.A2(n_82),
.B1(n_78),
.B2(n_75),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_79),
.A2(n_84),
.B(n_85),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_72),
.B(n_42),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_83),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_72),
.C(n_38),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_87),
.A2(n_89),
.B1(n_88),
.B2(n_71),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_81),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_92),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_93),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_94),
.A2(n_66),
.B1(n_7),
.B2(n_9),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_95),
.B(n_10),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_6),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_16),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_17),
.B(n_18),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_102),
.B(n_19),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_103),
.B(n_20),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_105),
.A2(n_99),
.B(n_26),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_25),
.B(n_27),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_32),
.B(n_33),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_34),
.Y(n_109)
);


endmodule