module real_jpeg_19403_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_0),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_1),
.A2(n_37),
.B1(n_38),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_1),
.A2(n_27),
.B1(n_29),
.B2(n_45),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_2),
.A2(n_27),
.B1(n_29),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_4),
.Y(n_65)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_6),
.A2(n_37),
.B1(n_38),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_6),
.A2(n_27),
.B1(n_29),
.B2(n_43),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_8),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_8),
.B(n_70),
.Y(n_106)
);

AOI21xp33_ASAP7_75t_L g128 ( 
.A1(n_8),
.A2(n_27),
.B(n_39),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_8),
.A2(n_37),
.B1(n_38),
.B2(n_66),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_8),
.A2(n_25),
.B1(n_31),
.B2(n_136),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_8),
.B(n_105),
.Y(n_149)
);

AOI21xp33_ASAP7_75t_L g166 ( 
.A1(n_8),
.A2(n_59),
.B(n_167),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_9),
.A2(n_54),
.B1(n_59),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_9),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_9),
.A2(n_27),
.B1(n_29),
.B2(n_62),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_9),
.A2(n_37),
.B1(n_38),
.B2(n_62),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_10),
.A2(n_65),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_10),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_10),
.A2(n_54),
.B1(n_59),
.B2(n_73),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_10),
.A2(n_37),
.B1(n_38),
.B2(n_73),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_10),
.A2(n_27),
.B1(n_29),
.B2(n_73),
.Y(n_136)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_12),
.A2(n_54),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_12),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_12),
.A2(n_60),
.B1(n_65),
.B2(n_74),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_12),
.A2(n_27),
.B1(n_29),
.B2(n_60),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_12),
.A2(n_37),
.B1(n_38),
.B2(n_60),
.Y(n_152)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_13),
.A2(n_37),
.B1(n_38),
.B2(n_55),
.Y(n_57)
);

OAI32xp33_ASAP7_75t_L g161 ( 
.A1(n_13),
.A2(n_38),
.A3(n_59),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_14),
.A2(n_37),
.B1(n_38),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_14),
.A2(n_50),
.B1(n_54),
.B2(n_59),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_14),
.A2(n_27),
.B1(n_29),
.B2(n_50),
.Y(n_154)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx3_ASAP7_75t_SL g38 ( 
.A(n_16),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_112),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_110),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_93),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_21),
.B(n_93),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_75),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_46),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_34),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_25),
.A2(n_28),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_25),
.A2(n_26),
.B1(n_90),
.B2(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_25),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_25),
.A2(n_91),
.B1(n_121),
.B2(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_25),
.A2(n_31),
.B1(n_124),
.B2(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_25),
.A2(n_91),
.B1(n_109),
.B2(n_154),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_27),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_27),
.A2(n_29),
.B1(n_39),
.B2(n_40),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_29),
.B(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_31),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_31),
.B(n_66),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_41),
.B1(n_42),
.B2(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_35),
.A2(n_41),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_35),
.A2(n_41),
.B1(n_132),
.B2(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_35),
.A2(n_41),
.B1(n_152),
.B2(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_35),
.A2(n_41),
.B1(n_49),
.B2(n_170),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_41),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_37),
.B(n_55),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_38),
.A2(n_40),
.B(n_66),
.C(n_128),
.Y(n_127)
);

CKINVDCx9p33_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_41),
.B(n_66),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_51),
.C(n_63),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_47),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_57),
.B1(n_58),
.B2(n_61),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_53),
.A2(n_57),
.B1(n_61),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_53),
.A2(n_57),
.B1(n_102),
.B2(n_166),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B(n_56),
.C(n_57),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_55),
.Y(n_56)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_59),
.B1(n_68),
.B2(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_64),
.B1(n_69),
.B2(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_54),
.B(n_66),
.Y(n_163)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_68),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_63),
.B(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_67),
.B1(n_70),
.B2(n_72),
.Y(n_63)
);

HAxp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_66),
.CON(n_64),
.SN(n_64)
);

O2A1O1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_65),
.A2(n_68),
.B(n_69),
.C(n_70),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_68),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_65),
.Y(n_74)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_72),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_86),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_83),
.B2(n_85),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_83),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_89),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_89),
.Y(n_97)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.C(n_98),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_94),
.B(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_106),
.C(n_107),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_100),
.B(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_106),
.A2(n_107),
.B1(n_108),
.B2(n_181),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_106),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_189),
.B(n_193),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_175),
.B(n_188),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_156),
.B(n_174),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_144),
.B(n_155),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_133),
.B(n_143),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_125),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_125),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_129),
.B2(n_130),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_129),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_138),
.B(n_142),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_137),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_146),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_153),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_151),
.C(n_153),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_158),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_164),
.B1(n_172),
.B2(n_173),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_159),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_161),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_163),
.Y(n_167)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_168),
.B1(n_169),
.B2(n_171),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_165),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_171),
.C(n_172),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_176),
.B(n_177),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_182),
.B2(n_183),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_185),
.C(n_186),
.Y(n_190)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_184),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_185),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_190),
.B(n_191),
.Y(n_193)
);


endmodule