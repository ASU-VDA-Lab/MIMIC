module real_jpeg_11939_n_16 (n_5, n_4, n_8, n_0, n_12, n_309, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_309;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;

BUFx2_ASAP7_75t_L g86 ( 
.A(n_0),
.Y(n_86)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_4),
.A2(n_62),
.B1(n_63),
.B2(n_66),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_4),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_4),
.A2(n_28),
.B1(n_30),
.B2(n_66),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_4),
.A2(n_35),
.B1(n_37),
.B2(n_66),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_4),
.A2(n_48),
.B1(n_52),
.B2(n_66),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_5),
.A2(n_62),
.B1(n_63),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_5),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_5),
.A2(n_28),
.B1(n_30),
.B2(n_165),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_5),
.A2(n_35),
.B1(n_37),
.B2(n_165),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_5),
.A2(n_48),
.B1(n_52),
.B2(n_165),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_6),
.A2(n_29),
.B1(n_35),
.B2(n_37),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_6),
.A2(n_29),
.B1(n_62),
.B2(n_63),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_6),
.A2(n_29),
.B1(n_48),
.B2(n_52),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_8),
.A2(n_35),
.B1(n_37),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_8),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_8),
.A2(n_48),
.B1(n_52),
.B2(n_56),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_8),
.A2(n_56),
.B1(n_62),
.B2(n_63),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_8),
.A2(n_28),
.B1(n_30),
.B2(n_56),
.Y(n_112)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

O2A1O1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_10),
.A2(n_59),
.B(n_62),
.C(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_10),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_10),
.A2(n_62),
.B1(n_63),
.B2(n_179),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_10),
.B(n_101),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_10),
.A2(n_35),
.B1(n_37),
.B2(n_179),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_10),
.A2(n_84),
.B1(n_87),
.B2(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_10),
.B(n_81),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_11),
.A2(n_62),
.B1(n_63),
.B2(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_11),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_11),
.A2(n_28),
.B1(n_30),
.B2(n_186),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_11),
.A2(n_35),
.B1(n_37),
.B2(n_186),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_11),
.A2(n_48),
.B1(n_52),
.B2(n_186),
.Y(n_265)
);

BUFx8_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_13),
.A2(n_28),
.B1(n_30),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_13),
.A2(n_43),
.B1(n_62),
.B2(n_63),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_13),
.A2(n_35),
.B1(n_37),
.B2(n_43),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_13),
.A2(n_43),
.B1(n_48),
.B2(n_52),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_14),
.A2(n_62),
.B1(n_63),
.B2(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_14),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_14),
.A2(n_28),
.B1(n_30),
.B2(n_140),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_14),
.A2(n_35),
.B1(n_37),
.B2(n_140),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_14),
.A2(n_48),
.B1(n_52),
.B2(n_140),
.Y(n_259)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_118),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_117),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_102),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_20),
.B(n_102),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_72),
.C(n_82),
.Y(n_20)
);

FAx1_ASAP7_75t_SL g304 ( 
.A(n_21),
.B(n_72),
.CI(n_82),
.CON(n_304),
.SN(n_304)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_57),
.B2(n_71),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_44),
.B2(n_45),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_24),
.B(n_45),
.C(n_57),
.Y(n_103)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B(n_40),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_27),
.A2(n_32),
.B1(n_79),
.B2(n_81),
.Y(n_78)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_28),
.A2(n_30),
.B1(n_34),
.B2(n_38),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_28),
.A2(n_30),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

HAxp5_ASAP7_75t_SL g228 ( 
.A(n_28),
.B(n_179),
.CON(n_228),
.SN(n_228)
);

OAI21xp33_ASAP7_75t_L g178 ( 
.A1(n_30),
.A2(n_60),
.B(n_179),
.Y(n_178)
);

NOR3xp33_ASAP7_75t_L g229 ( 
.A(n_30),
.B(n_35),
.C(n_38),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_31),
.A2(n_111),
.B(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_31),
.A2(n_33),
.B1(n_214),
.B2(n_216),
.Y(n_213)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_32),
.B(n_114),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_32),
.A2(n_41),
.B(n_112),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_32),
.A2(n_81),
.B1(n_182),
.B2(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_32),
.A2(n_81),
.B1(n_215),
.B2(n_228),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_39),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_33),
.A2(n_80),
.B(n_113),
.Y(n_136)
);

OA22x2_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_33)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_SL g226 ( 
.A1(n_34),
.A2(n_37),
.B(n_227),
.C(n_229),
.Y(n_226)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_35),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_37),
.B1(n_50),
.B2(n_51),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_37),
.B(n_249),
.Y(n_248)
);

INVxp33_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_42),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_44),
.A2(n_45),
.B1(n_110),
.B2(n_115),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_53),
.B(n_55),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_55),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_46),
.A2(n_53),
.B1(n_93),
.B2(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_46),
.A2(n_53),
.B1(n_234),
.B2(n_242),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_46),
.A2(n_53),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_46),
.A2(n_53),
.B1(n_242),
.B2(n_252),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_47),
.B(n_77),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_47),
.A2(n_75),
.B(n_135),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_47),
.B(n_179),
.Y(n_268)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_47)
);

CKINVDCx6p67_ASAP7_75t_R g52 ( 
.A(n_48),
.Y(n_52)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_50),
.B(n_52),
.C(n_179),
.Y(n_249)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_52),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_53),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_53),
.A2(n_55),
.B(n_94),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_53),
.Y(n_232)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_57),
.A2(n_71),
.B1(n_105),
.B2(n_116),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_61),
.B(n_67),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_58),
.A2(n_97),
.B1(n_184),
.B2(n_187),
.Y(n_183)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_61),
.Y(n_107)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_68),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_68),
.A2(n_101),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_68),
.A2(n_101),
.B1(n_139),
.B2(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_68),
.A2(n_101),
.B1(n_185),
.B2(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_72),
.A2(n_73),
.B(n_78),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_78),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_74),
.A2(n_232),
.B(n_233),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_112),
.Y(n_111)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_90),
.B(n_95),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_83),
.A2(n_95),
.B1(n_96),
.B2(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_83),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_83),
.A2(n_91),
.B1(n_92),
.B2(n_146),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_87),
.B(n_88),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_84),
.A2(n_157),
.B(n_159),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_84),
.A2(n_87),
.B1(n_257),
.B2(n_265),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_84),
.A2(n_128),
.B(n_259),
.Y(n_274)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_85),
.B(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_85),
.A2(n_86),
.B1(n_158),
.B2(n_175),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_85),
.A2(n_89),
.B(n_160),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_85),
.A2(n_86),
.B1(n_256),
.B2(n_258),
.Y(n_255)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_89),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_87),
.B(n_131),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_87),
.A2(n_129),
.B(n_176),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_87),
.B(n_179),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_90),
.B(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_98),
.B(n_100),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_97),
.A2(n_138),
.B(n_141),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_99),
.B(n_101),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_109),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_110),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_113),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_301),
.B(n_305),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_166),
.B(n_300),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_148),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_121),
.B(n_148),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_142),
.B2(n_147),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_122),
.B(n_143),
.C(n_144),
.Y(n_303)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_136),
.C(n_137),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_124),
.A2(n_125),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_132),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_126),
.A2(n_127),
.B1(n_132),
.B2(n_133),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_137),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_142),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_153),
.C(n_154),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_149),
.A2(n_150),
.B1(n_153),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_153),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_154),
.B(n_297),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_162),
.C(n_163),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_161),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_156),
.B(n_161),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_163),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_164),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_294),
.B(n_299),
.Y(n_166)
);

AOI221xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_203),
.B1(n_219),
.B2(n_293),
.C(n_309),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_192),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_169),
.B(n_192),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_188),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_170),
.B(n_189),
.C(n_190),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_180),
.C(n_183),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_171),
.A2(n_172),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_177),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_173),
.A2(n_174),
.B1(n_177),
.B2(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_177),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_180),
.B(n_183),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_196),
.C(n_202),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_202),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.C(n_200),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_198),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_199),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_206),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_217),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_204),
.B(n_217),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.C(n_209),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_205),
.B(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_207),
.B(n_209),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.C(n_213),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_213),
.B(n_236),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_292),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_287),
.B(n_291),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_243),
.B(n_286),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_238),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_223),
.B(n_238),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_235),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_231),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_225),
.B(n_231),
.C(n_235),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_230),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_226),
.B(n_230),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.C(n_241),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_239),
.B(n_283),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_240),
.B(n_241),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_281),
.B(n_285),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_271),
.B(n_280),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_260),
.B(n_270),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_255),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_255),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_250),
.B1(n_253),
.B2(n_254),
.Y(n_247)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_248),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_250),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_253),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_266),
.B(n_269),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_268),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_273),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_276),
.C(n_279),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_279),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_278),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_284),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_290),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_290),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_296),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_304),
.Y(n_306)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_304),
.Y(n_308)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);


endmodule