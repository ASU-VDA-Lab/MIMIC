module fake_jpeg_8805_n_235 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_235);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_235;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_34),
.B(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_44),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_27),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_21),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_33),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_41),
.C(n_35),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_40),
.C(n_38),
.Y(n_71)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_25),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_53),
.B(n_55),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_30),
.B1(n_27),
.B2(n_29),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_54),
.A2(n_56),
.B(n_22),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_36),
.A2(n_30),
.B1(n_29),
.B2(n_26),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_35),
.B(n_18),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_58),
.B(n_62),
.Y(n_83)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

CKINVDCx6p67_ASAP7_75t_R g84 ( 
.A(n_59),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_61),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_71),
.Y(n_92)
);

NAND2xp33_ASAP7_75t_SL g68 ( 
.A(n_49),
.B(n_22),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_68),
.A2(n_76),
.B(n_80),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_45),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_69),
.B(n_81),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_31),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_70),
.B(n_75),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_29),
.B1(n_21),
.B2(n_26),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_74),
.A2(n_24),
.B1(n_28),
.B2(n_48),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_62),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_51),
.A2(n_38),
.B1(n_19),
.B2(n_18),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_51),
.A2(n_19),
.B1(n_28),
.B2(n_24),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_40),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_65),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_L g87 ( 
.A1(n_52),
.A2(n_16),
.B(n_25),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_13),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_46),
.B(n_31),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_22),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_89),
.B(n_93),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_86),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_96),
.Y(n_129)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_86),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_97),
.B(n_98),
.Y(n_128)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

INVxp67_ASAP7_75t_SL g127 ( 
.A(n_99),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_100),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_79),
.B1(n_59),
.B2(n_61),
.Y(n_101)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_102),
.Y(n_126)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_105),
.Y(n_113)
);

AO22x1_ASAP7_75t_SL g106 ( 
.A1(n_68),
.A2(n_20),
.B1(n_32),
.B2(n_65),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_SL g131 ( 
.A1(n_106),
.A2(n_55),
.B(n_72),
.C(n_43),
.Y(n_131)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_82),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_111),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_70),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_97),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_115),
.B(n_117),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_91),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_119),
.A2(n_107),
.B(n_112),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_104),
.A2(n_71),
.B(n_73),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_134),
.B(n_43),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_72),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_130),
.B(n_132),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_131),
.A2(n_67),
.B1(n_64),
.B2(n_94),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_95),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_85),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_133),
.B(n_100),
.Y(n_147)
);

AND2x2_ASAP7_75t_SL g134 ( 
.A(n_106),
.B(n_57),
.Y(n_134)
);

OAI22x1_ASAP7_75t_L g135 ( 
.A1(n_131),
.A2(n_106),
.B1(n_103),
.B2(n_104),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_135),
.A2(n_136),
.B1(n_138),
.B2(n_131),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_115),
.B1(n_123),
.B2(n_101),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_133),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_137),
.B(n_140),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_103),
.B1(n_108),
.B2(n_99),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_130),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_147),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_141),
.B(n_142),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_116),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_132),
.A2(n_82),
.B1(n_93),
.B2(n_109),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_143),
.A2(n_154),
.B1(n_126),
.B2(n_113),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_144),
.B(n_149),
.Y(n_158)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_150),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_129),
.B(n_33),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_116),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_50),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_156),
.C(n_134),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_117),
.B(n_14),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_153),
.Y(n_168)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_124),
.B(n_110),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_124),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_128),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_135),
.B1(n_137),
.B2(n_122),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_167),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_131),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_169),
.C(n_172),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_113),
.Y(n_165)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_171),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_156),
.B(n_119),
.Y(n_169)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_170),
.Y(n_178)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_131),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_120),
.Y(n_173)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_173),
.Y(n_189)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_174),
.B(n_1),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_120),
.C(n_125),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_114),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_171),
.Y(n_176)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_176),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_160),
.Y(n_179)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_180),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_164),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_181),
.A2(n_187),
.B(n_191),
.Y(n_198)
);

XNOR2x1_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_149),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_158),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_1),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_161),
.A2(n_114),
.B1(n_94),
.B2(n_67),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_186),
.A2(n_190),
.B1(n_32),
.B2(n_3),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_175),
.A2(n_64),
.B1(n_44),
.B2(n_78),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_202),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_169),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_200),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_163),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_195),
.A2(n_187),
.B(n_178),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_197),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_162),
.C(n_172),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_168),
.C(n_33),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_66),
.C(n_44),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_203),
.Y(n_205)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_206),
.Y(n_218)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_198),
.Y(n_209)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_209),
.Y(n_219)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_210),
.A2(n_212),
.B1(n_186),
.B2(n_194),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_184),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_208),
.C(n_207),
.Y(n_214)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_199),
.Y(n_212)
);

NOR2x1_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_201),
.Y(n_213)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_213),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_215),
.C(n_208),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_202),
.Y(n_215)
);

NOR2xp67_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_189),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_216),
.A2(n_217),
.B(n_194),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_223),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_222),
.A2(n_213),
.B(n_219),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_176),
.C(n_211),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_196),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_224),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_2),
.C(n_4),
.Y(n_230)
);

AOI31xp67_ASAP7_75t_L g227 ( 
.A1(n_220),
.A2(n_183),
.A3(n_190),
.B(n_215),
.Y(n_227)
);

AOI322xp5_ASAP7_75t_L g229 ( 
.A1(n_227),
.A2(n_8),
.A3(n_13),
.B1(n_10),
.B2(n_9),
.C1(n_2),
.C2(n_6),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_229),
.B(n_230),
.Y(n_231)
);

AO221x1_ASAP7_75t_L g232 ( 
.A1(n_229),
.A2(n_226),
.B1(n_228),
.B2(n_32),
.C(n_6),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_232),
.A2(n_231),
.B1(n_4),
.B2(n_5),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_233),
.A2(n_2),
.B(n_4),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_234),
.B(n_5),
.Y(n_235)
);


endmodule