module fake_jpeg_23475_n_165 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_165);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_31),
.B(n_33),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_1),
.Y(n_33)
);

CKINVDCx9p33_ASAP7_75t_R g34 ( 
.A(n_19),
.Y(n_34)
);

INVx5_ASAP7_75t_SL g50 ( 
.A(n_34),
.Y(n_50)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_43),
.Y(n_53)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_20),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_1),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_16),
.B1(n_14),
.B2(n_25),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_46),
.A2(n_55),
.B1(n_65),
.B2(n_28),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_59),
.Y(n_73)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_32),
.A2(n_28),
.B1(n_16),
.B2(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_38),
.B(n_24),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_57),
.B(n_61),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_14),
.B1(n_24),
.B2(n_22),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_32),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_67),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_36),
.B(n_22),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_29),
.Y(n_64)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

AO22x1_ASAP7_75t_L g65 ( 
.A1(n_36),
.A2(n_17),
.B1(n_23),
.B2(n_18),
.Y(n_65)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_29),
.Y(n_68)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_71),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_39),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_28),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_76),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_79),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_53),
.B(n_39),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_52),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_46),
.B1(n_34),
.B2(n_70),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_45),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_81),
.B(n_87),
.Y(n_98)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_20),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_84),
.B(n_85),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_25),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_20),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_45),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_47),
.B(n_20),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_91),
.B(n_92),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_2),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_49),
.B(n_2),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_66),
.C(n_3),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_94),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_95),
.A2(n_99),
.B1(n_110),
.B2(n_75),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_70),
.B1(n_62),
.B2(n_51),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_106),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_66),
.C(n_55),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_101),
.A2(n_108),
.B(n_112),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_82),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_104),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

MAJx2_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_55),
.C(n_23),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_81),
.A2(n_51),
.B1(n_55),
.B2(n_63),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_79),
.C(n_74),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_93),
.B(n_88),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_113),
.A2(n_114),
.B(n_116),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_74),
.B(n_78),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_117),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_101),
.A2(n_78),
.B(n_89),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_89),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_120),
.Y(n_134)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_108),
.A2(n_97),
.B1(n_110),
.B2(n_106),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_123),
.A2(n_100),
.B1(n_103),
.B2(n_63),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_125),
.A2(n_126),
.B1(n_67),
.B2(n_102),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_85),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_127),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_128),
.A2(n_129),
.B(n_136),
.Y(n_143)
);

NOR2xp67_ASAP7_75t_SL g129 ( 
.A(n_114),
.B(n_85),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_131),
.A2(n_126),
.B1(n_40),
.B2(n_90),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_124),
.A2(n_83),
.B1(n_107),
.B2(n_23),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_133),
.A2(n_120),
.B1(n_121),
.B2(n_30),
.Y(n_144)
);

NAND3xp33_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_3),
.C(n_4),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_4),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_138),
.A2(n_136),
.B1(n_113),
.B2(n_125),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_130),
.B(n_118),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_141),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_122),
.C(n_116),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_142),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_122),
.C(n_115),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_145),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_134),
.B(n_4),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_146),
.A2(n_133),
.B(n_138),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

INVxp67_ASAP7_75t_SL g148 ( 
.A(n_147),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_128),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_152),
.B(n_140),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_141),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_155),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_149),
.B(n_143),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_157),
.C(n_158),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_150),
.A2(n_5),
.B(n_6),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_5),
.Y(n_158)
);

AO21x2_ASAP7_75t_L g160 ( 
.A1(n_154),
.A2(n_152),
.B(n_151),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_160),
.A2(n_18),
.B1(n_7),
.B2(n_12),
.Y(n_163)
);

AOI322xp5_ASAP7_75t_L g162 ( 
.A1(n_159),
.A2(n_151),
.A3(n_111),
.B1(n_40),
.B2(n_30),
.C1(n_18),
.C2(n_90),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g164 ( 
.A1(n_162),
.A2(n_163),
.B(n_161),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_160),
.Y(n_165)
);


endmodule