module fake_jpeg_19331_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_15),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_44),
.Y(n_59)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_28),
.B1(n_30),
.B2(n_33),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_52),
.A2(n_44),
.B1(n_35),
.B2(n_42),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_28),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_60),
.Y(n_66)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_23),
.Y(n_58)
);

AO21x1_ASAP7_75t_L g87 ( 
.A1(n_58),
.A2(n_42),
.B(n_41),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_23),
.Y(n_60)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_53),
.A2(n_30),
.B1(n_33),
.B2(n_44),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_64),
.A2(n_81),
.B1(n_92),
.B2(n_93),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_65),
.B(n_67),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_50),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_68),
.Y(n_124)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_72),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_58),
.C(n_47),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_71),
.B(n_37),
.C(n_23),
.Y(n_115)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_76),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_20),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_46),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_77),
.A2(n_83),
.B1(n_87),
.B2(n_89),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_43),
.B(n_26),
.C(n_21),
.Y(n_78)
);

OAI32xp33_ASAP7_75t_L g113 ( 
.A1(n_78),
.A2(n_22),
.A3(n_25),
.B1(n_26),
.B2(n_34),
.Y(n_113)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_79),
.Y(n_107)
);

BUFx4f_ASAP7_75t_SL g80 ( 
.A(n_61),
.Y(n_80)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_52),
.A2(n_44),
.B1(n_35),
.B2(n_43),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_35),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_85),
.Y(n_117)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_86),
.Y(n_112)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_61),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

BUFx4f_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_55),
.A2(n_30),
.B1(n_33),
.B2(n_44),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_48),
.A2(n_44),
.B1(n_20),
.B2(n_27),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_49),
.B(n_21),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_27),
.Y(n_125)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_96),
.A2(n_37),
.B1(n_36),
.B2(n_40),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_72),
.A2(n_35),
.B1(n_42),
.B2(n_41),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_97),
.A2(n_100),
.B1(n_106),
.B2(n_116),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_68),
.A2(n_35),
.B1(n_37),
.B2(n_22),
.Y(n_100)
);

CKINVDCx12_ASAP7_75t_R g101 ( 
.A(n_80),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_123),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_95),
.A2(n_42),
.B1(n_41),
.B2(n_22),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_103),
.A2(n_90),
.B1(n_96),
.B2(n_65),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_125),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_66),
.A2(n_37),
.B1(n_41),
.B2(n_36),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_114),
.A2(n_74),
.B1(n_84),
.B2(n_82),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_71),
.C(n_83),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_81),
.A2(n_34),
.B1(n_25),
.B2(n_18),
.Y(n_116)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_29),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_127),
.B(n_132),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_128),
.A2(n_138),
.B1(n_145),
.B2(n_149),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_131),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_83),
.C(n_69),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_109),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_133),
.B(n_141),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_78),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_139),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_136),
.A2(n_38),
.B1(n_32),
.B2(n_2),
.Y(n_188)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_102),
.A2(n_62),
.B1(n_70),
.B2(n_88),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_91),
.C(n_73),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_80),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_91),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_151),
.Y(n_177)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_102),
.A2(n_85),
.B1(n_40),
.B2(n_45),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_99),
.A2(n_18),
.B(n_29),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_147),
.A2(n_112),
.B(n_32),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_107),
.B(n_31),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_148),
.B(n_31),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_114),
.A2(n_40),
.B1(n_45),
.B2(n_73),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_105),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_153),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_108),
.B(n_104),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_106),
.A2(n_40),
.B1(n_45),
.B2(n_38),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_45),
.B1(n_119),
.B2(n_40),
.Y(n_181)
);

OAI21xp33_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_101),
.B(n_104),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_SL g201 ( 
.A1(n_156),
.A2(n_136),
.B(n_149),
.Y(n_201)
);

NOR2x1_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_107),
.Y(n_157)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_137),
.A2(n_112),
.B(n_118),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_158),
.A2(n_0),
.B(n_1),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_146),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_162),
.B(n_163),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_143),
.Y(n_163)
);

BUFx24_ASAP7_75t_SL g164 ( 
.A(n_140),
.Y(n_164)
);

BUFx24_ASAP7_75t_SL g204 ( 
.A(n_164),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_169),
.B(n_31),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_170),
.A2(n_32),
.B1(n_23),
.B2(n_19),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_127),
.A2(n_122),
.B1(n_121),
.B2(n_110),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_175),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_154),
.A2(n_122),
.B1(n_121),
.B2(n_110),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_134),
.A2(n_123),
.B1(n_117),
.B2(n_105),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_176),
.A2(n_181),
.B1(n_188),
.B2(n_0),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_144),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_133),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_130),
.B(n_117),
.Y(n_180)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_145),
.A2(n_119),
.B1(n_38),
.B2(n_11),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_182),
.A2(n_187),
.B1(n_152),
.B2(n_155),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_183),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_142),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_184),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_138),
.Y(n_185)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_128),
.A2(n_38),
.B1(n_11),
.B2(n_12),
.Y(n_187)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_189),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_129),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_190),
.B(n_175),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_192),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_131),
.C(n_151),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_210),
.C(n_218),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_134),
.Y(n_196)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_196),
.Y(n_235)
);

MAJx2_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_139),
.C(n_154),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_158),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_153),
.Y(n_198)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_198),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_201),
.A2(n_205),
.B(n_207),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_202),
.A2(n_203),
.B1(n_208),
.B2(n_215),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_160),
.A2(n_24),
.B1(n_32),
.B2(n_23),
.Y(n_203)
);

OA22x2_ASAP7_75t_L g207 ( 
.A1(n_166),
.A2(n_24),
.B1(n_19),
.B2(n_31),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_160),
.A2(n_24),
.B1(n_19),
.B2(n_31),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_159),
.Y(n_209)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_209),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_165),
.B(n_24),
.C(n_7),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_1),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_171),
.B(n_14),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_213),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_170),
.A2(n_13),
.B(n_11),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_214),
.A2(n_157),
.B(n_13),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_186),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_216),
.Y(n_230)
);

OA22x2_ASAP7_75t_L g217 ( 
.A1(n_167),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_217),
.A2(n_188),
.B(n_181),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_177),
.B(n_13),
.C(n_10),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_187),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_182),
.Y(n_231)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_183),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_220),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_197),
.B(n_177),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_223),
.B(n_225),
.Y(n_256)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_217),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_232),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_167),
.C(n_168),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_212),
.C(n_205),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_231),
.A2(n_237),
.B1(n_239),
.B2(n_214),
.Y(n_257)
);

INVx3_ASAP7_75t_SL g232 ( 
.A(n_206),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_240),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_195),
.Y(n_236)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_191),
.A2(n_185),
.B1(n_184),
.B2(n_178),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_194),
.B(n_210),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_174),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_240),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_243),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_200),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_246),
.B(n_227),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_234),
.B(n_199),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_258),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_239),
.A2(n_217),
.B(n_163),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_248),
.A2(n_243),
.B(n_217),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_264),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_259),
.C(n_261),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_226),
.A2(n_211),
.B1(n_193),
.B2(n_202),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_254),
.A2(n_257),
.B1(n_260),
.B2(n_232),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_230),
.B(n_193),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_173),
.C(n_174),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_235),
.A2(n_211),
.B1(n_173),
.B2(n_168),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_179),
.C(n_208),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_228),
.B(n_204),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_262),
.B(n_238),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_231),
.A2(n_203),
.B1(n_219),
.B2(n_179),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_242),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_223),
.B(n_207),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_222),
.B(n_207),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_266),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_222),
.B(n_207),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_267),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_278),
.Y(n_291)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_272),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_241),
.C(n_245),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_279),
.C(n_280),
.Y(n_297)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_250),
.Y(n_275)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_277),
.A2(n_256),
.B1(n_10),
.B2(n_9),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_244),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_251),
.B(n_236),
.C(n_224),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_224),
.C(n_221),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_221),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_282),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_283),
.A2(n_263),
.B(n_264),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_253),
.Y(n_296)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_287),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_268),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_293),
.Y(n_303)
);

BUFx24_ASAP7_75t_SL g293 ( 
.A(n_282),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_280),
.A2(n_266),
.B(n_265),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_276),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_279),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_273),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_296),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_281),
.A2(n_261),
.B1(n_256),
.B2(n_4),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_298),
.A2(n_276),
.B1(n_273),
.B2(n_9),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_299),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_270),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_300),
.B(n_304),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_308),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_274),
.C(n_270),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_307),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_7),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_9),
.C(n_3),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_288),
.C(n_299),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_312),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_292),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_309),
.A2(n_305),
.B1(n_290),
.B2(n_286),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_316),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_310),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_315),
.A2(n_287),
.B(n_4),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_303),
.A2(n_291),
.B(n_294),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_301),
.C(n_285),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_317),
.B(n_285),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_323),
.Y(n_327)
);

OAI21xp33_ASAP7_75t_L g324 ( 
.A1(n_319),
.A2(n_2),
.B(n_4),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_324),
.A2(n_325),
.B(n_5),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_SL g325 ( 
.A(n_313),
.B(n_5),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_326),
.B(n_328),
.C(n_315),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_318),
.Y(n_328)
);

INVxp33_ASAP7_75t_L g330 ( 
.A(n_329),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_318),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_R g332 ( 
.A(n_331),
.B(n_327),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_320),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_6),
.B(n_328),
.Y(n_334)
);


endmodule