module fake_jpeg_23970_n_27 (n_3, n_2, n_1, n_0, n_4, n_5, n_27);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_27;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

NAND2xp5_ASAP7_75t_L g6 ( 
.A(n_1),
.B(n_0),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_2),
.B(n_3),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_12),
.Y(n_18)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_13),
.A2(n_14),
.B(n_15),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_0),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_7),
.B(n_0),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_15),
.A2(n_8),
.B1(n_11),
.B2(n_10),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_16),
.A2(n_8),
.B(n_11),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_19),
.B(n_20),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_18),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_17),
.C(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_1),
.Y(n_25)
);

AOI31xp67_ASAP7_75t_L g24 ( 
.A1(n_22),
.A2(n_12),
.A3(n_10),
.B(n_4),
.Y(n_24)
);

NAND3xp33_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_25),
.C(n_5),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_26),
.A2(n_5),
.B(n_2),
.Y(n_27)
);


endmodule