module fake_netlist_5_2215_n_2265 (n_137, n_676, n_294, n_431, n_318, n_380, n_419, n_653, n_611, n_444, n_642, n_469, n_615, n_82, n_194, n_316, n_389, n_549, n_684, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_705, n_619, n_408, n_61, n_678, n_664, n_376, n_697, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_667, n_515, n_57, n_353, n_351, n_367, n_620, n_643, n_452, n_397, n_493, n_111, n_525, n_703, n_698, n_483, n_544, n_683, n_155, n_649, n_552, n_547, n_43, n_721, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_725, n_139, n_38, n_105, n_280, n_744, n_590, n_629, n_672, n_4, n_378, n_551, n_17, n_581, n_688, n_382, n_554, n_254, n_690, n_33, n_23, n_583, n_671, n_718, n_302, n_265, n_526, n_719, n_293, n_372, n_443, n_244, n_677, n_47, n_173, n_198, n_714, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_625, n_621, n_753, n_100, n_455, n_674, n_417, n_612, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_689, n_738, n_606, n_559, n_275, n_640, n_252, n_624, n_26, n_295, n_133, n_330, n_508, n_739, n_506, n_2, n_737, n_610, n_692, n_755, n_6, n_509, n_568, n_39, n_147, n_373, n_757, n_67, n_307, n_633, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_758, n_668, n_733, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_659, n_51, n_63, n_492, n_563, n_171, n_153, n_756, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_741, n_548, n_543, n_260, n_298, n_650, n_320, n_694, n_518, n_505, n_286, n_122, n_282, n_752, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_724, n_546, n_101, n_658, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_731, n_31, n_456, n_13, n_371, n_481, n_535, n_709, n_152, n_540, n_317, n_618, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_654, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_603, n_225, n_377, n_751, n_484, n_219, n_442, n_157, n_131, n_192, n_636, n_600, n_660, n_223, n_392, n_158, n_655, n_704, n_138, n_264, n_109, n_669, n_472, n_742, n_750, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_635, n_347, n_169, n_59, n_522, n_550, n_255, n_696, n_215, n_350, n_196, n_662, n_459, n_646, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_622, n_723, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_661, n_104, n_41, n_682, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_670, n_15, n_336, n_584, n_681, n_591, n_145, n_48, n_521, n_614, n_663, n_50, n_337, n_430, n_313, n_631, n_673, n_88, n_479, n_528, n_510, n_216, n_680, n_168, n_395, n_164, n_432, n_553, n_727, n_311, n_208, n_142, n_743, n_214, n_328, n_140, n_299, n_303, n_369, n_675, n_296, n_613, n_241, n_637, n_357, n_598, n_685, n_608, n_184, n_446, n_445, n_65, n_78, n_749, n_144, n_114, n_96, n_691, n_717, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_734, n_638, n_700, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_740, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_693, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_652, n_29, n_79, n_151, n_25, n_306, n_722, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_609, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_711, n_474, n_112, n_542, n_85, n_463, n_488, n_595, n_736, n_502, n_239, n_466, n_420, n_630, n_489, n_632, n_699, n_55, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_748, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_745, n_627, n_172, n_206, n_217, n_440, n_726, n_478, n_545, n_441, n_450, n_648, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_641, n_628, n_365, n_91, n_729, n_730, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_647, n_237, n_425, n_513, n_407, n_527, n_679, n_707, n_710, n_695, n_180, n_560, n_656, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_665, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_720, n_0, n_58, n_623, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_686, n_205, n_366, n_572, n_113, n_712, n_754, n_246, n_596, n_179, n_125, n_410, n_558, n_708, n_269, n_529, n_128, n_735, n_702, n_285, n_412, n_120, n_232, n_327, n_135, n_657, n_126, n_644, n_728, n_202, n_266, n_272, n_491, n_427, n_732, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_716, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_651, n_435, n_159, n_334, n_599, n_541, n_391, n_701, n_434, n_645, n_539, n_175, n_538, n_666, n_262, n_238, n_639, n_99, n_687, n_715, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_200, n_162, n_64, n_759, n_222, n_28, n_89, n_438, n_115, n_713, n_324, n_634, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_626, n_11, n_424, n_7, n_706, n_746, n_256, n_305, n_533, n_747, n_52, n_278, n_110, n_2265);

input n_137;
input n_676;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_653;
input n_611;
input n_444;
input n_642;
input n_469;
input n_615;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_684;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_705;
input n_619;
input n_408;
input n_61;
input n_678;
input n_664;
input n_376;
input n_697;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_667;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_643;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_703;
input n_698;
input n_483;
input n_544;
input n_683;
input n_155;
input n_649;
input n_552;
input n_547;
input n_43;
input n_721;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_725;
input n_139;
input n_38;
input n_105;
input n_280;
input n_744;
input n_590;
input n_629;
input n_672;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_688;
input n_382;
input n_554;
input n_254;
input n_690;
input n_33;
input n_23;
input n_583;
input n_671;
input n_718;
input n_302;
input n_265;
input n_526;
input n_719;
input n_293;
input n_372;
input n_443;
input n_244;
input n_677;
input n_47;
input n_173;
input n_198;
input n_714;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_625;
input n_621;
input n_753;
input n_100;
input n_455;
input n_674;
input n_417;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_689;
input n_738;
input n_606;
input n_559;
input n_275;
input n_640;
input n_252;
input n_624;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_739;
input n_506;
input n_2;
input n_737;
input n_610;
input n_692;
input n_755;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_757;
input n_67;
input n_307;
input n_633;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_758;
input n_668;
input n_733;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_659;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_756;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_741;
input n_548;
input n_543;
input n_260;
input n_298;
input n_650;
input n_320;
input n_694;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_752;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_724;
input n_546;
input n_101;
input n_658;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_731;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_709;
input n_152;
input n_540;
input n_317;
input n_618;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_654;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_603;
input n_225;
input n_377;
input n_751;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_636;
input n_600;
input n_660;
input n_223;
input n_392;
input n_158;
input n_655;
input n_704;
input n_138;
input n_264;
input n_109;
input n_669;
input n_472;
input n_742;
input n_750;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_635;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_696;
input n_215;
input n_350;
input n_196;
input n_662;
input n_459;
input n_646;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_723;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_661;
input n_104;
input n_41;
input n_682;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_670;
input n_15;
input n_336;
input n_584;
input n_681;
input n_591;
input n_145;
input n_48;
input n_521;
input n_614;
input n_663;
input n_50;
input n_337;
input n_430;
input n_313;
input n_631;
input n_673;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_680;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_727;
input n_311;
input n_208;
input n_142;
input n_743;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_675;
input n_296;
input n_613;
input n_241;
input n_637;
input n_357;
input n_598;
input n_685;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_749;
input n_144;
input n_114;
input n_96;
input n_691;
input n_717;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_734;
input n_638;
input n_700;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_740;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_693;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_652;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_722;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_609;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_711;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_736;
input n_502;
input n_239;
input n_466;
input n_420;
input n_630;
input n_489;
input n_632;
input n_699;
input n_55;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_748;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_745;
input n_627;
input n_172;
input n_206;
input n_217;
input n_440;
input n_726;
input n_478;
input n_545;
input n_441;
input n_450;
input n_648;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_641;
input n_628;
input n_365;
input n_91;
input n_729;
input n_730;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_647;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_679;
input n_707;
input n_710;
input n_695;
input n_180;
input n_560;
input n_656;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_665;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_720;
input n_0;
input n_58;
input n_623;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_686;
input n_205;
input n_366;
input n_572;
input n_113;
input n_712;
input n_754;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_708;
input n_269;
input n_529;
input n_128;
input n_735;
input n_702;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_657;
input n_126;
input n_644;
input n_728;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_732;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_716;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_651;
input n_435;
input n_159;
input n_334;
input n_599;
input n_541;
input n_391;
input n_701;
input n_434;
input n_645;
input n_539;
input n_175;
input n_538;
input n_666;
input n_262;
input n_238;
input n_639;
input n_99;
input n_687;
input n_715;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_200;
input n_162;
input n_64;
input n_759;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_713;
input n_324;
input n_634;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_626;
input n_11;
input n_424;
input n_7;
input n_706;
input n_746;
input n_256;
input n_305;
input n_533;
input n_747;
input n_52;
input n_278;
input n_110;

output n_2265;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_1508;
wire n_785;
wire n_2200;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_1780;
wire n_1488;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_1007;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_1939;
wire n_1806;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_1359;
wire n_1728;
wire n_1107;
wire n_2076;
wire n_2031;
wire n_1230;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_2203;
wire n_1243;
wire n_1016;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2144;
wire n_1778;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2085;
wire n_1669;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_897;
wire n_798;
wire n_1428;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_926;
wire n_2180;
wire n_2249;
wire n_1218;
wire n_1931;
wire n_1070;
wire n_777;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_1513;
wire n_1600;
wire n_845;
wire n_2235;
wire n_1862;
wire n_837;
wire n_1239;
wire n_1796;
wire n_1587;
wire n_1473;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_889;
wire n_973;
wire n_1700;
wire n_1585;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_2258;
wire n_1058;
wire n_1667;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_1385;
wire n_793;
wire n_2140;
wire n_1819;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_1072;
wire n_2218;
wire n_857;
wire n_832;
wire n_1319;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_847;
wire n_1393;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_1884;
wire n_1038;
wire n_1369;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_809;
wire n_870;
wire n_931;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_868;
wire n_914;
wire n_2120;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_1649;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_913;
wire n_1537;
wire n_865;
wire n_2227;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_1333;
wire n_1121;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_1624;
wire n_1510;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_1760;
wire n_936;
wire n_1500;
wire n_1090;
wire n_1832;
wire n_1851;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_959;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_1079;
wire n_2093;
wire n_1045;
wire n_1208;
wire n_2038;
wire n_2137;
wire n_1431;
wire n_1593;
wire n_1033;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_2029;
wire n_995;
wire n_2168;
wire n_1609;
wire n_1989;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_2048;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_1800;
wire n_1548;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_2081;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_1237;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_1823;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_860;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_1849;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_1351;
wire n_2240;
wire n_1205;
wire n_1044;
wire n_1209;
wire n_1552;
wire n_1435;
wire n_879;
wire n_2088;
wire n_824;
wire n_1645;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_1630;
wire n_2122;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_803;
wire n_1092;
wire n_1776;
wire n_2198;
wire n_2131;
wire n_2216;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_950;
wire n_1553;
wire n_1811;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_912;
wire n_968;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_1139;
wire n_885;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_1974;
wire n_2086;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_1179;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2123;
wire n_972;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_842;
wire n_984;
wire n_2082;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_896;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_2020;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_1149;
wire n_1671;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_1802;
wire n_849;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_830;
wire n_2098;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_939;
wire n_1088;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_1653;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_1465;
wire n_778;
wire n_1122;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_1174;
wire n_1371;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_1410;
wire n_1005;
wire n_1003;
wire n_2067;
wire n_1168;
wire n_2219;
wire n_2148;
wire n_937;
wire n_1427;
wire n_1584;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_1496;
wire n_1125;
wire n_1812;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_1533;
wire n_2224;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_1067;
wire n_1720;
wire n_2003;
wire n_766;
wire n_1457;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_872;
wire n_2012;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1184;
wire n_1011;
wire n_2184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_2023;
wire n_2213;
wire n_2211;
wire n_2095;
wire n_2103;
wire n_2160;
wire n_2228;
wire n_1602;
wire n_1178;
wire n_855;
wire n_1461;
wire n_850;
wire n_1999;
wire n_2065;
wire n_2136;
wire n_1372;
wire n_1273;
wire n_1822;
wire n_916;
wire n_1081;
wire n_1235;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_1120;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_825;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_1718;
wire n_986;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2239;
wire n_792;
wire n_1429;
wire n_1238;
wire n_812;
wire n_2104;
wire n_2057;
wire n_1772;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_1172;
wire n_1341;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_787;
wire n_1770;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1873;
wire n_1411;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2183;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_1589;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_1277;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_1546;
wire n_1337;
wire n_1495;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_1321;
wire n_1975;
wire n_2070;
wire n_1937;
wire n_2112;
wire n_1739;
wire n_1914;
wire n_2135;
wire n_1654;
wire n_1103;
wire n_1379;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_795;
wire n_2083;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2027;
wire n_1130;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_2049;
wire n_1493;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_1340;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_1138;
wire n_2044;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_1542;
wire n_1251;

INVx1_ASAP7_75t_L g760 ( 
.A(n_111),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_590),
.Y(n_761)
);

CKINVDCx20_ASAP7_75t_R g762 ( 
.A(n_99),
.Y(n_762)
);

INVx1_ASAP7_75t_SL g763 ( 
.A(n_227),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_497),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_574),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_756),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_727),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_445),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_591),
.Y(n_769)
);

CKINVDCx20_ASAP7_75t_R g770 ( 
.A(n_473),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_184),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_157),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_179),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_308),
.Y(n_774)
);

BUFx3_ASAP7_75t_L g775 ( 
.A(n_428),
.Y(n_775)
);

CKINVDCx20_ASAP7_75t_R g776 ( 
.A(n_194),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_499),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_322),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_292),
.Y(n_779)
);

CKINVDCx16_ASAP7_75t_R g780 ( 
.A(n_185),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_484),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_625),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_396),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_316),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_433),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_83),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_658),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_676),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_387),
.Y(n_789)
);

BUFx2_ASAP7_75t_R g790 ( 
.A(n_474),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_292),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_744),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_557),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_476),
.Y(n_794)
);

INVx1_ASAP7_75t_SL g795 ( 
.A(n_410),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_490),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_495),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_604),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_483),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_493),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_699),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_639),
.Y(n_802)
);

INVxp67_ASAP7_75t_L g803 ( 
.A(n_97),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_750),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_540),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_702),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_549),
.Y(n_807)
);

CKINVDCx20_ASAP7_75t_R g808 ( 
.A(n_406),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_281),
.Y(n_809)
);

BUFx5_ASAP7_75t_L g810 ( 
.A(n_675),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_226),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_524),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_522),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_370),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_109),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_475),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_226),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_446),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_152),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_254),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_196),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_28),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_417),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_333),
.Y(n_824)
);

INVxp67_ASAP7_75t_SL g825 ( 
.A(n_12),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_183),
.Y(n_826)
);

BUFx10_ASAP7_75t_L g827 ( 
.A(n_82),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_648),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_398),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_494),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_320),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_270),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_506),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_460),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_726),
.Y(n_835)
);

BUFx10_ASAP7_75t_L g836 ( 
.A(n_468),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_372),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_482),
.Y(n_838)
);

CKINVDCx20_ASAP7_75t_R g839 ( 
.A(n_244),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_136),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_372),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_517),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_62),
.Y(n_843)
);

BUFx3_ASAP7_75t_L g844 ( 
.A(n_740),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_82),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_754),
.Y(n_846)
);

INVx1_ASAP7_75t_SL g847 ( 
.A(n_43),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_43),
.Y(n_848)
);

CKINVDCx20_ASAP7_75t_R g849 ( 
.A(n_386),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_659),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_323),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_228),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_93),
.Y(n_853)
);

BUFx3_ASAP7_75t_L g854 ( 
.A(n_77),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_569),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_491),
.Y(n_856)
);

BUFx2_ASAP7_75t_L g857 ( 
.A(n_399),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_488),
.Y(n_858)
);

CKINVDCx20_ASAP7_75t_R g859 ( 
.A(n_736),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_560),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_106),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_757),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_732),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_507),
.Y(n_864)
);

CKINVDCx16_ASAP7_75t_R g865 ( 
.A(n_747),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_555),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_311),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_545),
.Y(n_868)
);

CKINVDCx20_ASAP7_75t_R g869 ( 
.A(n_125),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_496),
.Y(n_870)
);

CKINVDCx20_ASAP7_75t_R g871 ( 
.A(n_565),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_293),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_134),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_338),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_731),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_626),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_300),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_568),
.Y(n_878)
);

CKINVDCx20_ASAP7_75t_R g879 ( 
.A(n_577),
.Y(n_879)
);

BUFx10_ASAP7_75t_L g880 ( 
.A(n_263),
.Y(n_880)
);

CKINVDCx16_ASAP7_75t_R g881 ( 
.A(n_192),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_484),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_194),
.Y(n_883)
);

CKINVDCx20_ASAP7_75t_R g884 ( 
.A(n_176),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_501),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_237),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_497),
.Y(n_887)
);

CKINVDCx14_ASAP7_75t_R g888 ( 
.A(n_295),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_341),
.Y(n_889)
);

CKINVDCx20_ASAP7_75t_R g890 ( 
.A(n_101),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_624),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_462),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_495),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_153),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_743),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_694),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_16),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_715),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_665),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_236),
.Y(n_900)
);

INVx1_ASAP7_75t_SL g901 ( 
.A(n_615),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_471),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_415),
.Y(n_903)
);

BUFx5_ASAP7_75t_L g904 ( 
.A(n_723),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_36),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_608),
.Y(n_906)
);

CKINVDCx20_ASAP7_75t_R g907 ( 
.A(n_587),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_343),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_129),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_244),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_310),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_485),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_84),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_508),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_170),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_689),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_322),
.Y(n_917)
);

CKINVDCx20_ASAP7_75t_R g918 ( 
.A(n_430),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_710),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_396),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_201),
.Y(n_921)
);

BUFx8_ASAP7_75t_SL g922 ( 
.A(n_645),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_481),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_230),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_463),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_510),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_628),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_730),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_155),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_691),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_392),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_537),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_742),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_623),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_170),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_441),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_486),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_259),
.Y(n_938)
);

CKINVDCx20_ASAP7_75t_R g939 ( 
.A(n_3),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_228),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_746),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_187),
.Y(n_942)
);

CKINVDCx20_ASAP7_75t_R g943 ( 
.A(n_429),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_257),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_634),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_423),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_426),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_573),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_158),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_480),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_195),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_324),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_263),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_758),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_328),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_391),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_131),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_505),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_635),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_155),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_753),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_729),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_410),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_218),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_572),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_312),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_532),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_65),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_759),
.Y(n_969)
);

BUFx10_ASAP7_75t_L g970 ( 
.A(n_527),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_419),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_123),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_358),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_51),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_592),
.Y(n_975)
);

CKINVDCx20_ASAP7_75t_R g976 ( 
.A(n_128),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_257),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_479),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_333),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_594),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_324),
.Y(n_981)
);

CKINVDCx20_ASAP7_75t_R g982 ( 
.A(n_382),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_700),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_203),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_142),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_513),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_614),
.Y(n_987)
);

BUFx5_ASAP7_75t_L g988 ( 
.A(n_101),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_139),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_509),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_498),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_503),
.Y(n_992)
);

CKINVDCx14_ASAP7_75t_R g993 ( 
.A(n_535),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_489),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_91),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_610),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_384),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_361),
.Y(n_998)
);

BUFx5_ASAP7_75t_L g999 ( 
.A(n_636),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_552),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_533),
.Y(n_1001)
);

CKINVDCx20_ASAP7_75t_R g1002 ( 
.A(n_516),
.Y(n_1002)
);

INVx1_ASAP7_75t_SL g1003 ( 
.A(n_500),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_504),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_712),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_627),
.Y(n_1006)
);

INVxp67_ASAP7_75t_L g1007 ( 
.A(n_472),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_306),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_477),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_748),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_745),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_492),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_755),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_321),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_229),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_4),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_487),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_739),
.Y(n_1018)
);

CKINVDCx20_ASAP7_75t_R g1019 ( 
.A(n_332),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_393),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_582),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_749),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_232),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_603),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_356),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_35),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_656),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_98),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_561),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_455),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_660),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_456),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_705),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_317),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_41),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_99),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_558),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_383),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_453),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_502),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_143),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_60),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_242),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_239),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_288),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_602),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_469),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_250),
.Y(n_1048)
);

CKINVDCx16_ASAP7_75t_R g1049 ( 
.A(n_383),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_470),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_293),
.Y(n_1051)
);

HB1xp67_ASAP7_75t_L g1052 ( 
.A(n_299),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_709),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_53),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_579),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_159),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_19),
.Y(n_1057)
);

CKINVDCx20_ASAP7_75t_R g1058 ( 
.A(n_198),
.Y(n_1058)
);

BUFx5_ASAP7_75t_L g1059 ( 
.A(n_5),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_539),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_129),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_349),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_490),
.Y(n_1063)
);

CKINVDCx20_ASAP7_75t_R g1064 ( 
.A(n_633),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_377),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_734),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_737),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_275),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_752),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_222),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_416),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_567),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_316),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_103),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_344),
.Y(n_1075)
);

BUFx2_ASAP7_75t_SL g1076 ( 
.A(n_378),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_31),
.Y(n_1077)
);

CKINVDCx16_ASAP7_75t_R g1078 ( 
.A(n_599),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_500),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_751),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_455),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_311),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_595),
.Y(n_1083)
);

INVx1_ASAP7_75t_SL g1084 ( 
.A(n_211),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_19),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_478),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_741),
.Y(n_1087)
);

BUFx5_ASAP7_75t_L g1088 ( 
.A(n_169),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_407),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_168),
.Y(n_1090)
);

CKINVDCx20_ASAP7_75t_R g1091 ( 
.A(n_3),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_108),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_657),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_629),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_432),
.Y(n_1095)
);

INVxp67_ASAP7_75t_L g1096 ( 
.A(n_597),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_738),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_735),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_704),
.Y(n_1099)
);

INVx1_ASAP7_75t_SL g1100 ( 
.A(n_664),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_733),
.Y(n_1101)
);

CKINVDCx16_ASAP7_75t_R g1102 ( 
.A(n_780),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_922),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_806),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_988),
.Y(n_1105)
);

CKINVDCx20_ASAP7_75t_R g1106 ( 
.A(n_842),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_988),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_988),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1059),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_765),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1059),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1059),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1059),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_766),
.Y(n_1114)
);

CKINVDCx20_ASAP7_75t_R g1115 ( 
.A(n_846),
.Y(n_1115)
);

INVxp33_ASAP7_75t_SL g1116 ( 
.A(n_1052),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_767),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1059),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_859),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1088),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1088),
.Y(n_1121)
);

CKINVDCx20_ASAP7_75t_R g1122 ( 
.A(n_871),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_769),
.Y(n_1123)
);

NOR2xp67_ASAP7_75t_L g1124 ( 
.A(n_778),
.B(n_0),
.Y(n_1124)
);

CKINVDCx16_ASAP7_75t_R g1125 ( 
.A(n_881),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_879),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1088),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_778),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_764),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_764),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_764),
.Y(n_1131)
);

INVxp67_ASAP7_75t_L g1132 ( 
.A(n_857),
.Y(n_1132)
);

CKINVDCx20_ASAP7_75t_R g1133 ( 
.A(n_907),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_923),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_923),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_923),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_989),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_989),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_989),
.Y(n_1139)
);

CKINVDCx20_ASAP7_75t_R g1140 ( 
.A(n_969),
.Y(n_1140)
);

CKINVDCx20_ASAP7_75t_R g1141 ( 
.A(n_1002),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_782),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_788),
.Y(n_1143)
);

INVxp67_ASAP7_75t_SL g1144 ( 
.A(n_1060),
.Y(n_1144)
);

CKINVDCx20_ASAP7_75t_R g1145 ( 
.A(n_1064),
.Y(n_1145)
);

NAND2xp33_ASAP7_75t_R g1146 ( 
.A(n_962),
.B(n_0),
.Y(n_1146)
);

CKINVDCx20_ASAP7_75t_R g1147 ( 
.A(n_1066),
.Y(n_1147)
);

CKINVDCx20_ASAP7_75t_R g1148 ( 
.A(n_1080),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1041),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_888),
.B(n_1),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1041),
.Y(n_1151)
);

CKINVDCx20_ASAP7_75t_R g1152 ( 
.A(n_865),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1041),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_775),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_793),
.Y(n_1155)
);

CKINVDCx20_ASAP7_75t_R g1156 ( 
.A(n_1078),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_798),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_854),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_897),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_801),
.Y(n_1160)
);

CKINVDCx20_ASAP7_75t_R g1161 ( 
.A(n_993),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_1150),
.B(n_1049),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_1153),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1129),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1130),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1131),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1134),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1110),
.B(n_844),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1135),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1136),
.Y(n_1170)
);

OA21x2_ASAP7_75t_L g1171 ( 
.A1(n_1105),
.A2(n_1096),
.B(n_761),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_1114),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1137),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1138),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1139),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1149),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1151),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1117),
.B(n_1027),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_1154),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1108),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1107),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1109),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_1152),
.Y(n_1183)
);

CKINVDCx8_ASAP7_75t_R g1184 ( 
.A(n_1102),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_1111),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_1156),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1112),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_1113),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_1123),
.B(n_901),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1118),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1120),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1144),
.B(n_1056),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_1125),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1121),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_SL g1195 ( 
.A1(n_1116),
.A2(n_762),
.B1(n_776),
.B2(n_770),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1127),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_1128),
.Y(n_1197)
);

AND2x6_ASAP7_75t_L g1198 ( 
.A(n_1158),
.B(n_792),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_1159),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1142),
.B(n_1053),
.Y(n_1200)
);

INVx3_ASAP7_75t_L g1201 ( 
.A(n_1143),
.Y(n_1201)
);

INVx3_ASAP7_75t_L g1202 ( 
.A(n_1155),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1161),
.B(n_970),
.Y(n_1203)
);

BUFx6f_ASAP7_75t_L g1204 ( 
.A(n_1157),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1160),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1124),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1103),
.B(n_970),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1132),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1146),
.A2(n_813),
.B(n_805),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1189),
.B(n_1005),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1185),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1162),
.A2(n_1007),
.B1(n_803),
.B2(n_825),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1163),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1185),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_1188),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1182),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1187),
.Y(n_1217)
);

BUFx10_ASAP7_75t_L g1218 ( 
.A(n_1172),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_SL g1219 ( 
.A(n_1184),
.B(n_790),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1190),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1191),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_1199),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_1168),
.B(n_1104),
.Y(n_1223)
);

AOI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1192),
.A2(n_1115),
.B1(n_1119),
.B2(n_1106),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1178),
.B(n_1100),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1200),
.B(n_1122),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1199),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1208),
.B(n_827),
.Y(n_1228)
);

AND2x6_ASAP7_75t_L g1229 ( 
.A(n_1204),
.B(n_1017),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_1197),
.Y(n_1230)
);

INVx2_ASAP7_75t_SL g1231 ( 
.A(n_1193),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1181),
.Y(n_1232)
);

OR2x6_ASAP7_75t_L g1233 ( 
.A(n_1183),
.B(n_1076),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1180),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1201),
.B(n_1126),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1206),
.B(n_802),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_1194),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1209),
.B(n_804),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1202),
.B(n_1133),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1174),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_1179),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_1205),
.B(n_1207),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1196),
.B(n_807),
.Y(n_1243)
);

AND2x6_ASAP7_75t_L g1244 ( 
.A(n_1164),
.B(n_763),
.Y(n_1244)
);

INVxp33_ASAP7_75t_L g1245 ( 
.A(n_1195),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1165),
.Y(n_1246)
);

AND2x6_ASAP7_75t_L g1247 ( 
.A(n_1166),
.B(n_795),
.Y(n_1247)
);

AND2x6_ASAP7_75t_L g1248 ( 
.A(n_1167),
.B(n_847),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_1203),
.B(n_812),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1176),
.B(n_1169),
.Y(n_1250)
);

INVx4_ASAP7_75t_L g1251 ( 
.A(n_1171),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1170),
.B(n_823),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_1173),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_1175),
.B(n_1140),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_1186),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1177),
.B(n_835),
.Y(n_1256)
);

BUFx2_ASAP7_75t_L g1257 ( 
.A(n_1198),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1198),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1163),
.Y(n_1259)
);

INVx6_ASAP7_75t_L g1260 ( 
.A(n_1199),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_1172),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1185),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1193),
.Y(n_1263)
);

BUFx8_ASAP7_75t_L g1264 ( 
.A(n_1263),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1250),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1228),
.B(n_1141),
.Y(n_1266)
);

AOI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1210),
.A2(n_1147),
.B1(n_1148),
.B2(n_1145),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1225),
.B(n_787),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1240),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1232),
.Y(n_1270)
);

OR2x6_ASAP7_75t_L g1271 ( 
.A(n_1231),
.B(n_1233),
.Y(n_1271)
);

INVxp67_ASAP7_75t_L g1272 ( 
.A(n_1244),
.Y(n_1272)
);

BUFx2_ASAP7_75t_L g1273 ( 
.A(n_1255),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1246),
.Y(n_1274)
);

AND2x4_ASAP7_75t_L g1275 ( 
.A(n_1213),
.B(n_760),
.Y(n_1275)
);

OR2x6_ASAP7_75t_L g1276 ( 
.A(n_1260),
.B(n_920),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1216),
.B(n_828),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1217),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1237),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1237),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1220),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_1230),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1221),
.B(n_862),
.Y(n_1283)
);

AO22x2_ASAP7_75t_L g1284 ( 
.A1(n_1245),
.A2(n_1084),
.B1(n_1003),
.B2(n_838),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1223),
.B(n_836),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1259),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1253),
.Y(n_1287)
);

INVxp67_ASAP7_75t_L g1288 ( 
.A(n_1247),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1226),
.A2(n_855),
.B1(n_860),
.B2(n_850),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1253),
.Y(n_1290)
);

OAI221xp5_ASAP7_75t_L g1291 ( 
.A1(n_1236),
.A2(n_785),
.B1(n_794),
.B2(n_783),
.C(n_779),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1241),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1251),
.B(n_875),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1252),
.Y(n_1294)
);

BUFx8_ASAP7_75t_L g1295 ( 
.A(n_1229),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1218),
.B(n_836),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1211),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1214),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1262),
.Y(n_1299)
);

OAI221xp5_ASAP7_75t_L g1300 ( 
.A1(n_1256),
.A2(n_1095),
.B1(n_809),
.B2(n_814),
.C(n_799),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1261),
.Y(n_1301)
);

AO22x2_ASAP7_75t_L g1302 ( 
.A1(n_1249),
.A2(n_874),
.B1(n_909),
.B2(n_831),
.Y(n_1302)
);

OA22x2_ASAP7_75t_L g1303 ( 
.A1(n_1224),
.A2(n_771),
.B1(n_773),
.B2(n_768),
.Y(n_1303)
);

AO22x2_ASAP7_75t_L g1304 ( 
.A1(n_1219),
.A2(n_1242),
.B1(n_837),
.B2(n_848),
.Y(n_1304)
);

NAND2x1p5_ASAP7_75t_L g1305 ( 
.A(n_1222),
.B(n_898),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1215),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_SL g1307 ( 
.A1(n_1235),
.A2(n_839),
.B1(n_840),
.B2(n_808),
.Y(n_1307)
);

AND2x4_ASAP7_75t_L g1308 ( 
.A(n_1229),
.B(n_797),
.Y(n_1308)
);

OAI221xp5_ASAP7_75t_L g1309 ( 
.A1(n_1243),
.A2(n_819),
.B1(n_824),
.B2(n_817),
.C(n_816),
.Y(n_1309)
);

AND2x6_ASAP7_75t_L g1310 ( 
.A(n_1239),
.B(n_830),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1238),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1254),
.B(n_774),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1258),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1257),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1248),
.Y(n_1315)
);

AO22x2_ASAP7_75t_L g1316 ( 
.A1(n_1212),
.A2(n_942),
.B1(n_955),
.B2(n_924),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1250),
.Y(n_1317)
);

AO22x2_ASAP7_75t_L g1318 ( 
.A1(n_1212),
.A2(n_946),
.B1(n_972),
.B2(n_925),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1250),
.Y(n_1319)
);

INVx4_ASAP7_75t_L g1320 ( 
.A(n_1215),
.Y(n_1320)
);

AND2x2_ASAP7_75t_SL g1321 ( 
.A(n_1219),
.B(n_772),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1250),
.Y(n_1322)
);

AND2x4_ASAP7_75t_L g1323 ( 
.A(n_1213),
.B(n_834),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1234),
.Y(n_1324)
);

AO22x2_ASAP7_75t_L g1325 ( 
.A1(n_1212),
.A2(n_882),
.B1(n_953),
.B2(n_870),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1250),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1250),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_SL g1328 ( 
.A(n_1210),
.B(n_863),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1234),
.Y(n_1329)
);

OAI221xp5_ASAP7_75t_L g1330 ( 
.A1(n_1210),
.A2(n_867),
.B1(n_872),
.B2(n_858),
.C(n_852),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_SL g1331 ( 
.A(n_1210),
.B(n_1098),
.Y(n_1331)
);

AOI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1210),
.A2(n_868),
.B1(n_876),
.B2(n_866),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1210),
.B(n_899),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1250),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1250),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_SL g1336 ( 
.A(n_1210),
.B(n_1099),
.Y(n_1336)
);

AND2x6_ASAP7_75t_L g1337 ( 
.A(n_1223),
.B(n_885),
.Y(n_1337)
);

NAND2x1p5_ASAP7_75t_L g1338 ( 
.A(n_1227),
.B(n_941),
.Y(n_1338)
);

AO22x2_ASAP7_75t_L g1339 ( 
.A1(n_1212),
.A2(n_900),
.B1(n_937),
.B2(n_892),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_1260),
.Y(n_1340)
);

NAND2x1p5_ASAP7_75t_L g1341 ( 
.A(n_1227),
.B(n_945),
.Y(n_1341)
);

AO22x2_ASAP7_75t_L g1342 ( 
.A1(n_1212),
.A2(n_1036),
.B1(n_903),
.B2(n_887),
.Y(n_1342)
);

AO22x2_ASAP7_75t_L g1343 ( 
.A1(n_1212),
.A2(n_990),
.B1(n_1074),
.B2(n_963),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1250),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1210),
.B(n_948),
.Y(n_1345)
);

NAND2xp33_ASAP7_75t_L g1346 ( 
.A(n_1210),
.B(n_878),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1213),
.B(n_886),
.Y(n_1347)
);

AO22x2_ASAP7_75t_L g1348 ( 
.A1(n_1212),
.A2(n_921),
.B1(n_956),
.B2(n_914),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1250),
.Y(n_1349)
);

AOI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1210),
.A2(n_895),
.B1(n_896),
.B2(n_891),
.Y(n_1350)
);

INVxp67_ASAP7_75t_L g1351 ( 
.A(n_1228),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1250),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1250),
.Y(n_1353)
);

AO22x2_ASAP7_75t_L g1354 ( 
.A1(n_1212),
.A2(n_1045),
.B1(n_1054),
.B2(n_979),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1250),
.Y(n_1355)
);

OR2x6_ASAP7_75t_L g1356 ( 
.A(n_1231),
.B(n_786),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1250),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1210),
.B(n_1101),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1250),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1250),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1250),
.Y(n_1361)
);

INVxp67_ASAP7_75t_L g1362 ( 
.A(n_1228),
.Y(n_1362)
);

INVx4_ASAP7_75t_L g1363 ( 
.A(n_1215),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1250),
.Y(n_1364)
);

AO22x2_ASAP7_75t_L g1365 ( 
.A1(n_1212),
.A2(n_911),
.B1(n_917),
.B2(n_908),
.Y(n_1365)
);

NAND2xp33_ASAP7_75t_L g1366 ( 
.A(n_1210),
.B(n_906),
.Y(n_1366)
);

NAND2xp33_ASAP7_75t_SL g1367 ( 
.A(n_1315),
.B(n_849),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_SL g1368 ( 
.A(n_1351),
.B(n_916),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1333),
.B(n_965),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_SL g1370 ( 
.A(n_1362),
.B(n_919),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1345),
.B(n_975),
.Y(n_1371)
);

NAND2xp33_ASAP7_75t_SL g1372 ( 
.A(n_1301),
.B(n_861),
.Y(n_1372)
);

NAND2xp33_ASAP7_75t_SL g1373 ( 
.A(n_1314),
.B(n_869),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1312),
.B(n_926),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_SL g1375 ( 
.A(n_1285),
.B(n_927),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_SL g1376 ( 
.A(n_1265),
.B(n_928),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_SL g1377 ( 
.A(n_1317),
.B(n_930),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1319),
.B(n_880),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_SL g1379 ( 
.A(n_1322),
.B(n_933),
.Y(n_1379)
);

NAND2xp33_ASAP7_75t_SL g1380 ( 
.A(n_1282),
.B(n_884),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1268),
.B(n_986),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_SL g1382 ( 
.A(n_1326),
.B(n_934),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_SL g1383 ( 
.A(n_1327),
.B(n_954),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_SL g1384 ( 
.A(n_1334),
.B(n_959),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_SL g1385 ( 
.A(n_1335),
.B(n_961),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1344),
.B(n_880),
.Y(n_1386)
);

NAND2x1_ASAP7_75t_L g1387 ( 
.A(n_1313),
.B(n_792),
.Y(n_1387)
);

NAND2xp33_ASAP7_75t_SL g1388 ( 
.A(n_1296),
.B(n_889),
.Y(n_1388)
);

XNOR2xp5_ASAP7_75t_L g1389 ( 
.A(n_1267),
.B(n_890),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_SL g1390 ( 
.A(n_1349),
.B(n_1352),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1311),
.B(n_987),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1274),
.B(n_996),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_SL g1393 ( 
.A(n_1353),
.B(n_1355),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_SL g1394 ( 
.A(n_1357),
.B(n_967),
.Y(n_1394)
);

NAND2xp33_ASAP7_75t_SL g1395 ( 
.A(n_1266),
.B(n_912),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_SL g1396 ( 
.A(n_1359),
.B(n_980),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_SL g1397 ( 
.A(n_1360),
.B(n_1361),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_SL g1398 ( 
.A(n_1364),
.B(n_983),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_SL g1399 ( 
.A(n_1278),
.B(n_1006),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1272),
.B(n_918),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1281),
.B(n_1000),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1280),
.B(n_960),
.Y(n_1402)
);

NAND2xp33_ASAP7_75t_SL g1403 ( 
.A(n_1273),
.B(n_939),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_SL g1404 ( 
.A(n_1332),
.B(n_1011),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_SL g1405 ( 
.A(n_1350),
.B(n_1013),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_SL g1406 ( 
.A(n_1287),
.B(n_1018),
.Y(n_1406)
);

NAND2xp33_ASAP7_75t_SL g1407 ( 
.A(n_1320),
.B(n_1363),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_SL g1408 ( 
.A(n_1290),
.B(n_1021),
.Y(n_1408)
);

XNOR2xp5_ASAP7_75t_L g1409 ( 
.A(n_1307),
.B(n_943),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1324),
.B(n_1001),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_SL g1411 ( 
.A(n_1328),
.B(n_1024),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_SL g1412 ( 
.A(n_1331),
.B(n_1336),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_SL g1413 ( 
.A(n_1358),
.B(n_1029),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_SL g1414 ( 
.A(n_1289),
.B(n_1270),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_SL g1415 ( 
.A(n_1292),
.B(n_1031),
.Y(n_1415)
);

NAND2xp33_ASAP7_75t_SL g1416 ( 
.A(n_1294),
.B(n_976),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_SL g1417 ( 
.A(n_1269),
.B(n_1033),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_SL g1418 ( 
.A(n_1297),
.B(n_1037),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_SL g1419 ( 
.A(n_1298),
.B(n_1055),
.Y(n_1419)
);

NAND2xp33_ASAP7_75t_SL g1420 ( 
.A(n_1306),
.B(n_982),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_SL g1421 ( 
.A(n_1329),
.B(n_1067),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1288),
.B(n_1069),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1337),
.B(n_1046),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_SL g1424 ( 
.A(n_1277),
.B(n_1283),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_SL g1425 ( 
.A(n_1299),
.B(n_1083),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_SL g1426 ( 
.A(n_1286),
.B(n_1093),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_SL g1427 ( 
.A(n_1293),
.B(n_792),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_SL g1428 ( 
.A(n_1303),
.B(n_1072),
.Y(n_1428)
);

NAND2xp33_ASAP7_75t_SL g1429 ( 
.A(n_1308),
.B(n_1014),
.Y(n_1429)
);

NAND2xp33_ASAP7_75t_SL g1430 ( 
.A(n_1275),
.B(n_1019),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_SL g1431 ( 
.A(n_1323),
.B(n_1087),
.Y(n_1431)
);

NAND2xp33_ASAP7_75t_SL g1432 ( 
.A(n_1347),
.B(n_1023),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1356),
.B(n_777),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_SL g1434 ( 
.A(n_1305),
.B(n_1094),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1346),
.B(n_1097),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_SL g1436 ( 
.A(n_1340),
.B(n_810),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1366),
.B(n_932),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1284),
.B(n_781),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1310),
.B(n_1010),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_SL g1440 ( 
.A(n_1264),
.B(n_1295),
.Y(n_1440)
);

NAND2xp33_ASAP7_75t_SL g1441 ( 
.A(n_1304),
.B(n_1058),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_SL g1442 ( 
.A(n_1338),
.B(n_1341),
.Y(n_1442)
);

NAND2xp33_ASAP7_75t_SL g1443 ( 
.A(n_1310),
.B(n_1091),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_SL g1444 ( 
.A(n_1302),
.B(n_904),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_SL g1445 ( 
.A(n_1316),
.B(n_904),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1318),
.B(n_904),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_SL g1447 ( 
.A(n_1325),
.B(n_904),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_SL g1448 ( 
.A(n_1339),
.B(n_904),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_SL g1449 ( 
.A(n_1342),
.B(n_999),
.Y(n_1449)
);

AND2x4_ASAP7_75t_L g1450 ( 
.A(n_1271),
.B(n_964),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_SL g1451 ( 
.A(n_1343),
.B(n_999),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1348),
.B(n_1354),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_SL g1453 ( 
.A(n_1365),
.B(n_999),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_SL g1454 ( 
.A(n_1291),
.B(n_999),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1300),
.B(n_1022),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_SL g1456 ( 
.A(n_1309),
.B(n_999),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1276),
.B(n_784),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_SL g1458 ( 
.A(n_1330),
.B(n_789),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_SL g1459 ( 
.A(n_1321),
.B(n_791),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1333),
.B(n_796),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1333),
.B(n_800),
.Y(n_1461)
);

NAND2xp33_ASAP7_75t_SL g1462 ( 
.A(n_1315),
.B(n_815),
.Y(n_1462)
);

NAND2xp33_ASAP7_75t_SL g1463 ( 
.A(n_1315),
.B(n_818),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_SL g1464 ( 
.A(n_1321),
.B(n_820),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_SL g1465 ( 
.A(n_1321),
.B(n_821),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1321),
.B(n_822),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_SL g1467 ( 
.A(n_1321),
.B(n_826),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1321),
.B(n_829),
.Y(n_1468)
);

NAND2xp33_ASAP7_75t_SL g1469 ( 
.A(n_1315),
.B(n_832),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_SL g1470 ( 
.A(n_1321),
.B(n_833),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_SL g1471 ( 
.A(n_1321),
.B(n_841),
.Y(n_1471)
);

NAND2xp33_ASAP7_75t_SL g1472 ( 
.A(n_1315),
.B(n_843),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_SL g1473 ( 
.A(n_1321),
.B(n_845),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_SL g1474 ( 
.A(n_1321),
.B(n_851),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_1321),
.B(n_853),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_SL g1476 ( 
.A(n_1321),
.B(n_856),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_SL g1477 ( 
.A(n_1321),
.B(n_864),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_SL g1478 ( 
.A(n_1321),
.B(n_873),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1279),
.B(n_966),
.Y(n_1479)
);

NAND2xp33_ASAP7_75t_SL g1480 ( 
.A(n_1315),
.B(n_877),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_SL g1481 ( 
.A(n_1321),
.B(n_883),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_1321),
.B(n_893),
.Y(n_1482)
);

NAND2xp33_ASAP7_75t_SL g1483 ( 
.A(n_1315),
.B(n_894),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_SL g1484 ( 
.A(n_1321),
.B(n_902),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1321),
.B(n_905),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_SL g1486 ( 
.A(n_1321),
.B(n_910),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1285),
.B(n_915),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_SL g1488 ( 
.A(n_1321),
.B(n_929),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_SL g1489 ( 
.A(n_1321),
.B(n_931),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_SL g1490 ( 
.A(n_1321),
.B(n_935),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_SL g1491 ( 
.A(n_1321),
.B(n_936),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_SL g1492 ( 
.A(n_1321),
.B(n_938),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_SL g1493 ( 
.A(n_1321),
.B(n_940),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1285),
.B(n_944),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1279),
.B(n_968),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_SL g1496 ( 
.A(n_1321),
.B(n_947),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_SL g1497 ( 
.A(n_1321),
.B(n_949),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_SL g1498 ( 
.A(n_1321),
.B(n_950),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_1372),
.Y(n_1499)
);

CKINVDCx11_ASAP7_75t_R g1500 ( 
.A(n_1450),
.Y(n_1500)
);

BUFx2_ASAP7_75t_R g1501 ( 
.A(n_1440),
.Y(n_1501)
);

A2O1A1Ixp33_ASAP7_75t_L g1502 ( 
.A1(n_1391),
.A2(n_978),
.B(n_991),
.C(n_971),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1452),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1460),
.B(n_1461),
.Y(n_1504)
);

INVx3_ASAP7_75t_L g1505 ( 
.A(n_1402),
.Y(n_1505)
);

INVx2_ASAP7_75t_SL g1506 ( 
.A(n_1479),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1410),
.A2(n_1030),
.B(n_1028),
.Y(n_1507)
);

OAI22x1_ASAP7_75t_L g1508 ( 
.A1(n_1409),
.A2(n_952),
.B1(n_957),
.B2(n_951),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_SL g1509 ( 
.A1(n_1392),
.A2(n_913),
.B(n_811),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1495),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1495),
.Y(n_1511)
);

OAI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1414),
.A2(n_1039),
.B(n_1035),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1400),
.B(n_958),
.Y(n_1513)
);

OAI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1424),
.A2(n_1042),
.B(n_1040),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1412),
.A2(n_1073),
.B(n_1048),
.Y(n_1515)
);

AOI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1374),
.A2(n_1077),
.B(n_1075),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1390),
.Y(n_1517)
);

AOI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1376),
.A2(n_1081),
.B(n_1079),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1401),
.A2(n_1089),
.B(n_1082),
.Y(n_1519)
);

OAI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1369),
.A2(n_974),
.B(n_973),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1393),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1397),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_L g1523 ( 
.A1(n_1437),
.A2(n_1427),
.B(n_1387),
.Y(n_1523)
);

AOI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1371),
.A2(n_512),
.B(n_511),
.Y(n_1524)
);

OAI21x1_ASAP7_75t_L g1525 ( 
.A1(n_1435),
.A2(n_515),
.B(n_514),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1417),
.A2(n_519),
.B(n_518),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1381),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1455),
.Y(n_1528)
);

OA21x2_ASAP7_75t_L g1529 ( 
.A1(n_1444),
.A2(n_981),
.B(n_977),
.Y(n_1529)
);

INVx4_ASAP7_75t_L g1530 ( 
.A(n_1433),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1487),
.B(n_984),
.Y(n_1531)
);

OAI21x1_ASAP7_75t_L g1532 ( 
.A1(n_1421),
.A2(n_521),
.B(n_520),
.Y(n_1532)
);

AOI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1377),
.A2(n_525),
.B(n_523),
.Y(n_1533)
);

NAND2x1_ASAP7_75t_L g1534 ( 
.A(n_1439),
.B(n_526),
.Y(n_1534)
);

AO31x2_ASAP7_75t_L g1535 ( 
.A1(n_1423),
.A2(n_529),
.A3(n_530),
.B(n_528),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1375),
.A2(n_992),
.B1(n_994),
.B2(n_985),
.Y(n_1536)
);

A2O1A1Ixp33_ASAP7_75t_L g1537 ( 
.A1(n_1441),
.A2(n_997),
.B(n_998),
.C(n_995),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1426),
.A2(n_534),
.B(n_531),
.Y(n_1538)
);

INVx8_ASAP7_75t_L g1539 ( 
.A(n_1457),
.Y(n_1539)
);

BUFx12f_ASAP7_75t_L g1540 ( 
.A(n_1378),
.Y(n_1540)
);

AO21x2_ASAP7_75t_L g1541 ( 
.A1(n_1411),
.A2(n_538),
.B(n_536),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1494),
.A2(n_1008),
.B1(n_1009),
.B2(n_1004),
.Y(n_1542)
);

INVx2_ASAP7_75t_SL g1543 ( 
.A(n_1386),
.Y(n_1543)
);

NAND3x1_ASAP7_75t_L g1544 ( 
.A(n_1438),
.B(n_1016),
.C(n_1015),
.Y(n_1544)
);

NAND3xp33_ASAP7_75t_SL g1545 ( 
.A(n_1443),
.B(n_1020),
.C(n_1012),
.Y(n_1545)
);

INVx2_ASAP7_75t_SL g1546 ( 
.A(n_1428),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_L g1547 ( 
.A(n_1389),
.B(n_1459),
.Y(n_1547)
);

NAND2x1_ASAP7_75t_L g1548 ( 
.A(n_1407),
.B(n_541),
.Y(n_1548)
);

INVxp67_ASAP7_75t_SL g1549 ( 
.A(n_1379),
.Y(n_1549)
);

AO31x2_ASAP7_75t_L g1550 ( 
.A1(n_1445),
.A2(n_543),
.A3(n_544),
.B(n_542),
.Y(n_1550)
);

AOI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1382),
.A2(n_547),
.B(n_546),
.Y(n_1551)
);

OAI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1404),
.A2(n_1026),
.B(n_1025),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1446),
.Y(n_1553)
);

OAI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1415),
.A2(n_550),
.B(n_548),
.Y(n_1554)
);

AO31x2_ASAP7_75t_L g1555 ( 
.A1(n_1447),
.A2(n_553),
.A3(n_554),
.B(n_551),
.Y(n_1555)
);

BUFx10_ASAP7_75t_L g1556 ( 
.A(n_1403),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1464),
.B(n_1032),
.Y(n_1557)
);

OAI22x1_ASAP7_75t_L g1558 ( 
.A1(n_1465),
.A2(n_1038),
.B1(n_1043),
.B2(n_1034),
.Y(n_1558)
);

OAI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1405),
.A2(n_1047),
.B(n_1044),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1383),
.A2(n_559),
.B(n_556),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1466),
.B(n_1050),
.Y(n_1561)
);

INVx2_ASAP7_75t_SL g1562 ( 
.A(n_1436),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1467),
.B(n_1051),
.Y(n_1563)
);

AO21x2_ASAP7_75t_L g1564 ( 
.A1(n_1413),
.A2(n_563),
.B(n_562),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1448),
.Y(n_1565)
);

AO31x2_ASAP7_75t_L g1566 ( 
.A1(n_1449),
.A2(n_566),
.A3(n_570),
.B(n_564),
.Y(n_1566)
);

BUFx3_ASAP7_75t_L g1567 ( 
.A(n_1380),
.Y(n_1567)
);

AO31x2_ASAP7_75t_L g1568 ( 
.A1(n_1451),
.A2(n_1453),
.A3(n_1454),
.B(n_1456),
.Y(n_1568)
);

OAI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1418),
.A2(n_575),
.B(n_571),
.Y(n_1569)
);

NOR2xp67_ASAP7_75t_SL g1570 ( 
.A(n_1442),
.B(n_1434),
.Y(n_1570)
);

NAND2xp33_ASAP7_75t_L g1571 ( 
.A(n_1399),
.B(n_1086),
.Y(n_1571)
);

INVxp67_ASAP7_75t_SL g1572 ( 
.A(n_1384),
.Y(n_1572)
);

OAI21x1_ASAP7_75t_L g1573 ( 
.A1(n_1419),
.A2(n_578),
.B(n_576),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1373),
.B(n_1057),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_L g1575 ( 
.A(n_1468),
.B(n_1061),
.Y(n_1575)
);

AOI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1385),
.A2(n_581),
.B(n_580),
.Y(n_1576)
);

INVxp67_ASAP7_75t_SL g1577 ( 
.A(n_1394),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1470),
.B(n_1062),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1395),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1471),
.B(n_1063),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_SL g1581 ( 
.A(n_1388),
.B(n_1065),
.Y(n_1581)
);

AO22x2_ASAP7_75t_L g1582 ( 
.A1(n_1473),
.A2(n_1474),
.B1(n_1476),
.B2(n_1475),
.Y(n_1582)
);

O2A1O1Ixp33_ASAP7_75t_L g1583 ( 
.A1(n_1477),
.A2(n_1070),
.B(n_1071),
.C(n_1068),
.Y(n_1583)
);

BUFx3_ASAP7_75t_L g1584 ( 
.A(n_1420),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1431),
.Y(n_1585)
);

INVx3_ASAP7_75t_L g1586 ( 
.A(n_1462),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1396),
.A2(n_1090),
.B1(n_1092),
.B2(n_1085),
.Y(n_1587)
);

AOI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1398),
.A2(n_584),
.B(n_583),
.Y(n_1588)
);

AOI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1367),
.A2(n_586),
.B1(n_588),
.B2(n_585),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1425),
.A2(n_593),
.B(n_589),
.Y(n_1590)
);

BUFx3_ASAP7_75t_L g1591 ( 
.A(n_1463),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1478),
.B(n_2),
.Y(n_1592)
);

OAI21xp5_ASAP7_75t_L g1593 ( 
.A1(n_1481),
.A2(n_598),
.B(n_596),
.Y(n_1593)
);

OAI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1482),
.A2(n_601),
.B(n_600),
.Y(n_1594)
);

OAI21x1_ASAP7_75t_L g1595 ( 
.A1(n_1406),
.A2(n_606),
.B(n_605),
.Y(n_1595)
);

OAI21x1_ASAP7_75t_L g1596 ( 
.A1(n_1408),
.A2(n_609),
.B(n_607),
.Y(n_1596)
);

AO31x2_ASAP7_75t_L g1597 ( 
.A1(n_1469),
.A2(n_1472),
.A3(n_1483),
.B(n_1480),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1484),
.B(n_1485),
.Y(n_1598)
);

AOI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1368),
.A2(n_1370),
.B(n_1422),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1486),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1517),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1522),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_1540),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1521),
.Y(n_1604)
);

OR2x6_ASAP7_75t_L g1605 ( 
.A(n_1539),
.B(n_1488),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1504),
.B(n_1489),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1528),
.Y(n_1607)
);

INVx3_ASAP7_75t_L g1608 ( 
.A(n_1539),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1547),
.A2(n_1492),
.B1(n_1493),
.B2(n_1491),
.Y(n_1609)
);

INVx3_ASAP7_75t_L g1610 ( 
.A(n_1530),
.Y(n_1610)
);

NAND2x1p5_ASAP7_75t_L g1611 ( 
.A(n_1505),
.B(n_1490),
.Y(n_1611)
);

AO32x2_ASAP7_75t_L g1612 ( 
.A1(n_1542),
.A2(n_1546),
.A3(n_1587),
.B1(n_1536),
.B2(n_1506),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1527),
.Y(n_1613)
);

OAI21x1_ASAP7_75t_L g1614 ( 
.A1(n_1526),
.A2(n_1497),
.B(n_1496),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_1499),
.Y(n_1615)
);

AO21x2_ASAP7_75t_L g1616 ( 
.A1(n_1512),
.A2(n_1498),
.B(n_1458),
.Y(n_1616)
);

AOI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1598),
.A2(n_1429),
.B1(n_1416),
.B2(n_1430),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1510),
.Y(n_1618)
);

CKINVDCx20_ASAP7_75t_R g1619 ( 
.A(n_1500),
.Y(n_1619)
);

OAI21xp5_ASAP7_75t_L g1620 ( 
.A1(n_1599),
.A2(n_1432),
.B(n_612),
.Y(n_1620)
);

BUFx2_ASAP7_75t_L g1621 ( 
.A(n_1503),
.Y(n_1621)
);

NAND2x1p5_ASAP7_75t_L g1622 ( 
.A(n_1543),
.B(n_616),
.Y(n_1622)
);

OAI21x1_ASAP7_75t_L g1623 ( 
.A1(n_1532),
.A2(n_613),
.B(n_611),
.Y(n_1623)
);

AOI221xp5_ASAP7_75t_L g1624 ( 
.A1(n_1508),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.C(n_9),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_R g1625 ( 
.A(n_1545),
.B(n_617),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1511),
.Y(n_1626)
);

OAI21x1_ASAP7_75t_L g1627 ( 
.A1(n_1569),
.A2(n_1573),
.B(n_1538),
.Y(n_1627)
);

OA21x2_ASAP7_75t_L g1628 ( 
.A1(n_1507),
.A2(n_619),
.B(n_618),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1553),
.Y(n_1629)
);

AND2x4_ASAP7_75t_SL g1630 ( 
.A(n_1556),
.B(n_620),
.Y(n_1630)
);

BUFx2_ASAP7_75t_L g1631 ( 
.A(n_1567),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1575),
.A2(n_1578),
.B1(n_1579),
.B2(n_1584),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1565),
.Y(n_1633)
);

AOI21xp33_ASAP7_75t_L g1634 ( 
.A1(n_1583),
.A2(n_10),
.B(n_11),
.Y(n_1634)
);

INVxp67_ASAP7_75t_L g1635 ( 
.A(n_1600),
.Y(n_1635)
);

OAI21x1_ASAP7_75t_L g1636 ( 
.A1(n_1554),
.A2(n_622),
.B(n_621),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1592),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_1637)
);

INVx1_ASAP7_75t_SL g1638 ( 
.A(n_1501),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1568),
.Y(n_1639)
);

BUFx8_ASAP7_75t_SL g1640 ( 
.A(n_1591),
.Y(n_1640)
);

OAI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1595),
.A2(n_1596),
.B(n_1525),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1585),
.Y(n_1642)
);

OR2x6_ASAP7_75t_L g1643 ( 
.A(n_1548),
.B(n_630),
.Y(n_1643)
);

OAI21x1_ASAP7_75t_SL g1644 ( 
.A1(n_1509),
.A2(n_632),
.B(n_631),
.Y(n_1644)
);

BUFx2_ASAP7_75t_L g1645 ( 
.A(n_1529),
.Y(n_1645)
);

OAI21x1_ASAP7_75t_L g1646 ( 
.A1(n_1524),
.A2(n_638),
.B(n_637),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1586),
.B(n_640),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1562),
.Y(n_1648)
);

OAI21x1_ASAP7_75t_L g1649 ( 
.A1(n_1534),
.A2(n_642),
.B(n_641),
.Y(n_1649)
);

OR2x6_ASAP7_75t_L g1650 ( 
.A(n_1582),
.B(n_643),
.Y(n_1650)
);

OAI21x1_ASAP7_75t_L g1651 ( 
.A1(n_1593),
.A2(n_646),
.B(n_644),
.Y(n_1651)
);

OA21x2_ASAP7_75t_L g1652 ( 
.A1(n_1594),
.A2(n_649),
.B(n_647),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1549),
.A2(n_20),
.B1(n_17),
.B2(n_18),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1561),
.B(n_21),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1550),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1580),
.B(n_22),
.Y(n_1656)
);

AOI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1572),
.A2(n_651),
.B(n_650),
.Y(n_1657)
);

OAI21x1_ASAP7_75t_L g1658 ( 
.A1(n_1533),
.A2(n_653),
.B(n_652),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_1558),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1577),
.B(n_22),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1550),
.Y(n_1661)
);

OAI21x1_ASAP7_75t_L g1662 ( 
.A1(n_1551),
.A2(n_655),
.B(n_654),
.Y(n_1662)
);

OAI21x1_ASAP7_75t_L g1663 ( 
.A1(n_1560),
.A2(n_1588),
.B(n_1576),
.Y(n_1663)
);

OAI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1557),
.A2(n_662),
.B(n_661),
.Y(n_1664)
);

OAI21x1_ASAP7_75t_L g1665 ( 
.A1(n_1590),
.A2(n_666),
.B(n_663),
.Y(n_1665)
);

OAI21x1_ASAP7_75t_L g1666 ( 
.A1(n_1514),
.A2(n_668),
.B(n_667),
.Y(n_1666)
);

OAI21x1_ASAP7_75t_L g1667 ( 
.A1(n_1515),
.A2(n_1516),
.B(n_1518),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1555),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1531),
.B(n_23),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1597),
.B(n_669),
.Y(n_1670)
);

OAI21x1_ASAP7_75t_L g1671 ( 
.A1(n_1589),
.A2(n_1563),
.B(n_1559),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1520),
.B(n_24),
.Y(n_1672)
);

OAI21x1_ASAP7_75t_L g1673 ( 
.A1(n_1552),
.A2(n_671),
.B(n_670),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1555),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1502),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1570),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1537),
.B(n_24),
.Y(n_1677)
);

AOI21x1_ASAP7_75t_L g1678 ( 
.A1(n_1581),
.A2(n_673),
.B(n_672),
.Y(n_1678)
);

OAI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1571),
.A2(n_677),
.B(n_674),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1574),
.B(n_25),
.Y(n_1680)
);

INVx2_ASAP7_75t_SL g1681 ( 
.A(n_1566),
.Y(n_1681)
);

AO31x2_ASAP7_75t_L g1682 ( 
.A1(n_1535),
.A2(n_1566),
.A3(n_1564),
.B(n_1541),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1544),
.Y(n_1683)
);

OAI21x1_ASAP7_75t_L g1684 ( 
.A1(n_1523),
.A2(n_679),
.B(n_678),
.Y(n_1684)
);

AOI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1547),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_1685)
);

NAND2x1p5_ASAP7_75t_L g1686 ( 
.A(n_1505),
.B(n_684),
.Y(n_1686)
);

OA21x2_ASAP7_75t_L g1687 ( 
.A1(n_1519),
.A2(n_681),
.B(n_680),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1517),
.Y(n_1688)
);

OAI21x1_ASAP7_75t_L g1689 ( 
.A1(n_1523),
.A2(n_683),
.B(n_682),
.Y(n_1689)
);

OA21x2_ASAP7_75t_L g1690 ( 
.A1(n_1519),
.A2(n_686),
.B(n_685),
.Y(n_1690)
);

AOI221xp5_ASAP7_75t_L g1691 ( 
.A1(n_1513),
.A2(n_30),
.B1(n_27),
.B2(n_29),
.C(n_31),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1547),
.A2(n_32),
.B1(n_29),
.B2(n_30),
.Y(n_1692)
);

OA21x2_ASAP7_75t_L g1693 ( 
.A1(n_1519),
.A2(n_688),
.B(n_687),
.Y(n_1693)
);

AOI221xp5_ASAP7_75t_L g1694 ( 
.A1(n_1513),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.C(n_35),
.Y(n_1694)
);

INVx3_ASAP7_75t_L g1695 ( 
.A(n_1540),
.Y(n_1695)
);

NAND2x1p5_ASAP7_75t_L g1696 ( 
.A(n_1505),
.B(n_690),
.Y(n_1696)
);

INVx6_ASAP7_75t_L g1697 ( 
.A(n_1540),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1613),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1601),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1602),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1604),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1654),
.B(n_37),
.Y(n_1702)
);

OAI21x1_ASAP7_75t_L g1703 ( 
.A1(n_1627),
.A2(n_693),
.B(n_692),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1688),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1606),
.B(n_38),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1642),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1607),
.Y(n_1707)
);

HB1xp67_ASAP7_75t_L g1708 ( 
.A(n_1621),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1629),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1633),
.Y(n_1710)
);

AND2x4_ASAP7_75t_L g1711 ( 
.A(n_1608),
.B(n_695),
.Y(n_1711)
);

OAI21x1_ASAP7_75t_L g1712 ( 
.A1(n_1641),
.A2(n_697),
.B(n_696),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1626),
.Y(n_1713)
);

AOI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1672),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_1714)
);

AND2x4_ASAP7_75t_L g1715 ( 
.A(n_1610),
.B(n_698),
.Y(n_1715)
);

NAND2x1p5_ASAP7_75t_L g1716 ( 
.A(n_1631),
.B(n_701),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1635),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_1640),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1618),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1676),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1648),
.Y(n_1721)
);

OA21x2_ASAP7_75t_L g1722 ( 
.A1(n_1655),
.A2(n_706),
.B(n_703),
.Y(n_1722)
);

INVx3_ASAP7_75t_L g1723 ( 
.A(n_1697),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1660),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1656),
.B(n_40),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1677),
.Y(n_1726)
);

OAI21xp33_ASAP7_75t_L g1727 ( 
.A1(n_1669),
.A2(n_42),
.B(n_44),
.Y(n_1727)
);

OAI21x1_ASAP7_75t_L g1728 ( 
.A1(n_1684),
.A2(n_708),
.B(n_707),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1639),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1675),
.Y(n_1730)
);

AOI21x1_ASAP7_75t_L g1731 ( 
.A1(n_1674),
.A2(n_713),
.B(n_711),
.Y(n_1731)
);

OAI211xp5_ASAP7_75t_L g1732 ( 
.A1(n_1624),
.A2(n_1691),
.B(n_1694),
.C(n_1685),
.Y(n_1732)
);

AOI21x1_ASAP7_75t_L g1733 ( 
.A1(n_1645),
.A2(n_716),
.B(n_714),
.Y(n_1733)
);

NAND2x1_ASAP7_75t_L g1734 ( 
.A(n_1643),
.B(n_717),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1611),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1695),
.B(n_718),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1689),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1612),
.Y(n_1738)
);

INVx2_ASAP7_75t_SL g1739 ( 
.A(n_1615),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1680),
.Y(n_1740)
);

OAI222xp33_ASAP7_75t_L g1741 ( 
.A1(n_1692),
.A2(n_47),
.B1(n_49),
.B2(n_45),
.C1(n_46),
.C2(n_48),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_1619),
.Y(n_1742)
);

INVx2_ASAP7_75t_SL g1743 ( 
.A(n_1603),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1670),
.Y(n_1744)
);

AOI21x1_ASAP7_75t_L g1745 ( 
.A1(n_1661),
.A2(n_720),
.B(n_719),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1632),
.B(n_48),
.Y(n_1746)
);

OAI21x1_ASAP7_75t_L g1747 ( 
.A1(n_1663),
.A2(n_722),
.B(n_721),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1668),
.Y(n_1748)
);

BUFx6f_ASAP7_75t_L g1749 ( 
.A(n_1605),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1647),
.Y(n_1750)
);

OAI21xp5_ASAP7_75t_L g1751 ( 
.A1(n_1620),
.A2(n_50),
.B(n_51),
.Y(n_1751)
);

INVx3_ASAP7_75t_L g1752 ( 
.A(n_1630),
.Y(n_1752)
);

INVx3_ASAP7_75t_L g1753 ( 
.A(n_1622),
.Y(n_1753)
);

INVx2_ASAP7_75t_SL g1754 ( 
.A(n_1638),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1678),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1617),
.B(n_52),
.Y(n_1756)
);

AND2x4_ASAP7_75t_L g1757 ( 
.A(n_1683),
.B(n_724),
.Y(n_1757)
);

NAND2xp33_ASAP7_75t_R g1758 ( 
.A(n_1742),
.B(n_1625),
.Y(n_1758)
);

INVxp67_ASAP7_75t_L g1759 ( 
.A(n_1708),
.Y(n_1759)
);

AND2x4_ASAP7_75t_L g1760 ( 
.A(n_1750),
.B(n_1643),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_R g1761 ( 
.A(n_1752),
.B(n_1659),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1724),
.B(n_1609),
.Y(n_1762)
);

INVxp67_ASAP7_75t_L g1763 ( 
.A(n_1717),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1707),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1744),
.B(n_1650),
.Y(n_1765)
);

NAND2xp33_ASAP7_75t_R g1766 ( 
.A(n_1718),
.B(n_1652),
.Y(n_1766)
);

OR2x6_ASAP7_75t_L g1767 ( 
.A(n_1716),
.B(n_1686),
.Y(n_1767)
);

NAND2xp33_ASAP7_75t_R g1768 ( 
.A(n_1723),
.B(n_1687),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1699),
.Y(n_1769)
);

INVxp67_ASAP7_75t_L g1770 ( 
.A(n_1721),
.Y(n_1770)
);

CKINVDCx16_ASAP7_75t_R g1771 ( 
.A(n_1739),
.Y(n_1771)
);

BUFx3_ASAP7_75t_L g1772 ( 
.A(n_1743),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_R g1773 ( 
.A(n_1753),
.B(n_1681),
.Y(n_1773)
);

NAND2xp33_ASAP7_75t_R g1774 ( 
.A(n_1757),
.B(n_1690),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1726),
.B(n_1637),
.Y(n_1775)
);

OR2x6_ASAP7_75t_L g1776 ( 
.A(n_1734),
.B(n_1696),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1709),
.Y(n_1777)
);

INVxp67_ASAP7_75t_L g1778 ( 
.A(n_1740),
.Y(n_1778)
);

NAND2xp33_ASAP7_75t_R g1779 ( 
.A(n_1756),
.B(n_1693),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1749),
.B(n_1649),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_R g1781 ( 
.A(n_1754),
.B(n_725),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1746),
.B(n_1705),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1701),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_1749),
.B(n_1614),
.Y(n_1784)
);

AND2x4_ASAP7_75t_L g1785 ( 
.A(n_1735),
.B(n_1657),
.Y(n_1785)
);

XNOR2xp5_ASAP7_75t_L g1786 ( 
.A(n_1736),
.B(n_1653),
.Y(n_1786)
);

AND2x4_ASAP7_75t_L g1787 ( 
.A(n_1711),
.B(n_1658),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1702),
.B(n_1634),
.Y(n_1788)
);

NAND2xp33_ASAP7_75t_R g1789 ( 
.A(n_1715),
.B(n_1628),
.Y(n_1789)
);

NAND2xp33_ASAP7_75t_R g1790 ( 
.A(n_1725),
.B(n_1664),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_L g1791 ( 
.A(n_1698),
.B(n_1616),
.Y(n_1791)
);

AND2x4_ASAP7_75t_L g1792 ( 
.A(n_1719),
.B(n_1662),
.Y(n_1792)
);

AND2x4_ASAP7_75t_L g1793 ( 
.A(n_1700),
.B(n_1665),
.Y(n_1793)
);

NOR2x1_ASAP7_75t_L g1794 ( 
.A(n_1720),
.B(n_1679),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1764),
.Y(n_1795)
);

OAI22xp5_ASAP7_75t_L g1796 ( 
.A1(n_1762),
.A2(n_1732),
.B1(n_1714),
.B2(n_1751),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1782),
.B(n_1704),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_SL g1798 ( 
.A(n_1771),
.B(n_1741),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1763),
.B(n_1706),
.Y(n_1799)
);

CKINVDCx16_ASAP7_75t_R g1800 ( 
.A(n_1761),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1769),
.Y(n_1801)
);

BUFx2_ASAP7_75t_L g1802 ( 
.A(n_1773),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1759),
.B(n_1710),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1783),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1778),
.B(n_1713),
.Y(n_1805)
);

INVxp67_ASAP7_75t_SL g1806 ( 
.A(n_1791),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1788),
.B(n_1738),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1770),
.B(n_1729),
.Y(n_1808)
);

INVx3_ASAP7_75t_L g1809 ( 
.A(n_1765),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1777),
.B(n_1727),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1792),
.Y(n_1811)
);

INVx1_ASAP7_75t_SL g1812 ( 
.A(n_1772),
.Y(n_1812)
);

NOR2x1_ASAP7_75t_L g1813 ( 
.A(n_1794),
.B(n_1730),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1784),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1793),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1780),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1785),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1775),
.B(n_1748),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1760),
.B(n_1787),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1767),
.B(n_1755),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1767),
.B(n_1682),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1776),
.Y(n_1822)
);

AND2x2_ASAP7_75t_SL g1823 ( 
.A(n_1790),
.B(n_1722),
.Y(n_1823)
);

HB1xp67_ASAP7_75t_L g1824 ( 
.A(n_1779),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1776),
.Y(n_1825)
);

INVxp67_ASAP7_75t_L g1826 ( 
.A(n_1758),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1786),
.B(n_1733),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1766),
.B(n_1682),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1781),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1768),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1774),
.B(n_1671),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1789),
.B(n_1733),
.Y(n_1832)
);

INVx2_ASAP7_75t_SL g1833 ( 
.A(n_1812),
.Y(n_1833)
);

AOI22xp33_ASAP7_75t_L g1834 ( 
.A1(n_1796),
.A2(n_1644),
.B1(n_1667),
.B2(n_1673),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1795),
.Y(n_1835)
);

NOR2x1_ASAP7_75t_L g1836 ( 
.A(n_1813),
.B(n_1722),
.Y(n_1836)
);

BUFx6f_ASAP7_75t_L g1837 ( 
.A(n_1802),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1806),
.B(n_1737),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1801),
.Y(n_1839)
);

AOI33xp33_ASAP7_75t_L g1840 ( 
.A1(n_1827),
.A2(n_56),
.A3(n_58),
.B1(n_54),
.B2(n_55),
.B3(n_57),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1805),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1824),
.B(n_1747),
.Y(n_1842)
);

AOI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1817),
.A2(n_1651),
.B1(n_1666),
.B2(n_1728),
.Y(n_1843)
);

AOI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1817),
.A2(n_1646),
.B1(n_1712),
.B2(n_1703),
.Y(n_1844)
);

NAND4xp25_ASAP7_75t_L g1845 ( 
.A(n_1799),
.B(n_58),
.C(n_56),
.D(n_57),
.Y(n_1845)
);

INVx1_ASAP7_75t_SL g1846 ( 
.A(n_1829),
.Y(n_1846)
);

NOR2x1_ASAP7_75t_L g1847 ( 
.A(n_1830),
.B(n_1731),
.Y(n_1847)
);

AND2x4_ASAP7_75t_L g1848 ( 
.A(n_1814),
.B(n_1816),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1808),
.Y(n_1849)
);

OAI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1826),
.A2(n_1745),
.B1(n_1636),
.B2(n_1623),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1797),
.B(n_59),
.Y(n_1851)
);

INVx1_ASAP7_75t_SL g1852 ( 
.A(n_1819),
.Y(n_1852)
);

AOI21xp5_ASAP7_75t_L g1853 ( 
.A1(n_1823),
.A2(n_59),
.B(n_60),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1803),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1822),
.A2(n_64),
.B1(n_61),
.B2(n_63),
.Y(n_1855)
);

BUFx3_ASAP7_75t_L g1856 ( 
.A(n_1809),
.Y(n_1856)
);

AND2x2_ASAP7_75t_SL g1857 ( 
.A(n_1800),
.B(n_65),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_SL g1858 ( 
.A(n_1825),
.B(n_728),
.Y(n_1858)
);

INVx1_ASAP7_75t_SL g1859 ( 
.A(n_1820),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1811),
.B(n_66),
.Y(n_1860)
);

AOI221xp5_ASAP7_75t_L g1861 ( 
.A1(n_1810),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.C(n_70),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1815),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1821),
.Y(n_1863)
);

INVx3_ASAP7_75t_L g1864 ( 
.A(n_1828),
.Y(n_1864)
);

AOI22xp33_ASAP7_75t_L g1865 ( 
.A1(n_1832),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1818),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1831),
.B(n_71),
.Y(n_1867)
);

HB1xp67_ASAP7_75t_L g1868 ( 
.A(n_1824),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1807),
.B(n_73),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1807),
.B(n_73),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1807),
.B(n_74),
.Y(n_1871)
);

AOI221xp5_ASAP7_75t_L g1872 ( 
.A1(n_1796),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.C(n_78),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1804),
.Y(n_1873)
);

AOI22xp33_ASAP7_75t_SL g1874 ( 
.A1(n_1798),
.A2(n_79),
.B1(n_76),
.B2(n_78),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1807),
.B(n_80),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1795),
.Y(n_1876)
);

HB1xp67_ASAP7_75t_L g1877 ( 
.A(n_1824),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1795),
.Y(n_1878)
);

NOR2xp33_ASAP7_75t_L g1879 ( 
.A(n_1826),
.B(n_81),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1795),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1864),
.B(n_85),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1868),
.B(n_86),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1835),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1877),
.B(n_87),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1866),
.B(n_87),
.Y(n_1885)
);

AND2x4_ASAP7_75t_L g1886 ( 
.A(n_1856),
.B(n_88),
.Y(n_1886)
);

INVx4_ASAP7_75t_R g1887 ( 
.A(n_1833),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1876),
.Y(n_1888)
);

NOR2xp67_ASAP7_75t_L g1889 ( 
.A(n_1863),
.B(n_89),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1839),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1852),
.B(n_90),
.Y(n_1891)
);

AND2x4_ASAP7_75t_L g1892 ( 
.A(n_1848),
.B(n_91),
.Y(n_1892)
);

INVx3_ASAP7_75t_L g1893 ( 
.A(n_1837),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1878),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1880),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1841),
.B(n_92),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1849),
.B(n_94),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1854),
.B(n_94),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_SL g1899 ( 
.A(n_1857),
.B(n_95),
.Y(n_1899)
);

OR2x2_ASAP7_75t_L g1900 ( 
.A(n_1873),
.B(n_96),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1862),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1846),
.B(n_100),
.Y(n_1902)
);

OAI32xp33_ASAP7_75t_L g1903 ( 
.A1(n_1845),
.A2(n_104),
.A3(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_1903)
);

OR3x2_ASAP7_75t_L g1904 ( 
.A(n_1867),
.B(n_104),
.C(n_105),
.Y(n_1904)
);

OR2x2_ASAP7_75t_L g1905 ( 
.A(n_1838),
.B(n_107),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1842),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1836),
.Y(n_1907)
);

INVx2_ASAP7_75t_SL g1908 ( 
.A(n_1860),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1869),
.B(n_109),
.Y(n_1909)
);

OR2x2_ASAP7_75t_L g1910 ( 
.A(n_1851),
.B(n_110),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1870),
.B(n_110),
.Y(n_1911)
);

INVx1_ASAP7_75t_SL g1912 ( 
.A(n_1871),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1875),
.B(n_112),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1847),
.Y(n_1914)
);

AND2x4_ASAP7_75t_L g1915 ( 
.A(n_1853),
.B(n_112),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1879),
.B(n_113),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1850),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1865),
.B(n_114),
.Y(n_1918)
);

OR2x2_ASAP7_75t_L g1919 ( 
.A(n_1834),
.B(n_115),
.Y(n_1919)
);

NOR2xp33_ASAP7_75t_SL g1920 ( 
.A(n_1874),
.B(n_116),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1872),
.B(n_116),
.Y(n_1921)
);

BUFx2_ASAP7_75t_L g1922 ( 
.A(n_1861),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1858),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1843),
.B(n_1855),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1844),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1859),
.B(n_117),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1835),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1839),
.Y(n_1928)
);

OR2x2_ASAP7_75t_L g1929 ( 
.A(n_1864),
.B(n_118),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1835),
.Y(n_1930)
);

INVx1_ASAP7_75t_SL g1931 ( 
.A(n_1837),
.Y(n_1931)
);

OR2x2_ASAP7_75t_L g1932 ( 
.A(n_1864),
.B(n_119),
.Y(n_1932)
);

HB1xp67_ASAP7_75t_L g1933 ( 
.A(n_1868),
.Y(n_1933)
);

NAND3xp33_ASAP7_75t_L g1934 ( 
.A(n_1872),
.B(n_120),
.C(n_121),
.Y(n_1934)
);

NOR2x1_ASAP7_75t_L g1935 ( 
.A(n_1836),
.B(n_122),
.Y(n_1935)
);

NAND4xp25_ASAP7_75t_L g1936 ( 
.A(n_1840),
.B(n_126),
.C(n_124),
.D(n_125),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1859),
.B(n_124),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1839),
.Y(n_1938)
);

AND2x4_ASAP7_75t_L g1939 ( 
.A(n_1856),
.B(n_127),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1835),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1859),
.B(n_130),
.Y(n_1941)
);

INVxp67_ASAP7_75t_L g1942 ( 
.A(n_1868),
.Y(n_1942)
);

CKINVDCx8_ASAP7_75t_R g1943 ( 
.A(n_1886),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1883),
.Y(n_1944)
);

AO221x2_ASAP7_75t_L g1945 ( 
.A1(n_1934),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.C(n_135),
.Y(n_1945)
);

OAI22xp33_ASAP7_75t_L g1946 ( 
.A1(n_1922),
.A2(n_140),
.B1(n_137),
.B2(n_138),
.Y(n_1946)
);

CKINVDCx5p33_ASAP7_75t_R g1947 ( 
.A(n_1931),
.Y(n_1947)
);

CKINVDCx5p33_ASAP7_75t_R g1948 ( 
.A(n_1893),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1942),
.B(n_138),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1917),
.B(n_141),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1906),
.B(n_141),
.Y(n_1951)
);

INVx2_ASAP7_75t_SL g1952 ( 
.A(n_1887),
.Y(n_1952)
);

INVxp67_ASAP7_75t_L g1953 ( 
.A(n_1935),
.Y(n_1953)
);

AO221x2_ASAP7_75t_L g1954 ( 
.A1(n_1904),
.A2(n_145),
.B1(n_147),
.B2(n_144),
.C(n_146),
.Y(n_1954)
);

NOR2x1_ASAP7_75t_L g1955 ( 
.A(n_1907),
.B(n_145),
.Y(n_1955)
);

AO221x2_ASAP7_75t_L g1956 ( 
.A1(n_1924),
.A2(n_148),
.B1(n_150),
.B2(n_147),
.C(n_149),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1888),
.B(n_146),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1894),
.B(n_149),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1895),
.B(n_150),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1927),
.B(n_151),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1930),
.Y(n_1961)
);

CKINVDCx5p33_ASAP7_75t_R g1962 ( 
.A(n_1939),
.Y(n_1962)
);

NAND2xp33_ASAP7_75t_SL g1963 ( 
.A(n_1902),
.B(n_153),
.Y(n_1963)
);

INVx2_ASAP7_75t_SL g1964 ( 
.A(n_1908),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1940),
.Y(n_1965)
);

NOR2x1_ASAP7_75t_L g1966 ( 
.A(n_1914),
.B(n_154),
.Y(n_1966)
);

OR2x2_ASAP7_75t_L g1967 ( 
.A(n_1901),
.B(n_156),
.Y(n_1967)
);

OAI22xp33_ASAP7_75t_L g1968 ( 
.A1(n_1936),
.A2(n_1920),
.B1(n_1919),
.B2(n_1921),
.Y(n_1968)
);

NOR2xp33_ASAP7_75t_SL g1969 ( 
.A(n_1889),
.B(n_156),
.Y(n_1969)
);

NAND2xp33_ASAP7_75t_SL g1970 ( 
.A(n_1891),
.B(n_157),
.Y(n_1970)
);

INVxp67_ASAP7_75t_L g1971 ( 
.A(n_1905),
.Y(n_1971)
);

INVx3_ASAP7_75t_L g1972 ( 
.A(n_1890),
.Y(n_1972)
);

INVxp67_ASAP7_75t_L g1973 ( 
.A(n_1885),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1928),
.B(n_1938),
.Y(n_1974)
);

AOI221xp5_ASAP7_75t_L g1975 ( 
.A1(n_1903),
.A2(n_162),
.B1(n_160),
.B2(n_161),
.C(n_163),
.Y(n_1975)
);

AO221x2_ASAP7_75t_L g1976 ( 
.A1(n_1918),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.C(n_167),
.Y(n_1976)
);

AO221x2_ASAP7_75t_L g1977 ( 
.A1(n_1898),
.A2(n_1923),
.B1(n_1915),
.B2(n_1912),
.C(n_1882),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_1892),
.Y(n_1978)
);

AOI22xp5_ASAP7_75t_SL g1979 ( 
.A1(n_1884),
.A2(n_173),
.B1(n_174),
.B2(n_172),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1897),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1881),
.B(n_1929),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1932),
.B(n_171),
.Y(n_1982)
);

CKINVDCx5p33_ASAP7_75t_R g1983 ( 
.A(n_1926),
.Y(n_1983)
);

NAND2xp33_ASAP7_75t_SL g1984 ( 
.A(n_1937),
.B(n_1941),
.Y(n_1984)
);

AO221x2_ASAP7_75t_L g1985 ( 
.A1(n_1916),
.A2(n_178),
.B1(n_175),
.B2(n_177),
.C(n_179),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1900),
.Y(n_1986)
);

INVx3_ASAP7_75t_L g1987 ( 
.A(n_1896),
.Y(n_1987)
);

OAI22xp33_ASAP7_75t_L g1988 ( 
.A1(n_1910),
.A2(n_1911),
.B1(n_1913),
.B2(n_1909),
.Y(n_1988)
);

NOR2x1_ASAP7_75t_L g1989 ( 
.A(n_1935),
.B(n_180),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1933),
.B(n_180),
.Y(n_1990)
);

OR2x2_ASAP7_75t_L g1991 ( 
.A(n_1906),
.B(n_181),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1933),
.B(n_182),
.Y(n_1992)
);

NOR2xp67_ASAP7_75t_L g1993 ( 
.A(n_1907),
.B(n_184),
.Y(n_1993)
);

NOR2x1_ASAP7_75t_L g1994 ( 
.A(n_1935),
.B(n_186),
.Y(n_1994)
);

AOI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1922),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.Y(n_1995)
);

NAND2xp33_ASAP7_75t_R g1996 ( 
.A(n_1922),
.B(n_190),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_SL g1997 ( 
.A(n_1925),
.B(n_191),
.Y(n_1997)
);

NOR4xp25_ASAP7_75t_SL g1998 ( 
.A(n_1907),
.B(n_193),
.C(n_191),
.D(n_192),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1933),
.B(n_193),
.Y(n_1999)
);

NOR2xp33_ASAP7_75t_SL g2000 ( 
.A(n_1899),
.B(n_197),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1933),
.B(n_199),
.Y(n_2001)
);

NAND2xp33_ASAP7_75t_R g2002 ( 
.A(n_1922),
.B(n_200),
.Y(n_2002)
);

INVx1_ASAP7_75t_SL g2003 ( 
.A(n_1952),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1977),
.B(n_201),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1972),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1944),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1986),
.B(n_1987),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1961),
.Y(n_2008)
);

INVx4_ASAP7_75t_L g2009 ( 
.A(n_1947),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1980),
.B(n_202),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1964),
.B(n_203),
.Y(n_2011)
);

AOI22xp33_ASAP7_75t_L g2012 ( 
.A1(n_1954),
.A2(n_1968),
.B1(n_1945),
.B2(n_1956),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_SL g2013 ( 
.A(n_1969),
.B(n_204),
.Y(n_2013)
);

AOI22xp33_ASAP7_75t_L g2014 ( 
.A1(n_1945),
.A2(n_206),
.B1(n_204),
.B2(n_205),
.Y(n_2014)
);

INVx1_ASAP7_75t_SL g2015 ( 
.A(n_1984),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1965),
.Y(n_2016)
);

AOI22xp33_ASAP7_75t_L g2017 ( 
.A1(n_1976),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1951),
.B(n_207),
.Y(n_2018)
);

OR2x2_ASAP7_75t_L g2019 ( 
.A(n_1981),
.B(n_208),
.Y(n_2019)
);

INVx1_ASAP7_75t_SL g2020 ( 
.A(n_1983),
.Y(n_2020)
);

INVx1_ASAP7_75t_SL g2021 ( 
.A(n_1970),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1950),
.B(n_209),
.Y(n_2022)
);

OAI21x1_ASAP7_75t_SL g2023 ( 
.A1(n_1955),
.A2(n_210),
.B(n_211),
.Y(n_2023)
);

INVx1_ASAP7_75t_SL g2024 ( 
.A(n_1963),
.Y(n_2024)
);

OAI21x1_ASAP7_75t_L g2025 ( 
.A1(n_1974),
.A2(n_212),
.B(n_213),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1967),
.Y(n_2026)
);

INVx1_ASAP7_75t_SL g2027 ( 
.A(n_1948),
.Y(n_2027)
);

OR2x2_ASAP7_75t_L g2028 ( 
.A(n_1991),
.B(n_212),
.Y(n_2028)
);

AOI22xp33_ASAP7_75t_L g2029 ( 
.A1(n_1976),
.A2(n_216),
.B1(n_214),
.B2(n_215),
.Y(n_2029)
);

OAI21x1_ASAP7_75t_L g2030 ( 
.A1(n_1966),
.A2(n_1992),
.B(n_1990),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1957),
.B(n_217),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1943),
.Y(n_2032)
);

INVxp67_ASAP7_75t_L g2033 ( 
.A(n_2002),
.Y(n_2033)
);

BUFx3_ASAP7_75t_L g2034 ( 
.A(n_1962),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1958),
.B(n_219),
.Y(n_2035)
);

NOR2xp33_ASAP7_75t_SL g2036 ( 
.A(n_1989),
.B(n_220),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1959),
.B(n_220),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1960),
.B(n_221),
.Y(n_2038)
);

INVxp67_ASAP7_75t_L g2039 ( 
.A(n_1994),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1999),
.B(n_223),
.Y(n_2040)
);

AND3x2_ASAP7_75t_L g2041 ( 
.A(n_1975),
.B(n_224),
.C(n_225),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1978),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_2001),
.B(n_229),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1949),
.B(n_231),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1982),
.Y(n_2045)
);

AND4x1_ASAP7_75t_L g2046 ( 
.A(n_1995),
.B(n_235),
.C(n_233),
.D(n_234),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1988),
.B(n_1997),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1985),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1979),
.Y(n_2049)
);

HB1xp67_ASAP7_75t_L g2050 ( 
.A(n_1946),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1998),
.B(n_238),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1944),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_1952),
.B(n_240),
.Y(n_2053)
);

INVx1_ASAP7_75t_SL g2054 ( 
.A(n_1952),
.Y(n_2054)
);

INVx1_ASAP7_75t_SL g2055 ( 
.A(n_1952),
.Y(n_2055)
);

NOR2xp33_ASAP7_75t_L g2056 ( 
.A(n_1973),
.B(n_241),
.Y(n_2056)
);

OR2x2_ASAP7_75t_L g2057 ( 
.A(n_1971),
.B(n_243),
.Y(n_2057)
);

AND3x1_ASAP7_75t_L g2058 ( 
.A(n_2000),
.B(n_245),
.C(n_246),
.Y(n_2058)
);

OR2x2_ASAP7_75t_L g2059 ( 
.A(n_1971),
.B(n_247),
.Y(n_2059)
);

BUFx2_ASAP7_75t_L g2060 ( 
.A(n_1952),
.Y(n_2060)
);

AOI22xp33_ASAP7_75t_L g2061 ( 
.A1(n_1954),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.Y(n_2061)
);

NOR2xp67_ASAP7_75t_L g2062 ( 
.A(n_1953),
.B(n_249),
.Y(n_2062)
);

NOR2x1_ASAP7_75t_L g2063 ( 
.A(n_1993),
.B(n_251),
.Y(n_2063)
);

INVx1_ASAP7_75t_SL g2064 ( 
.A(n_1952),
.Y(n_2064)
);

NOR2xp33_ASAP7_75t_L g2065 ( 
.A(n_1973),
.B(n_252),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1944),
.Y(n_2066)
);

HB1xp67_ASAP7_75t_L g2067 ( 
.A(n_1953),
.Y(n_2067)
);

AOI22xp33_ASAP7_75t_L g2068 ( 
.A1(n_1954),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.Y(n_2068)
);

INVx1_ASAP7_75t_SL g2069 ( 
.A(n_1952),
.Y(n_2069)
);

AND3x1_ASAP7_75t_L g2070 ( 
.A(n_2000),
.B(n_256),
.C(n_258),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_1973),
.B(n_258),
.Y(n_2071)
);

INVx1_ASAP7_75t_SL g2072 ( 
.A(n_1952),
.Y(n_2072)
);

NAND2x1p5_ASAP7_75t_L g2073 ( 
.A(n_1952),
.B(n_260),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_1952),
.B(n_261),
.Y(n_2074)
);

NAND3xp33_ASAP7_75t_L g2075 ( 
.A(n_1996),
.B(n_262),
.C(n_264),
.Y(n_2075)
);

AOI222xp33_ASAP7_75t_L g2076 ( 
.A1(n_1968),
.A2(n_267),
.B1(n_269),
.B2(n_265),
.C1(n_266),
.C2(n_268),
.Y(n_2076)
);

INVx2_ASAP7_75t_SL g2077 ( 
.A(n_2060),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2006),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2039),
.B(n_271),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2008),
.Y(n_2080)
);

AOI221x1_ASAP7_75t_SL g2081 ( 
.A1(n_2048),
.A2(n_274),
.B1(n_272),
.B2(n_273),
.C(n_275),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2016),
.Y(n_2082)
);

AOI21xp33_ASAP7_75t_L g2083 ( 
.A1(n_2015),
.A2(n_276),
.B(n_277),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_2052),
.Y(n_2084)
);

NAND4xp25_ASAP7_75t_L g2085 ( 
.A(n_2012),
.B(n_279),
.C(n_280),
.D(n_278),
.Y(n_2085)
);

AND2x2_ASAP7_75t_L g2086 ( 
.A(n_2003),
.B(n_2054),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_2067),
.B(n_278),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_2055),
.B(n_282),
.Y(n_2088)
);

AOI32xp33_ASAP7_75t_L g2089 ( 
.A1(n_2058),
.A2(n_285),
.A3(n_283),
.B1(n_284),
.B2(n_286),
.Y(n_2089)
);

A2O1A1Ixp33_ASAP7_75t_L g2090 ( 
.A1(n_2033),
.A2(n_285),
.B(n_283),
.C(n_284),
.Y(n_2090)
);

A2O1A1Ixp33_ASAP7_75t_L g2091 ( 
.A1(n_2075),
.A2(n_289),
.B(n_287),
.C(n_288),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_2064),
.B(n_289),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_2004),
.B(n_290),
.Y(n_2093)
);

AOI21xp33_ASAP7_75t_L g2094 ( 
.A1(n_2076),
.A2(n_291),
.B(n_294),
.Y(n_2094)
);

AOI22xp33_ASAP7_75t_SL g2095 ( 
.A1(n_2050),
.A2(n_296),
.B1(n_294),
.B2(n_295),
.Y(n_2095)
);

AOI21xp33_ASAP7_75t_SL g2096 ( 
.A1(n_2013),
.A2(n_296),
.B(n_297),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_2049),
.B(n_298),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_SL g2098 ( 
.A(n_2009),
.B(n_2032),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_2069),
.B(n_2072),
.Y(n_2099)
);

NOR5xp2_ASAP7_75t_SL g2100 ( 
.A(n_2070),
.B(n_303),
.C(n_301),
.D(n_302),
.E(n_304),
.Y(n_2100)
);

AND2x4_ASAP7_75t_L g2101 ( 
.A(n_2007),
.B(n_301),
.Y(n_2101)
);

INVxp67_ASAP7_75t_L g2102 ( 
.A(n_2036),
.Y(n_2102)
);

AO21x1_ASAP7_75t_L g2103 ( 
.A1(n_2047),
.A2(n_303),
.B(n_304),
.Y(n_2103)
);

AND2x4_ASAP7_75t_L g2104 ( 
.A(n_2026),
.B(n_2066),
.Y(n_2104)
);

OAI21xp33_ASAP7_75t_L g2105 ( 
.A1(n_2017),
.A2(n_305),
.B(n_306),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_2005),
.Y(n_2106)
);

AOI21xp33_ASAP7_75t_L g2107 ( 
.A1(n_2021),
.A2(n_307),
.B(n_308),
.Y(n_2107)
);

NOR2xp67_ASAP7_75t_L g2108 ( 
.A(n_2062),
.B(n_309),
.Y(n_2108)
);

INVx1_ASAP7_75t_SL g2109 ( 
.A(n_2024),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2045),
.B(n_313),
.Y(n_2110)
);

OAI21xp33_ASAP7_75t_SL g2111 ( 
.A1(n_2030),
.A2(n_314),
.B(n_315),
.Y(n_2111)
);

INVx1_ASAP7_75t_SL g2112 ( 
.A(n_2020),
.Y(n_2112)
);

OA21x2_ASAP7_75t_L g2113 ( 
.A1(n_2010),
.A2(n_318),
.B(n_319),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2057),
.Y(n_2114)
);

OAI21xp5_ASAP7_75t_SL g2115 ( 
.A1(n_2041),
.A2(n_325),
.B(n_326),
.Y(n_2115)
);

OAI22xp5_ASAP7_75t_L g2116 ( 
.A1(n_2029),
.A2(n_329),
.B1(n_327),
.B2(n_328),
.Y(n_2116)
);

OAI211xp5_ASAP7_75t_L g2117 ( 
.A1(n_2061),
.A2(n_331),
.B(n_329),
.C(n_330),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2059),
.Y(n_2118)
);

OAI21xp33_ASAP7_75t_L g2119 ( 
.A1(n_2068),
.A2(n_334),
.B(n_335),
.Y(n_2119)
);

NAND4xp25_ASAP7_75t_L g2120 ( 
.A(n_2014),
.B(n_336),
.C(n_334),
.D(n_335),
.Y(n_2120)
);

INVx1_ASAP7_75t_SL g2121 ( 
.A(n_2027),
.Y(n_2121)
);

OR2x2_ASAP7_75t_L g2122 ( 
.A(n_2019),
.B(n_337),
.Y(n_2122)
);

INVx3_ASAP7_75t_L g2123 ( 
.A(n_2034),
.Y(n_2123)
);

HB1xp67_ASAP7_75t_L g2124 ( 
.A(n_2025),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_2056),
.B(n_339),
.Y(n_2125)
);

AO22x1_ASAP7_75t_L g2126 ( 
.A1(n_2063),
.A2(n_342),
.B1(n_340),
.B2(n_341),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_2065),
.B(n_340),
.Y(n_2127)
);

NOR2xp33_ASAP7_75t_L g2128 ( 
.A(n_2042),
.B(n_342),
.Y(n_2128)
);

NAND3xp33_ASAP7_75t_L g2129 ( 
.A(n_2046),
.B(n_343),
.C(n_345),
.Y(n_2129)
);

AOI221xp5_ASAP7_75t_L g2130 ( 
.A1(n_2023),
.A2(n_347),
.B1(n_345),
.B2(n_346),
.C(n_348),
.Y(n_2130)
);

NAND3xp33_ASAP7_75t_L g2131 ( 
.A(n_2051),
.B(n_350),
.C(n_351),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_2086),
.B(n_2073),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2078),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2080),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_2099),
.B(n_2053),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2082),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2084),
.Y(n_2137)
);

NOR2xp33_ASAP7_75t_L g2138 ( 
.A(n_2123),
.B(n_2071),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_2109),
.B(n_2040),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_2077),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2112),
.B(n_2121),
.Y(n_2141)
);

NOR2x1_ASAP7_75t_L g2142 ( 
.A(n_2108),
.B(n_2028),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_2103),
.B(n_2043),
.Y(n_2143)
);

OAI22xp5_ASAP7_75t_L g2144 ( 
.A1(n_2129),
.A2(n_2031),
.B1(n_2037),
.B2(n_2035),
.Y(n_2144)
);

NOR2xp33_ASAP7_75t_L g2145 ( 
.A(n_2098),
.B(n_2022),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_2124),
.B(n_2011),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2114),
.B(n_2118),
.Y(n_2147)
);

CKINVDCx5p33_ASAP7_75t_R g2148 ( 
.A(n_2100),
.Y(n_2148)
);

AOI22xp33_ASAP7_75t_L g2149 ( 
.A1(n_2094),
.A2(n_2044),
.B1(n_2038),
.B2(n_2018),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2101),
.Y(n_2150)
);

HB1xp67_ASAP7_75t_L g2151 ( 
.A(n_2102),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2104),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_2106),
.B(n_2074),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2088),
.B(n_352),
.Y(n_2154)
);

HB1xp67_ASAP7_75t_L g2155 ( 
.A(n_2113),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_2111),
.B(n_352),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_SL g2157 ( 
.A(n_2089),
.B(n_353),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_2092),
.B(n_354),
.Y(n_2158)
);

NOR2xp33_ASAP7_75t_L g2159 ( 
.A(n_2110),
.B(n_355),
.Y(n_2159)
);

NOR2xp33_ASAP7_75t_L g2160 ( 
.A(n_2093),
.B(n_357),
.Y(n_2160)
);

OAI22xp5_ASAP7_75t_L g2161 ( 
.A1(n_2115),
.A2(n_359),
.B1(n_357),
.B2(n_358),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_2095),
.B(n_360),
.Y(n_2162)
);

NAND2xp33_ASAP7_75t_L g2163 ( 
.A(n_2090),
.B(n_362),
.Y(n_2163)
);

OAI221xp5_ASAP7_75t_L g2164 ( 
.A1(n_2081),
.A2(n_364),
.B1(n_362),
.B2(n_363),
.C(n_365),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2126),
.B(n_363),
.Y(n_2165)
);

HB1xp67_ASAP7_75t_L g2166 ( 
.A(n_2142),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2151),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_2132),
.B(n_2135),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2147),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2155),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2133),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2134),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2136),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2137),
.Y(n_2174)
);

INVx2_ASAP7_75t_SL g2175 ( 
.A(n_2150),
.Y(n_2175)
);

NOR2xp33_ASAP7_75t_L g2176 ( 
.A(n_2148),
.B(n_2097),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_2140),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_2153),
.B(n_2128),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2152),
.Y(n_2179)
);

INVx2_ASAP7_75t_SL g2180 ( 
.A(n_2154),
.Y(n_2180)
);

HB1xp67_ASAP7_75t_L g2181 ( 
.A(n_2139),
.Y(n_2181)
);

INVxp67_ASAP7_75t_L g2182 ( 
.A(n_2143),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2146),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2158),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2156),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2165),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2144),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_2138),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2160),
.Y(n_2189)
);

INVx2_ASAP7_75t_SL g2190 ( 
.A(n_2157),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_2145),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_2162),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2159),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2161),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_2164),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2163),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2149),
.Y(n_2197)
);

INVx8_ASAP7_75t_L g2198 ( 
.A(n_2141),
.Y(n_2198)
);

OAI321xp33_ASAP7_75t_L g2199 ( 
.A1(n_2182),
.A2(n_2085),
.A3(n_2120),
.B1(n_2105),
.B2(n_2116),
.C(n_2119),
.Y(n_2199)
);

AND4x1_ASAP7_75t_L g2200 ( 
.A(n_2176),
.B(n_2131),
.C(n_2091),
.D(n_2130),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_2168),
.B(n_2087),
.Y(n_2201)
);

OR3x1_ASAP7_75t_L g2202 ( 
.A(n_2167),
.B(n_2083),
.C(n_2107),
.Y(n_2202)
);

NAND3xp33_ASAP7_75t_SL g2203 ( 
.A(n_2166),
.B(n_2096),
.C(n_2117),
.Y(n_2203)
);

AOI211xp5_ASAP7_75t_L g2204 ( 
.A1(n_2196),
.A2(n_2187),
.B(n_2197),
.C(n_2190),
.Y(n_2204)
);

OAI211xp5_ASAP7_75t_SL g2205 ( 
.A1(n_2186),
.A2(n_2125),
.B(n_2127),
.C(n_2079),
.Y(n_2205)
);

XNOR2x1_ASAP7_75t_L g2206 ( 
.A(n_2195),
.B(n_2122),
.Y(n_2206)
);

AOI221x1_ASAP7_75t_L g2207 ( 
.A1(n_2170),
.A2(n_367),
.B1(n_365),
.B2(n_366),
.C(n_368),
.Y(n_2207)
);

NOR3xp33_ASAP7_75t_L g2208 ( 
.A(n_2185),
.B(n_369),
.C(n_370),
.Y(n_2208)
);

NOR4xp25_ASAP7_75t_L g2209 ( 
.A(n_2192),
.B(n_374),
.C(n_371),
.D(n_373),
.Y(n_2209)
);

NOR3xp33_ASAP7_75t_L g2210 ( 
.A(n_2191),
.B(n_371),
.C(n_373),
.Y(n_2210)
);

NOR4xp25_ASAP7_75t_L g2211 ( 
.A(n_2175),
.B(n_2179),
.C(n_2194),
.D(n_2177),
.Y(n_2211)
);

AOI21xp5_ASAP7_75t_L g2212 ( 
.A1(n_2198),
.A2(n_375),
.B(n_376),
.Y(n_2212)
);

AOI221xp5_ASAP7_75t_L g2213 ( 
.A1(n_2181),
.A2(n_381),
.B1(n_379),
.B2(n_380),
.C(n_382),
.Y(n_2213)
);

NOR3xp33_ASAP7_75t_L g2214 ( 
.A(n_2188),
.B(n_380),
.C(n_381),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_2178),
.B(n_384),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_2180),
.B(n_385),
.Y(n_2216)
);

HB1xp67_ASAP7_75t_L g2217 ( 
.A(n_2169),
.Y(n_2217)
);

AOI311xp33_ASAP7_75t_L g2218 ( 
.A1(n_2183),
.A2(n_390),
.A3(n_388),
.B(n_389),
.C(n_391),
.Y(n_2218)
);

BUFx2_ASAP7_75t_L g2219 ( 
.A(n_2184),
.Y(n_2219)
);

AOI211xp5_ASAP7_75t_L g2220 ( 
.A1(n_2193),
.A2(n_397),
.B(n_394),
.C(n_395),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_SL g2221 ( 
.A(n_2189),
.B(n_394),
.Y(n_2221)
);

OAI22xp5_ASAP7_75t_L g2222 ( 
.A1(n_2202),
.A2(n_2172),
.B1(n_2173),
.B2(n_2171),
.Y(n_2222)
);

NAND2xp33_ASAP7_75t_L g2223 ( 
.A(n_2218),
.B(n_2174),
.Y(n_2223)
);

OAI211xp5_ASAP7_75t_SL g2224 ( 
.A1(n_2204),
.A2(n_402),
.B(n_400),
.C(n_401),
.Y(n_2224)
);

NAND3xp33_ASAP7_75t_L g2225 ( 
.A(n_2200),
.B(n_403),
.C(n_404),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2219),
.Y(n_2226)
);

AOI21xp33_ASAP7_75t_SL g2227 ( 
.A1(n_2206),
.A2(n_2209),
.B(n_2210),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_2215),
.B(n_405),
.Y(n_2228)
);

AOI21xp33_ASAP7_75t_SL g2229 ( 
.A1(n_2214),
.A2(n_405),
.B(n_406),
.Y(n_2229)
);

AOI221xp5_ASAP7_75t_L g2230 ( 
.A1(n_2199),
.A2(n_409),
.B1(n_407),
.B2(n_408),
.C(n_411),
.Y(n_2230)
);

AOI22xp33_ASAP7_75t_L g2231 ( 
.A1(n_2201),
.A2(n_2205),
.B1(n_2217),
.B2(n_2208),
.Y(n_2231)
);

OAI211xp5_ASAP7_75t_SL g2232 ( 
.A1(n_2213),
.A2(n_414),
.B(n_412),
.C(n_413),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2216),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2212),
.B(n_418),
.Y(n_2234)
);

OAI21xp33_ASAP7_75t_SL g2235 ( 
.A1(n_2221),
.A2(n_420),
.B(n_421),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_2207),
.B(n_422),
.Y(n_2236)
);

O2A1O1Ixp33_ASAP7_75t_L g2237 ( 
.A1(n_2220),
.A2(n_427),
.B(n_424),
.C(n_425),
.Y(n_2237)
);

AOI211x1_ASAP7_75t_SL g2238 ( 
.A1(n_2203),
.A2(n_435),
.B(n_431),
.C(n_434),
.Y(n_2238)
);

AOI221xp5_ASAP7_75t_L g2239 ( 
.A1(n_2211),
.A2(n_438),
.B1(n_436),
.B2(n_437),
.C(n_439),
.Y(n_2239)
);

NOR4xp75_ASAP7_75t_L g2240 ( 
.A(n_2222),
.B(n_443),
.C(n_440),
.D(n_442),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2226),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2228),
.Y(n_2242)
);

NAND4xp75_ASAP7_75t_L g2243 ( 
.A(n_2239),
.B(n_447),
.C(n_444),
.D(n_445),
.Y(n_2243)
);

NOR2x1_ASAP7_75t_L g2244 ( 
.A(n_2225),
.B(n_447),
.Y(n_2244)
);

NOR2x1_ASAP7_75t_L g2245 ( 
.A(n_2236),
.B(n_448),
.Y(n_2245)
);

NAND4xp75_ASAP7_75t_L g2246 ( 
.A(n_2230),
.B(n_451),
.C(n_449),
.D(n_450),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_2231),
.B(n_451),
.Y(n_2247)
);

OR2x6_ASAP7_75t_L g2248 ( 
.A(n_2234),
.B(n_452),
.Y(n_2248)
);

NOR2xp67_ASAP7_75t_L g2249 ( 
.A(n_2235),
.B(n_2227),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2233),
.Y(n_2250)
);

AOI22xp5_ASAP7_75t_L g2251 ( 
.A1(n_2223),
.A2(n_454),
.B1(n_452),
.B2(n_453),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_SL g2252 ( 
.A(n_2249),
.B(n_2229),
.Y(n_2252)
);

OAI21xp5_ASAP7_75t_SL g2253 ( 
.A1(n_2251),
.A2(n_2224),
.B(n_2238),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_2245),
.B(n_2247),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2254),
.Y(n_2255)
);

OAI221xp5_ASAP7_75t_L g2256 ( 
.A1(n_2253),
.A2(n_2241),
.B1(n_2244),
.B2(n_2250),
.C(n_2237),
.Y(n_2256)
);

NOR4xp25_ASAP7_75t_L g2257 ( 
.A(n_2252),
.B(n_2242),
.C(n_2232),
.D(n_2240),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2255),
.Y(n_2258)
);

OAI22xp5_ASAP7_75t_SL g2259 ( 
.A1(n_2258),
.A2(n_2248),
.B1(n_2256),
.B2(n_2257),
.Y(n_2259)
);

AOI31xp33_ASAP7_75t_L g2260 ( 
.A1(n_2259),
.A2(n_2248),
.A3(n_2243),
.B(n_2246),
.Y(n_2260)
);

AOI22xp5_ASAP7_75t_L g2261 ( 
.A1(n_2260),
.A2(n_459),
.B1(n_457),
.B2(n_458),
.Y(n_2261)
);

OAI22x1_ASAP7_75t_L g2262 ( 
.A1(n_2261),
.A2(n_463),
.B1(n_461),
.B2(n_462),
.Y(n_2262)
);

INVx1_ASAP7_75t_SL g2263 ( 
.A(n_2262),
.Y(n_2263)
);

OAI221xp5_ASAP7_75t_R g2264 ( 
.A1(n_2263),
.A2(n_466),
.B1(n_464),
.B2(n_465),
.C(n_467),
.Y(n_2264)
);

AOI211xp5_ASAP7_75t_L g2265 ( 
.A1(n_2264),
.A2(n_468),
.B(n_465),
.C(n_467),
.Y(n_2265)
);


endmodule