module fake_jpeg_22201_n_204 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_38),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g36 ( 
.A(n_32),
.B(n_1),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_37),
.C(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_2),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_2),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_18),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_45),
.B(n_52),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_41),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_46),
.Y(n_69)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_29),
.B1(n_34),
.B2(n_27),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_49),
.A2(n_51),
.B1(n_31),
.B2(n_47),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_29),
.B1(n_27),
.B2(n_24),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVxp67_ASAP7_75t_SL g71 ( 
.A(n_56),
.Y(n_71)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_30),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_62),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_22),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_64),
.B(n_18),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_66),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_63),
.A2(n_36),
.B(n_24),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_68),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_36),
.C(n_22),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_83),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_80),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_36),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_87),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_47),
.A2(n_38),
.B1(n_16),
.B2(n_19),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_75),
.A2(n_93),
.B1(n_26),
.B2(n_23),
.Y(n_111)
);

NOR2x1_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_16),
.Y(n_77)
);

NOR2x1_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_33),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_19),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_78),
.B(n_20),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_13),
.Y(n_102)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_55),
.A2(n_31),
.B1(n_21),
.B2(n_28),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_85),
.Y(n_103)
);

FAx1_ASAP7_75t_SL g86 ( 
.A(n_65),
.B(n_59),
.CI(n_45),
.CON(n_86),
.SN(n_86)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_86),
.B(n_58),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_25),
.Y(n_87)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_50),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

AO21x2_ASAP7_75t_L g93 ( 
.A1(n_52),
.A2(n_25),
.B(n_26),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_50),
.B1(n_53),
.B2(n_58),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_94),
.A2(n_93),
.B1(n_72),
.B2(n_84),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_95),
.A2(n_114),
.B(n_70),
.Y(n_121)
);

NOR3xp33_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_28),
.C(n_21),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_112),
.Y(n_124)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_102),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_100),
.B(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_69),
.B(n_20),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_113),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_108),
.A2(n_111),
.B1(n_93),
.B2(n_81),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_74),
.B(n_58),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_68),
.Y(n_123)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_33),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_3),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_33),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_86),
.Y(n_129)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_116),
.B(n_3),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_118),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_106),
.A2(n_116),
.B1(n_103),
.B2(n_95),
.Y(n_120)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

AO21x1_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_126),
.B(n_105),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_123),
.A2(n_134),
.B(n_137),
.Y(n_150)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_132),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_110),
.C(n_105),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_133),
.C(n_137),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_129),
.B(n_131),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_108),
.A2(n_72),
.B1(n_81),
.B2(n_93),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_104),
.B(n_112),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_101),
.B(n_76),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_84),
.C(n_67),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_82),
.B1(n_67),
.B2(n_53),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_78),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_136),
.Y(n_139)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_117),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_138),
.B(n_144),
.Y(n_166)
);

NAND3xp33_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_108),
.C(n_99),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_143),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_114),
.C(n_105),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_123),
.B(n_121),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_117),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_146),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_131),
.B(n_100),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_151),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_134),
.B1(n_111),
.B2(n_118),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_127),
.C(n_133),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_119),
.B(n_102),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_128),
.Y(n_153)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_153),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_128),
.Y(n_155)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_164),
.C(n_168),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_162),
.A2(n_165),
.B1(n_167),
.B2(n_4),
.Y(n_180)
);

BUFx12_ASAP7_75t_L g163 ( 
.A(n_154),
.Y(n_163)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_163),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_122),
.C(n_136),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_142),
.A2(n_124),
.B1(n_122),
.B2(n_94),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_132),
.C(n_91),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_91),
.C(n_90),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_26),
.C(n_23),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_156),
.A2(n_152),
.B(n_150),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_172),
.A2(n_179),
.B(n_161),
.Y(n_184)
);

AOI322xp5_ASAP7_75t_L g173 ( 
.A1(n_166),
.A2(n_152),
.A3(n_146),
.B1(n_140),
.B2(n_139),
.C1(n_153),
.C2(n_145),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_175),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_168),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_176),
.Y(n_183)
);

AOI322xp5_ASAP7_75t_L g175 ( 
.A1(n_158),
.A2(n_140),
.A3(n_138),
.B1(n_150),
.B2(n_147),
.C1(n_151),
.C2(n_119),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_90),
.C(n_92),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_177),
.A2(n_180),
.B(n_5),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_23),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_5),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_157),
.A2(n_3),
.B(n_4),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_179),
.B(n_159),
.Y(n_181)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_171),
.B(n_163),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_187),
.C(n_188),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_184),
.A2(n_185),
.B1(n_177),
.B2(n_170),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_170),
.A2(n_163),
.B(n_12),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_190),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_174),
.C(n_178),
.Y(n_190)
);

BUFx24_ASAP7_75t_SL g192 ( 
.A(n_181),
.Y(n_192)
);

AO21x1_ASAP7_75t_L g195 ( 
.A1(n_192),
.A2(n_193),
.B(n_182),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_11),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_195),
.B(n_15),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_191),
.A2(n_194),
.B1(n_190),
.B2(n_14),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_197),
.Y(n_201)
);

AOI322xp5_ASAP7_75t_L g198 ( 
.A1(n_191),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_13),
.C1(n_15),
.C2(n_192),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_198),
.B(n_7),
.C(n_8),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_200),
.Y(n_203)
);

AO21x1_ASAP7_75t_L g202 ( 
.A1(n_201),
.A2(n_196),
.B(n_198),
.Y(n_202)
);

FAx1_ASAP7_75t_SL g204 ( 
.A(n_202),
.B(n_9),
.CI(n_203),
.CON(n_204),
.SN(n_204)
);


endmodule