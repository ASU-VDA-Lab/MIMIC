module real_jpeg_22289_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_342, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_342;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_0),
.A2(n_27),
.B1(n_29),
.B2(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_0),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_0),
.A2(n_23),
.B1(n_25),
.B2(n_115),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_0),
.A2(n_47),
.B1(n_48),
.B2(n_115),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_0),
.A2(n_41),
.B1(n_42),
.B2(n_115),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_1),
.A2(n_23),
.B1(n_25),
.B2(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_1),
.A2(n_47),
.B1(n_48),
.B2(n_58),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_1),
.A2(n_41),
.B1(n_42),
.B2(n_58),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_1),
.A2(n_27),
.B1(n_29),
.B2(n_58),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_2),
.A2(n_27),
.B1(n_29),
.B2(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_2),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_2),
.A2(n_47),
.B1(n_48),
.B2(n_117),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_2),
.A2(n_41),
.B1(n_42),
.B2(n_117),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_2),
.A2(n_23),
.B1(n_25),
.B2(n_117),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_3),
.A2(n_24),
.B1(n_41),
.B2(n_42),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_3),
.A2(n_24),
.B1(n_27),
.B2(n_29),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_3),
.A2(n_24),
.B1(n_47),
.B2(n_48),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_4),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_4),
.B(n_26),
.Y(n_149)
);

AOI21xp33_ASAP7_75t_L g170 ( 
.A1(n_4),
.A2(n_14),
.B(n_48),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_4),
.A2(n_41),
.B1(n_42),
.B2(n_120),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_4),
.A2(n_94),
.B1(n_99),
.B2(n_179),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_4),
.B(n_76),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_4),
.B(n_29),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g211 ( 
.A1(n_4),
.A2(n_29),
.B(n_207),
.Y(n_211)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_6),
.A2(n_23),
.B1(n_25),
.B2(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_6),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_6),
.A2(n_27),
.B1(n_29),
.B2(n_122),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_6),
.A2(n_41),
.B1(n_42),
.B2(n_122),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_6),
.A2(n_47),
.B1(n_48),
.B2(n_122),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_7),
.B(n_47),
.Y(n_95)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_7),
.Y(n_99)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_7),
.Y(n_180)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_9),
.A2(n_23),
.B1(n_25),
.B2(n_32),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_9),
.A2(n_27),
.B1(n_29),
.B2(n_32),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_9),
.A2(n_32),
.B1(n_47),
.B2(n_48),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_9),
.A2(n_32),
.B1(n_41),
.B2(n_42),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_11),
.A2(n_23),
.B1(n_25),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_11),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_11),
.A2(n_41),
.B1(n_42),
.B2(n_56),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_11),
.A2(n_47),
.B1(n_48),
.B2(n_56),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_11),
.A2(n_27),
.B1(n_29),
.B2(n_56),
.Y(n_272)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_12),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_14),
.A2(n_41),
.B(n_45),
.C(n_46),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_41),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_14),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_46)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_15),
.Y(n_44)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.C(n_339),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_82),
.B(n_337),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_35),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_20),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_30),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_21),
.A2(n_54),
.B(n_255),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_26),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_22),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_22),
.A2(n_26),
.B(n_33),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_23),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_23),
.A2(n_26),
.B(n_28),
.C(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_28),
.Y(n_34)
);

HAxp5_ASAP7_75t_SL g119 ( 
.A(n_23),
.B(n_120),
.CON(n_119),
.SN(n_119)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_26),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_26),
.B(n_31),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_26),
.A2(n_33),
.B1(n_119),
.B2(n_121),
.Y(n_118)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_27),
.A2(n_34),
.B1(n_119),
.B2(n_126),
.Y(n_125)
);

AOI32xp33_ASAP7_75t_L g206 ( 
.A1(n_27),
.A2(n_41),
.A3(n_66),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_28),
.B(n_29),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_29),
.A2(n_64),
.B(n_65),
.C(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_29),
.B(n_65),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_30),
.A2(n_55),
.B(n_59),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_33),
.A2(n_79),
.B(n_80),
.Y(n_78)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_36),
.B(n_338),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_74),
.C(n_78),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_37),
.A2(n_38),
.B1(n_333),
.B2(n_335),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_52),
.C(n_60),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_39),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_39),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_39),
.A2(n_60),
.B1(n_61),
.B2(n_313),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_46),
.B(n_50),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_40),
.A2(n_50),
.B(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_40),
.A2(n_46),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_40),
.A2(n_46),
.B1(n_174),
.B2(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_40),
.A2(n_46),
.B1(n_195),
.B2(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_40),
.A2(n_214),
.B(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_40),
.A2(n_46),
.B1(n_102),
.B2(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_40),
.A2(n_110),
.B(n_247),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_42),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_42),
.A2(n_49),
.B(n_120),
.C(n_170),
.Y(n_169)
);

NAND2xp33_ASAP7_75t_SL g208 ( 
.A(n_42),
.B(n_65),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_46),
.A2(n_102),
.B(n_103),
.Y(n_101)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_46),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_46),
.B(n_120),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_47),
.B(n_184),
.Y(n_183)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_51),
.B(n_111),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_52),
.A2(n_53),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_59),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_54),
.A2(n_59),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_54),
.A2(n_59),
.B1(n_133),
.B2(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_54),
.A2(n_81),
.B(n_301),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_57),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_68),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_63),
.A2(n_69),
.B(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_64),
.A2(n_70),
.B1(n_114),
.B2(n_116),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_64),
.A2(n_70),
.B1(n_152),
.B2(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_64),
.B(n_73),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_64),
.A2(n_68),
.B(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_64),
.A2(n_70),
.B1(n_272),
.B2(n_293),
.Y(n_292)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_67),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_69),
.A2(n_76),
.B(n_77),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_69),
.A2(n_76),
.B1(n_151),
.B2(n_153),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_69),
.A2(n_77),
.B(n_258),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_69),
.A2(n_258),
.B(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_74),
.A2(n_75),
.B1(n_78),
.B2(n_334),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_78),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_330),
.B(n_336),
.Y(n_82)
);

OAI321xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_306),
.A3(n_325),
.B1(n_328),
.B2(n_329),
.C(n_342),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_285),
.B(n_305),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_263),
.B(n_284),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_154),
.B(n_238),
.C(n_262),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_138),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_88),
.B(n_138),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_123),
.B2(n_137),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_107),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_91),
.B(n_107),
.C(n_137),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_101),
.B2(n_106),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_92),
.B(n_106),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_96),
.B(n_97),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_94),
.A2(n_96),
.B1(n_99),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_94),
.A2(n_163),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_94),
.A2(n_166),
.B(n_197),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_94),
.A2(n_180),
.B(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_95),
.B(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_95),
.A2(n_162),
.B1(n_164),
.B2(n_165),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_95),
.A2(n_98),
.B(n_199),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_99),
.A2(n_128),
.B(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_99),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_99),
.B(n_120),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_101),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_103),
.B(n_229),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_104),
.B(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.C(n_118),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_108),
.A2(n_109),
.B1(n_112),
.B2(n_113),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_114),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_116),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_118),
.B(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_121),
.Y(n_132)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_129),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_124),
.B(n_130),
.C(n_135),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_127),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_134),
.B2(n_135),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.C(n_143),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_139),
.B(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_149),
.C(n_150),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_145),
.A2(n_146),
.B1(n_149),
.B2(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_147),
.B(n_197),
.Y(n_245)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_149),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_150),
.B(n_224),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_237),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_232),
.B(n_236),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_219),
.B(n_231),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_201),
.B(n_218),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_187),
.B(n_200),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_175),
.B(n_186),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_167),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_167),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_171),
.B2(n_172),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_169),
.B(n_171),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_181),
.B(n_185),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_178),
.Y(n_185)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_180),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_188),
.B(n_189),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_196),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_194),
.C(n_196),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_199),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_203),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_209),
.B1(n_216),
.B2(n_217),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_204),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_206),
.Y(n_230)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_209),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_212),
.B1(n_213),
.B2(n_215),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_210),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_215),
.C(n_216),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_220),
.B(n_221),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_226),
.B2(n_227),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_228),
.C(n_230),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_233),
.B(n_234),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_239),
.B(n_240),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_260),
.B2(n_261),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_248),
.B2(n_249),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_249),
.C(n_261),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_246),
.Y(n_269)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_252),
.B2(n_259),
.Y(n_249)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_250),
.Y(n_259)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_256),
.B2(n_257),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_257),
.C(n_259),
.Y(n_283)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_260),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_264),
.B(n_265),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_283),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_276),
.B2(n_277),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_277),
.C(n_283),
.Y(n_286)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_269),
.B(n_273),
.C(n_275),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_271),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_281),
.B2(n_282),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_278),
.A2(n_279),
.B1(n_300),
.B2(n_302),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_278),
.A2(n_296),
.B(n_300),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_281),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_281),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_286),
.B(n_287),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_303),
.B2(n_304),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_295),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_290),
.B(n_295),
.C(n_304),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B(n_294),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_292),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_293),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_308),
.C(n_317),
.Y(n_307)
);

FAx1_ASAP7_75t_SL g327 ( 
.A(n_294),
.B(n_308),
.CI(n_317),
.CON(n_327),
.SN(n_327)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_300),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_303),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_318),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_307),
.B(n_318),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_309),
.A2(n_310),
.B1(n_320),
.B2(n_323),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_310),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_313),
.C(n_315),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_310),
.B(n_323),
.C(n_324),
.Y(n_331)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_324),
.Y(n_318)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_320),
.Y(n_323)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_326),
.B(n_327),
.Y(n_328)
);

BUFx24_ASAP7_75t_SL g341 ( 
.A(n_327),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_332),
.Y(n_336)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_333),
.Y(n_335)
);


endmodule