module fake_ariane_1078_n_7467 (n_913, n_1681, n_1486, n_1507, n_589, n_1174, n_1469, n_691, n_1353, n_1355, n_423, n_1383, n_603, n_373, n_1250, n_1169, n_789, n_850, n_610, n_245, n_96, n_319, n_49, n_1436, n_690, n_416, n_1109, n_1430, n_525, n_187, n_1463, n_1238, n_1515, n_817, n_924, n_781, n_1566, n_189, n_717, n_72, n_952, n_864, n_1096, n_1379, n_57, n_1706, n_117, n_524, n_1214, n_634, n_1246, n_1138, n_214, n_764, n_1503, n_462, n_1196, n_1181, n_32, n_410, n_1187, n_1131, n_1225, n_737, n_137, n_1298, n_1366, n_232, n_52, n_568, n_1088, n_77, n_1424, n_766, n_1457, n_377, n_1682, n_520, n_870, n_1453, n_279, n_945, n_958, n_813, n_419, n_146, n_270, n_338, n_995, n_285, n_1184, n_202, n_1535, n_500, n_665, n_754, n_903, n_871, n_1073, n_239, n_402, n_1277, n_54, n_829, n_1062, n_339, n_738, n_1690, n_672, n_740, n_1283, n_167, n_1018, n_69, n_259, n_953, n_1364, n_143, n_1224, n_1425, n_625, n_557, n_1107, n_1688, n_989, n_242, n_645, n_331, n_559, n_267, n_495, n_350, n_381, n_795, n_721, n_1084, n_1276, n_200, n_1428, n_1284, n_1241, n_821, n_561, n_770, n_1514, n_1528, n_507, n_486, n_901, n_569, n_1145, n_971, n_787, n_1650, n_31, n_1519, n_1195, n_1522, n_518, n_1207, n_222, n_786, n_1404, n_868, n_1542, n_1314, n_1512, n_1539, n_884, n_1415, n_1034, n_1652, n_1676, n_1085, n_277, n_1636, n_432, n_293, n_823, n_620, n_93, n_1074, n_859, n_108, n_587, n_693, n_863, n_303, n_1254, n_929, n_206, n_352, n_899, n_1703, n_611, n_1295, n_238, n_365, n_1013, n_1495, n_1637, n_136, n_334, n_192, n_661, n_300, n_533, n_104, n_438, n_1560, n_1654, n_1548, n_16, n_440, n_273, n_1396, n_1230, n_612, n_333, n_376, n_512, n_1597, n_1544, n_579, n_844, n_1012, n_1267, n_1354, n_149, n_1213, n_237, n_780, n_1021, n_1443, n_491, n_1465, n_1595, n_1142, n_1140, n_705, n_570, n_260, n_942, n_1437, n_7, n_1378, n_461, n_1121, n_1416, n_209, n_490, n_1461, n_17, n_1391, n_225, n_1599, n_1006, n_575, n_546, n_503, n_1112, n_700, n_1159, n_772, n_1216, n_1245, n_1669, n_1675, n_676, n_42, n_1594, n_680, n_287, n_302, n_380, n_1585, n_1432, n_94, n_4, n_249, n_1108, n_355, n_212, n_65, n_123, n_444, n_851, n_1590, n_1351, n_1274, n_257, n_652, n_475, n_135, n_947, n_930, n_1260, n_1179, n_468, n_102, n_182, n_696, n_1442, n_482, n_798, n_577, n_407, n_1691, n_27, n_916, n_1386, n_912, n_460, n_1555, n_366, n_762, n_1253, n_1468, n_1661, n_555, n_804, n_1656, n_1382, n_966, n_992, n_955, n_1182, n_794, n_78, n_1692, n_1562, n_514, n_418, n_1376, n_513, n_288, n_179, n_1292, n_1178, n_1435, n_1026, n_1506, n_1610, n_306, n_92, n_203, n_436, n_150, n_324, n_669, n_931, n_1491, n_619, n_337, n_437, n_111, n_21, n_274, n_967, n_1083, n_1418, n_746, n_1357, n_292, n_1079, n_1389, n_615, n_1139, n_76, n_517, n_1312, n_0, n_824, n_428, n_159, n_892, n_959, n_30, n_1399, n_1101, n_1567, n_1343, n_563, n_144, n_990, n_1623, n_867, n_1226, n_944, n_749, n_815, n_542, n_1340, n_470, n_1240, n_1087, n_632, n_477, n_650, n_425, n_1433, n_1155, n_1071, n_712, n_976, n_909, n_1392, n_767, n_1680, n_964, n_1627, n_382, n_489, n_80, n_251, n_974, n_506, n_799, n_1147, n_397, n_471, n_351, n_965, n_155, n_934, n_1447, n_1220, n_356, n_698, n_1674, n_124, n_307, n_1209, n_1020, n_1563, n_646, n_1633, n_34, n_404, n_172, n_1058, n_347, n_1042, n_183, n_1234, n_479, n_1578, n_1455, n_299, n_836, n_1279, n_564, n_133, n_66, n_205, n_1029, n_1247, n_760, n_522, n_1568, n_20, n_1483, n_1363, n_367, n_1111, n_970, n_1689, n_713, n_1255, n_1646, n_598, n_345, n_1237, n_927, n_261, n_1095, n_370, n_706, n_286, n_1401, n_1419, n_1531, n_776, n_424, n_1651, n_85, n_130, n_1387, n_466, n_1263, n_346, n_348, n_552, n_670, n_379, n_138, n_162, n_264, n_441, n_1032, n_1217, n_1496, n_637, n_1592, n_73, n_327, n_1259, n_1177, n_1231, n_980, n_1618, n_905, n_207, n_720, n_926, n_41, n_194, n_1163, n_186, n_1384, n_145, n_59, n_1501, n_1173, n_1068, n_1198, n_1570, n_487, n_1518, n_1456, n_90, n_1648, n_1413, n_855, n_158, n_808, n_1365, n_553, n_1439, n_814, n_578, n_1665, n_1287, n_405, n_1611, n_120, n_320, n_1414, n_1134, n_1484, n_647, n_1423, n_481, n_600, n_1053, n_1609, n_529, n_502, n_218, n_1467, n_247, n_1304, n_1608, n_1105, n_547, n_439, n_604, n_677, n_478, n_703, n_1349, n_1061, n_326, n_681, n_227, n_874, n_1278, n_707, n_11, n_129, n_126, n_983, n_590, n_699, n_727, n_301, n_545, n_1015, n_1377, n_1162, n_536, n_1614, n_325, n_1602, n_688, n_636, n_427, n_1098, n_1490, n_442, n_777, n_1553, n_1080, n_920, n_1086, n_1092, n_986, n_1104, n_729, n_887, n_1122, n_1205, n_1408, n_163, n_1693, n_1132, n_390, n_1156, n_501, n_314, n_1120, n_1202, n_627, n_1188, n_1498, n_1371, n_233, n_957, n_388, n_1402, n_1242, n_1607, n_1489, n_1218, n_221, n_321, n_86, n_1586, n_861, n_1543, n_1431, n_877, n_1119, n_1666, n_1500, n_616, n_1055, n_1395, n_1346, n_1189, n_1089, n_281, n_262, n_1502, n_1523, n_1478, n_735, n_297, n_1005, n_527, n_46, n_84, n_1294, n_1667, n_845, n_888, n_1649, n_1677, n_1297, n_178, n_551, n_417, n_1708, n_70, n_343, n_1222, n_582, n_755, n_1097, n_1219, n_710, n_534, n_1460, n_1239, n_278, n_560, n_890, n_842, n_148, n_451, n_745, n_1572, n_61, n_742, n_1081, n_1373, n_1388, n_1266, n_1540, n_769, n_13, n_1372, n_476, n_832, n_55, n_535, n_744, n_982, n_915, n_215, n_1075, n_454, n_298, n_1331, n_1529, n_1227, n_655, n_403, n_1007, n_1580, n_1319, n_657, n_837, n_812, n_606, n_951, n_862, n_1700, n_659, n_1332, n_509, n_666, n_430, n_1206, n_722, n_1508, n_1532, n_1171, n_1030, n_785, n_1309, n_999, n_1338, n_1342, n_456, n_852, n_1394, n_704, n_1060, n_1044, n_521, n_873, n_1301, n_1243, n_1400, n_342, n_1466, n_1513, n_1527, n_358, n_608, n_1538, n_1037, n_1329, n_317, n_1545, n_134, n_1257, n_1480, n_1668, n_1605, n_1078, n_266, n_157, n_1161, n_811, n_624, n_791, n_876, n_618, n_1191, n_736, n_1025, n_1215, n_241, n_1449, n_687, n_797, n_480, n_1327, n_1475, n_211, n_642, n_97, n_408, n_1406, n_595, n_1405, n_602, n_592, n_1499, n_854, n_1318, n_393, n_1632, n_474, n_805, n_295, n_1658, n_190, n_1072, n_695, n_1526, n_1305, n_64, n_180, n_730, n_386, n_1596, n_1281, n_516, n_1137, n_1258, n_197, n_640, n_463, n_1476, n_1524, n_943, n_1118, n_678, n_651, n_1293, n_961, n_469, n_1046, n_726, n_1123, n_1657, n_878, n_771, n_1321, n_752, n_71, n_1488, n_985, n_421, n_1330, n_906, n_1180, n_1697, n_283, n_806, n_1350, n_1556, n_649, n_1561, n_374, n_1352, n_643, n_1492, n_226, n_1441, n_682, n_36, n_1616, n_819, n_586, n_1324, n_1429, n_686, n_605, n_1154, n_584, n_1557, n_1130, n_1450, n_349, n_756, n_1016, n_1149, n_1505, n_979, n_1642, n_2, n_897, n_949, n_1493, n_515, n_807, n_891, n_885, n_1659, n_198, n_1208, n_396, n_802, n_23, n_1151, n_554, n_960, n_1256, n_87, n_714, n_790, n_354, n_140, n_725, n_1577, n_151, n_1448, n_28, n_1009, n_230, n_1133, n_154, n_883, n_142, n_473, n_801, n_1286, n_818, n_1685, n_779, n_594, n_1397, n_35, n_1052, n_272, n_1333, n_1306, n_833, n_1426, n_879, n_1117, n_38, n_422, n_1269, n_1303, n_1547, n_1438, n_1541, n_597, n_75, n_1047, n_95, n_1472, n_1593, n_1050, n_566, n_152, n_169, n_106, n_1201, n_1288, n_173, n_858, n_1185, n_335, n_1035, n_1143, n_344, n_426, n_433, n_398, n_62, n_210, n_1090, n_1367, n_166, n_253, n_928, n_1153, n_271, n_465, n_825, n_1103, n_732, n_1565, n_1192, n_128, n_224, n_82, n_894, n_1380, n_1624, n_420, n_1291, n_562, n_748, n_510, n_1045, n_256, n_1160, n_1023, n_988, n_330, n_914, n_400, n_689, n_1116, n_282, n_328, n_368, n_467, n_1511, n_1422, n_644, n_1197, n_276, n_497, n_1165, n_1641, n_168, n_81, n_538, n_1517, n_576, n_843, n_511, n_455, n_429, n_588, n_638, n_1307, n_1128, n_1671, n_1417, n_1048, n_775, n_667, n_1049, n_14, n_869, n_141, n_846, n_1398, n_1356, n_1341, n_1504, n_1440, n_1370, n_1603, n_305, n_312, n_56, n_60, n_728, n_413, n_715, n_889, n_1066, n_1549, n_935, n_685, n_911, n_361, n_89, n_623, n_1403, n_1065, n_453, n_1534, n_74, n_810, n_19, n_40, n_1290, n_181, n_617, n_543, n_1362, n_1559, n_236, n_601, n_683, n_565, n_628, n_1300, n_743, n_1194, n_1647, n_1546, n_1420, n_907, n_1454, n_660, n_464, n_962, n_941, n_1210, n_847, n_747, n_1622, n_1135, n_918, n_107, n_639, n_452, n_673, n_1038, n_414, n_571, n_1521, n_1694, n_6, n_284, n_593, n_1695, n_1164, n_37, n_58, n_609, n_1193, n_1345, n_613, n_1022, n_1336, n_1033, n_409, n_171, n_519, n_384, n_1166, n_1056, n_526, n_1040, n_674, n_1158, n_316, n_125, n_1444, n_820, n_43, n_872, n_1653, n_254, n_1157, n_1584, n_234, n_848, n_1664, n_280, n_629, n_161, n_532, n_763, n_99, n_540, n_216, n_692, n_5, n_984, n_1687, n_223, n_1552, n_750, n_834, n_1612, n_800, n_1606, n_395, n_621, n_1587, n_213, n_67, n_1014, n_724, n_1427, n_1481, n_493, n_1311, n_1589, n_114, n_1100, n_585, n_875, n_1617, n_827, n_697, n_622, n_1626, n_1335, n_296, n_880, n_793, n_1175, n_132, n_751, n_1027, n_1070, n_1621, n_739, n_1485, n_1028, n_1221, n_530, n_792, n_1262, n_580, n_1579, n_494, n_434, n_975, n_229, n_394, n_923, n_1645, n_1124, n_1381, n_1494, n_932, n_1183, n_1326, n_981, n_1110, n_243, n_1407, n_185, n_1204, n_1554, n_994, n_1360, n_973, n_268, n_972, n_164, n_184, n_856, n_1248, n_1176, n_1564, n_1054, n_508, n_118, n_121, n_1679, n_353, n_1678, n_1482, n_1361, n_1601, n_1057, n_191, n_978, n_1011, n_1520, n_1509, n_828, n_322, n_1411, n_1359, n_558, n_116, n_39, n_653, n_1445, n_1317, n_783, n_556, n_1127, n_170, n_1536, n_1471, n_160, n_119, n_1008, n_332, n_581, n_294, n_1024, n_830, n_176, n_987, n_936, n_1620, n_1385, n_1525, n_541, n_499, n_788, n_12, n_908, n_1036, n_341, n_1270, n_109, n_1167, n_1272, n_549, n_591, n_969, n_919, n_1663, n_50, n_1625, n_318, n_1458, n_103, n_244, n_679, n_1630, n_220, n_663, n_443, n_1412, n_1550, n_528, n_1358, n_1200, n_387, n_406, n_826, n_139, n_391, n_940, n_1537, n_1077, n_607, n_956, n_445, n_765, n_122, n_1268, n_385, n_917, n_1271, n_372, n_15, n_1530, n_631, n_399, n_1170, n_1261, n_702, n_857, n_898, n_363, n_968, n_1067, n_1235, n_1323, n_1462, n_1064, n_633, n_900, n_1446, n_1282, n_1701, n_1093, n_1551, n_1285, n_193, n_733, n_761, n_731, n_336, n_315, n_311, n_1452, n_1573, n_8, n_668, n_758, n_1106, n_47, n_153, n_18, n_648, n_784, n_269, n_816, n_1322, n_1473, n_835, n_446, n_1076, n_1348, n_753, n_701, n_1003, n_1125, n_309, n_1344, n_115, n_1390, n_401, n_485, n_504, n_483, n_435, n_1141, n_1629, n_291, n_1640, n_822, n_1094, n_840, n_1459, n_1510, n_1099, n_839, n_79, n_3, n_759, n_567, n_91, n_240, n_369, n_44, n_1575, n_1172, n_614, n_1212, n_831, n_778, n_48, n_1619, n_188, n_323, n_550, n_1315, n_1660, n_997, n_635, n_694, n_1643, n_1320, n_1113, n_248, n_1152, n_921, n_1615, n_1236, n_228, n_1265, n_1576, n_1470, n_671, n_1533, n_1, n_1409, n_1148, n_1588, n_1684, n_1673, n_1334, n_654, n_1275, n_488, n_904, n_505, n_88, n_1696, n_498, n_1059, n_684, n_1039, n_539, n_1150, n_977, n_449, n_392, n_1628, n_1289, n_1497, n_459, n_1136, n_458, n_1190, n_1600, n_1144, n_383, n_838, n_1558, n_1316, n_175, n_950, n_1017, n_711, n_734, n_723, n_1393, n_658, n_630, n_1369, n_53, n_362, n_310, n_709, n_24, n_809, n_1686, n_235, n_881, n_1019, n_1477, n_662, n_641, n_910, n_290, n_741, n_939, n_1410, n_371, n_199, n_217, n_1114, n_1325, n_708, n_308, n_1223, n_201, n_572, n_1199, n_865, n_10, n_1273, n_1041, n_993, n_948, n_922, n_1004, n_448, n_1347, n_860, n_1043, n_255, n_450, n_896, n_1479, n_1613, n_902, n_1031, n_1638, n_853, n_716, n_1571, n_1698, n_196, n_1337, n_774, n_933, n_596, n_954, n_1168, n_219, n_1310, n_231, n_656, n_492, n_574, n_252, n_664, n_1591, n_1229, n_1683, n_68, n_415, n_63, n_1280, n_544, n_1516, n_1186, n_1705, n_599, n_768, n_1091, n_537, n_1063, n_25, n_991, n_83, n_389, n_1670, n_1707, n_1126, n_195, n_938, n_1328, n_895, n_110, n_304, n_1639, n_583, n_1302, n_1000, n_313, n_626, n_378, n_1581, n_98, n_946, n_757, n_375, n_113, n_1655, n_33, n_1146, n_1634, n_1203, n_998, n_1699, n_1598, n_472, n_937, n_1474, n_265, n_1583, n_1604, n_208, n_1631, n_1702, n_156, n_174, n_275, n_100, n_1375, n_147, n_204, n_1232, n_996, n_1211, n_1368, n_963, n_1264, n_51, n_1082, n_496, n_866, n_26, n_246, n_925, n_1313, n_1001, n_1115, n_1339, n_1002, n_1644, n_105, n_1051, n_719, n_131, n_263, n_1102, n_360, n_1129, n_1252, n_250, n_1464, n_1296, n_773, n_165, n_1010, n_882, n_1249, n_101, n_803, n_329, n_718, n_1434, n_340, n_1569, n_289, n_9, n_112, n_45, n_548, n_523, n_1662, n_457, n_1299, n_177, n_782, n_364, n_258, n_431, n_1228, n_1244, n_411, n_484, n_849, n_22, n_29, n_357, n_412, n_1251, n_447, n_1421, n_1233, n_1574, n_1672, n_1635, n_1704, n_893, n_1582, n_841, n_886, n_1069, n_359, n_1308, n_573, n_796, n_127, n_531, n_1374, n_1451, n_1487, n_675, n_7467);

input n_913;
input n_1681;
input n_1486;
input n_1507;
input n_589;
input n_1174;
input n_1469;
input n_691;
input n_1353;
input n_1355;
input n_423;
input n_1383;
input n_603;
input n_373;
input n_1250;
input n_1169;
input n_789;
input n_850;
input n_610;
input n_245;
input n_96;
input n_319;
input n_49;
input n_1436;
input n_690;
input n_416;
input n_1109;
input n_1430;
input n_525;
input n_187;
input n_1463;
input n_1238;
input n_1515;
input n_817;
input n_924;
input n_781;
input n_1566;
input n_189;
input n_717;
input n_72;
input n_952;
input n_864;
input n_1096;
input n_1379;
input n_57;
input n_1706;
input n_117;
input n_524;
input n_1214;
input n_634;
input n_1246;
input n_1138;
input n_214;
input n_764;
input n_1503;
input n_462;
input n_1196;
input n_1181;
input n_32;
input n_410;
input n_1187;
input n_1131;
input n_1225;
input n_737;
input n_137;
input n_1298;
input n_1366;
input n_232;
input n_52;
input n_568;
input n_1088;
input n_77;
input n_1424;
input n_766;
input n_1457;
input n_377;
input n_1682;
input n_520;
input n_870;
input n_1453;
input n_279;
input n_945;
input n_958;
input n_813;
input n_419;
input n_146;
input n_270;
input n_338;
input n_995;
input n_285;
input n_1184;
input n_202;
input n_1535;
input n_500;
input n_665;
input n_754;
input n_903;
input n_871;
input n_1073;
input n_239;
input n_402;
input n_1277;
input n_54;
input n_829;
input n_1062;
input n_339;
input n_738;
input n_1690;
input n_672;
input n_740;
input n_1283;
input n_167;
input n_1018;
input n_69;
input n_259;
input n_953;
input n_1364;
input n_143;
input n_1224;
input n_1425;
input n_625;
input n_557;
input n_1107;
input n_1688;
input n_989;
input n_242;
input n_645;
input n_331;
input n_559;
input n_267;
input n_495;
input n_350;
input n_381;
input n_795;
input n_721;
input n_1084;
input n_1276;
input n_200;
input n_1428;
input n_1284;
input n_1241;
input n_821;
input n_561;
input n_770;
input n_1514;
input n_1528;
input n_507;
input n_486;
input n_901;
input n_569;
input n_1145;
input n_971;
input n_787;
input n_1650;
input n_31;
input n_1519;
input n_1195;
input n_1522;
input n_518;
input n_1207;
input n_222;
input n_786;
input n_1404;
input n_868;
input n_1542;
input n_1314;
input n_1512;
input n_1539;
input n_884;
input n_1415;
input n_1034;
input n_1652;
input n_1676;
input n_1085;
input n_277;
input n_1636;
input n_432;
input n_293;
input n_823;
input n_620;
input n_93;
input n_1074;
input n_859;
input n_108;
input n_587;
input n_693;
input n_863;
input n_303;
input n_1254;
input n_929;
input n_206;
input n_352;
input n_899;
input n_1703;
input n_611;
input n_1295;
input n_238;
input n_365;
input n_1013;
input n_1495;
input n_1637;
input n_136;
input n_334;
input n_192;
input n_661;
input n_300;
input n_533;
input n_104;
input n_438;
input n_1560;
input n_1654;
input n_1548;
input n_16;
input n_440;
input n_273;
input n_1396;
input n_1230;
input n_612;
input n_333;
input n_376;
input n_512;
input n_1597;
input n_1544;
input n_579;
input n_844;
input n_1012;
input n_1267;
input n_1354;
input n_149;
input n_1213;
input n_237;
input n_780;
input n_1021;
input n_1443;
input n_491;
input n_1465;
input n_1595;
input n_1142;
input n_1140;
input n_705;
input n_570;
input n_260;
input n_942;
input n_1437;
input n_7;
input n_1378;
input n_461;
input n_1121;
input n_1416;
input n_209;
input n_490;
input n_1461;
input n_17;
input n_1391;
input n_225;
input n_1599;
input n_1006;
input n_575;
input n_546;
input n_503;
input n_1112;
input n_700;
input n_1159;
input n_772;
input n_1216;
input n_1245;
input n_1669;
input n_1675;
input n_676;
input n_42;
input n_1594;
input n_680;
input n_287;
input n_302;
input n_380;
input n_1585;
input n_1432;
input n_94;
input n_4;
input n_249;
input n_1108;
input n_355;
input n_212;
input n_65;
input n_123;
input n_444;
input n_851;
input n_1590;
input n_1351;
input n_1274;
input n_257;
input n_652;
input n_475;
input n_135;
input n_947;
input n_930;
input n_1260;
input n_1179;
input n_468;
input n_102;
input n_182;
input n_696;
input n_1442;
input n_482;
input n_798;
input n_577;
input n_407;
input n_1691;
input n_27;
input n_916;
input n_1386;
input n_912;
input n_460;
input n_1555;
input n_366;
input n_762;
input n_1253;
input n_1468;
input n_1661;
input n_555;
input n_804;
input n_1656;
input n_1382;
input n_966;
input n_992;
input n_955;
input n_1182;
input n_794;
input n_78;
input n_1692;
input n_1562;
input n_514;
input n_418;
input n_1376;
input n_513;
input n_288;
input n_179;
input n_1292;
input n_1178;
input n_1435;
input n_1026;
input n_1506;
input n_1610;
input n_306;
input n_92;
input n_203;
input n_436;
input n_150;
input n_324;
input n_669;
input n_931;
input n_1491;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_967;
input n_1083;
input n_1418;
input n_746;
input n_1357;
input n_292;
input n_1079;
input n_1389;
input n_615;
input n_1139;
input n_76;
input n_517;
input n_1312;
input n_0;
input n_824;
input n_428;
input n_159;
input n_892;
input n_959;
input n_30;
input n_1399;
input n_1101;
input n_1567;
input n_1343;
input n_563;
input n_144;
input n_990;
input n_1623;
input n_867;
input n_1226;
input n_944;
input n_749;
input n_815;
input n_542;
input n_1340;
input n_470;
input n_1240;
input n_1087;
input n_632;
input n_477;
input n_650;
input n_425;
input n_1433;
input n_1155;
input n_1071;
input n_712;
input n_976;
input n_909;
input n_1392;
input n_767;
input n_1680;
input n_964;
input n_1627;
input n_382;
input n_489;
input n_80;
input n_251;
input n_974;
input n_506;
input n_799;
input n_1147;
input n_397;
input n_471;
input n_351;
input n_965;
input n_155;
input n_934;
input n_1447;
input n_1220;
input n_356;
input n_698;
input n_1674;
input n_124;
input n_307;
input n_1209;
input n_1020;
input n_1563;
input n_646;
input n_1633;
input n_34;
input n_404;
input n_172;
input n_1058;
input n_347;
input n_1042;
input n_183;
input n_1234;
input n_479;
input n_1578;
input n_1455;
input n_299;
input n_836;
input n_1279;
input n_564;
input n_133;
input n_66;
input n_205;
input n_1029;
input n_1247;
input n_760;
input n_522;
input n_1568;
input n_20;
input n_1483;
input n_1363;
input n_367;
input n_1111;
input n_970;
input n_1689;
input n_713;
input n_1255;
input n_1646;
input n_598;
input n_345;
input n_1237;
input n_927;
input n_261;
input n_1095;
input n_370;
input n_706;
input n_286;
input n_1401;
input n_1419;
input n_1531;
input n_776;
input n_424;
input n_1651;
input n_85;
input n_130;
input n_1387;
input n_466;
input n_1263;
input n_346;
input n_348;
input n_552;
input n_670;
input n_379;
input n_138;
input n_162;
input n_264;
input n_441;
input n_1032;
input n_1217;
input n_1496;
input n_637;
input n_1592;
input n_73;
input n_327;
input n_1259;
input n_1177;
input n_1231;
input n_980;
input n_1618;
input n_905;
input n_207;
input n_720;
input n_926;
input n_41;
input n_194;
input n_1163;
input n_186;
input n_1384;
input n_145;
input n_59;
input n_1501;
input n_1173;
input n_1068;
input n_1198;
input n_1570;
input n_487;
input n_1518;
input n_1456;
input n_90;
input n_1648;
input n_1413;
input n_855;
input n_158;
input n_808;
input n_1365;
input n_553;
input n_1439;
input n_814;
input n_578;
input n_1665;
input n_1287;
input n_405;
input n_1611;
input n_120;
input n_320;
input n_1414;
input n_1134;
input n_1484;
input n_647;
input n_1423;
input n_481;
input n_600;
input n_1053;
input n_1609;
input n_529;
input n_502;
input n_218;
input n_1467;
input n_247;
input n_1304;
input n_1608;
input n_1105;
input n_547;
input n_439;
input n_604;
input n_677;
input n_478;
input n_703;
input n_1349;
input n_1061;
input n_326;
input n_681;
input n_227;
input n_874;
input n_1278;
input n_707;
input n_11;
input n_129;
input n_126;
input n_983;
input n_590;
input n_699;
input n_727;
input n_301;
input n_545;
input n_1015;
input n_1377;
input n_1162;
input n_536;
input n_1614;
input n_325;
input n_1602;
input n_688;
input n_636;
input n_427;
input n_1098;
input n_1490;
input n_442;
input n_777;
input n_1553;
input n_1080;
input n_920;
input n_1086;
input n_1092;
input n_986;
input n_1104;
input n_729;
input n_887;
input n_1122;
input n_1205;
input n_1408;
input n_163;
input n_1693;
input n_1132;
input n_390;
input n_1156;
input n_501;
input n_314;
input n_1120;
input n_1202;
input n_627;
input n_1188;
input n_1498;
input n_1371;
input n_233;
input n_957;
input n_388;
input n_1402;
input n_1242;
input n_1607;
input n_1489;
input n_1218;
input n_221;
input n_321;
input n_86;
input n_1586;
input n_861;
input n_1543;
input n_1431;
input n_877;
input n_1119;
input n_1666;
input n_1500;
input n_616;
input n_1055;
input n_1395;
input n_1346;
input n_1189;
input n_1089;
input n_281;
input n_262;
input n_1502;
input n_1523;
input n_1478;
input n_735;
input n_297;
input n_1005;
input n_527;
input n_46;
input n_84;
input n_1294;
input n_1667;
input n_845;
input n_888;
input n_1649;
input n_1677;
input n_1297;
input n_178;
input n_551;
input n_417;
input n_1708;
input n_70;
input n_343;
input n_1222;
input n_582;
input n_755;
input n_1097;
input n_1219;
input n_710;
input n_534;
input n_1460;
input n_1239;
input n_278;
input n_560;
input n_890;
input n_842;
input n_148;
input n_451;
input n_745;
input n_1572;
input n_61;
input n_742;
input n_1081;
input n_1373;
input n_1388;
input n_1266;
input n_1540;
input n_769;
input n_13;
input n_1372;
input n_476;
input n_832;
input n_55;
input n_535;
input n_744;
input n_982;
input n_915;
input n_215;
input n_1075;
input n_454;
input n_298;
input n_1331;
input n_1529;
input n_1227;
input n_655;
input n_403;
input n_1007;
input n_1580;
input n_1319;
input n_657;
input n_837;
input n_812;
input n_606;
input n_951;
input n_862;
input n_1700;
input n_659;
input n_1332;
input n_509;
input n_666;
input n_430;
input n_1206;
input n_722;
input n_1508;
input n_1532;
input n_1171;
input n_1030;
input n_785;
input n_1309;
input n_999;
input n_1338;
input n_1342;
input n_456;
input n_852;
input n_1394;
input n_704;
input n_1060;
input n_1044;
input n_521;
input n_873;
input n_1301;
input n_1243;
input n_1400;
input n_342;
input n_1466;
input n_1513;
input n_1527;
input n_358;
input n_608;
input n_1538;
input n_1037;
input n_1329;
input n_317;
input n_1545;
input n_134;
input n_1257;
input n_1480;
input n_1668;
input n_1605;
input n_1078;
input n_266;
input n_157;
input n_1161;
input n_811;
input n_624;
input n_791;
input n_876;
input n_618;
input n_1191;
input n_736;
input n_1025;
input n_1215;
input n_241;
input n_1449;
input n_687;
input n_797;
input n_480;
input n_1327;
input n_1475;
input n_211;
input n_642;
input n_97;
input n_408;
input n_1406;
input n_595;
input n_1405;
input n_602;
input n_592;
input n_1499;
input n_854;
input n_1318;
input n_393;
input n_1632;
input n_474;
input n_805;
input n_295;
input n_1658;
input n_190;
input n_1072;
input n_695;
input n_1526;
input n_1305;
input n_64;
input n_180;
input n_730;
input n_386;
input n_1596;
input n_1281;
input n_516;
input n_1137;
input n_1258;
input n_197;
input n_640;
input n_463;
input n_1476;
input n_1524;
input n_943;
input n_1118;
input n_678;
input n_651;
input n_1293;
input n_961;
input n_469;
input n_1046;
input n_726;
input n_1123;
input n_1657;
input n_878;
input n_771;
input n_1321;
input n_752;
input n_71;
input n_1488;
input n_985;
input n_421;
input n_1330;
input n_906;
input n_1180;
input n_1697;
input n_283;
input n_806;
input n_1350;
input n_1556;
input n_649;
input n_1561;
input n_374;
input n_1352;
input n_643;
input n_1492;
input n_226;
input n_1441;
input n_682;
input n_36;
input n_1616;
input n_819;
input n_586;
input n_1324;
input n_1429;
input n_686;
input n_605;
input n_1154;
input n_584;
input n_1557;
input n_1130;
input n_1450;
input n_349;
input n_756;
input n_1016;
input n_1149;
input n_1505;
input n_979;
input n_1642;
input n_2;
input n_897;
input n_949;
input n_1493;
input n_515;
input n_807;
input n_891;
input n_885;
input n_1659;
input n_198;
input n_1208;
input n_396;
input n_802;
input n_23;
input n_1151;
input n_554;
input n_960;
input n_1256;
input n_87;
input n_714;
input n_790;
input n_354;
input n_140;
input n_725;
input n_1577;
input n_151;
input n_1448;
input n_28;
input n_1009;
input n_230;
input n_1133;
input n_154;
input n_883;
input n_142;
input n_473;
input n_801;
input n_1286;
input n_818;
input n_1685;
input n_779;
input n_594;
input n_1397;
input n_35;
input n_1052;
input n_272;
input n_1333;
input n_1306;
input n_833;
input n_1426;
input n_879;
input n_1117;
input n_38;
input n_422;
input n_1269;
input n_1303;
input n_1547;
input n_1438;
input n_1541;
input n_597;
input n_75;
input n_1047;
input n_95;
input n_1472;
input n_1593;
input n_1050;
input n_566;
input n_152;
input n_169;
input n_106;
input n_1201;
input n_1288;
input n_173;
input n_858;
input n_1185;
input n_335;
input n_1035;
input n_1143;
input n_344;
input n_426;
input n_433;
input n_398;
input n_62;
input n_210;
input n_1090;
input n_1367;
input n_166;
input n_253;
input n_928;
input n_1153;
input n_271;
input n_465;
input n_825;
input n_1103;
input n_732;
input n_1565;
input n_1192;
input n_128;
input n_224;
input n_82;
input n_894;
input n_1380;
input n_1624;
input n_420;
input n_1291;
input n_562;
input n_748;
input n_510;
input n_1045;
input n_256;
input n_1160;
input n_1023;
input n_988;
input n_330;
input n_914;
input n_400;
input n_689;
input n_1116;
input n_282;
input n_328;
input n_368;
input n_467;
input n_1511;
input n_1422;
input n_644;
input n_1197;
input n_276;
input n_497;
input n_1165;
input n_1641;
input n_168;
input n_81;
input n_538;
input n_1517;
input n_576;
input n_843;
input n_511;
input n_455;
input n_429;
input n_588;
input n_638;
input n_1307;
input n_1128;
input n_1671;
input n_1417;
input n_1048;
input n_775;
input n_667;
input n_1049;
input n_14;
input n_869;
input n_141;
input n_846;
input n_1398;
input n_1356;
input n_1341;
input n_1504;
input n_1440;
input n_1370;
input n_1603;
input n_305;
input n_312;
input n_56;
input n_60;
input n_728;
input n_413;
input n_715;
input n_889;
input n_1066;
input n_1549;
input n_935;
input n_685;
input n_911;
input n_361;
input n_89;
input n_623;
input n_1403;
input n_1065;
input n_453;
input n_1534;
input n_74;
input n_810;
input n_19;
input n_40;
input n_1290;
input n_181;
input n_617;
input n_543;
input n_1362;
input n_1559;
input n_236;
input n_601;
input n_683;
input n_565;
input n_628;
input n_1300;
input n_743;
input n_1194;
input n_1647;
input n_1546;
input n_1420;
input n_907;
input n_1454;
input n_660;
input n_464;
input n_962;
input n_941;
input n_1210;
input n_847;
input n_747;
input n_1622;
input n_1135;
input n_918;
input n_107;
input n_639;
input n_452;
input n_673;
input n_1038;
input n_414;
input n_571;
input n_1521;
input n_1694;
input n_6;
input n_284;
input n_593;
input n_1695;
input n_1164;
input n_37;
input n_58;
input n_609;
input n_1193;
input n_1345;
input n_613;
input n_1022;
input n_1336;
input n_1033;
input n_409;
input n_171;
input n_519;
input n_384;
input n_1166;
input n_1056;
input n_526;
input n_1040;
input n_674;
input n_1158;
input n_316;
input n_125;
input n_1444;
input n_820;
input n_43;
input n_872;
input n_1653;
input n_254;
input n_1157;
input n_1584;
input n_234;
input n_848;
input n_1664;
input n_280;
input n_629;
input n_161;
input n_532;
input n_763;
input n_99;
input n_540;
input n_216;
input n_692;
input n_5;
input n_984;
input n_1687;
input n_223;
input n_1552;
input n_750;
input n_834;
input n_1612;
input n_800;
input n_1606;
input n_395;
input n_621;
input n_1587;
input n_213;
input n_67;
input n_1014;
input n_724;
input n_1427;
input n_1481;
input n_493;
input n_1311;
input n_1589;
input n_114;
input n_1100;
input n_585;
input n_875;
input n_1617;
input n_827;
input n_697;
input n_622;
input n_1626;
input n_1335;
input n_296;
input n_880;
input n_793;
input n_1175;
input n_132;
input n_751;
input n_1027;
input n_1070;
input n_1621;
input n_739;
input n_1485;
input n_1028;
input n_1221;
input n_530;
input n_792;
input n_1262;
input n_580;
input n_1579;
input n_494;
input n_434;
input n_975;
input n_229;
input n_394;
input n_923;
input n_1645;
input n_1124;
input n_1381;
input n_1494;
input n_932;
input n_1183;
input n_1326;
input n_981;
input n_1110;
input n_243;
input n_1407;
input n_185;
input n_1204;
input n_1554;
input n_994;
input n_1360;
input n_973;
input n_268;
input n_972;
input n_164;
input n_184;
input n_856;
input n_1248;
input n_1176;
input n_1564;
input n_1054;
input n_508;
input n_118;
input n_121;
input n_1679;
input n_353;
input n_1678;
input n_1482;
input n_1361;
input n_1601;
input n_1057;
input n_191;
input n_978;
input n_1011;
input n_1520;
input n_1509;
input n_828;
input n_322;
input n_1411;
input n_1359;
input n_558;
input n_116;
input n_39;
input n_653;
input n_1445;
input n_1317;
input n_783;
input n_556;
input n_1127;
input n_170;
input n_1536;
input n_1471;
input n_160;
input n_119;
input n_1008;
input n_332;
input n_581;
input n_294;
input n_1024;
input n_830;
input n_176;
input n_987;
input n_936;
input n_1620;
input n_1385;
input n_1525;
input n_541;
input n_499;
input n_788;
input n_12;
input n_908;
input n_1036;
input n_341;
input n_1270;
input n_109;
input n_1167;
input n_1272;
input n_549;
input n_591;
input n_969;
input n_919;
input n_1663;
input n_50;
input n_1625;
input n_318;
input n_1458;
input n_103;
input n_244;
input n_679;
input n_1630;
input n_220;
input n_663;
input n_443;
input n_1412;
input n_1550;
input n_528;
input n_1358;
input n_1200;
input n_387;
input n_406;
input n_826;
input n_139;
input n_391;
input n_940;
input n_1537;
input n_1077;
input n_607;
input n_956;
input n_445;
input n_765;
input n_122;
input n_1268;
input n_385;
input n_917;
input n_1271;
input n_372;
input n_15;
input n_1530;
input n_631;
input n_399;
input n_1170;
input n_1261;
input n_702;
input n_857;
input n_898;
input n_363;
input n_968;
input n_1067;
input n_1235;
input n_1323;
input n_1462;
input n_1064;
input n_633;
input n_900;
input n_1446;
input n_1282;
input n_1701;
input n_1093;
input n_1551;
input n_1285;
input n_193;
input n_733;
input n_761;
input n_731;
input n_336;
input n_315;
input n_311;
input n_1452;
input n_1573;
input n_8;
input n_668;
input n_758;
input n_1106;
input n_47;
input n_153;
input n_18;
input n_648;
input n_784;
input n_269;
input n_816;
input n_1322;
input n_1473;
input n_835;
input n_446;
input n_1076;
input n_1348;
input n_753;
input n_701;
input n_1003;
input n_1125;
input n_309;
input n_1344;
input n_115;
input n_1390;
input n_401;
input n_485;
input n_504;
input n_483;
input n_435;
input n_1141;
input n_1629;
input n_291;
input n_1640;
input n_822;
input n_1094;
input n_840;
input n_1459;
input n_1510;
input n_1099;
input n_839;
input n_79;
input n_3;
input n_759;
input n_567;
input n_91;
input n_240;
input n_369;
input n_44;
input n_1575;
input n_1172;
input n_614;
input n_1212;
input n_831;
input n_778;
input n_48;
input n_1619;
input n_188;
input n_323;
input n_550;
input n_1315;
input n_1660;
input n_997;
input n_635;
input n_694;
input n_1643;
input n_1320;
input n_1113;
input n_248;
input n_1152;
input n_921;
input n_1615;
input n_1236;
input n_228;
input n_1265;
input n_1576;
input n_1470;
input n_671;
input n_1533;
input n_1;
input n_1409;
input n_1148;
input n_1588;
input n_1684;
input n_1673;
input n_1334;
input n_654;
input n_1275;
input n_488;
input n_904;
input n_505;
input n_88;
input n_1696;
input n_498;
input n_1059;
input n_684;
input n_1039;
input n_539;
input n_1150;
input n_977;
input n_449;
input n_392;
input n_1628;
input n_1289;
input n_1497;
input n_459;
input n_1136;
input n_458;
input n_1190;
input n_1600;
input n_1144;
input n_383;
input n_838;
input n_1558;
input n_1316;
input n_175;
input n_950;
input n_1017;
input n_711;
input n_734;
input n_723;
input n_1393;
input n_658;
input n_630;
input n_1369;
input n_53;
input n_362;
input n_310;
input n_709;
input n_24;
input n_809;
input n_1686;
input n_235;
input n_881;
input n_1019;
input n_1477;
input n_662;
input n_641;
input n_910;
input n_290;
input n_741;
input n_939;
input n_1410;
input n_371;
input n_199;
input n_217;
input n_1114;
input n_1325;
input n_708;
input n_308;
input n_1223;
input n_201;
input n_572;
input n_1199;
input n_865;
input n_10;
input n_1273;
input n_1041;
input n_993;
input n_948;
input n_922;
input n_1004;
input n_448;
input n_1347;
input n_860;
input n_1043;
input n_255;
input n_450;
input n_896;
input n_1479;
input n_1613;
input n_902;
input n_1031;
input n_1638;
input n_853;
input n_716;
input n_1571;
input n_1698;
input n_196;
input n_1337;
input n_774;
input n_933;
input n_596;
input n_954;
input n_1168;
input n_219;
input n_1310;
input n_231;
input n_656;
input n_492;
input n_574;
input n_252;
input n_664;
input n_1591;
input n_1229;
input n_1683;
input n_68;
input n_415;
input n_63;
input n_1280;
input n_544;
input n_1516;
input n_1186;
input n_1705;
input n_599;
input n_768;
input n_1091;
input n_537;
input n_1063;
input n_25;
input n_991;
input n_83;
input n_389;
input n_1670;
input n_1707;
input n_1126;
input n_195;
input n_938;
input n_1328;
input n_895;
input n_110;
input n_304;
input n_1639;
input n_583;
input n_1302;
input n_1000;
input n_313;
input n_626;
input n_378;
input n_1581;
input n_98;
input n_946;
input n_757;
input n_375;
input n_113;
input n_1655;
input n_33;
input n_1146;
input n_1634;
input n_1203;
input n_998;
input n_1699;
input n_1598;
input n_472;
input n_937;
input n_1474;
input n_265;
input n_1583;
input n_1604;
input n_208;
input n_1631;
input n_1702;
input n_156;
input n_174;
input n_275;
input n_100;
input n_1375;
input n_147;
input n_204;
input n_1232;
input n_996;
input n_1211;
input n_1368;
input n_963;
input n_1264;
input n_51;
input n_1082;
input n_496;
input n_866;
input n_26;
input n_246;
input n_925;
input n_1313;
input n_1001;
input n_1115;
input n_1339;
input n_1002;
input n_1644;
input n_105;
input n_1051;
input n_719;
input n_131;
input n_263;
input n_1102;
input n_360;
input n_1129;
input n_1252;
input n_250;
input n_1464;
input n_1296;
input n_773;
input n_165;
input n_1010;
input n_882;
input n_1249;
input n_101;
input n_803;
input n_329;
input n_718;
input n_1434;
input n_340;
input n_1569;
input n_289;
input n_9;
input n_112;
input n_45;
input n_548;
input n_523;
input n_1662;
input n_457;
input n_1299;
input n_177;
input n_782;
input n_364;
input n_258;
input n_431;
input n_1228;
input n_1244;
input n_411;
input n_484;
input n_849;
input n_22;
input n_29;
input n_357;
input n_412;
input n_1251;
input n_447;
input n_1421;
input n_1233;
input n_1574;
input n_1672;
input n_1635;
input n_1704;
input n_893;
input n_1582;
input n_841;
input n_886;
input n_1069;
input n_359;
input n_1308;
input n_573;
input n_796;
input n_127;
input n_531;
input n_1374;
input n_1451;
input n_1487;
input n_675;

output n_7467;

wire n_3527;
wire n_2752;
wire n_4474;
wire n_7329;
wire n_4030;
wire n_7029;
wire n_6790;
wire n_4770;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_6603;
wire n_2679;
wire n_6557;
wire n_5402;
wire n_6581;
wire n_2182;
wire n_5553;
wire n_6002;
wire n_7277;
wire n_2680;
wire n_3264;
wire n_5717;
wire n_2993;
wire n_4283;
wire n_2879;
wire n_4403;
wire n_4962;
wire n_2002;
wire n_2729;
wire n_4302;
wire n_5791;
wire n_7127;
wire n_4547;
wire n_5090;
wire n_3765;
wire n_5302;
wire n_2376;
wire n_2790;
wire n_2207;
wire n_7053;
wire n_5712;
wire n_3954;
wire n_6297;
wire n_4982;
wire n_2042;
wire n_5479;
wire n_2646;
wire n_2653;
wire n_4610;
wire n_6058;
wire n_3115;
wire n_4028;
wire n_5263;
wire n_5565;
wire n_6358;
wire n_6293;
wire n_2482;
wire n_7001;
wire n_6129;
wire n_2554;
wire n_4321;
wire n_1985;
wire n_5590;
wire n_2621;
wire n_6524;
wire n_4853;
wire n_1909;
wire n_5229;
wire n_6313;
wire n_7464;
wire n_4260;
wire n_3348;
wire n_3261;
wire n_1761;
wire n_7368;
wire n_2807;
wire n_6664;
wire n_7428;
wire n_4512;
wire n_6190;
wire n_4132;
wire n_7373;
wire n_2390;
wire n_6891;
wire n_4500;
wire n_2322;
wire n_2663;
wire n_5481;
wire n_6539;
wire n_4824;
wire n_5340;
wire n_3545;
wire n_6797;
wire n_7392;
wire n_4741;
wire n_4143;
wire n_4273;
wire n_4136;
wire n_3144;
wire n_2359;
wire n_5896;
wire n_7338;
wire n_4567;
wire n_5833;
wire n_6249;
wire n_6887;
wire n_6253;
wire n_6128;
wire n_3552;
wire n_2950;
wire n_6197;
wire n_7200;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_5589;
wire n_3015;
wire n_5744;
wire n_3870;
wire n_6808;
wire n_3749;
wire n_5691;
wire n_3482;
wire n_6295;
wire n_5403;
wire n_1900;
wire n_6096;
wire n_4268;
wire n_6338;
wire n_6992;
wire n_3960;
wire n_2433;
wire n_3975;
wire n_5830;
wire n_2004;
wire n_4018;
wire n_3325;
wire n_6681;
wire n_4227;
wire n_5158;
wire n_5152;
wire n_1917;
wire n_2456;
wire n_5092;
wire n_1924;
wire n_6542;
wire n_1811;
wire n_6161;
wire n_3612;
wire n_4505;
wire n_6452;
wire n_1840;
wire n_5247;
wire n_5464;
wire n_7306;
wire n_4476;
wire n_6740;
wire n_6978;
wire n_2956;
wire n_5210;
wire n_7215;
wire n_2382;
wire n_7379;
wire n_7441;
wire n_5292;
wire n_1918;
wire n_7438;
wire n_4119;
wire n_4443;
wire n_4000;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_6136;
wire n_3458;
wire n_5843;
wire n_7108;
wire n_3511;
wire n_2077;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_6156;
wire n_4908;
wire n_3754;
wire n_5060;
wire n_7162;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_7331;
wire n_5913;
wire n_4530;
wire n_2245;
wire n_5614;
wire n_5391;
wire n_5452;
wire n_3359;
wire n_3841;
wire n_5249;
wire n_3900;
wire n_3413;
wire n_5076;
wire n_3539;
wire n_5757;
wire n_6872;
wire n_6644;
wire n_5062;
wire n_2134;
wire n_3862;
wire n_4912;
wire n_4226;
wire n_4311;
wire n_3284;
wire n_5046;
wire n_6236;
wire n_7104;
wire n_3506;
wire n_4827;
wire n_6801;
wire n_1842;
wire n_4993;
wire n_7397;
wire n_3678;
wire n_7205;
wire n_2791;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_6563;
wire n_5968;
wire n_3549;
wire n_3914;
wire n_6398;
wire n_5586;
wire n_7461;
wire n_2611;
wire n_5468;
wire n_3029;
wire n_4745;
wire n_2398;
wire n_4233;
wire n_4791;
wire n_5971;
wire n_6319;
wire n_7224;
wire n_6966;
wire n_5056;
wire n_2015;
wire n_7259;
wire n_5984;
wire n_5204;
wire n_6705;
wire n_6724;
wire n_2877;
wire n_7307;
wire n_6776;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_2161;
wire n_6624;
wire n_6710;
wire n_1787;
wire n_6883;
wire n_3172;
wire n_4033;
wire n_2659;
wire n_3747;
wire n_6553;
wire n_4905;
wire n_4508;
wire n_5897;
wire n_4045;
wire n_4894;
wire n_3651;
wire n_1812;
wire n_6261;
wire n_6659;
wire n_7351;
wire n_3614;
wire n_7256;
wire n_2257;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_6893;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_3559;
wire n_5778;
wire n_7021;
wire n_5179;
wire n_2435;
wire n_6337;
wire n_5680;
wire n_1932;
wire n_6210;
wire n_1780;
wire n_2825;
wire n_5685;
wire n_5974;
wire n_5723;
wire n_5922;
wire n_6378;
wire n_5549;
wire n_2388;
wire n_2273;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_3700;
wire n_4307;
wire n_2795;
wire n_6044;
wire n_1841;
wire n_6206;
wire n_2954;
wire n_4438;
wire n_6538;
wire n_3814;
wire n_6996;
wire n_5831;
wire n_4367;
wire n_5134;
wire n_2467;
wire n_7231;
wire n_4195;
wire n_7007;
wire n_6579;
wire n_5091;
wire n_4866;
wire n_7230;
wire n_2019;
wire n_5708;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_5454;
wire n_4254;
wire n_3438;
wire n_2625;
wire n_5373;
wire n_7403;
wire n_6665;
wire n_3147;
wire n_3661;
wire n_7168;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_2649;
wire n_6033;
wire n_6461;
wire n_6860;
wire n_2919;
wire n_7322;
wire n_6060;
wire n_3108;
wire n_5788;
wire n_5983;
wire n_6709;
wire n_2632;
wire n_5557;
wire n_6914;
wire n_4314;
wire n_2980;
wire n_5951;
wire n_1728;
wire n_4315;
wire n_5647;
wire n_6117;
wire n_7287;
wire n_3239;
wire n_2631;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_4857;
wire n_3087;
wire n_6009;
wire n_7221;
wire n_4637;
wire n_5523;
wire n_2697;
wire n_1817;
wire n_3704;
wire n_6382;
wire n_2677;
wire n_4296;
wire n_2483;
wire n_5088;
wire n_6615;
wire n_7294;
wire n_6192;
wire n_5773;
wire n_7414;
wire n_5392;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_3589;
wire n_6418;
wire n_1743;
wire n_6263;
wire n_1943;
wire n_6731;
wire n_5138;
wire n_4588;
wire n_6048;
wire n_7185;
wire n_5149;
wire n_3054;
wire n_4970;
wire n_5280;
wire n_6234;
wire n_4153;
wire n_1868;
wire n_5052;
wire n_3601;
wire n_5137;
wire n_7141;
wire n_2373;
wire n_3881;
wire n_6224;
wire n_5089;
wire n_5775;
wire n_2099;
wire n_3759;
wire n_3323;
wire n_4643;
wire n_6142;
wire n_2617;
wire n_6119;
wire n_6619;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_6759;
wire n_6903;
wire n_3466;
wire n_7416;
wire n_2074;
wire n_5031;
wire n_6768;
wire n_7092;
wire n_7233;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_5082;
wire n_4788;
wire n_2067;
wire n_4555;
wire n_5230;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_7191;
wire n_2117;
wire n_6189;
wire n_5796;
wire n_5296;
wire n_5398;
wire n_1906;
wire n_6761;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_1828;
wire n_7202;
wire n_3335;
wire n_5960;
wire n_3007;
wire n_2267;
wire n_7445;
wire n_5858;
wire n_5985;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_3370;
wire n_3949;
wire n_2286;
wire n_5192;
wire n_4247;
wire n_5051;
wire n_5336;
wire n_3036;
wire n_2783;
wire n_4583;
wire n_6366;
wire n_6304;
wire n_4292;
wire n_2118;
wire n_7176;
wire n_5552;
wire n_6074;
wire n_3764;
wire n_4773;
wire n_1760;
wire n_5028;
wire n_3025;
wire n_3051;
wire n_2802;
wire n_2125;
wire n_5123;
wire n_4974;
wire n_6689;
wire n_2861;
wire n_4344;
wire n_5242;
wire n_3130;
wire n_4856;
wire n_2618;
wire n_7096;
wire n_4216;
wire n_2707;
wire n_5596;
wire n_6482;
wire n_2849;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_6335;
wire n_5742;
wire n_5127;
wire n_4313;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_3713;
wire n_6229;
wire n_1863;
wire n_5933;
wire n_5536;
wire n_4798;
wire n_7293;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_5810;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_7144;
wire n_2190;
wire n_3931;
wire n_2516;
wire n_4991;
wire n_7316;
wire n_3070;
wire n_5818;
wire n_3275;
wire n_5198;
wire n_3245;
wire n_2894;
wire n_2452;
wire n_4182;
wire n_2827;
wire n_3214;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5539;
wire n_5009;
wire n_3710;
wire n_1844;
wire n_6943;
wire n_1957;
wire n_1953;
wire n_6631;
wire n_5889;
wire n_7151;
wire n_3944;
wire n_5632;
wire n_4729;
wire n_6728;
wire n_1793;
wire n_4446;
wire n_4662;
wire n_5613;
wire n_4800;
wire n_7075;
wire n_5427;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_6770;
wire n_5450;
wire n_6508;
wire n_2821;
wire n_3696;
wire n_4781;
wire n_6031;
wire n_3531;
wire n_5124;
wire n_4237;
wire n_5297;
wire n_4828;
wire n_3333;
wire n_4652;
wire n_4114;
wire n_7105;
wire n_7013;
wire n_3135;
wire n_4925;
wire n_5719;
wire n_7254;
wire n_2448;
wire n_2211;
wire n_5904;
wire n_6628;
wire n_5318;
wire n_5374;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_6456;
wire n_7407;
wire n_3277;
wire n_4863;
wire n_1766;
wire n_5463;
wire n_2978;
wire n_6328;
wire n_6929;
wire n_4859;
wire n_4568;
wire n_3617;
wire n_6012;
wire n_2958;
wire n_1714;
wire n_4429;
wire n_5435;
wire n_6484;
wire n_3340;
wire n_5053;
wire n_7182;
wire n_5476;
wire n_5483;
wire n_5511;
wire n_3486;
wire n_6639;
wire n_2457;
wire n_2992;
wire n_6124;
wire n_3197;
wire n_7423;
wire n_3256;
wire n_1878;
wire n_7375;
wire n_7076;
wire n_6344;
wire n_6435;
wire n_3646;
wire n_5829;
wire n_2520;
wire n_7419;
wire n_6600;
wire n_7010;
wire n_5881;
wire n_3864;
wire n_4694;
wire n_4664;
wire n_6201;
wire n_3450;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_5073;
wire n_6555;
wire n_4306;
wire n_6360;
wire n_6735;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_3266;
wire n_3102;
wire n_6803;
wire n_4288;
wire n_3452;
wire n_4098;
wire n_2691;
wire n_5894;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_2991;
wire n_5419;
wire n_4289;
wire n_4972;
wire n_2723;
wire n_6036;
wire n_7346;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_5165;
wire n_2850;
wire n_1874;
wire n_5077;
wire n_6102;
wire n_3780;
wire n_6650;
wire n_6573;
wire n_6904;
wire n_3753;
wire n_6329;
wire n_7385;
wire n_6244;
wire n_4846;
wire n_6204;
wire n_2295;
wire n_5225;
wire n_7295;
wire n_4076;
wire n_7148;
wire n_3142;
wire n_7169;
wire n_3129;
wire n_3495;
wire n_3843;
wire n_6756;
wire n_4805;
wire n_2606;
wire n_2386;
wire n_5826;
wire n_4822;
wire n_6946;
wire n_5931;
wire n_1829;
wire n_4635;
wire n_5532;
wire n_7311;
wire n_3740;
wire n_6804;
wire n_5441;
wire n_6179;
wire n_2417;
wire n_6059;
wire n_1815;
wire n_7039;
wire n_2911;
wire n_3313;
wire n_2354;
wire n_6427;
wire n_4281;
wire n_3945;
wire n_5994;
wire n_3726;
wire n_4419;
wire n_5405;
wire n_5365;
wire n_3560;
wire n_3345;
wire n_5772;
wire n_6442;
wire n_6188;
wire n_3421;
wire n_3548;
wire n_4906;
wire n_6846;
wire n_4630;
wire n_6840;
wire n_6645;
wire n_4829;
wire n_6749;
wire n_6915;
wire n_2612;
wire n_5259;
wire n_3236;
wire n_1995;
wire n_7455;
wire n_5921;
wire n_6247;
wire n_1849;
wire n_4966;
wire n_2250;
wire n_6104;
wire n_3321;
wire n_4188;
wire n_2001;
wire n_6205;
wire n_2506;
wire n_2413;
wire n_4825;
wire n_3715;
wire n_2610;
wire n_2626;
wire n_7315;
wire n_2892;
wire n_6939;
wire n_2605;
wire n_2804;
wire n_5884;
wire n_5006;
wire n_4882;
wire n_3206;
wire n_5728;
wire n_3475;
wire n_4878;
wire n_2070;
wire n_6706;
wire n_7431;
wire n_3842;
wire n_4202;
wire n_6909;
wire n_2044;
wire n_5679;
wire n_6487;
wire n_3886;
wire n_2619;
wire n_5141;
wire n_3098;
wire n_6627;
wire n_4503;
wire n_7253;
wire n_5208;
wire n_5113;
wire n_3987;
wire n_5205;
wire n_4249;
wire n_3160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_7452;
wire n_6551;
wire n_3386;
wire n_3921;
wire n_2177;
wire n_6516;
wire n_2766;
wire n_4196;
wire n_7318;
wire n_2613;
wire n_7411;
wire n_7326;
wire n_5667;
wire n_2647;
wire n_5508;
wire n_5105;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_5879;
wire n_6500;
wire n_5027;
wire n_2343;
wire n_3380;
wire n_5688;
wire n_2826;
wire n_5825;
wire n_1921;
wire n_6630;
wire n_5629;
wire n_5759;
wire n_2411;
wire n_4631;
wire n_6798;
wire n_5999;
wire n_2110;
wire n_6421;
wire n_5377;
wire n_6180;
wire n_3822;
wire n_4355;
wire n_7453;
wire n_3818;
wire n_5599;
wire n_3587;
wire n_2608;
wire n_6004;
wire n_1948;
wire n_6652;
wire n_7183;
wire n_4155;
wire n_4278;
wire n_4710;
wire n_1959;
wire n_6275;
wire n_6395;
wire n_3497;
wire n_6403;
wire n_4542;
wire n_5451;
wire n_6578;
wire n_3243;
wire n_4326;
wire n_2121;
wire n_3865;
wire n_6350;
wire n_5460;
wire n_4685;
wire n_3927;
wire n_6141;
wire n_2068;
wire n_3595;
wire n_6875;
wire n_7189;
wire n_4060;
wire n_6194;
wire n_2459;
wire n_3396;
wire n_5517;
wire n_5807;
wire n_5426;
wire n_6475;
wire n_4093;
wire n_5693;
wire n_5695;
wire n_4123;
wire n_4294;
wire n_1940;
wire n_3683;
wire n_6502;
wire n_6944;
wire n_4452;
wire n_3887;
wire n_3195;
wire n_5587;
wire n_4722;
wire n_6318;
wire n_6805;
wire n_3048;
wire n_3339;
wire n_4126;
wire n_4164;
wire n_5030;
wire n_7240;
wire n_2963;
wire n_5674;
wire n_2561;
wire n_5584;
wire n_3168;
wire n_5320;
wire n_4079;
wire n_1749;
wire n_6075;
wire n_6559;
wire n_4088;
wire n_2669;
wire n_3911;
wire n_6068;
wire n_3802;
wire n_4366;
wire n_6248;
wire n_6541;
wire n_5125;
wire n_4922;
wire n_6066;
wire n_6080;
wire n_4733;
wire n_1814;
wire n_7219;
wire n_2441;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_6150;
wire n_6638;
wire n_7063;
wire n_7402;
wire n_6351;
wire n_4935;
wire n_4509;
wire n_2073;
wire n_7382;
wire n_4004;
wire n_5238;
wire n_3630;
wire n_1910;
wire n_5906;
wire n_2189;
wire n_5732;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_2602;
wire n_5780;
wire n_2931;
wire n_3433;
wire n_5556;
wire n_6006;
wire n_3597;
wire n_6474;
wire n_5743;
wire n_6481;
wire n_1956;
wire n_4111;
wire n_5633;
wire n_3786;
wire n_6022;
wire n_6991;
wire n_2828;
wire n_7434;
wire n_5950;
wire n_1715;
wire n_4204;
wire n_3553;
wire n_5323;
wire n_6744;
wire n_3645;
wire n_5705;
wire n_6927;
wire n_7335;
wire n_4996;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_6116;
wire n_3550;
wire n_5510;
wire n_4785;
wire n_2870;
wire n_1893;
wire n_1805;
wire n_4068;
wire n_5440;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_3610;
wire n_2443;
wire n_5011;
wire n_6757;
wire n_3279;
wire n_5513;
wire n_5875;
wire n_4262;
wire n_2923;
wire n_2843;
wire n_3714;
wire n_4832;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_6485;
wire n_5848;
wire n_5834;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_5784;
wire n_3125;
wire n_5128;
wire n_2356;
wire n_5618;
wire n_6495;
wire n_6209;
wire n_4672;
wire n_2564;
wire n_3558;
wire n_3034;
wire n_3502;
wire n_4053;
wire n_7413;
wire n_3963;
wire n_3091;
wire n_6274;
wire n_5157;
wire n_4496;
wire n_2518;
wire n_4596;
wire n_5178;
wire n_3105;
wire n_6237;
wire n_4628;
wire n_6802;
wire n_7343;
wire n_5982;
wire n_1775;
wire n_7109;
wire n_4083;
wire n_2794;
wire n_6155;
wire n_2901;
wire n_3940;
wire n_6809;
wire n_6099;
wire n_3225;
wire n_3621;
wire n_5529;
wire n_3473;
wire n_6349;
wire n_3680;
wire n_6716;
wire n_3565;
wire n_6905;
wire n_5388;
wire n_5824;
wire n_5354;
wire n_2453;
wire n_3331;
wire n_1788;
wire n_6203;
wire n_2138;
wire n_6407;
wire n_3040;
wire n_4230;
wire n_6899;
wire n_6413;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_7070;
wire n_2000;
wire n_5276;
wire n_4037;
wire n_3804;
wire n_4659;
wire n_3211;
wire n_7299;
wire n_5196;
wire n_2440;
wire n_2096;
wire n_2556;
wire n_2215;
wire n_3847;
wire n_6960;
wire n_4073;
wire n_7249;
wire n_5763;
wire n_3633;
wire n_6061;
wire n_2584;
wire n_4001;
wire n_5701;
wire n_7002;
wire n_6273;
wire n_7094;
wire n_7396;
wire n_3111;
wire n_1813;
wire n_2997;
wire n_7018;
wire n_6746;
wire n_3258;
wire n_3691;
wire n_2252;
wire n_6174;
wire n_6545;
wire n_6763;
wire n_1996;
wire n_2009;
wire n_5907;
wire n_4339;
wire n_7297;
wire n_6013;
wire n_6182;
wire n_6754;
wire n_4690;
wire n_2987;
wire n_6279;
wire n_5895;
wire n_2651;
wire n_2445;
wire n_2733;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_3316;
wire n_4023;
wire n_4253;
wire n_3632;
wire n_2522;
wire n_4064;
wire n_6131;
wire n_3351;
wire n_5478;
wire n_6113;
wire n_3457;
wire n_5384;
wire n_6477;
wire n_2324;
wire n_6575;
wire n_5283;
wire n_3454;
wire n_5961;
wire n_2139;
wire n_2521;
wire n_5686;
wire n_6391;
wire n_2740;
wire n_1991;
wire n_7140;
wire n_4066;
wire n_6252;
wire n_6426;
wire n_4681;
wire n_3303;
wire n_6592;
wire n_4414;
wire n_2541;
wire n_5094;
wire n_3232;
wire n_3768;
wire n_4295;
wire n_4100;
wire n_6668;
wire n_2372;
wire n_2105;
wire n_3445;
wire n_1806;
wire n_4087;
wire n_4473;
wire n_4619;
wire n_6670;
wire n_5371;
wire n_2290;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_5350;
wire n_3265;
wire n_3018;
wire n_1875;
wire n_6962;
wire n_2429;
wire n_6779;
wire n_5286;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_5676;
wire n_5949;
wire n_5040;
wire n_6901;
wire n_4266;
wire n_6336;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_6503;
wire n_6049;
wire n_5885;
wire n_3628;
wire n_7100;
wire n_4777;
wire n_7243;
wire n_5243;
wire n_3941;
wire n_1915;
wire n_7415;
wire n_5399;
wire n_2846;
wire n_3371;
wire n_4918;
wire n_5856;
wire n_3872;
wire n_5760;
wire n_4415;
wire n_5110;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_1777;
wire n_3366;
wire n_6998;
wire n_7395;
wire n_5844;
wire n_6298;
wire n_3441;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_6609;
wire n_2545;
wire n_2513;
wire n_4408;
wire n_2115;
wire n_2017;
wire n_1810;
wire n_4976;
wire n_6525;
wire n_3555;
wire n_5938;
wire n_7274;
wire n_3534;
wire n_4548;
wire n_2670;
wire n_6494;
wire n_3556;
wire n_4574;
wire n_2644;
wire n_6132;
wire n_4557;
wire n_3071;
wire n_2148;
wire n_5548;
wire n_6974;
wire n_4663;
wire n_5840;
wire n_6882;
wire n_3296;
wire n_3762;
wire n_3794;
wire n_4624;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_6498;
wire n_6562;
wire n_3293;
wire n_4902;
wire n_4686;
wire n_2384;
wire n_3707;
wire n_3895;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_5917;
wire n_6965;
wire n_2058;
wire n_3231;
wire n_1846;
wire n_4161;
wire n_6168;
wire n_5304;
wire n_5437;
wire n_6963;
wire n_6951;
wire n_3058;
wire n_5355;
wire n_2047;
wire n_3398;
wire n_3709;
wire n_6284;
wire n_3592;
wire n_5321;
wire n_7454;
wire n_2536;
wire n_3399;
wire n_4772;
wire n_6931;
wire n_6521;
wire n_5915;
wire n_7276;
wire n_6379;
wire n_7085;
wire n_6306;
wire n_4120;
wire n_6834;
wire n_2880;
wire n_4716;
wire n_3722;
wire n_4654;
wire n_5116;
wire n_3771;
wire n_7225;
wire n_3158;
wire n_3221;
wire n_2316;
wire n_2830;
wire n_5500;
wire n_4622;
wire n_4757;
wire n_1871;
wire n_6471;
wire n_6949;
wire n_5669;
wire n_5672;
wire n_4016;
wire n_3334;
wire n_5621;
wire n_6760;
wire n_2940;
wire n_3427;
wire n_3162;
wire n_5569;
wire n_4591;
wire n_5966;
wire n_5515;
wire n_6589;
wire n_3083;
wire n_4570;
wire n_7014;
wire n_2491;
wire n_1931;
wire n_5559;
wire n_2259;
wire n_5337;
wire n_5059;
wire n_4655;
wire n_7459;
wire n_1820;
wire n_7160;
wire n_7324;
wire n_6046;
wire n_7054;
wire n_4493;
wire n_6055;
wire n_7161;
wire n_1808;
wire n_6364;
wire n_6091;
wire n_6348;
wire n_4896;
wire n_4851;
wire n_6848;
wire n_2479;
wire n_6788;
wire n_6144;
wire n_5528;
wire n_5605;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_6896;
wire n_2484;
wire n_5753;
wire n_5358;
wire n_4901;
wire n_3480;
wire n_7201;
wire n_4213;
wire n_4127;
wire n_6221;
wire n_2500;
wire n_2334;
wire n_5467;
wire n_7241;
wire n_3181;
wire n_5493;
wire n_1916;
wire n_6285;
wire n_4602;
wire n_1713;
wire n_2818;
wire n_4900;
wire n_3578;
wire n_2537;
wire n_3745;
wire n_6748;
wire n_7430;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_5901;
wire n_2837;
wire n_2446;
wire n_6582;
wire n_4116;
wire n_5360;
wire n_7269;
wire n_7047;
wire n_2671;
wire n_2702;
wire n_6937;
wire n_4363;
wire n_3561;
wire n_1839;
wire n_4103;
wire n_2529;
wire n_2374;
wire n_5439;
wire n_6115;
wire n_3154;
wire n_3938;
wire n_2278;
wire n_6272;
wire n_7067;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_5250;
wire n_4416;
wire n_6607;
wire n_4439;
wire n_4985;
wire n_3382;
wire n_7117;
wire n_3930;
wire n_3808;
wire n_5471;
wire n_2248;
wire n_4660;
wire n_3081;
wire n_6446;
wire n_5497;
wire n_5519;
wire n_6071;
wire n_2579;
wire n_1961;
wire n_6849;
wire n_2960;
wire n_3270;
wire n_6807;
wire n_2844;
wire n_1979;
wire n_6616;
wire n_6719;
wire n_4814;
wire n_6178;
wire n_6677;
wire n_2221;
wire n_5502;
wire n_2317;
wire n_2838;
wire n_1736;
wire n_2200;
wire n_7302;
wire n_2781;
wire n_6191;
wire n_2442;
wire n_7238;
wire n_6862;
wire n_3657;
wire n_5706;
wire n_2634;
wire n_2746;
wire n_7292;
wire n_5098;
wire n_6000;
wire n_6774;
wire n_6443;
wire n_5145;
wire n_6072;
wire n_2878;
wire n_7248;
wire n_3830;
wire n_3252;
wire n_6647;
wire n_5466;
wire n_6941;
wire n_7239;
wire n_6552;
wire n_3315;
wire n_6094;
wire n_3523;
wire n_3999;
wire n_7112;
wire n_3420;
wire n_3859;
wire n_5213;
wire n_3474;
wire n_5738;
wire n_2458;
wire n_5592;
wire n_5620;
wire n_3150;
wire n_5491;
wire n_4831;
wire n_4782;
wire n_2859;
wire n_5216;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_5953;
wire n_5703;
wire n_6886;
wire n_7078;
wire n_4597;
wire n_4546;
wire n_5187;
wire n_7006;
wire n_4031;
wire n_5119;
wire n_4147;
wire n_3073;
wire n_6531;
wire n_3571;
wire n_4576;
wire n_7354;
wire n_6098;
wire n_5995;
wire n_3297;
wire n_5148;
wire n_3003;
wire n_6726;
wire n_6983;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_5330;
wire n_6935;
wire n_2899;
wire n_6984;
wire n_6778;
wire n_6897;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5526;
wire n_5202;
wire n_3817;
wire n_6345;
wire n_6386;
wire n_3728;
wire n_2722;
wire n_6596;
wire n_5107;
wire n_7165;
wire n_4680;
wire n_5067;
wire n_6830;
wire n_2685;
wire n_2061;
wire n_5987;
wire n_2512;
wire n_1790;
wire n_2788;
wire n_6642;
wire n_6291;
wire n_6510;
wire n_5264;
wire n_2595;
wire n_3084;
wire n_6781;
wire n_4593;
wire n_7123;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_3554;
wire n_6509;
wire n_2717;
wire n_6376;
wire n_2981;
wire n_4995;
wire n_5873;
wire n_6514;
wire n_4498;
wire n_6741;
wire n_6434;
wire n_5741;
wire n_2743;
wire n_2969;
wire n_3429;
wire n_2466;
wire n_6593;
wire n_3758;
wire n_6690;
wire n_5423;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_4109;
wire n_1935;
wire n_3777;
wire n_1872;
wire n_3767;
wire n_6056;
wire n_5926;
wire n_5866;
wire n_3692;
wire n_3234;
wire n_2216;
wire n_2426;
wire n_6947;
wire n_4850;
wire n_3716;
wire n_7157;
wire n_2926;
wire n_4937;
wire n_5574;
wire n_3391;
wire n_5877;
wire n_6375;
wire n_4786;
wire n_6042;
wire n_5203;
wire n_7091;
wire n_4354;
wire n_6429;
wire n_4235;
wire n_3159;
wire n_6315;
wire n_2855;
wire n_2848;
wire n_6775;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_6970;
wire n_6948;
wire n_3460;
wire n_5155;
wire n_2202;
wire n_2952;
wire n_3530;
wire n_6133;
wire n_6920;
wire n_2693;
wire n_7409;
wire n_5408;
wire n_5812;
wire n_5540;
wire n_7381;
wire n_5804;
wire n_3240;
wire n_5066;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_7087;
wire n_5130;
wire n_4175;
wire n_6241;
wire n_5200;
wire n_3393;
wire n_2836;
wire n_2864;
wire n_4456;
wire n_1717;
wire n_5992;
wire n_2172;
wire n_2601;
wire n_2365;
wire n_1880;
wire n_5684;
wire n_7228;
wire n_5981;
wire n_1855;
wire n_6632;
wire n_2333;
wire n_3629;
wire n_4948;
wire n_5413;
wire n_1903;
wire n_2147;
wire n_6623;
wire n_4020;
wire n_5111;
wire n_5150;
wire n_2224;
wire n_6933;
wire n_1970;
wire n_3724;
wire n_3287;
wire n_2167;
wire n_3046;
wire n_2293;
wire n_2921;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_5444;
wire n_3257;
wire n_5737;
wire n_3730;
wire n_5615;
wire n_3979;
wire n_6908;
wire n_5097;
wire n_2695;
wire n_7084;
wire n_2598;
wire n_3727;
wire n_6083;
wire n_6537;
wire n_4003;
wire n_1832;
wire n_6390;
wire n_2302;
wire n_6799;
wire n_3014;
wire n_2294;
wire n_6278;
wire n_2274;
wire n_7195;
wire n_5640;
wire n_3342;
wire n_2895;
wire n_6101;
wire n_7298;
wire n_3796;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_5550;
wire n_3375;
wire n_2768;
wire n_3760;
wire n_5661;
wire n_4975;
wire n_3515;
wire n_2363;
wire n_5306;
wire n_5905;
wire n_6112;
wire n_2728;
wire n_2025;
wire n_3744;
wire n_5457;
wire n_5159;
wire n_4022;
wire n_7115;
wire n_2495;
wire n_4336;
wire n_5314;
wire n_5231;
wire n_5064;
wire n_2223;
wire n_6412;
wire n_6271;
wire n_7235;
wire n_2511;
wire n_6572;
wire n_3981;
wire n_7271;
wire n_2681;
wire n_7222;
wire n_2535;
wire n_3031;
wire n_6930;
wire n_2335;
wire n_5482;
wire n_3215;
wire n_3138;
wire n_2860;
wire n_2041;
wire n_1933;
wire n_6584;
wire n_4494;
wire n_6387;
wire n_4201;
wire n_6470;
wire n_7206;
wire n_5287;
wire n_4719;
wire n_5651;
wire n_3577;
wire n_6625;
wire n_4074;
wire n_7383;
wire n_3994;
wire n_4636;
wire n_4983;
wire n_3185;
wire n_6826;
wire n_2662;
wire n_4386;
wire n_6341;
wire n_6374;
wire n_3917;
wire n_5623;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_5524;
wire n_2296;
wire n_5735;
wire n_6363;
wire n_6588;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_4225;
wire n_6811;
wire n_6687;
wire n_4658;
wire n_7135;
wire n_6037;
wire n_4186;
wire n_2241;
wire n_6865;
wire n_7211;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_2531;
wire n_7132;
wire n_3377;
wire n_6722;
wire n_6420;
wire n_4907;
wire n_3961;
wire n_5153;
wire n_2059;
wire n_4713;
wire n_5787;
wire n_6911;
wire n_7129;
wire n_7080;
wire n_3374;
wire n_4870;
wire n_6981;
wire n_4818;
wire n_7436;
wire n_7020;
wire n_5935;
wire n_6696;
wire n_4916;
wire n_5967;
wire n_6095;
wire n_4323;
wire n_6045;
wire n_1899;
wire n_5934;
wire n_5376;
wire n_3508;
wire n_6300;
wire n_6653;
wire n_6372;
wire n_4129;
wire n_7120;
wire n_5488;
wire n_6900;
wire n_5727;
wire n_3599;
wire n_6660;
wire n_5988;
wire n_6424;
wire n_5646;
wire n_7448;
wire n_4480;
wire n_5711;
wire n_3734;
wire n_6787;
wire n_5832;
wire n_6254;
wire n_7460;
wire n_3401;
wire n_7142;
wire n_6423;
wire n_6526;
wire n_3542;
wire n_3263;
wire n_5891;
wire n_2523;
wire n_1945;
wire n_2418;
wire n_5328;
wire n_3819;
wire n_3222;
wire n_1740;
wire n_4616;
wire n_5016;
wire n_6011;
wire n_7465;
wire n_5470;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_6176;
wire n_1963;
wire n_3868;
wire n_6222;
wire n_2218;
wire n_2593;
wire n_6969;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_6587;
wire n_6688;
wire n_6505;
wire n_5362;
wire n_2754;
wire n_4580;
wire n_6762;
wire n_3611;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_6987;
wire n_3995;
wire n_3908;
wire n_6453;
wire n_6308;
wire n_3892;
wire n_7449;
wire n_3501;
wire n_3216;
wire n_3568;
wire n_2555;
wire n_2708;
wire n_6187;
wire n_6597;
wire n_4844;
wire n_6220;
wire n_4049;
wire n_2661;
wire n_2470;
wire n_3551;
wire n_5037;
wire n_7305;
wire n_5650;
wire n_5729;
wire n_5581;
wire n_4677;
wire n_5189;
wire n_4525;
wire n_6149;
wire n_3364;
wire n_2643;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_4369;
wire n_3826;
wire n_5648;
wire n_2266;
wire n_6439;
wire n_4324;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_6547;
wire n_7177;
wire n_5160;
wire n_1719;
wire n_2742;
wire n_3671;
wire n_2366;
wire n_5762;
wire n_1753;
wire n_5484;
wire n_1895;
wire n_7353;
wire n_4104;
wire n_3791;
wire n_6478;
wire n_2008;
wire n_4989;
wire n_5874;
wire n_3064;
wire n_3199;
wire n_2127;
wire n_7050;
wire n_3151;
wire n_6906;
wire n_3016;
wire n_2460;
wire n_6739;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_4528;
wire n_2772;
wire n_5385;
wire n_1747;
wire n_3990;
wire n_5622;
wire n_5635;
wire n_4069;
wire n_3582;
wire n_4280;
wire n_1867;
wire n_6034;
wire n_5609;
wire n_3993;
wire n_3459;
wire n_2576;
wire n_4811;
wire n_2696;
wire n_5595;
wire n_5256;
wire n_4779;
wire n_5910;
wire n_2140;
wire n_2157;
wire n_1966;
wire n_5380;
wire n_3735;
wire n_7410;
wire n_6422;
wire n_3656;
wire n_4524;
wire n_2831;
wire n_3069;
wire n_4657;
wire n_5568;
wire n_5941;
wire n_4891;
wire n_2629;
wire n_3369;
wire n_1954;
wire n_6604;
wire n_3964;
wire n_6611;
wire n_5364;
wire n_3302;
wire n_5597;
wire n_2486;
wire n_1897;
wire n_6999;
wire n_5469;
wire n_2137;
wire n_3685;
wire n_6019;
wire n_6440;
wire n_4977;
wire n_2492;
wire n_6976;
wire n_7234;
wire n_2939;
wire n_3425;
wire n_4876;
wire n_5021;
wire n_2900;
wire n_2912;
wire n_5936;
wire n_3813;
wire n_5312;
wire n_2622;
wire n_3447;
wire n_6784;
wire n_1757;
wire n_1950;
wire n_2264;
wire n_5928;
wire n_2032;
wire n_2090;
wire n_3124;
wire n_3811;
wire n_4200;
wire n_2249;
wire n_5785;
wire n_3411;
wire n_5222;
wire n_6165;
wire n_3463;
wire n_2785;
wire n_4938;
wire n_2574;
wire n_2364;
wire n_6114;
wire n_1856;
wire n_2928;
wire n_5505;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_5504;
wire n_7348;
wire n_4118;
wire n_6829;
wire n_3857;
wire n_3110;
wire n_4239;
wire n_3157;
wire n_2730;
wire n_6464;
wire n_5129;
wire n_7320;
wire n_4704;
wire n_2720;
wire n_5494;
wire n_5970;
wire n_2405;
wire n_6838;
wire n_2700;
wire n_6368;
wire n_2416;
wire n_2064;
wire n_3640;
wire n_5663;
wire n_5161;
wire n_6640;
wire n_7155;
wire n_6166;
wire n_4744;
wire n_5378;
wire n_5626;
wire n_4706;
wire n_3879;
wire n_2022;
wire n_4343;
wire n_6850;
wire n_2408;
wire n_4764;
wire n_5389;
wire n_4990;
wire n_2986;
wire n_2454;
wire n_6550;
wire n_6656;
wire n_6972;
wire n_3591;
wire n_2760;
wire n_4919;
wire n_7043;
wire n_3317;
wire n_7266;
wire n_5653;
wire n_4835;
wire n_4420;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_5266;
wire n_4559;
wire n_4742;
wire n_5038;
wire n_3566;
wire n_5800;
wire n_4372;
wire n_5396;
wire n_4097;
wire n_4162;
wire n_5766;
wire n_5293;
wire n_4790;
wire n_7035;
wire n_4173;
wire n_5309;
wire n_6047;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_7442;
wire n_4727;
wire n_6568;
wire n_3654;
wire n_5627;
wire n_3783;
wire n_4008;
wire n_2158;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_7153;
wire n_6258;
wire n_2173;
wire n_3982;
wire n_7350;
wire n_3647;
wire n_7314;
wire n_6026;
wire n_3973;
wire n_4799;
wire n_5882;
wire n_6700;
wire n_7136;
wire n_4534;
wire n_5636;
wire n_4960;
wire n_5707;
wire n_5594;
wire n_3738;
wire n_5697;
wire n_2020;
wire n_5606;
wire n_6727;
wire n_2310;
wire n_5911;
wire n_7340;
wire n_3600;
wire n_7303;
wire n_6139;
wire n_7399;
wire n_5382;
wire n_4327;
wire n_7387;
wire n_3190;
wire n_3027;
wire n_6454;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_3733;
wire n_3967;
wire n_6333;
wire n_7004;
wire n_4370;
wire n_5638;
wire n_4816;
wire n_4091;
wire n_5058;
wire n_3096;
wire n_7207;
wire n_4166;
wire n_2777;
wire n_5356;
wire n_7167;
wire n_2234;
wire n_5849;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_5841;
wire n_7146;
wire n_7030;
wire n_4478;
wire n_2935;
wire n_4246;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_4061;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_4754;
wire n_4375;
wire n_2396;
wire n_3368;
wire n_3117;
wire n_4684;
wire n_3384;
wire n_5279;
wire n_7159;
wire n_2592;
wire n_3490;
wire n_7280;
wire n_5043;
wire n_7339;
wire n_4241;
wire n_3113;
wire n_2751;
wire n_4183;
wire n_1968;
wire n_5645;
wire n_5020;
wire n_6455;
wire n_2842;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_3720;
wire n_6183;
wire n_6107;
wire n_6476;
wire n_5232;
wire n_2560;
wire n_4256;
wire n_5035;
wire n_3037;
wire n_5453;
wire n_4333;
wire n_5339;
wire n_6003;
wire n_5443;
wire n_2007;
wire n_3363;
wire n_6636;
wire n_1803;
wire n_3522;
wire n_4455;
wire n_3241;
wire n_3899;
wire n_6554;
wire n_5631;
wire n_3481;
wire n_6994;
wire n_7401;
wire n_5101;
wire n_6020;
wire n_2236;
wire n_6185;
wire n_7321;
wire n_4457;
wire n_2150;
wire n_6785;
wire n_1816;
wire n_2803;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_6870;
wire n_3305;
wire n_6643;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_6695;
wire n_3354;
wire n_5608;
wire n_6501;
wire n_2204;
wire n_2040;
wire n_6466;
wire n_2151;
wire n_2455;
wire n_3437;
wire n_6467;
wire n_2231;
wire n_4212;
wire n_4584;
wire n_7188;
wire n_5702;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_2406;
wire n_4477;
wire n_5806;
wire n_4110;
wire n_5182;
wire n_4217;
wire n_5277;
wire n_6507;
wire n_1942;
wire n_6618;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_6213;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_3969;
wire n_6873;
wire n_2282;
wire n_4605;
wire n_3873;
wire n_4649;
wire n_5747;
wire n_7101;
wire n_2428;
wire n_6063;
wire n_2858;
wire n_3076;
wire n_3410;
wire n_5415;
wire n_7261;
wire n_4592;
wire n_4999;
wire n_6993;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_1858;
wire n_2589;
wire n_4086;
wire n_6767;
wire n_4656;
wire n_4862;
wire n_5687;
wire n_6558;
wire n_6755;
wire n_6153;
wire n_3536;
wire n_1721;
wire n_7263;
wire n_3782;
wire n_6608;
wire n_6202;
wire n_6780;
wire n_3594;
wire n_5383;
wire n_2385;
wire n_6635;
wire n_7245;
wire n_7310;
wire n_6359;
wire n_5690;
wire n_1980;
wire n_5740;
wire n_7093;
wire n_4177;
wire n_2501;
wire n_1998;
wire n_5029;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_3855;
wire n_7418;
wire n_6353;
wire n_2985;
wire n_5218;
wire n_2630;
wire n_6577;
wire n_2028;
wire n_3114;
wire n_2092;
wire n_6082;
wire n_3622;
wire n_2817;
wire n_2773;
wire n_2402;
wire n_3047;
wire n_3163;
wire n_5361;
wire n_7312;
wire n_6105;
wire n_5512;
wire n_2808;
wire n_2344;
wire n_3520;
wire n_2392;
wire n_3272;
wire n_3122;
wire n_5898;
wire n_7113;
wire n_6548;
wire n_5923;
wire n_3687;
wire n_2787;
wire n_6657;
wire n_5617;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_5946;
wire n_2676;
wire n_7282;
wire n_2770;
wire n_4550;
wire n_4347;
wire n_5193;
wire n_4933;
wire n_4144;
wire n_5514;
wire n_5611;
wire n_3278;
wire n_2375;
wire n_5579;
wire n_4167;
wire n_6380;
wire n_3608;
wire n_4895;
wire n_6163;
wire n_7170;
wire n_4726;
wire n_5573;
wire n_5143;
wire n_5836;
wire n_1755;
wire n_5188;
wire n_6674;
wire n_5049;
wire n_2212;
wire n_6331;
wire n_5308;
wire n_4434;
wire n_5068;
wire n_6493;
wire n_7363;
wire n_7281;
wire n_5739;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_6023;
wire n_3829;
wire n_4510;
wire n_5057;
wire n_6196;
wire n_5425;
wire n_5273;
wire n_5839;
wire n_2469;
wire n_2358;
wire n_1710;
wire n_3546;
wire n_2355;
wire n_5887;
wire n_3068;
wire n_6321;
wire n_5683;
wire n_3002;
wire n_7192;
wire n_5248;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_4156;
wire n_1727;
wire n_3693;
wire n_5880;
wire n_3132;
wire n_5002;
wire n_5487;
wire n_5649;
wire n_5531;
wire n_3681;
wire n_5666;
wire n_3970;
wire n_2351;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_6824;
wire n_6954;
wire n_6450;
wire n_6995;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_4579;
wire n_6347;
wire n_6496;
wire n_4776;
wire n_2704;
wire n_6745;
wire n_3729;
wire n_6698;
wire n_4471;
wire n_6968;
wire n_7377;
wire n_4392;
wire n_3103;
wire n_6064;
wire n_2048;
wire n_3028;
wire n_4691;
wire n_3148;
wire n_3775;
wire n_5682;
wire n_5461;
wire n_7296;
wire n_3966;
wire n_4397;
wire n_6164;
wire n_3616;
wire n_4753;
wire n_4803;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_5730;
wire n_6292;
wire n_6743;
wire n_4165;
wire n_2056;
wire n_5754;
wire n_2852;
wire n_2515;
wire n_6330;
wire n_7178;
wire n_1941;
wire n_7045;
wire n_3637;
wire n_4893;
wire n_2240;
wire n_4258;
wire n_5756;
wire n_2917;
wire n_3194;
wire n_2432;
wire n_2085;
wire n_5033;
wire n_6015;
wire n_6408;
wire n_4232;
wire n_5075;
wire n_2097;
wire n_3461;
wire n_7300;
wire n_2297;
wire n_6861;
wire n_4203;
wire n_5789;
wire n_5400;
wire n_5347;
wire n_2957;
wire n_1983;
wire n_4767;
wire n_4569;
wire n_6528;
wire n_3820;
wire n_5144;
wire n_6895;
wire n_3072;
wire n_2961;
wire n_4468;
wire n_5509;
wire n_1923;
wire n_3848;
wire n_7400;
wire n_3631;
wire n_7393;
wire n_6590;
wire n_6523;
wire n_5169;
wire n_4885;
wire n_4698;
wire n_3674;
wire n_5349;
wire n_6472;
wire n_3763;
wire n_6389;
wire n_3499;
wire n_5534;
wire n_1821;
wire n_3910;
wire n_3947;
wire n_5183;
wire n_2585;
wire n_3361;
wire n_2995;
wire n_6073;
wire n_4533;
wire n_4287;
wire n_3228;
wire n_2164;
wire n_1732;
wire n_2678;
wire n_6869;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_4556;
wire n_6137;
wire n_2205;
wire n_2183;
wire n_1724;
wire n_3088;
wire n_2080;
wire n_5254;
wire n_3590;
wire n_5079;
wire n_2761;
wire n_2357;
wire n_4520;
wire n_2421;
wire n_3295;
wire n_5751;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_6885;
wire n_5039;
wire n_1818;
wire n_6580;
wire n_6613;
wire n_4265;
wire n_6404;
wire n_6120;
wire n_3557;
wire n_2269;
wire n_4612;
wire n_5997;
wire n_5375;
wire n_5438;
wire n_7150;
wire n_6530;
wire n_6602;
wire n_4149;
wire n_1827;
wire n_4958;
wire n_6135;
wire n_1752;
wire n_2361;
wire n_4538;
wire n_3030;
wire n_3505;
wire n_5563;
wire n_3075;
wire n_2239;
wire n_6942;
wire n_6892;
wire n_4730;
wire n_7357;
wire n_6782;
wire n_4421;
wire n_6230;
wire n_2464;
wire n_3697;
wire n_2304;
wire n_2514;
wire n_6977;
wire n_7229;
wire n_7336;
wire n_5932;
wire n_6598;
wire n_6795;
wire n_6121;
wire n_3430;
wire n_5919;
wire n_2063;
wire n_3489;
wire n_5012;
wire n_6614;
wire n_6506;
wire n_2079;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_3484;
wire n_6001;
wire n_4971;
wire n_2095;
wire n_5664;
wire n_2738;
wire n_6406;
wire n_5890;
wire n_2590;
wire n_4661;
wire n_2797;
wire n_3041;
wire n_5823;
wire n_2208;
wire n_2423;
wire n_5422;
wire n_5944;
wire n_6989;
wire n_6299;
wire n_7424;
wire n_5246;
wire n_4376;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_4305;
wire n_2037;
wire n_2953;
wire n_2823;
wire n_7273;
wire n_3684;
wire n_5725;
wire n_5404;
wire n_4834;
wire n_5332;
wire n_7149;
wire n_2866;
wire n_7116;
wire n_3153;
wire n_2346;
wire n_4692;
wire n_3268;
wire n_2559;
wire n_5616;
wire n_4259;
wire n_5870;
wire n_2030;
wire n_6053;
wire n_6233;
wire n_4299;
wire n_5625;
wire n_6758;
wire n_2407;
wire n_5367;
wire n_2243;
wire n_6629;
wire n_5288;
wire n_2694;
wire n_6356;
wire n_5601;
wire n_3742;
wire n_4965;
wire n_1837;
wire n_7033;
wire n_4178;
wire n_6010;
wire n_2006;
wire n_4953;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_7147;
wire n_5294;
wire n_5570;
wire n_6411;
wire n_2731;
wire n_3703;
wire n_5411;
wire n_5670;
wire n_5265;
wire n_5955;
wire n_2123;
wire n_2238;
wire n_4802;
wire n_4793;
wire n_6032;
wire n_5733;
wire n_3435;
wire n_2380;
wire n_4897;
wire n_6918;
wire n_1745;
wire n_4674;
wire n_4796;
wire n_7138;
wire n_6401;
wire n_7279;
wire n_5184;
wire n_2750;
wire n_2547;
wire n_4575;
wire n_3665;
wire n_3063;
wire n_3281;
wire n_7137;
wire n_3535;
wire n_5061;
wire n_2288;
wire n_3858;
wire n_4653;
wire n_4589;
wire n_7124;
wire n_5978;
wire n_6853;
wire n_3220;
wire n_4581;
wire n_6008;
wire n_4625;
wire n_7098;
wire n_6181;
wire n_2107;
wire n_5070;
wire n_4845;
wire n_4148;
wire n_3679;
wire n_5575;
wire n_6654;
wire n_4968;
wire n_6907;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_4038;
wire n_3856;
wire n_5316;
wire n_2735;
wire n_4214;
wire n_1888;
wire n_5290;
wire n_2109;
wire n_2709;
wire n_3419;
wire n_7323;
wire n_5048;
wire n_2233;
wire n_5363;
wire n_5665;
wire n_6517;
wire n_4892;
wire n_6339;
wire n_1936;
wire n_3890;
wire n_6170;
wire n_7247;
wire n_6394;
wire n_5607;
wire n_2782;
wire n_3929;
wire n_4353;
wire n_2201;
wire n_4950;
wire n_6504;
wire n_4176;
wire n_4124;
wire n_4431;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_5462;
wire n_6814;
wire n_7216;
wire n_4488;
wire n_5278;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_5214;
wire n_3756;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_5845;
wire n_4608;
wire n_6691;
wire n_3948;
wire n_4839;
wire n_5969;
wire n_1765;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_2332;
wire n_2391;
wire n_6343;
wire n_6005;
wire n_2060;
wire n_3883;
wire n_6686;
wire n_4032;
wire n_2571;
wire n_6437;
wire n_5736;
wire n_4929;
wire n_2874;
wire n_6029;
wire n_6536;
wire n_6684;
wire n_4117;
wire n_6025;
wire n_3049;
wire n_3634;
wire n_5436;
wire n_2341;
wire n_6697;
wire n_3066;
wire n_2045;
wire n_6085;
wire n_3913;
wire n_5341;
wire n_2575;
wire n_3739;
wire n_5140;
wire n_2942;
wire n_6062;
wire n_1771;
wire n_4541;
wire n_6715;
wire n_3271;
wire n_3164;
wire n_3861;
wire n_5096;
wire n_2043;
wire n_6771;
wire n_4171;
wire n_5847;
wire n_7204;
wire n_7022;
wire n_6383;
wire n_4815;
wire n_4665;
wire n_5639;
wire n_6877;
wire n_7308;
wire n_4884;
wire n_3580;
wire n_4276;
wire n_5268;
wire n_5050;
wire n_5240;
wire n_5503;
wire n_5718;
wire n_7208;
wire n_1876;
wire n_1830;
wire n_5001;
wire n_6567;
wire n_5658;
wire n_4174;
wire n_6868;
wire n_7290;
wire n_5131;
wire n_6813;
wire n_5546;
wire n_6294;
wire n_5174;
wire n_2145;
wire n_4801;
wire n_6079;
wire n_6260;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_5289;
wire n_6520;
wire n_3119;
wire n_6671;
wire n_4740;
wire n_4394;
wire n_5544;
wire n_6444;
wire n_6637;
wire n_6729;
wire n_5660;
wire n_6958;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_5541;
wire n_6314;
wire n_5610;
wire n_2810;
wire n_6703;
wire n_1884;
wire n_4378;
wire n_5166;
wire n_2683;
wire n_6065;
wire n_7265;
wire n_4180;
wire n_4459;
wire n_6878;
wire n_3624;
wire n_6725;
wire n_5808;
wire n_6527;
wire n_4594;
wire n_7289;
wire n_2748;
wire n_4642;
wire n_6913;
wire n_7242;
wire n_6533;
wire n_7164;
wire n_2925;
wire n_1750;
wire n_3544;
wire n_6845;
wire n_5300;
wire n_2072;
wire n_3852;
wire n_5233;
wire n_5381;
wire n_5770;
wire n_5710;
wire n_2628;
wire n_7389;
wire n_3219;
wire n_5333;
wire n_5799;
wire n_6265;
wire n_4914;
wire n_3510;
wire n_7046;
wire n_4587;
wire n_3688;
wire n_5008;
wire n_3871;
wire n_3757;
wire n_2219;
wire n_6148;
wire n_2100;
wire n_3666;
wire n_5538;
wire n_6357;
wire n_3479;
wire n_5499;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_6522;
wire n_4285;
wire n_7097;
wire n_7000;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_3741;
wire n_5582;
wire n_2567;
wire n_2557;
wire n_1908;
wire n_5675;
wire n_2755;
wire n_5109;
wire n_6713;
wire n_2066;
wire n_5281;
wire n_2762;
wire n_6087;
wire n_2220;
wire n_7342;
wire n_7044;
wire n_6108;
wire n_6100;
wire n_6800;
wire n_7364;
wire n_6866;
wire n_7114;
wire n_6373;
wire n_4433;
wire n_2829;
wire n_7332;
wire n_5862;
wire n_1914;
wire n_2253;
wire n_5886;
wire n_6415;
wire n_6783;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_5285;
wire n_2328;
wire n_2434;
wire n_3936;
wire n_5564;
wire n_2261;
wire n_3082;
wire n_5162;
wire n_5442;
wire n_2473;
wire n_5802;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_6340;
wire n_3867;
wire n_3397;
wire n_6103;
wire n_6392;
wire n_6513;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_6720;
wire n_5883;
wire n_3078;
wire n_6078;
wire n_3971;
wire n_5630;
wire n_6666;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_2113;
wire n_6815;
wire n_6207;
wire n_6381;
wire n_3711;
wire n_5054;
wire n_6571;
wire n_3171;
wire n_5929;
wire n_5394;
wire n_4751;
wire n_4242;
wire n_5975;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_2812;
wire n_3300;
wire n_7061;
wire n_7066;
wire n_5496;
wire n_3104;
wire n_7174;
wire n_4122;
wire n_6661;
wire n_2132;
wire n_4522;
wire n_5991;
wire n_4952;
wire n_6967;
wire n_4426;
wire n_5956;
wire n_5699;
wire n_4362;
wire n_3267;
wire n_6017;
wire n_3946;
wire n_5920;
wire n_2112;
wire n_2640;
wire n_6125;
wire n_5000;
wire n_4634;
wire n_4932;
wire n_1795;
wire n_2237;
wire n_2983;
wire n_5211;
wire n_4089;
wire n_3513;
wire n_3498;
wire n_5132;
wire n_2350;
wire n_6414;
wire n_5535;
wire n_4506;
wire n_6097;
wire n_6057;
wire n_6936;
wire n_4728;
wire n_7171;
wire n_1886;
wire n_4346;
wire n_7003;
wire n_2187;
wire n_2481;
wire n_3863;
wire n_6302;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_6922;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_3332;
wire n_6432;
wire n_2055;
wire n_2998;
wire n_7366;
wire n_4359;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_4447;
wire n_2937;
wire n_4293;
wire n_6880;
wire n_5176;
wire n_6223;
wire n_4039;
wire n_5793;
wire n_6926;
wire n_1798;
wire n_3057;
wire n_5761;
wire n_6699;
wire n_3983;
wire n_3318;
wire n_7232;
wire n_3385;
wire n_3773;
wire n_3494;
wire n_6957;
wire n_5074;
wire n_3939;
wire n_3788;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_6694;
wire n_3260;
wire n_2496;
wire n_3349;
wire n_6449;
wire n_4348;
wire n_7422;
wire n_3139;
wire n_3801;
wire n_5681;
wire n_2338;
wire n_5261;
wire n_3636;
wire n_6591;
wire n_7466;
wire n_3653;
wire n_3823;
wire n_3403;
wire n_2057;
wire n_6594;
wire n_6342;
wire n_6195;
wire n_2716;
wire n_6441;
wire n_7158;
wire n_2944;
wire n_3439;
wire n_2780;
wire n_4084;
wire n_4240;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_2774;
wire n_6354;
wire n_2799;
wire n_5748;
wire n_4393;
wire n_6662;
wire n_3984;
wire n_4389;
wire n_6433;
wire n_1763;
wire n_6200;
wire n_5641;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_1859;
wire n_3426;
wire n_2660;
wire n_6902;
wire n_4615;
wire n_3044;
wire n_3492;
wire n_7197;
wire n_3737;
wire n_6369;
wire n_5657;
wire n_3579;
wire n_2379;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_5244;
wire n_5765;
wire n_5114;
wire n_4551;
wire n_4521;
wire n_6956;
wire n_2284;
wire n_6451;
wire n_3005;
wire n_5420;
wire n_6497;
wire n_2283;
wire n_5206;
wire n_2526;
wire n_1711;
wire n_4387;
wire n_3186;
wire n_2508;
wire n_6701;
wire n_2594;
wire n_5298;
wire n_3417;
wire n_3626;
wire n_4598;
wire n_4464;
wire n_5106;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_2119;
wire n_2493;
wire n_5080;
wire n_4565;
wire n_7032;
wire n_3392;
wire n_1800;
wire n_7198;
wire n_6884;
wire n_5081;
wire n_6921;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_6106;
wire n_6876;
wire n_3512;
wire n_1860;
wire n_1734;
wire n_4552;
wire n_7193;
wire n_6287;
wire n_2840;
wire n_6172;
wire n_4482;
wire n_5957;
wire n_4172;
wire n_4040;
wire n_3024;
wire n_5567;
wire n_5406;
wire n_6362;
wire n_4328;
wire n_1854;
wire n_5191;
wire n_1729;
wire n_6067;
wire n_2893;
wire n_6833;
wire n_4940;
wire n_3161;
wire n_2389;
wire n_2280;
wire n_7126;
wire n_5867;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_6430;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_6296;
wire n_4112;
wire n_5602;
wire n_2035;
wire n_4928;
wire n_7196;
wire n_2614;
wire n_7360;
wire n_5428;
wire n_6325;
wire n_2494;
wire n_4865;
wire n_6678;
wire n_2128;
wire n_4071;
wire n_6564;
wire n_7268;
wire n_4436;
wire n_5822;
wire n_5786;
wire n_3586;
wire n_5817;
wire n_4160;
wire n_6109;
wire n_6385;
wire n_5798;
wire n_4137;
wire n_5417;
wire n_4545;
wire n_4758;
wire n_4840;
wire n_5713;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_4535;
wire n_4385;
wire n_3748;
wire n_4731;
wire n_2337;
wire n_7073;
wire n_1786;
wire n_6309;
wire n_3732;
wire n_1804;
wire n_6519;
wire n_4671;
wire n_2272;
wire n_5571;
wire n_4766;
wire n_5989;
wire n_4558;
wire n_1769;
wire n_7349;
wire n_1929;
wire n_4319;
wire n_6585;
wire n_2929;
wire n_4358;
wire n_7122;
wire n_4874;
wire n_2656;
wire n_4904;
wire n_1997;
wire n_1733;
wire n_6490;
wire n_4651;
wire n_3167;
wire n_4748;
wire n_1807;
wire n_2857;
wire n_1784;
wire n_4618;
wire n_6721;
wire n_3787;
wire n_4025;
wire n_3050;
wire n_3919;
wire n_5506;
wire n_5475;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_5908;
wire n_5431;
wire n_5100;
wire n_2383;
wire n_2764;
wire n_1822;
wire n_7019;
wire n_5315;
wire n_2633;
wire n_3708;
wire n_5752;
wire n_2907;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_5746;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_3718;
wire n_6685;
wire n_3390;
wire n_2298;
wire n_4666;
wire n_3140;
wire n_2320;
wire n_4082;
wire n_3976;
wire n_2813;
wire n_2546;
wire n_3381;
wire n_7347;
wire n_3736;
wire n_4466;
wire n_6016;
wire n_3955;
wire n_5366;
wire n_5322;
wire n_1864;
wire n_5414;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_6971;
wire n_3336;
wire n_5903;
wire n_7199;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_5151;
wire n_3605;
wire n_5307;
wire n_2170;
wire n_4721;
wire n_6549;
wire n_5003;
wire n_3840;
wire n_6540;
wire n_7166;
wire n_2198;
wire n_6658;
wire n_5369;
wire n_6683;
wire n_3067;
wire n_3809;
wire n_4921;
wire n_1852;
wire n_5912;
wire n_5745;
wire n_6086;
wire n_4377;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_5803;
wire n_6327;
wire n_5593;
wire n_5270;
wire n_5853;
wire n_6171;
wire n_3468;
wire n_5779;
wire n_1877;
wire n_7213;
wire n_4301;
wire n_5313;
wire n_2133;
wire n_6820;
wire n_2497;
wire n_5446;
wire n_7107;
wire n_4561;
wire n_3291;
wire n_7456;
wire n_7369;
wire n_2578;
wire n_2475;
wire n_7250;
wire n_4715;
wire n_6157;
wire n_2715;
wire n_2665;
wire n_4879;
wire n_5044;
wire n_3755;
wire n_4536;
wire n_6676;
wire n_4304;
wire n_4927;
wire n_4078;
wire n_5459;
wire n_1801;
wire n_2854;
wire n_4418;
wire n_3341;
wire n_4125;
wire n_5390;
wire n_5351;
wire n_5267;
wire n_5024;
wire n_7012;
wire n_3043;
wire n_2747;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_4151;
wire n_2845;
wire n_4412;
wire n_2036;
wire n_6923;
wire n_3358;
wire n_6704;
wire n_2003;
wire n_2533;
wire n_7406;
wire n_4682;
wire n_6673;
wire n_2419;
wire n_2330;
wire n_6534;
wire n_5078;
wire n_4810;
wire n_6162;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_3289;
wire n_1955;
wire n_6127;
wire n_6246;
wire n_5005;
wire n_6126;
wire n_7372;
wire n_7427;
wire n_6151;
wire n_6828;
wire n_6841;
wire n_5207;
wire n_2658;
wire n_5624;
wire n_3620;
wire n_4601;
wire n_4518;
wire n_2767;
wire n_5474;
wire n_7009;
wire n_3376;
wire n_7371;
wire n_3123;
wire n_5447;
wire n_2692;
wire n_7463;
wire n_1960;
wire n_4102;
wire n_4308;
wire n_5700;
wire n_5755;
wire n_2862;
wire n_4325;
wire n_2645;
wire n_2553;
wire n_4711;
wire n_6889;
wire n_2749;
wire n_5962;
wire n_4413;
wire n_3307;
wire n_3251;
wire n_1885;
wire n_3288;
wire n_2833;
wire n_6723;
wire n_7398;
wire n_3723;
wire n_4135;
wire n_6154;
wire n_5223;
wire n_5662;
wire n_3880;
wire n_5801;
wire n_3904;
wire n_6054;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_7011;
wire n_3405;
wire n_2313;
wire n_6393;
wire n_7074;
wire n_5465;
wire n_3532;
wire n_5154;
wire n_5721;
wire n_2609;
wire n_6184;
wire n_1767;
wire n_3131;
wire n_4138;
wire n_7083;
wire n_1973;
wire n_2882;
wire n_7143;
wire n_2303;
wire n_4384;
wire n_4639;
wire n_4577;
wire n_6312;
wire n_2154;
wire n_1986;
wire n_6711;
wire n_2624;
wire n_6818;
wire n_6438;
wire n_2054;
wire n_1857;
wire n_3926;
wire n_4481;
wire n_5087;
wire n_2938;
wire n_7209;
wire n_2498;
wire n_6193;
wire n_3992;
wire n_7330;
wire n_6007;
wire n_6734;
wire n_6535;
wire n_1772;
wire n_6879;
wire n_3106;
wire n_6208;
wire n_7190;
wire n_2881;
wire n_6303;
wire n_3092;
wire n_6014;
wire n_4270;
wire n_4620;
wire n_5397;
wire n_6255;
wire n_6457;
wire n_4924;
wire n_4044;
wire n_6270;
wire n_2305;
wire n_5996;
wire n_5566;
wire n_3304;
wire n_7288;
wire n_4388;
wire n_7362;
wire n_7082;
wire n_7237;
wire n_3247;
wire n_7131;
wire n_6276;
wire n_4406;
wire n_2180;
wire n_4271;
wire n_7042;
wire n_2809;
wire n_5652;
wire n_5805;
wire n_7304;
wire n_6266;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_3785;
wire n_5492;
wire n_2465;
wire n_5501;
wire n_6934;
wire n_7386;
wire n_2972;
wire n_7391;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_3178;
wire n_7023;
wire n_2251;
wire n_5758;
wire n_5842;
wire n_3100;
wire n_3721;
wire n_7404;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_6147;
wire n_5692;
wire n_6765;
wire n_4973;
wire n_4792;
wire n_3537;
wire n_4402;
wire n_2487;
wire n_5473;
wire n_1834;
wire n_2534;
wire n_6352;
wire n_2941;
wire n_4286;
wire n_3638;
wire n_6211;
wire n_3576;
wire n_5562;
wire n_4858;
wire n_6093;
wire n_5370;
wire n_7378;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_5458;
wire n_2387;
wire n_4318;
wire n_5227;
wire n_5902;
wire n_2510;
wire n_6402;
wire n_3570;
wire n_3227;
wire n_5359;
wire n_4673;
wire n_2793;
wire n_5282;
wire n_6764;
wire n_2639;
wire n_7016;
wire n_4738;
wire n_2603;
wire n_5386;
wire n_6215;
wire n_4554;
wire n_4526;
wire n_4105;
wire n_3663;
wire n_6955;
wire n_5952;
wire n_7180;
wire n_2086;
wire n_1926;
wire n_6569;
wire n_1720;
wire n_2966;
wire n_2409;
wire n_3431;
wire n_3355;
wire n_7031;
wire n_1738;
wire n_5716;
wire n_3897;
wire n_7103;
wire n_6605;
wire n_1735;
wire n_5888;
wire n_4005;
wire n_4181;
wire n_2543;
wire n_2321;
wire n_2597;
wire n_6832;
wire n_5980;
wire n_4092;
wire n_4875;
wire n_4255;
wire n_2758;
wire n_6544;
wire n_6469;
wire n_5036;
wire n_6332;
wire n_2186;
wire n_5790;
wire n_7130;
wire n_6680;
wire n_4647;
wire n_3575;
wire n_6310;
wire n_2471;
wire n_7134;
wire n_3042;
wire n_1937;
wire n_4142;
wire n_5118;
wire n_5485;
wire n_5525;
wire n_7102;
wire n_6259;
wire n_3004;
wire n_4849;
wire n_5271;
wire n_2039;
wire n_7133;
wire n_6289;
wire n_3838;
wire n_6651;
wire n_4059;
wire n_6565;
wire n_5194;
wire n_5445;
wire n_2734;
wire n_5948;
wire n_7227;
wire n_4499;
wire n_4504;
wire n_3598;
wire n_4917;
wire n_2420;
wire n_6836;
wire n_3273;
wire n_2918;
wire n_6595;
wire n_6186;
wire n_1865;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_1792;
wire n_5628;
wire n_5245;
wire n_2062;
wire n_4489;
wire n_2153;
wire n_5329;
wire n_5472;
wire n_6035;
wire n_1754;
wire n_7236;
wire n_4833;
wire n_3394;
wire n_6405;
wire n_2235;
wire n_5850;
wire n_6786;
wire n_4564;
wire n_1848;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_3581;
wire n_5072;
wire n_3778;
wire n_6769;
wire n_6844;
wire n_4322;
wire n_6361;
wire n_2260;
wire n_4080;
wire n_2206;
wire n_6766;
wire n_4185;
wire n_5940;
wire n_3001;
wire n_5260;
wire n_6751;
wire n_4981;
wire n_6232;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_7457;
wire n_5372;
wire n_6736;
wire n_4507;
wire n_4756;
wire n_5860;
wire n_2422;
wire n_6416;
wire n_2933;
wire n_3387;
wire n_6214;
wire n_3952;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_7049;
wire n_6945;
wire n_6143;
wire n_2736;
wire n_6491;
wire n_3825;
wire n_4198;
wire n_7172;
wire n_2339;
wire n_6225;
wire n_2532;
wire n_4373;
wire n_1866;
wire n_2664;
wire n_4154;
wire n_7344;
wire n_5859;
wire n_6447;
wire n_4390;
wire n_1782;
wire n_4107;
wire n_2519;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_7325;
wire n_2360;
wire n_4453;
wire n_6219;
wire n_6175;
wire n_6445;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_3032;
wire n_5612;
wire n_4886;
wire n_6198;
wire n_5172;
wire n_6499;
wire n_1982;
wire n_5311;
wire n_5164;
wire n_4964;
wire n_4700;
wire n_6842;
wire n_4002;
wire n_7361;
wire n_1742;
wire n_4679;
wire n_6397;
wire n_3815;
wire n_6827;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_2982;
wire n_5495;
wire n_6281;
wire n_4483;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_5547;
wire n_4693;
wire n_6822;
wire n_5121;
wire n_4956;
wire n_2869;
wire n_5379;
wire n_7079;
wire n_4487;
wire n_5878;
wire n_2674;
wire n_5820;
wire n_1737;
wire n_7309;
wire n_7119;
wire n_3026;
wire n_7184;
wire n_2979;
wire n_4329;
wire n_5291;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_3902;
wire n_3244;
wire n_1779;
wire n_3112;
wire n_2562;
wire n_2051;
wire n_3196;
wire n_5964;
wire n_2673;
wire n_6076;
wire n_4678;
wire n_5301;
wire n_5126;
wire n_6732;
wire n_2548;
wire n_3488;
wire n_2381;
wire n_2744;
wire n_6817;
wire n_1967;
wire n_5776;
wire n_2179;
wire n_3779;
wire n_6982;
wire n_7291;
wire n_2275;
wire n_7435;
wire n_4606;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_5603;
wire n_1891;
wire n_6560;
wire n_6634;
wire n_5348;
wire n_4868;
wire n_7017;
wire n_4072;
wire n_2792;
wire n_4465;
wire n_2596;
wire n_5217;
wire n_3986;
wire n_5558;
wire n_3725;
wire n_4026;
wire n_4245;
wire n_5520;
wire n_2524;
wire n_3894;
wire n_5909;
wire n_4852;
wire n_3202;
wire n_4290;
wire n_4945;
wire n_5750;
wire n_1725;
wire n_5654;
wire n_2318;
wire n_2819;
wire n_1722;
wire n_2229;
wire n_6400;
wire n_3547;
wire n_4014;
wire n_2551;
wire n_2255;
wire n_5554;
wire n_3045;
wire n_5135;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_6655;
wire n_1905;
wire n_5448;
wire n_2573;
wire n_6480;
wire n_5837;
wire n_2336;
wire n_5412;
wire n_3249;
wire n_3483;
wire n_6621;
wire n_6851;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_2915;
wire n_7420;
wire n_4869;
wire n_3213;
wire n_5533;
wire n_4047;
wire n_1796;
wire n_2719;
wire n_2876;
wire n_4063;
wire n_5224;
wire n_2778;
wire n_6226;
wire n_3033;
wire n_1981;
wire n_2824;
wire n_5327;
wire n_4417;
wire n_2089;
wire n_6283;
wire n_4688;
wire n_7156;
wire n_4939;
wire n_5900;
wire n_7319;
wire n_3619;
wire n_6158;
wire n_4013;
wire n_3434;
wire n_4342;
wire n_6819;
wire n_4903;
wire n_6122;
wire n_2131;
wire n_3853;
wire n_4382;
wire n_4085;
wire n_2509;
wire n_6898;
wire n_6570;
wire n_5486;
wire n_2135;
wire n_7260;
wire n_6894;
wire n_4475;
wire n_6843;
wire n_5432;
wire n_5851;
wire n_6317;
wire n_6928;
wire n_6707;
wire n_7244;
wire n_4626;
wire n_4997;
wire n_5065;
wire n_6806;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_6835;
wire n_7286;
wire n_2436;
wire n_3517;
wire n_6269;
wire n_2461;
wire n_3719;
wire n_7154;
wire n_3526;
wire n_3888;
wire n_3198;
wire n_1853;
wire n_5295;
wire n_6088;
wire n_1999;
wire n_7194;
wire n_4841;
wire n_4683;
wire n_5173;
wire n_2873;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_5655;
wire n_3383;
wire n_1835;
wire n_5855;
wire n_7175;
wire n_3965;
wire n_3905;
wire n_7163;
wire n_3797;
wire n_1836;
wire n_7027;
wire n_3416;
wire n_4600;
wire n_5861;
wire n_6964;
wire n_3943;
wire n_3145;
wire n_5749;
wire n_6320;
wire n_6316;
wire n_7068;
wire n_2908;
wire n_4106;
wire n_2156;
wire n_2323;
wire n_4549;
wire n_7327;
wire n_1746;
wire n_6610;
wire n_5998;
wire n_4702;
wire n_5102;
wire n_4954;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_6752;
wire n_6959;
wire n_6250;
wire n_3283;
wire n_4331;
wire n_7317;
wire n_4159;
wire n_3451;
wire n_4734;
wire n_6675;
wire n_2832;
wire n_5827;
wire n_2370;
wire n_1944;
wire n_7384;
wire n_2914;
wire n_5656;
wire n_7218;
wire n_1988;
wire n_5678;
wire n_6561;
wire n_6858;
wire n_5865;
wire n_6050;
wire n_1718;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_2539;
wire n_5555;
wire n_2078;
wire n_4809;
wire n_7152;
wire n_4012;
wire n_2049;
wire n_5212;
wire n_4760;
wire n_6823;
wire n_3606;
wire n_7062;
wire n_7090;
wire n_2232;
wire n_1847;
wire n_5815;
wire n_4320;
wire n_5084;
wire n_7223;
wire n_5251;
wire n_5965;
wire n_4980;
wire n_3324;
wire n_2192;
wire n_6796;
wire n_5407;
wire n_2988;
wire n_4560;
wire n_3230;
wire n_3793;
wire n_5042;
wire n_7055;
wire n_6024;
wire n_4768;
wire n_1889;
wire n_6090;
wire n_5368;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_3607;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_7388;
wire n_1751;
wire n_7056;
wire n_7437;
wire n_6489;
wire n_5310;
wire n_2769;
wire n_4987;
wire n_6714;
wire n_3013;
wire n_4572;
wire n_7417;
wire n_2739;
wire n_3962;
wire n_4988;
wire n_7446;
wire n_6038;
wire n_2902;
wire n_6030;
wire n_6245;
wire n_4360;
wire n_6620;
wire n_6791;
wire n_4540;
wire n_6821;
wire n_2094;
wire n_5588;
wire n_3854;
wire n_6583;
wire n_2349;
wire n_3652;
wire n_3449;
wire n_3089;
wire n_4854;
wire n_5477;
wire n_2727;
wire n_5234;
wire n_6890;
wire n_6988;
wire n_5871;
wire n_4747;
wire n_3472;
wire n_2527;
wire n_6052;
wire n_7257;
wire n_3126;
wire n_2759;
wire n_6973;
wire n_5007;
wire n_4881;
wire n_2038;
wire n_6488;
wire n_3958;
wire n_4495;
wire n_4737;
wire n_1838;
wire n_4357;
wire n_2806;
wire n_4502;
wire n_3191;
wire n_1716;
wire n_7005;
wire n_5334;
wire n_3562;
wire n_2281;
wire n_7081;
wire n_5253;
wire n_3588;
wire n_6280;
wire n_3280;
wire n_4115;
wire n_5274;
wire n_6399;
wire n_5418;
wire n_5019;
wire n_5939;
wire n_1819;
wire n_3095;
wire n_7341;
wire n_5792;
wire n_3698;
wire n_4513;
wire n_4775;
wire n_6256;
wire n_2620;
wire n_1833;
wire n_7264;
wire n_2499;
wire n_2549;
wire n_6648;
wire n_6649;
wire n_3093;
wire n_2970;
wire n_6910;
wire n_3885;
wire n_4264;
wire n_5954;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_6431;
wire n_3250;
wire n_4223;
wire n_3538;
wire n_3915;
wire n_3839;
wire n_7285;
wire n_5490;
wire n_5694;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_6324;
wire n_5489;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_4206;
wire n_2415;
wire n_4099;
wire n_3120;
wire n_6512;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_5342;
wire n_4794;
wire n_4843;
wire n_5580;
wire n_5215;
wire n_3937;
wire n_4763;
wire n_6243;
wire n_5795;
wire n_5715;
wire n_4170;
wire n_5561;
wire n_2462;
wire n_7051;
wire n_6773;
wire n_2155;
wire n_6231;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_3604;
wire n_5430;
wire n_6041;
wire n_5659;
wire n_6859;
wire n_4272;
wire n_5195;
wire n_3176;
wire n_3792;
wire n_6323;
wire n_5720;
wire n_4267;
wire n_2083;
wire n_5598;
wire n_2753;
wire n_3021;
wire n_4352;
wire n_2712;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_2898;
wire n_1825;
wire n_6912;
wire n_3567;
wire n_7425;
wire n_2682;
wire n_5854;
wire n_5958;
wire n_5585;
wire n_5112;
wire n_5326;
wire n_5783;
wire n_6837;
wire n_6747;
wire n_2903;
wire n_5303;
wire n_3812;
wire n_3127;
wire n_6916;
wire n_1731;
wire n_2378;
wire n_5530;
wire n_6718;
wire n_5809;
wire n_2213;
wire n_7121;
wire n_6410;
wire n_6473;
wire n_4056;
wire n_4806;
wire n_5993;
wire n_4015;
wire n_6574;
wire n_2924;
wire n_6492;
wire n_4445;
wire n_4462;
wire n_5299;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_2142;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_3170;
wire n_2311;
wire n_6857;
wire n_2287;
wire n_3415;
wire n_6975;
wire n_3464;
wire n_6290;
wire n_3414;
wire n_6646;
wire n_4234;
wire n_3467;
wire n_5821;
wire n_3179;
wire n_6622;
wire n_5522;
wire n_4836;
wire n_3889;
wire n_5262;
wire n_3262;
wire n_5319;
wire n_3699;
wire n_6118;
wire n_2120;
wire n_7125;
wire n_6028;
wire n_6663;
wire n_6532;
wire n_3816;
wire n_3528;
wire n_6267;
wire n_6682;
wire n_4207;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_4725;
wire n_2312;
wire n_7203;
wire n_1826;
wire n_5943;
wire n_6556;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_6216;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_7128;
wire n_5335;
wire n_6365;
wire n_7111;
wire n_2801;
wire n_4334;
wire n_5284;
wire n_4978;
wire n_5771;
wire n_3246;
wire n_3299;
wire n_1869;
wire n_3623;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_6950;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_5516;
wire n_7284;
wire n_3615;
wire n_7057;
wire n_1802;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_3200;
wire n_6167;
wire n_3642;
wire n_2146;
wire n_4274;
wire n_5583;
wire n_3276;
wire n_7064;
wire n_5433;
wire n_3682;
wire n_5429;
wire n_7278;
wire n_6772;
wire n_7088;
wire n_5698;
wire n_5731;
wire n_4007;
wire n_1879;
wire n_6159;
wire n_2129;
wire n_5857;
wire n_7048;
wire n_6617;
wire n_5120;
wire n_3572;
wire n_2975;
wire n_2399;
wire n_3471;
wire n_4075;
wire n_2932;
wire n_2027;
wire n_6217;
wire n_3118;
wire n_5560;
wire n_4441;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_5455;
wire n_6777;
wire n_6742;
wire n_7447;
wire n_5209;
wire n_6307;
wire n_5704;
wire n_4458;
wire n_2159;
wire n_4889;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_3618;
wire n_5916;
wire n_3705;
wire n_3022;
wire n_1709;
wire n_6479;
wire n_5099;
wire n_3286;
wire n_5781;
wire n_5619;
wire n_2023;
wire n_3974;
wire n_7365;
wire n_3443;
wire n_3988;
wire n_2599;
wire n_5022;
wire n_6370;
wire n_2075;
wire n_1726;
wire n_2031;
wire n_3761;
wire n_3996;
wire n_7275;
wire n_5353;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_6856;
wire n_3009;
wire n_7095;
wire n_7390;
wire n_6140;
wire n_6111;
wire n_5219;
wire n_3951;
wire n_5518;
wire n_3035;
wire n_4261;
wire n_7037;
wire n_1823;
wire n_6240;
wire n_5236;
wire n_4236;
wire n_3942;
wire n_3023;
wire n_2254;
wire n_3290;
wire n_6693;
wire n_6712;
wire n_3957;
wire n_3418;
wire n_6465;
wire n_5673;
wire n_5814;
wire n_6586;
wire n_7058;
wire n_5103;
wire n_4648;
wire n_2214;
wire n_6730;
wire n_6367;
wire n_2256;
wire n_3326;
wire n_6069;
wire n_2732;
wire n_1883;
wire n_6515;
wire n_4094;
wire n_2776;
wire n_6077;
wire n_3224;
wire n_1969;
wire n_5671;
wire n_7429;
wire n_6940;
wire n_2949;
wire n_7008;
wire n_6468;
wire n_4269;
wire n_1927;
wire n_7139;
wire n_3803;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_7432;
wire n_2124;
wire n_1894;
wire n_4913;
wire n_2449;
wire n_4428;
wire n_6483;
wire n_4463;
wire n_5357;
wire n_7173;
wire n_3648;
wire n_6576;
wire n_6810;
wire n_1975;
wire n_5421;
wire n_4396;
wire n_1990;
wire n_6708;
wire n_6667;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_6040;
wire n_1890;
wire n_6847;
wire n_6305;
wire n_4034;
wire n_4228;
wire n_7251;
wire n_3166;
wire n_7356;
wire n_3649;
wire n_7412;
wire n_3065;
wire n_7212;
wire n_5045;
wire n_5237;
wire n_7060;
wire n_3924;
wire n_3997;
wire n_3564;
wire n_5769;
wire n_2637;
wire n_6750;
wire n_7444;
wire n_3795;
wire n_4931;
wire n_2306;
wire n_2071;
wire n_7426;
wire n_3953;
wire n_4400;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_5434;
wire n_6855;
wire n_5181;
wire n_6239;
wire n_3208;
wire n_5768;
wire n_6199;
wire n_2737;
wire n_3282;
wire n_2916;
wire n_7252;
wire n_5963;
wire n_4424;
wire n_4351;
wire n_6543;
wire n_4192;
wire n_1748;
wire n_6789;
wire n_5972;
wire n_3400;
wire n_7065;
wire n_6177;
wire n_2581;
wire n_5937;
wire n_1783;
wire n_5146;
wire n_7367;
wire n_7267;
wire n_7405;
wire n_4646;
wire n_4221;
wire n_3650;
wire n_6825;
wire n_1993;
wire n_6460;
wire n_4035;
wire n_6952;
wire n_3670;
wire n_6173;
wire n_2540;
wire n_4190;
wire n_3060;
wire n_6218;
wire n_6486;
wire n_2984;
wire n_4009;
wire n_2489;
wire n_5013;
wire n_4145;
wire n_6852;
wire n_5577;
wire n_5872;
wire n_6692;
wire n_5017;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_7220;
wire n_2106;
wire n_5976;
wire n_4717;
wire n_6888;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_2091;
wire n_4312;
wire n_5424;
wire n_3789;
wire n_7270;
wire n_4750;
wire n_2348;
wire n_1873;
wire n_2667;
wire n_2725;
wire n_3746;
wire n_6626;
wire n_4537;
wire n_5838;
wire n_7034;
wire n_3694;
wire n_6854;
wire n_6793;
wire n_5456;
wire n_3893;
wire n_4847;
wire n_5846;
wire n_2307;
wire n_3702;
wire n_5930;
wire n_1984;
wire n_3453;
wire n_6980;
wire n_7040;
wire n_5345;
wire n_2815;
wire n_4427;
wire n_7458;
wire n_1824;
wire n_4065;
wire n_4705;
wire n_6794;
wire n_2945;
wire n_1971;
wire n_3543;
wire n_7179;
wire n_3448;
wire n_1776;
wire n_7433;
wire n_4279;
wire n_2936;
wire n_3609;
wire n_4330;
wire n_6334;
wire n_6257;
wire n_4152;
wire n_6874;
wire n_5537;
wire n_2698;
wire n_5572;
wire n_4783;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_2789;
wire n_5409;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_5142;
wire n_6355;
wire n_7015;
wire n_6039;
wire n_6286;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_7226;
wire n_1987;
wire n_7217;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_6377;
wire n_5401;
wire n_4595;
wire n_7272;
wire n_2352;
wire n_5201;
wire n_5816;
wire n_5551;
wire n_5416;
wire n_4404;
wire n_2377;
wire n_2652;
wire n_5498;
wire n_5543;
wire n_4054;
wire n_6018;
wire n_6021;
wire n_4617;
wire n_2477;
wire n_4611;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_5797;
wire n_6511;
wire n_4732;
wire n_2076;
wire n_2203;
wire n_5942;
wire n_5764;
wire n_4969;
wire n_5252;
wire n_5777;
wire n_4641;
wire n_5063;
wire n_4399;
wire n_6867;
wire n_4140;
wire n_5171;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_7255;
wire n_3309;
wire n_7181;
wire n_2796;
wire n_5393;
wire n_4817;
wire n_6863;
wire n_7352;
wire n_7355;
wire n_2136;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_7328;
wire n_2771;
wire n_6322;
wire n_7359;
wire n_2403;
wire n_2947;
wire n_5643;
wire n_3769;
wire n_4437;
wire n_6419;
wire n_3055;
wire n_4070;
wire n_5346;
wire n_7283;
wire n_7089;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_4139;
wire n_4769;
wire n_6130;
wire n_5868;
wire n_6417;
wire n_7145;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_2713;
wire n_1965;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_6979;
wire n_5986;
wire n_6932;
wire n_2934;
wire n_7258;
wire n_5104;
wire n_6961;
wire n_6792;
wire n_2210;
wire n_4368;
wire n_5794;
wire n_3141;
wire n_2053;
wire n_5272;
wire n_3476;
wire n_6919;
wire n_4430;
wire n_6123;
wire n_3238;
wire n_2450;
wire n_5338;
wire n_7440;
wire n_6831;
wire n_1773;
wire n_3175;
wire n_4544;
wire n_2666;
wire n_5578;
wire n_4191;
wire n_4409;
wire n_2401;
wire n_3255;
wire n_2588;
wire n_5722;
wire n_5811;
wire n_7072;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_3509;
wire n_5395;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_6458;
wire n_6986;
wire n_3456;
wire n_4532;
wire n_5863;
wire n_6633;
wire n_3790;
wire n_7118;
wire n_6152;
wire n_5734;
wire n_2566;
wire n_5095;
wire n_3101;
wire n_3662;
wire n_6169;
wire n_5774;
wire n_7069;
wire n_5199;
wire n_6546;
wire n_4257;
wire n_4282;
wire n_4341;
wire n_6925;
wire n_7186;
wire n_4027;
wire n_4309;
wire n_4650;
wire n_5480;
wire n_6428;
wire n_6924;
wire n_3077;
wire n_4944;
wire n_6425;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_4994;
wire n_5977;
wire n_3533;
wire n_5175;
wire n_7246;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_3409;
wire n_4381;
wire n_3583;
wire n_4316;
wire n_7301;
wire n_4860;
wire n_4469;
wire n_3540;
wire n_4930;
wire n_5352;
wire n_7262;
wire n_5959;
wire n_3563;
wire n_5945;
wire n_1739;
wire n_3310;
wire n_2642;
wire n_4423;
wire n_3689;
wire n_1789;
wire n_6301;
wire n_2174;
wire n_5668;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_4703;
wire n_6282;
wire n_4934;
wire n_2638;
wire n_2046;
wire n_7059;
wire n_6985;
wire n_1756;
wire n_4350;
wire n_5600;
wire n_6737;
wire n_2340;
wire n_4804;
wire n_2444;
wire n_4888;
wire n_5767;
wire n_6459;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_2199;
wire n_6384;
wire n_4669;
wire n_5228;
wire n_2600;
wire n_7443;
wire n_3436;
wire n_5973;
wire n_1962;
wire n_3806;
wire n_4759;
wire n_5869;
wire n_5914;
wire n_2114;
wire n_6753;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_4887;
wire n_3751;
wire n_3402;
wire n_6448;
wire n_5186;
wire n_4585;
wire n_1785;
wire n_3406;
wire n_3664;
wire n_4218;
wire n_4687;
wire n_7077;
wire n_3686;
wire n_4720;
wire n_2889;
wire n_6043;
wire n_6268;
wire n_2141;
wire n_1758;
wire n_5604;
wire n_3470;
wire n_5221;
wire n_7024;
wire n_6145;
wire n_2865;
wire n_5925;
wire n_6529;
wire n_5591;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_7214;
wire n_2572;
wire n_4490;
wire n_3677;
wire n_5387;
wire n_3292;
wire n_6311;
wire n_3989;
wire n_4644;
wire n_4752;
wire n_4746;
wire n_4131;
wire n_5449;
wire n_4215;
wire n_2488;
wire n_6134;
wire n_4158;
wire n_6812;
wire n_3079;
wire n_5190;
wire n_6733;
wire n_3269;
wire n_5325;
wire n_4231;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_6262;
wire n_4926;
wire n_2050;
wire n_6938;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_5876;
wire n_5344;
wire n_2550;
wire n_3177;
wire n_6160;
wire n_4667;
wire n_5813;
wire n_6235;
wire n_6212;
wire n_3440;
wire n_6816;
wire n_3658;
wire n_7374;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_2542;
wire n_5892;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_7110;
wire n_5714;
wire n_2169;
wire n_6953;
wire n_6089;
wire n_5634;
wire n_5133;
wire n_5305;
wire n_5990;
wire n_2175;
wire n_7086;
wire n_5689;
wire n_4578;
wire n_5644;
wire n_3644;
wire n_2176;
wire n_3059;
wire n_6138;
wire n_1922;
wire n_4877;
wire n_2065;
wire n_7038;
wire n_4470;
wire n_4187;
wire n_1904;
wire n_4998;
wire n_5576;
wire n_2395;
wire n_2868;
wire n_7345;
wire n_4057;
wire n_6070;
wire n_5852;
wire n_5918;
wire n_2724;
wire n_2258;
wire n_7041;
wire n_6717;
wire n_6881;
wire n_3328;
wire n_2012;
wire n_3182;
wire n_6871;
wire n_2967;
wire n_5343;
wire n_6672;
wire n_6518;
wire n_7334;
wire n_4021;
wire n_6396;
wire n_7028;
wire n_3379;
wire n_4379;
wire n_5947;
wire n_6242;
wire n_6601;
wire n_2268;
wire n_3469;
wire n_2835;
wire n_5835;
wire n_2111;
wire n_3743;
wire n_5542;
wire n_2948;
wire n_5015;
wire n_3099;
wire n_5527;
wire n_2897;
wire n_4812;
wire n_4497;
wire n_6606;
wire n_2583;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_1770;
wire n_4472;
wire n_2699;
wire n_5819;
wire n_3901;
wire n_5180;
wire n_2973;
wire n_5893;
wire n_2710;
wire n_6092;
wire n_6462;
wire n_2505;
wire n_4519;
wire n_5025;
wire n_2397;
wire n_7333;
wire n_3878;
wire n_4197;
wire n_6669;
wire n_2721;
wire n_1892;
wire n_6251;
wire n_2615;
wire n_4787;
wire n_7337;
wire n_4310;
wire n_4566;
wire n_3933;
wire n_5726;
wire n_7439;
wire n_4371;
wire n_1902;
wire n_5828;
wire n_2784;
wire n_7210;
wire n_3898;
wire n_6228;
wire n_6702;
wire n_7358;
wire n_4749;
wire n_5924;
wire n_1845;
wire n_5545;
wire n_2104;
wire n_2552;
wire n_5083;
wire n_3253;
wire n_2088;
wire n_6997;
wire n_4238;
wire n_6371;
wire n_2005;
wire n_7187;
wire n_2108;
wire n_3824;
wire n_2246;
wire n_7313;
wire n_5899;
wire n_3846;
wire n_5122;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_6641;
wire n_3845;
wire n_6463;
wire n_3203;
wire n_4986;
wire n_4668;
wire n_6264;
wire n_5782;
wire n_4168;
wire n_7036;
wire n_4298;
wire n_7370;
wire n_4743;
wire n_1781;
wire n_4250;
wire n_3143;
wire n_3690;
wire n_3229;
wire n_5864;
wire n_2188;
wire n_2430;
wire n_2504;
wire n_5637;
wire n_4211;
wire n_6084;
wire n_3094;
wire n_5185;
wire n_2964;
wire n_5032;
wire n_6990;
wire n_5034;
wire n_3312;
wire n_7071;
wire n_2451;
wire n_2913;
wire n_6288;
wire n_1862;
wire n_3752;
wire n_3672;
wire n_7380;
wire n_2839;
wire n_3237;
wire n_4128;
wire n_4036;
wire n_5269;
wire n_3655;
wire n_2955;
wire n_5709;
wire n_1764;
wire n_4807;
wire n_6277;
wire n_5115;
wire n_7376;
wire n_1723;
wire n_3918;
wire n_5324;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_6409;
wire n_4095;
wire n_5927;
wire n_4485;
wire n_6388;
wire n_3593;
wire n_6839;
wire n_5163;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_1896;
wire n_6864;
wire n_4890;
wire n_2485;
wire n_6679;
wire n_6051;
wire n_2563;
wire n_4224;
wire n_1799;
wire n_5507;
wire n_4573;
wire n_4943;
wire n_2875;
wire n_6599;
wire n_3519;
wire n_2209;
wire n_4042;
wire n_7099;
wire n_4244;
wire n_1928;
wire n_5642;
wire n_4708;
wire n_4883;
wire n_6227;
wire n_4553;
wire n_7052;
wire n_6738;
wire n_5226;
wire n_2081;
wire n_6566;
wire n_1794;
wire n_5696;
wire n_3053;
wire n_5014;
wire n_7106;
wire n_6346;
wire n_3772;
wire n_7408;
wire n_2891;
wire n_4335;
wire n_7026;
wire n_3128;
wire n_6146;
wire n_5677;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_7394;
wire n_4516;
wire n_5235;
wire n_6436;
wire n_2798;
wire n_7450;
wire n_3217;
wire n_6081;
wire n_5724;
wire n_3821;
wire n_3201;
wire n_7462;
wire n_3503;
wire n_5979;
wire n_6027;
wire n_1870;
wire n_4467;
wire n_5521;
wire n_2654;
wire n_3935;
wire n_7421;
wire n_1861;
wire n_2319;
wire n_2965;
wire n_4955;
wire n_5410;
wire n_1989;
wire n_2689;
wire n_6110;
wire n_1762;
wire n_6238;
wire n_7025;
wire n_3798;
wire n_3080;
wire n_5241;
wire n_4248;
wire n_2228;
wire n_4645;
wire n_5331;
wire n_3308;
wire n_6326;
wire n_3204;
wire n_7451;
wire n_4134;
wire n_5018;
wire n_6917;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_1730;
wire n_6612;
wire n_5258;

INVx1_ASAP7_75t_L g1709 ( 
.A(n_445),
.Y(n_1709)
);

CKINVDCx5p33_ASAP7_75t_R g1710 ( 
.A(n_1414),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_890),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_1296),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_306),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1262),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1482),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_1458),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_1536),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_654),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_126),
.Y(n_1719)
);

BUFx3_ASAP7_75t_L g1720 ( 
.A(n_1474),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1645),
.Y(n_1721)
);

INVx2_ASAP7_75t_SL g1722 ( 
.A(n_914),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_890),
.Y(n_1723)
);

CKINVDCx5p33_ASAP7_75t_R g1724 ( 
.A(n_676),
.Y(n_1724)
);

CKINVDCx14_ASAP7_75t_R g1725 ( 
.A(n_228),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_592),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_1550),
.Y(n_1727)
);

BUFx10_ASAP7_75t_L g1728 ( 
.A(n_1623),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_194),
.Y(n_1729)
);

CKINVDCx5p33_ASAP7_75t_R g1730 ( 
.A(n_1219),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1698),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_790),
.Y(n_1732)
);

CKINVDCx16_ASAP7_75t_R g1733 ( 
.A(n_1667),
.Y(n_1733)
);

INVxp67_ASAP7_75t_SL g1734 ( 
.A(n_523),
.Y(n_1734)
);

BUFx10_ASAP7_75t_L g1735 ( 
.A(n_476),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1073),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_474),
.Y(n_1737)
);

CKINVDCx20_ASAP7_75t_R g1738 ( 
.A(n_1358),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_1061),
.Y(n_1739)
);

BUFx3_ASAP7_75t_L g1740 ( 
.A(n_1017),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_1512),
.Y(n_1741)
);

INVxp67_ASAP7_75t_L g1742 ( 
.A(n_616),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_1563),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_1137),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_1244),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_1174),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_1226),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_839),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_1630),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_1643),
.Y(n_1750)
);

INVx2_ASAP7_75t_SL g1751 ( 
.A(n_500),
.Y(n_1751)
);

BUFx6f_ASAP7_75t_L g1752 ( 
.A(n_1125),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1049),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_350),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_1460),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_1578),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_1268),
.Y(n_1757)
);

BUFx6f_ASAP7_75t_L g1758 ( 
.A(n_791),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_1547),
.Y(n_1759)
);

CKINVDCx14_ASAP7_75t_R g1760 ( 
.A(n_323),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1327),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_1451),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_161),
.Y(n_1763)
);

INVx1_ASAP7_75t_SL g1764 ( 
.A(n_606),
.Y(n_1764)
);

INVx1_ASAP7_75t_SL g1765 ( 
.A(n_244),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_563),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_1646),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_1463),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1411),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_44),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_331),
.Y(n_1771)
);

CKINVDCx5p33_ASAP7_75t_R g1772 ( 
.A(n_361),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_792),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1469),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_1597),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1589),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_128),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_498),
.Y(n_1778)
);

CKINVDCx20_ASAP7_75t_R g1779 ( 
.A(n_218),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_550),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_517),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_1200),
.Y(n_1782)
);

CKINVDCx5p33_ASAP7_75t_R g1783 ( 
.A(n_1702),
.Y(n_1783)
);

CKINVDCx20_ASAP7_75t_R g1784 ( 
.A(n_676),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_977),
.Y(n_1785)
);

BUFx3_ASAP7_75t_L g1786 ( 
.A(n_1118),
.Y(n_1786)
);

CKINVDCx5p33_ASAP7_75t_R g1787 ( 
.A(n_427),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_175),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_775),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_1422),
.Y(n_1790)
);

INVx3_ASAP7_75t_L g1791 ( 
.A(n_1484),
.Y(n_1791)
);

CKINVDCx5p33_ASAP7_75t_R g1792 ( 
.A(n_1670),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1602),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_867),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_1346),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1493),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1688),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1342),
.Y(n_1798)
);

BUFx3_ASAP7_75t_L g1799 ( 
.A(n_231),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_1334),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_582),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_1222),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1542),
.Y(n_1803)
);

CKINVDCx5p33_ASAP7_75t_R g1804 ( 
.A(n_1491),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_1398),
.Y(n_1805)
);

BUFx10_ASAP7_75t_L g1806 ( 
.A(n_323),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1468),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_290),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1499),
.Y(n_1809)
);

CKINVDCx5p33_ASAP7_75t_R g1810 ( 
.A(n_343),
.Y(n_1810)
);

CKINVDCx20_ASAP7_75t_R g1811 ( 
.A(n_413),
.Y(n_1811)
);

CKINVDCx5p33_ASAP7_75t_R g1812 ( 
.A(n_348),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_30),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_1112),
.Y(n_1814)
);

CKINVDCx20_ASAP7_75t_R g1815 ( 
.A(n_195),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1348),
.Y(n_1816)
);

CKINVDCx5p33_ASAP7_75t_R g1817 ( 
.A(n_1592),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_574),
.Y(n_1818)
);

CKINVDCx5p33_ASAP7_75t_R g1819 ( 
.A(n_1194),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_647),
.Y(n_1820)
);

CKINVDCx5p33_ASAP7_75t_R g1821 ( 
.A(n_1494),
.Y(n_1821)
);

CKINVDCx5p33_ASAP7_75t_R g1822 ( 
.A(n_294),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_304),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_294),
.Y(n_1824)
);

INVx1_ASAP7_75t_SL g1825 ( 
.A(n_1276),
.Y(n_1825)
);

BUFx3_ASAP7_75t_L g1826 ( 
.A(n_1205),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1333),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_447),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_1197),
.Y(n_1829)
);

CKINVDCx5p33_ASAP7_75t_R g1830 ( 
.A(n_1616),
.Y(n_1830)
);

CKINVDCx20_ASAP7_75t_R g1831 ( 
.A(n_1178),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1675),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_437),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_520),
.Y(n_1834)
);

CKINVDCx5p33_ASAP7_75t_R g1835 ( 
.A(n_1660),
.Y(n_1835)
);

CKINVDCx5p33_ASAP7_75t_R g1836 ( 
.A(n_1671),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_893),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1700),
.Y(n_1838)
);

INVx1_ASAP7_75t_SL g1839 ( 
.A(n_1707),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_771),
.Y(n_1840)
);

CKINVDCx5p33_ASAP7_75t_R g1841 ( 
.A(n_1190),
.Y(n_1841)
);

CKINVDCx5p33_ASAP7_75t_R g1842 ( 
.A(n_812),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_1518),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_986),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_1048),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_639),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_1485),
.Y(n_1847)
);

CKINVDCx5p33_ASAP7_75t_R g1848 ( 
.A(n_1640),
.Y(n_1848)
);

CKINVDCx5p33_ASAP7_75t_R g1849 ( 
.A(n_526),
.Y(n_1849)
);

CKINVDCx20_ASAP7_75t_R g1850 ( 
.A(n_441),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_81),
.Y(n_1851)
);

CKINVDCx5p33_ASAP7_75t_R g1852 ( 
.A(n_551),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_144),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_1607),
.Y(n_1854)
);

BUFx3_ASAP7_75t_L g1855 ( 
.A(n_243),
.Y(n_1855)
);

CKINVDCx5p33_ASAP7_75t_R g1856 ( 
.A(n_1042),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_599),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_223),
.Y(n_1858)
);

CKINVDCx14_ASAP7_75t_R g1859 ( 
.A(n_1520),
.Y(n_1859)
);

BUFx10_ASAP7_75t_L g1860 ( 
.A(n_1673),
.Y(n_1860)
);

CKINVDCx5p33_ASAP7_75t_R g1861 ( 
.A(n_1477),
.Y(n_1861)
);

CKINVDCx5p33_ASAP7_75t_R g1862 ( 
.A(n_109),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_161),
.Y(n_1863)
);

CKINVDCx14_ASAP7_75t_R g1864 ( 
.A(n_153),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_1701),
.Y(n_1865)
);

CKINVDCx5p33_ASAP7_75t_R g1866 ( 
.A(n_1516),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1040),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1588),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_1523),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_550),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_811),
.Y(n_1871)
);

CKINVDCx5p33_ASAP7_75t_R g1872 ( 
.A(n_1526),
.Y(n_1872)
);

BUFx10_ASAP7_75t_L g1873 ( 
.A(n_487),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1245),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1591),
.Y(n_1875)
);

CKINVDCx5p33_ASAP7_75t_R g1876 ( 
.A(n_199),
.Y(n_1876)
);

CKINVDCx5p33_ASAP7_75t_R g1877 ( 
.A(n_1247),
.Y(n_1877)
);

BUFx5_ASAP7_75t_L g1878 ( 
.A(n_1652),
.Y(n_1878)
);

CKINVDCx5p33_ASAP7_75t_R g1879 ( 
.A(n_949),
.Y(n_1879)
);

CKINVDCx20_ASAP7_75t_R g1880 ( 
.A(n_282),
.Y(n_1880)
);

BUFx10_ASAP7_75t_L g1881 ( 
.A(n_1177),
.Y(n_1881)
);

CKINVDCx5p33_ASAP7_75t_R g1882 ( 
.A(n_1445),
.Y(n_1882)
);

CKINVDCx5p33_ASAP7_75t_R g1883 ( 
.A(n_1560),
.Y(n_1883)
);

BUFx5_ASAP7_75t_L g1884 ( 
.A(n_314),
.Y(n_1884)
);

CKINVDCx5p33_ASAP7_75t_R g1885 ( 
.A(n_1598),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1188),
.Y(n_1886)
);

CKINVDCx5p33_ASAP7_75t_R g1887 ( 
.A(n_384),
.Y(n_1887)
);

CKINVDCx5p33_ASAP7_75t_R g1888 ( 
.A(n_1225),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_1436),
.Y(n_1889)
);

CKINVDCx20_ASAP7_75t_R g1890 ( 
.A(n_545),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_1092),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1507),
.Y(n_1892)
);

CKINVDCx16_ASAP7_75t_R g1893 ( 
.A(n_154),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1427),
.Y(n_1894)
);

CKINVDCx5p33_ASAP7_75t_R g1895 ( 
.A(n_1223),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_554),
.Y(n_1896)
);

CKINVDCx5p33_ASAP7_75t_R g1897 ( 
.A(n_1168),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_575),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1228),
.Y(n_1899)
);

CKINVDCx5p33_ASAP7_75t_R g1900 ( 
.A(n_1462),
.Y(n_1900)
);

INVx4_ASAP7_75t_R g1901 ( 
.A(n_401),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_509),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_34),
.Y(n_1903)
);

CKINVDCx5p33_ASAP7_75t_R g1904 ( 
.A(n_1254),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1641),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_1539),
.Y(n_1906)
);

CKINVDCx5p33_ASAP7_75t_R g1907 ( 
.A(n_616),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_1666),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_40),
.Y(n_1909)
);

CKINVDCx5p33_ASAP7_75t_R g1910 ( 
.A(n_45),
.Y(n_1910)
);

CKINVDCx5p33_ASAP7_75t_R g1911 ( 
.A(n_1448),
.Y(n_1911)
);

CKINVDCx20_ASAP7_75t_R g1912 ( 
.A(n_889),
.Y(n_1912)
);

CKINVDCx5p33_ASAP7_75t_R g1913 ( 
.A(n_891),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_988),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_835),
.Y(n_1915)
);

BUFx3_ASAP7_75t_L g1916 ( 
.A(n_81),
.Y(n_1916)
);

CKINVDCx5p33_ASAP7_75t_R g1917 ( 
.A(n_331),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_477),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1095),
.Y(n_1919)
);

CKINVDCx5p33_ASAP7_75t_R g1920 ( 
.A(n_1030),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_1613),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_394),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_97),
.Y(n_1923)
);

CKINVDCx5p33_ASAP7_75t_R g1924 ( 
.A(n_710),
.Y(n_1924)
);

CKINVDCx5p33_ASAP7_75t_R g1925 ( 
.A(n_1420),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_832),
.Y(n_1926)
);

CKINVDCx5p33_ASAP7_75t_R g1927 ( 
.A(n_542),
.Y(n_1927)
);

CKINVDCx20_ASAP7_75t_R g1928 ( 
.A(n_397),
.Y(n_1928)
);

CKINVDCx20_ASAP7_75t_R g1929 ( 
.A(n_1403),
.Y(n_1929)
);

INVx4_ASAP7_75t_R g1930 ( 
.A(n_511),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1452),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_940),
.Y(n_1932)
);

CKINVDCx16_ASAP7_75t_R g1933 ( 
.A(n_1453),
.Y(n_1933)
);

CKINVDCx5p33_ASAP7_75t_R g1934 ( 
.A(n_845),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1017),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_922),
.Y(n_1936)
);

CKINVDCx5p33_ASAP7_75t_R g1937 ( 
.A(n_1237),
.Y(n_1937)
);

CKINVDCx5p33_ASAP7_75t_R g1938 ( 
.A(n_729),
.Y(n_1938)
);

INVx2_ASAP7_75t_SL g1939 ( 
.A(n_281),
.Y(n_1939)
);

CKINVDCx5p33_ASAP7_75t_R g1940 ( 
.A(n_1404),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_663),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_1389),
.Y(n_1942)
);

CKINVDCx5p33_ASAP7_75t_R g1943 ( 
.A(n_955),
.Y(n_1943)
);

CKINVDCx20_ASAP7_75t_R g1944 ( 
.A(n_420),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_533),
.Y(n_1945)
);

CKINVDCx5p33_ASAP7_75t_R g1946 ( 
.A(n_1035),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_178),
.Y(n_1947)
);

CKINVDCx5p33_ASAP7_75t_R g1948 ( 
.A(n_1631),
.Y(n_1948)
);

CKINVDCx5p33_ASAP7_75t_R g1949 ( 
.A(n_1019),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_871),
.Y(n_1950)
);

BUFx3_ASAP7_75t_L g1951 ( 
.A(n_361),
.Y(n_1951)
);

BUFx6f_ASAP7_75t_L g1952 ( 
.A(n_1545),
.Y(n_1952)
);

CKINVDCx5p33_ASAP7_75t_R g1953 ( 
.A(n_116),
.Y(n_1953)
);

CKINVDCx5p33_ASAP7_75t_R g1954 ( 
.A(n_1246),
.Y(n_1954)
);

CKINVDCx5p33_ASAP7_75t_R g1955 ( 
.A(n_1196),
.Y(n_1955)
);

BUFx2_ASAP7_75t_L g1956 ( 
.A(n_1191),
.Y(n_1956)
);

CKINVDCx5p33_ASAP7_75t_R g1957 ( 
.A(n_1426),
.Y(n_1957)
);

CKINVDCx5p33_ASAP7_75t_R g1958 ( 
.A(n_481),
.Y(n_1958)
);

CKINVDCx5p33_ASAP7_75t_R g1959 ( 
.A(n_1551),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1326),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1647),
.Y(n_1961)
);

CKINVDCx16_ASAP7_75t_R g1962 ( 
.A(n_496),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_228),
.Y(n_1963)
);

BUFx6f_ASAP7_75t_L g1964 ( 
.A(n_1156),
.Y(n_1964)
);

CKINVDCx5p33_ASAP7_75t_R g1965 ( 
.A(n_1025),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1173),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_892),
.Y(n_1967)
);

CKINVDCx5p33_ASAP7_75t_R g1968 ( 
.A(n_1205),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_198),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1428),
.Y(n_1970)
);

INVxp67_ASAP7_75t_L g1971 ( 
.A(n_1400),
.Y(n_1971)
);

CKINVDCx5p33_ASAP7_75t_R g1972 ( 
.A(n_836),
.Y(n_1972)
);

CKINVDCx5p33_ASAP7_75t_R g1973 ( 
.A(n_664),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_376),
.Y(n_1974)
);

INVx1_ASAP7_75t_SL g1975 ( 
.A(n_1705),
.Y(n_1975)
);

CKINVDCx5p33_ASAP7_75t_R g1976 ( 
.A(n_1590),
.Y(n_1976)
);

INVxp67_ASAP7_75t_SL g1977 ( 
.A(n_680),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_1568),
.Y(n_1978)
);

CKINVDCx5p33_ASAP7_75t_R g1979 ( 
.A(n_1549),
.Y(n_1979)
);

CKINVDCx5p33_ASAP7_75t_R g1980 ( 
.A(n_1556),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_991),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_209),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1681),
.Y(n_1983)
);

CKINVDCx5p33_ASAP7_75t_R g1984 ( 
.A(n_1522),
.Y(n_1984)
);

CKINVDCx5p33_ASAP7_75t_R g1985 ( 
.A(n_711),
.Y(n_1985)
);

CKINVDCx5p33_ASAP7_75t_R g1986 ( 
.A(n_628),
.Y(n_1986)
);

CKINVDCx5p33_ASAP7_75t_R g1987 ( 
.A(n_883),
.Y(n_1987)
);

CKINVDCx5p33_ASAP7_75t_R g1988 ( 
.A(n_1661),
.Y(n_1988)
);

CKINVDCx5p33_ASAP7_75t_R g1989 ( 
.A(n_1500),
.Y(n_1989)
);

CKINVDCx5p33_ASAP7_75t_R g1990 ( 
.A(n_1689),
.Y(n_1990)
);

BUFx6f_ASAP7_75t_L g1991 ( 
.A(n_97),
.Y(n_1991)
);

CKINVDCx20_ASAP7_75t_R g1992 ( 
.A(n_1208),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_1283),
.Y(n_1993)
);

CKINVDCx20_ASAP7_75t_R g1994 ( 
.A(n_1473),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_949),
.Y(n_1995)
);

INVx1_ASAP7_75t_SL g1996 ( 
.A(n_789),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1464),
.Y(n_1997)
);

INVx4_ASAP7_75t_R g1998 ( 
.A(n_1092),
.Y(n_1998)
);

CKINVDCx5p33_ASAP7_75t_R g1999 ( 
.A(n_1605),
.Y(n_1999)
);

CKINVDCx5p33_ASAP7_75t_R g2000 ( 
.A(n_287),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_190),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_266),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_1119),
.Y(n_2003)
);

CKINVDCx5p33_ASAP7_75t_R g2004 ( 
.A(n_855),
.Y(n_2004)
);

CKINVDCx5p33_ASAP7_75t_R g2005 ( 
.A(n_1087),
.Y(n_2005)
);

CKINVDCx20_ASAP7_75t_R g2006 ( 
.A(n_1650),
.Y(n_2006)
);

CKINVDCx5p33_ASAP7_75t_R g2007 ( 
.A(n_56),
.Y(n_2007)
);

CKINVDCx5p33_ASAP7_75t_R g2008 ( 
.A(n_947),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1638),
.Y(n_2009)
);

CKINVDCx5p33_ASAP7_75t_R g2010 ( 
.A(n_1626),
.Y(n_2010)
);

CKINVDCx5p33_ASAP7_75t_R g2011 ( 
.A(n_788),
.Y(n_2011)
);

CKINVDCx5p33_ASAP7_75t_R g2012 ( 
.A(n_744),
.Y(n_2012)
);

CKINVDCx5p33_ASAP7_75t_R g2013 ( 
.A(n_1524),
.Y(n_2013)
);

CKINVDCx5p33_ASAP7_75t_R g2014 ( 
.A(n_1488),
.Y(n_2014)
);

CKINVDCx5p33_ASAP7_75t_R g2015 ( 
.A(n_1418),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1697),
.Y(n_2016)
);

CKINVDCx20_ASAP7_75t_R g2017 ( 
.A(n_365),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1027),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1684),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1209),
.Y(n_2020)
);

CKINVDCx5p33_ASAP7_75t_R g2021 ( 
.A(n_168),
.Y(n_2021)
);

BUFx6f_ASAP7_75t_L g2022 ( 
.A(n_1421),
.Y(n_2022)
);

CKINVDCx5p33_ASAP7_75t_R g2023 ( 
.A(n_644),
.Y(n_2023)
);

CKINVDCx5p33_ASAP7_75t_R g2024 ( 
.A(n_1699),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_774),
.Y(n_2025)
);

INVx3_ASAP7_75t_L g2026 ( 
.A(n_462),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_374),
.Y(n_2027)
);

INVx2_ASAP7_75t_SL g2028 ( 
.A(n_1297),
.Y(n_2028)
);

INVx1_ASAP7_75t_SL g2029 ( 
.A(n_1627),
.Y(n_2029)
);

CKINVDCx5p33_ASAP7_75t_R g2030 ( 
.A(n_643),
.Y(n_2030)
);

CKINVDCx5p33_ASAP7_75t_R g2031 ( 
.A(n_411),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1628),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_398),
.Y(n_2033)
);

INVx1_ASAP7_75t_SL g2034 ( 
.A(n_712),
.Y(n_2034)
);

CKINVDCx5p33_ASAP7_75t_R g2035 ( 
.A(n_1347),
.Y(n_2035)
);

BUFx6f_ASAP7_75t_L g2036 ( 
.A(n_572),
.Y(n_2036)
);

CKINVDCx5p33_ASAP7_75t_R g2037 ( 
.A(n_1147),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_358),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_179),
.Y(n_2039)
);

CKINVDCx5p33_ASAP7_75t_R g2040 ( 
.A(n_297),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1555),
.Y(n_2041)
);

CKINVDCx5p33_ASAP7_75t_R g2042 ( 
.A(n_665),
.Y(n_2042)
);

CKINVDCx5p33_ASAP7_75t_R g2043 ( 
.A(n_1446),
.Y(n_2043)
);

INVxp67_ASAP7_75t_L g2044 ( 
.A(n_1046),
.Y(n_2044)
);

CKINVDCx5p33_ASAP7_75t_R g2045 ( 
.A(n_155),
.Y(n_2045)
);

CKINVDCx5p33_ASAP7_75t_R g2046 ( 
.A(n_1189),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_382),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1413),
.Y(n_2048)
);

CKINVDCx5p33_ASAP7_75t_R g2049 ( 
.A(n_503),
.Y(n_2049)
);

CKINVDCx5p33_ASAP7_75t_R g2050 ( 
.A(n_430),
.Y(n_2050)
);

CKINVDCx5p33_ASAP7_75t_R g2051 ( 
.A(n_1572),
.Y(n_2051)
);

CKINVDCx5p33_ASAP7_75t_R g2052 ( 
.A(n_1668),
.Y(n_2052)
);

CKINVDCx5p33_ASAP7_75t_R g2053 ( 
.A(n_558),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_104),
.Y(n_2054)
);

CKINVDCx5p33_ASAP7_75t_R g2055 ( 
.A(n_903),
.Y(n_2055)
);

CKINVDCx5p33_ASAP7_75t_R g2056 ( 
.A(n_1558),
.Y(n_2056)
);

BUFx3_ASAP7_75t_L g2057 ( 
.A(n_885),
.Y(n_2057)
);

CKINVDCx5p33_ASAP7_75t_R g2058 ( 
.A(n_115),
.Y(n_2058)
);

CKINVDCx5p33_ASAP7_75t_R g2059 ( 
.A(n_1620),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1199),
.Y(n_2060)
);

CKINVDCx5p33_ASAP7_75t_R g2061 ( 
.A(n_1271),
.Y(n_2061)
);

CKINVDCx5p33_ASAP7_75t_R g2062 ( 
.A(n_1595),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1386),
.Y(n_2063)
);

CKINVDCx5p33_ASAP7_75t_R g2064 ( 
.A(n_271),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1148),
.Y(n_2065)
);

CKINVDCx5p33_ASAP7_75t_R g2066 ( 
.A(n_1309),
.Y(n_2066)
);

CKINVDCx5p33_ASAP7_75t_R g2067 ( 
.A(n_1125),
.Y(n_2067)
);

CKINVDCx5p33_ASAP7_75t_R g2068 ( 
.A(n_337),
.Y(n_2068)
);

CKINVDCx5p33_ASAP7_75t_R g2069 ( 
.A(n_1240),
.Y(n_2069)
);

CKINVDCx5p33_ASAP7_75t_R g2070 ( 
.A(n_562),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1201),
.Y(n_2071)
);

INVxp67_ASAP7_75t_L g2072 ( 
.A(n_1583),
.Y(n_2072)
);

CKINVDCx5p33_ASAP7_75t_R g2073 ( 
.A(n_1055),
.Y(n_2073)
);

CKINVDCx5p33_ASAP7_75t_R g2074 ( 
.A(n_1655),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_975),
.Y(n_2075)
);

INVxp67_ASAP7_75t_L g2076 ( 
.A(n_1041),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_167),
.Y(n_2077)
);

BUFx3_ASAP7_75t_L g2078 ( 
.A(n_1168),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_489),
.Y(n_2079)
);

BUFx10_ASAP7_75t_L g2080 ( 
.A(n_1490),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_475),
.Y(n_2081)
);

CKINVDCx5p33_ASAP7_75t_R g2082 ( 
.A(n_1202),
.Y(n_2082)
);

BUFx2_ASAP7_75t_L g2083 ( 
.A(n_1136),
.Y(n_2083)
);

CKINVDCx5p33_ASAP7_75t_R g2084 ( 
.A(n_1678),
.Y(n_2084)
);

BUFx5_ASAP7_75t_L g2085 ( 
.A(n_1483),
.Y(n_2085)
);

CKINVDCx5p33_ASAP7_75t_R g2086 ( 
.A(n_1541),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1625),
.Y(n_2087)
);

CKINVDCx5p33_ASAP7_75t_R g2088 ( 
.A(n_1471),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_286),
.Y(n_2089)
);

CKINVDCx5p33_ASAP7_75t_R g2090 ( 
.A(n_1314),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1294),
.Y(n_2091)
);

CKINVDCx5p33_ASAP7_75t_R g2092 ( 
.A(n_919),
.Y(n_2092)
);

CKINVDCx5p33_ASAP7_75t_R g2093 ( 
.A(n_1259),
.Y(n_2093)
);

CKINVDCx5p33_ASAP7_75t_R g2094 ( 
.A(n_1683),
.Y(n_2094)
);

CKINVDCx5p33_ASAP7_75t_R g2095 ( 
.A(n_1708),
.Y(n_2095)
);

CKINVDCx5p33_ASAP7_75t_R g2096 ( 
.A(n_1574),
.Y(n_2096)
);

INVxp67_ASAP7_75t_L g2097 ( 
.A(n_1163),
.Y(n_2097)
);

CKINVDCx5p33_ASAP7_75t_R g2098 ( 
.A(n_1457),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_520),
.Y(n_2099)
);

CKINVDCx5p33_ASAP7_75t_R g2100 ( 
.A(n_1120),
.Y(n_2100)
);

CKINVDCx16_ASAP7_75t_R g2101 ( 
.A(n_1142),
.Y(n_2101)
);

BUFx6f_ASAP7_75t_L g2102 ( 
.A(n_1561),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_574),
.Y(n_2103)
);

BUFx10_ASAP7_75t_L g2104 ( 
.A(n_1515),
.Y(n_2104)
);

INVxp33_ASAP7_75t_SL g2105 ( 
.A(n_160),
.Y(n_2105)
);

CKINVDCx5p33_ASAP7_75t_R g2106 ( 
.A(n_393),
.Y(n_2106)
);

INVx1_ASAP7_75t_SL g2107 ( 
.A(n_1063),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_637),
.Y(n_2108)
);

CKINVDCx20_ASAP7_75t_R g2109 ( 
.A(n_289),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_239),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1009),
.Y(n_2111)
);

CKINVDCx5p33_ASAP7_75t_R g2112 ( 
.A(n_1528),
.Y(n_2112)
);

CKINVDCx20_ASAP7_75t_R g2113 ( 
.A(n_346),
.Y(n_2113)
);

CKINVDCx5p33_ASAP7_75t_R g2114 ( 
.A(n_1633),
.Y(n_2114)
);

CKINVDCx5p33_ASAP7_75t_R g2115 ( 
.A(n_1079),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1618),
.Y(n_2116)
);

CKINVDCx5p33_ASAP7_75t_R g2117 ( 
.A(n_950),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1225),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1304),
.Y(n_2119)
);

CKINVDCx5p33_ASAP7_75t_R g2120 ( 
.A(n_928),
.Y(n_2120)
);

CKINVDCx5p33_ASAP7_75t_R g2121 ( 
.A(n_1466),
.Y(n_2121)
);

BUFx2_ASAP7_75t_L g2122 ( 
.A(n_1280),
.Y(n_2122)
);

CKINVDCx5p33_ASAP7_75t_R g2123 ( 
.A(n_95),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_773),
.Y(n_2124)
);

CKINVDCx5p33_ASAP7_75t_R g2125 ( 
.A(n_1119),
.Y(n_2125)
);

CKINVDCx20_ASAP7_75t_R g2126 ( 
.A(n_1621),
.Y(n_2126)
);

CKINVDCx5p33_ASAP7_75t_R g2127 ( 
.A(n_555),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1486),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1467),
.Y(n_2129)
);

CKINVDCx5p33_ASAP7_75t_R g2130 ( 
.A(n_338),
.Y(n_2130)
);

CKINVDCx5p33_ASAP7_75t_R g2131 ( 
.A(n_715),
.Y(n_2131)
);

CKINVDCx5p33_ASAP7_75t_R g2132 ( 
.A(n_1614),
.Y(n_2132)
);

CKINVDCx5p33_ASAP7_75t_R g2133 ( 
.A(n_192),
.Y(n_2133)
);

CKINVDCx5p33_ASAP7_75t_R g2134 ( 
.A(n_450),
.Y(n_2134)
);

CKINVDCx5p33_ASAP7_75t_R g2135 ( 
.A(n_1257),
.Y(n_2135)
);

CKINVDCx5p33_ASAP7_75t_R g2136 ( 
.A(n_671),
.Y(n_2136)
);

CKINVDCx5p33_ASAP7_75t_R g2137 ( 
.A(n_827),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1601),
.Y(n_2138)
);

CKINVDCx5p33_ASAP7_75t_R g2139 ( 
.A(n_1557),
.Y(n_2139)
);

CKINVDCx5p33_ASAP7_75t_R g2140 ( 
.A(n_1510),
.Y(n_2140)
);

CKINVDCx20_ASAP7_75t_R g2141 ( 
.A(n_1264),
.Y(n_2141)
);

CKINVDCx5p33_ASAP7_75t_R g2142 ( 
.A(n_58),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_154),
.Y(n_2143)
);

BUFx2_ASAP7_75t_L g2144 ( 
.A(n_1529),
.Y(n_2144)
);

CKINVDCx5p33_ASAP7_75t_R g2145 ( 
.A(n_1180),
.Y(n_2145)
);

CKINVDCx5p33_ASAP7_75t_R g2146 ( 
.A(n_634),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_782),
.Y(n_2147)
);

BUFx2_ASAP7_75t_L g2148 ( 
.A(n_833),
.Y(n_2148)
);

CKINVDCx5p33_ASAP7_75t_R g2149 ( 
.A(n_551),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_196),
.Y(n_2150)
);

CKINVDCx5p33_ASAP7_75t_R g2151 ( 
.A(n_721),
.Y(n_2151)
);

CKINVDCx5p33_ASAP7_75t_R g2152 ( 
.A(n_1069),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_250),
.Y(n_2153)
);

CKINVDCx5p33_ASAP7_75t_R g2154 ( 
.A(n_1656),
.Y(n_2154)
);

CKINVDCx5p33_ASAP7_75t_R g2155 ( 
.A(n_1552),
.Y(n_2155)
);

CKINVDCx5p33_ASAP7_75t_R g2156 ( 
.A(n_679),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_14),
.Y(n_2157)
);

CKINVDCx5p33_ASAP7_75t_R g2158 ( 
.A(n_943),
.Y(n_2158)
);

CKINVDCx16_ASAP7_75t_R g2159 ( 
.A(n_1214),
.Y(n_2159)
);

CKINVDCx5p33_ASAP7_75t_R g2160 ( 
.A(n_696),
.Y(n_2160)
);

CKINVDCx5p33_ASAP7_75t_R g2161 ( 
.A(n_213),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1612),
.Y(n_2162)
);

CKINVDCx5p33_ASAP7_75t_R g2163 ( 
.A(n_429),
.Y(n_2163)
);

CKINVDCx5p33_ASAP7_75t_R g2164 ( 
.A(n_1672),
.Y(n_2164)
);

CKINVDCx5p33_ASAP7_75t_R g2165 ( 
.A(n_1694),
.Y(n_2165)
);

CKINVDCx5p33_ASAP7_75t_R g2166 ( 
.A(n_303),
.Y(n_2166)
);

CKINVDCx5p33_ASAP7_75t_R g2167 ( 
.A(n_215),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_943),
.Y(n_2168)
);

CKINVDCx5p33_ASAP7_75t_R g2169 ( 
.A(n_1182),
.Y(n_2169)
);

CKINVDCx5p33_ASAP7_75t_R g2170 ( 
.A(n_1380),
.Y(n_2170)
);

INVx2_ASAP7_75t_SL g2171 ( 
.A(n_779),
.Y(n_2171)
);

CKINVDCx5p33_ASAP7_75t_R g2172 ( 
.A(n_590),
.Y(n_2172)
);

CKINVDCx5p33_ASAP7_75t_R g2173 ( 
.A(n_1540),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_564),
.Y(n_2174)
);

CKINVDCx5p33_ASAP7_75t_R g2175 ( 
.A(n_1393),
.Y(n_2175)
);

CKINVDCx5p33_ASAP7_75t_R g2176 ( 
.A(n_1209),
.Y(n_2176)
);

CKINVDCx5p33_ASAP7_75t_R g2177 ( 
.A(n_1489),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_690),
.Y(n_2178)
);

BUFx10_ASAP7_75t_L g2179 ( 
.A(n_354),
.Y(n_2179)
);

INVxp67_ASAP7_75t_L g2180 ( 
.A(n_629),
.Y(n_2180)
);

CKINVDCx5p33_ASAP7_75t_R g2181 ( 
.A(n_1222),
.Y(n_2181)
);

CKINVDCx5p33_ASAP7_75t_R g2182 ( 
.A(n_922),
.Y(n_2182)
);

BUFx3_ASAP7_75t_L g2183 ( 
.A(n_904),
.Y(n_2183)
);

BUFx5_ASAP7_75t_L g2184 ( 
.A(n_1455),
.Y(n_2184)
);

CKINVDCx5p33_ASAP7_75t_R g2185 ( 
.A(n_967),
.Y(n_2185)
);

CKINVDCx20_ASAP7_75t_R g2186 ( 
.A(n_273),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_784),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_367),
.Y(n_2188)
);

CKINVDCx5p33_ASAP7_75t_R g2189 ( 
.A(n_1573),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_885),
.Y(n_2190)
);

CKINVDCx5p33_ASAP7_75t_R g2191 ( 
.A(n_271),
.Y(n_2191)
);

CKINVDCx5p33_ASAP7_75t_R g2192 ( 
.A(n_1513),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_182),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_908),
.Y(n_2194)
);

CKINVDCx5p33_ASAP7_75t_R g2195 ( 
.A(n_292),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_443),
.Y(n_2196)
);

CKINVDCx5p33_ASAP7_75t_R g2197 ( 
.A(n_675),
.Y(n_2197)
);

CKINVDCx5p33_ASAP7_75t_R g2198 ( 
.A(n_716),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_857),
.Y(n_2199)
);

CKINVDCx5p33_ASAP7_75t_R g2200 ( 
.A(n_1387),
.Y(n_2200)
);

CKINVDCx5p33_ASAP7_75t_R g2201 ( 
.A(n_698),
.Y(n_2201)
);

CKINVDCx5p33_ASAP7_75t_R g2202 ( 
.A(n_1504),
.Y(n_2202)
);

CKINVDCx5p33_ASAP7_75t_R g2203 ( 
.A(n_565),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1481),
.Y(n_2204)
);

CKINVDCx5p33_ASAP7_75t_R g2205 ( 
.A(n_1210),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_275),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_262),
.Y(n_2207)
);

BUFx3_ASAP7_75t_L g2208 ( 
.A(n_1703),
.Y(n_2208)
);

CKINVDCx20_ASAP7_75t_R g2209 ( 
.A(n_45),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1311),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_483),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1417),
.Y(n_2212)
);

CKINVDCx5p33_ASAP7_75t_R g2213 ( 
.A(n_444),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_283),
.Y(n_2214)
);

CKINVDCx5p33_ASAP7_75t_R g2215 ( 
.A(n_1498),
.Y(n_2215)
);

CKINVDCx5p33_ASAP7_75t_R g2216 ( 
.A(n_1330),
.Y(n_2216)
);

INVx2_ASAP7_75t_SL g2217 ( 
.A(n_1098),
.Y(n_2217)
);

CKINVDCx5p33_ASAP7_75t_R g2218 ( 
.A(n_870),
.Y(n_2218)
);

CKINVDCx20_ASAP7_75t_R g2219 ( 
.A(n_1459),
.Y(n_2219)
);

CKINVDCx5p33_ASAP7_75t_R g2220 ( 
.A(n_1048),
.Y(n_2220)
);

CKINVDCx5p33_ASAP7_75t_R g2221 ( 
.A(n_1476),
.Y(n_2221)
);

CKINVDCx5p33_ASAP7_75t_R g2222 ( 
.A(n_778),
.Y(n_2222)
);

CKINVDCx5p33_ASAP7_75t_R g2223 ( 
.A(n_1439),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1559),
.Y(n_2224)
);

CKINVDCx5p33_ASAP7_75t_R g2225 ( 
.A(n_1116),
.Y(n_2225)
);

INVx3_ASAP7_75t_L g2226 ( 
.A(n_1352),
.Y(n_2226)
);

CKINVDCx5p33_ASAP7_75t_R g2227 ( 
.A(n_894),
.Y(n_2227)
);

CKINVDCx5p33_ASAP7_75t_R g2228 ( 
.A(n_807),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_839),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1095),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_770),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1450),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_742),
.Y(n_2233)
);

CKINVDCx5p33_ASAP7_75t_R g2234 ( 
.A(n_275),
.Y(n_2234)
);

CKINVDCx5p33_ASAP7_75t_R g2235 ( 
.A(n_1044),
.Y(n_2235)
);

CKINVDCx5p33_ASAP7_75t_R g2236 ( 
.A(n_772),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_122),
.Y(n_2237)
);

CKINVDCx5p33_ASAP7_75t_R g2238 ( 
.A(n_1685),
.Y(n_2238)
);

CKINVDCx5p33_ASAP7_75t_R g2239 ( 
.A(n_423),
.Y(n_2239)
);

INVx2_ASAP7_75t_SL g2240 ( 
.A(n_1097),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1171),
.Y(n_2241)
);

CKINVDCx5p33_ASAP7_75t_R g2242 ( 
.A(n_76),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_844),
.Y(n_2243)
);

CKINVDCx5p33_ASAP7_75t_R g2244 ( 
.A(n_1074),
.Y(n_2244)
);

CKINVDCx5p33_ASAP7_75t_R g2245 ( 
.A(n_19),
.Y(n_2245)
);

CKINVDCx5p33_ASAP7_75t_R g2246 ( 
.A(n_792),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1527),
.Y(n_2247)
);

CKINVDCx5p33_ASAP7_75t_R g2248 ( 
.A(n_1435),
.Y(n_2248)
);

CKINVDCx20_ASAP7_75t_R g2249 ( 
.A(n_353),
.Y(n_2249)
);

CKINVDCx20_ASAP7_75t_R g2250 ( 
.A(n_220),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_526),
.Y(n_2251)
);

CKINVDCx5p33_ASAP7_75t_R g2252 ( 
.A(n_1525),
.Y(n_2252)
);

INVx2_ASAP7_75t_SL g2253 ( 
.A(n_582),
.Y(n_2253)
);

CKINVDCx5p33_ASAP7_75t_R g2254 ( 
.A(n_1370),
.Y(n_2254)
);

CKINVDCx5p33_ASAP7_75t_R g2255 ( 
.A(n_1281),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1609),
.Y(n_2256)
);

CKINVDCx5p33_ASAP7_75t_R g2257 ( 
.A(n_1312),
.Y(n_2257)
);

CKINVDCx5p33_ASAP7_75t_R g2258 ( 
.A(n_1135),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_437),
.Y(n_2259)
);

INVx1_ASAP7_75t_SL g2260 ( 
.A(n_1047),
.Y(n_2260)
);

CKINVDCx5p33_ASAP7_75t_R g2261 ( 
.A(n_17),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_365),
.Y(n_2262)
);

CKINVDCx20_ASAP7_75t_R g2263 ( 
.A(n_807),
.Y(n_2263)
);

CKINVDCx5p33_ASAP7_75t_R g2264 ( 
.A(n_963),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_1170),
.Y(n_2265)
);

BUFx8_ASAP7_75t_SL g2266 ( 
.A(n_672),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1437),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1567),
.Y(n_2268)
);

CKINVDCx5p33_ASAP7_75t_R g2269 ( 
.A(n_1084),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_1503),
.Y(n_2270)
);

CKINVDCx5p33_ASAP7_75t_R g2271 ( 
.A(n_1128),
.Y(n_2271)
);

CKINVDCx20_ASAP7_75t_R g2272 ( 
.A(n_1041),
.Y(n_2272)
);

CKINVDCx5p33_ASAP7_75t_R g2273 ( 
.A(n_951),
.Y(n_2273)
);

CKINVDCx20_ASAP7_75t_R g2274 ( 
.A(n_1335),
.Y(n_2274)
);

CKINVDCx5p33_ASAP7_75t_R g2275 ( 
.A(n_1021),
.Y(n_2275)
);

CKINVDCx5p33_ASAP7_75t_R g2276 ( 
.A(n_1565),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_1606),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1669),
.Y(n_2278)
);

CKINVDCx20_ASAP7_75t_R g2279 ( 
.A(n_854),
.Y(n_2279)
);

CKINVDCx5p33_ASAP7_75t_R g2280 ( 
.A(n_446),
.Y(n_2280)
);

CKINVDCx20_ASAP7_75t_R g2281 ( 
.A(n_57),
.Y(n_2281)
);

BUFx8_ASAP7_75t_SL g2282 ( 
.A(n_1665),
.Y(n_2282)
);

CKINVDCx5p33_ASAP7_75t_R g2283 ( 
.A(n_1022),
.Y(n_2283)
);

CKINVDCx5p33_ASAP7_75t_R g2284 ( 
.A(n_879),
.Y(n_2284)
);

CKINVDCx5p33_ASAP7_75t_R g2285 ( 
.A(n_846),
.Y(n_2285)
);

CKINVDCx5p33_ASAP7_75t_R g2286 ( 
.A(n_1193),
.Y(n_2286)
);

CKINVDCx5p33_ASAP7_75t_R g2287 ( 
.A(n_1088),
.Y(n_2287)
);

CKINVDCx5p33_ASAP7_75t_R g2288 ( 
.A(n_1198),
.Y(n_2288)
);

BUFx6f_ASAP7_75t_L g2289 ( 
.A(n_1082),
.Y(n_2289)
);

INVx2_ASAP7_75t_SL g2290 ( 
.A(n_1206),
.Y(n_2290)
);

CKINVDCx5p33_ASAP7_75t_R g2291 ( 
.A(n_579),
.Y(n_2291)
);

CKINVDCx5p33_ASAP7_75t_R g2292 ( 
.A(n_36),
.Y(n_2292)
);

CKINVDCx5p33_ASAP7_75t_R g2293 ( 
.A(n_942),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_1581),
.Y(n_2294)
);

INVx1_ASAP7_75t_SL g2295 ( 
.A(n_1682),
.Y(n_2295)
);

CKINVDCx5p33_ASAP7_75t_R g2296 ( 
.A(n_240),
.Y(n_2296)
);

CKINVDCx5p33_ASAP7_75t_R g2297 ( 
.A(n_1251),
.Y(n_2297)
);

CKINVDCx5p33_ASAP7_75t_R g2298 ( 
.A(n_1480),
.Y(n_2298)
);

HB1xp67_ASAP7_75t_L g2299 ( 
.A(n_1569),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_507),
.Y(n_2300)
);

BUFx10_ASAP7_75t_L g2301 ( 
.A(n_1047),
.Y(n_2301)
);

CKINVDCx5p33_ASAP7_75t_R g2302 ( 
.A(n_1217),
.Y(n_2302)
);

CKINVDCx5p33_ASAP7_75t_R g2303 ( 
.A(n_706),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_1570),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_1706),
.Y(n_2305)
);

CKINVDCx5p33_ASAP7_75t_R g2306 ( 
.A(n_613),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_1461),
.Y(n_2307)
);

INVx1_ASAP7_75t_SL g2308 ( 
.A(n_1663),
.Y(n_2308)
);

CKINVDCx5p33_ASAP7_75t_R g2309 ( 
.A(n_566),
.Y(n_2309)
);

CKINVDCx5p33_ASAP7_75t_R g2310 ( 
.A(n_401),
.Y(n_2310)
);

CKINVDCx5p33_ASAP7_75t_R g2311 ( 
.A(n_1186),
.Y(n_2311)
);

BUFx10_ASAP7_75t_L g2312 ( 
.A(n_190),
.Y(n_2312)
);

CKINVDCx20_ASAP7_75t_R g2313 ( 
.A(n_306),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_1636),
.Y(n_2314)
);

CKINVDCx5p33_ASAP7_75t_R g2315 ( 
.A(n_89),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_1132),
.Y(n_2316)
);

CKINVDCx5p33_ASAP7_75t_R g2317 ( 
.A(n_1564),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_1644),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_151),
.Y(n_2319)
);

CKINVDCx5p33_ASAP7_75t_R g2320 ( 
.A(n_667),
.Y(n_2320)
);

CKINVDCx20_ASAP7_75t_R g2321 ( 
.A(n_115),
.Y(n_2321)
);

CKINVDCx20_ASAP7_75t_R g2322 ( 
.A(n_1440),
.Y(n_2322)
);

CKINVDCx5p33_ASAP7_75t_R g2323 ( 
.A(n_803),
.Y(n_2323)
);

INVx2_ASAP7_75t_SL g2324 ( 
.A(n_407),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_1229),
.Y(n_2325)
);

CKINVDCx20_ASAP7_75t_R g2326 ( 
.A(n_1128),
.Y(n_2326)
);

CKINVDCx5p33_ASAP7_75t_R g2327 ( 
.A(n_1456),
.Y(n_2327)
);

CKINVDCx20_ASAP7_75t_R g2328 ( 
.A(n_643),
.Y(n_2328)
);

CKINVDCx5p33_ASAP7_75t_R g2329 ( 
.A(n_1349),
.Y(n_2329)
);

INVx2_ASAP7_75t_SL g2330 ( 
.A(n_1676),
.Y(n_2330)
);

HB1xp67_ASAP7_75t_L g2331 ( 
.A(n_1216),
.Y(n_2331)
);

CKINVDCx5p33_ASAP7_75t_R g2332 ( 
.A(n_1548),
.Y(n_2332)
);

CKINVDCx5p33_ASAP7_75t_R g2333 ( 
.A(n_1175),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_581),
.Y(n_2334)
);

CKINVDCx5p33_ASAP7_75t_R g2335 ( 
.A(n_867),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_1508),
.Y(n_2336)
);

CKINVDCx5p33_ASAP7_75t_R g2337 ( 
.A(n_1063),
.Y(n_2337)
);

CKINVDCx5p33_ASAP7_75t_R g2338 ( 
.A(n_1664),
.Y(n_2338)
);

CKINVDCx20_ASAP7_75t_R g2339 ( 
.A(n_797),
.Y(n_2339)
);

INVx1_ASAP7_75t_SL g2340 ( 
.A(n_597),
.Y(n_2340)
);

CKINVDCx5p33_ASAP7_75t_R g2341 ( 
.A(n_118),
.Y(n_2341)
);

CKINVDCx5p33_ASAP7_75t_R g2342 ( 
.A(n_264),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_408),
.Y(n_2343)
);

CKINVDCx5p33_ASAP7_75t_R g2344 ( 
.A(n_1343),
.Y(n_2344)
);

CKINVDCx5p33_ASAP7_75t_R g2345 ( 
.A(n_372),
.Y(n_2345)
);

CKINVDCx5p33_ASAP7_75t_R g2346 ( 
.A(n_1180),
.Y(n_2346)
);

CKINVDCx5p33_ASAP7_75t_R g2347 ( 
.A(n_214),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_1025),
.Y(n_2348)
);

BUFx3_ASAP7_75t_L g2349 ( 
.A(n_1337),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_1492),
.Y(n_2350)
);

HB1xp67_ASAP7_75t_L g2351 ( 
.A(n_820),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_1057),
.Y(n_2352)
);

INVx1_ASAP7_75t_SL g2353 ( 
.A(n_1161),
.Y(n_2353)
);

CKINVDCx5p33_ASAP7_75t_R g2354 ( 
.A(n_608),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_773),
.Y(n_2355)
);

CKINVDCx5p33_ASAP7_75t_R g2356 ( 
.A(n_214),
.Y(n_2356)
);

CKINVDCx5p33_ASAP7_75t_R g2357 ( 
.A(n_1067),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_1224),
.Y(n_2358)
);

CKINVDCx5p33_ASAP7_75t_R g2359 ( 
.A(n_187),
.Y(n_2359)
);

CKINVDCx5p33_ASAP7_75t_R g2360 ( 
.A(n_1635),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_322),
.Y(n_2361)
);

INVx2_ASAP7_75t_SL g2362 ( 
.A(n_1321),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_515),
.Y(n_2363)
);

CKINVDCx5p33_ASAP7_75t_R g2364 ( 
.A(n_626),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_524),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_811),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_1429),
.Y(n_2367)
);

CKINVDCx16_ASAP7_75t_R g2368 ( 
.A(n_368),
.Y(n_2368)
);

CKINVDCx5p33_ASAP7_75t_R g2369 ( 
.A(n_157),
.Y(n_2369)
);

CKINVDCx5p33_ASAP7_75t_R g2370 ( 
.A(n_928),
.Y(n_2370)
);

CKINVDCx5p33_ASAP7_75t_R g2371 ( 
.A(n_801),
.Y(n_2371)
);

BUFx3_ASAP7_75t_L g2372 ( 
.A(n_1307),
.Y(n_2372)
);

CKINVDCx5p33_ASAP7_75t_R g2373 ( 
.A(n_585),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_900),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_926),
.Y(n_2375)
);

CKINVDCx5p33_ASAP7_75t_R g2376 ( 
.A(n_441),
.Y(n_2376)
);

CKINVDCx5p33_ASAP7_75t_R g2377 ( 
.A(n_1454),
.Y(n_2377)
);

CKINVDCx5p33_ASAP7_75t_R g2378 ( 
.A(n_1662),
.Y(n_2378)
);

CKINVDCx5p33_ASAP7_75t_R g2379 ( 
.A(n_876),
.Y(n_2379)
);

INVx1_ASAP7_75t_SL g2380 ( 
.A(n_153),
.Y(n_2380)
);

CKINVDCx5p33_ASAP7_75t_R g2381 ( 
.A(n_1585),
.Y(n_2381)
);

CKINVDCx5p33_ASAP7_75t_R g2382 ( 
.A(n_545),
.Y(n_2382)
);

CKINVDCx5p33_ASAP7_75t_R g2383 ( 
.A(n_55),
.Y(n_2383)
);

CKINVDCx5p33_ASAP7_75t_R g2384 ( 
.A(n_1692),
.Y(n_2384)
);

CKINVDCx5p33_ASAP7_75t_R g2385 ( 
.A(n_1475),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_314),
.Y(n_2386)
);

CKINVDCx5p33_ASAP7_75t_R g2387 ( 
.A(n_281),
.Y(n_2387)
);

CKINVDCx20_ASAP7_75t_R g2388 ( 
.A(n_1208),
.Y(n_2388)
);

CKINVDCx5p33_ASAP7_75t_R g2389 ( 
.A(n_682),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_961),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_462),
.Y(n_2391)
);

BUFx2_ASAP7_75t_L g2392 ( 
.A(n_999),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_1632),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_1537),
.Y(n_2394)
);

CKINVDCx20_ASAP7_75t_R g2395 ( 
.A(n_700),
.Y(n_2395)
);

INVx1_ASAP7_75t_SL g2396 ( 
.A(n_1546),
.Y(n_2396)
);

CKINVDCx5p33_ASAP7_75t_R g2397 ( 
.A(n_524),
.Y(n_2397)
);

CKINVDCx5p33_ASAP7_75t_R g2398 ( 
.A(n_1123),
.Y(n_2398)
);

BUFx2_ASAP7_75t_SL g2399 ( 
.A(n_336),
.Y(n_2399)
);

CKINVDCx5p33_ASAP7_75t_R g2400 ( 
.A(n_210),
.Y(n_2400)
);

CKINVDCx5p33_ASAP7_75t_R g2401 ( 
.A(n_531),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_267),
.Y(n_2402)
);

CKINVDCx20_ASAP7_75t_R g2403 ( 
.A(n_1374),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_552),
.Y(n_2404)
);

BUFx3_ASAP7_75t_L g2405 ( 
.A(n_1691),
.Y(n_2405)
);

INVx1_ASAP7_75t_SL g2406 ( 
.A(n_484),
.Y(n_2406)
);

CKINVDCx5p33_ASAP7_75t_R g2407 ( 
.A(n_1176),
.Y(n_2407)
);

INVx2_ASAP7_75t_SL g2408 ( 
.A(n_929),
.Y(n_2408)
);

BUFx10_ASAP7_75t_L g2409 ( 
.A(n_1230),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_1278),
.Y(n_2410)
);

CKINVDCx5p33_ASAP7_75t_R g2411 ( 
.A(n_721),
.Y(n_2411)
);

CKINVDCx5p33_ASAP7_75t_R g2412 ( 
.A(n_1213),
.Y(n_2412)
);

CKINVDCx5p33_ASAP7_75t_R g2413 ( 
.A(n_803),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_240),
.Y(n_2414)
);

HB1xp67_ASAP7_75t_L g2415 ( 
.A(n_463),
.Y(n_2415)
);

INVx2_ASAP7_75t_L g2416 ( 
.A(n_1069),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_991),
.Y(n_2417)
);

CKINVDCx5p33_ASAP7_75t_R g2418 ( 
.A(n_1291),
.Y(n_2418)
);

CKINVDCx5p33_ASAP7_75t_R g2419 ( 
.A(n_1449),
.Y(n_2419)
);

CKINVDCx5p33_ASAP7_75t_R g2420 ( 
.A(n_999),
.Y(n_2420)
);

CKINVDCx5p33_ASAP7_75t_R g2421 ( 
.A(n_1509),
.Y(n_2421)
);

CKINVDCx5p33_ASAP7_75t_R g2422 ( 
.A(n_764),
.Y(n_2422)
);

CKINVDCx20_ASAP7_75t_R g2423 ( 
.A(n_1178),
.Y(n_2423)
);

CKINVDCx5p33_ASAP7_75t_R g2424 ( 
.A(n_768),
.Y(n_2424)
);

CKINVDCx5p33_ASAP7_75t_R g2425 ( 
.A(n_369),
.Y(n_2425)
);

CKINVDCx5p33_ASAP7_75t_R g2426 ( 
.A(n_470),
.Y(n_2426)
);

CKINVDCx16_ASAP7_75t_R g2427 ( 
.A(n_200),
.Y(n_2427)
);

CKINVDCx5p33_ASAP7_75t_R g2428 ( 
.A(n_670),
.Y(n_2428)
);

CKINVDCx5p33_ASAP7_75t_R g2429 ( 
.A(n_1014),
.Y(n_2429)
);

INVx2_ASAP7_75t_L g2430 ( 
.A(n_56),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_873),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_1014),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_951),
.Y(n_2433)
);

INVx2_ASAP7_75t_SL g2434 ( 
.A(n_1502),
.Y(n_2434)
);

CKINVDCx5p33_ASAP7_75t_R g2435 ( 
.A(n_1423),
.Y(n_2435)
);

CKINVDCx5p33_ASAP7_75t_R g2436 ( 
.A(n_1519),
.Y(n_2436)
);

CKINVDCx5p33_ASAP7_75t_R g2437 ( 
.A(n_1185),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_732),
.Y(n_2438)
);

BUFx5_ASAP7_75t_L g2439 ( 
.A(n_704),
.Y(n_2439)
);

BUFx10_ASAP7_75t_L g2440 ( 
.A(n_960),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_1183),
.Y(n_2441)
);

CKINVDCx20_ASAP7_75t_R g2442 ( 
.A(n_859),
.Y(n_2442)
);

CKINVDCx5p33_ASAP7_75t_R g2443 ( 
.A(n_1535),
.Y(n_2443)
);

CKINVDCx5p33_ASAP7_75t_R g2444 ( 
.A(n_1704),
.Y(n_2444)
);

INVx1_ASAP7_75t_SL g2445 ( 
.A(n_1110),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_43),
.Y(n_2446)
);

CKINVDCx5p33_ASAP7_75t_R g2447 ( 
.A(n_635),
.Y(n_2447)
);

CKINVDCx5p33_ASAP7_75t_R g2448 ( 
.A(n_146),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_264),
.Y(n_2449)
);

BUFx2_ASAP7_75t_L g2450 ( 
.A(n_1194),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_444),
.Y(n_2451)
);

CKINVDCx5p33_ASAP7_75t_R g2452 ( 
.A(n_583),
.Y(n_2452)
);

CKINVDCx14_ASAP7_75t_R g2453 ( 
.A(n_1596),
.Y(n_2453)
);

BUFx10_ASAP7_75t_L g2454 ( 
.A(n_1629),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_1339),
.Y(n_2455)
);

CKINVDCx5p33_ASAP7_75t_R g2456 ( 
.A(n_491),
.Y(n_2456)
);

CKINVDCx5p33_ASAP7_75t_R g2457 ( 
.A(n_812),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_776),
.Y(n_2458)
);

CKINVDCx5p33_ASAP7_75t_R g2459 ( 
.A(n_1198),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_485),
.Y(n_2460)
);

CKINVDCx20_ASAP7_75t_R g2461 ( 
.A(n_1114),
.Y(n_2461)
);

CKINVDCx5p33_ASAP7_75t_R g2462 ( 
.A(n_1506),
.Y(n_2462)
);

CKINVDCx5p33_ASAP7_75t_R g2463 ( 
.A(n_913),
.Y(n_2463)
);

BUFx5_ASAP7_75t_L g2464 ( 
.A(n_910),
.Y(n_2464)
);

CKINVDCx5p33_ASAP7_75t_R g2465 ( 
.A(n_1686),
.Y(n_2465)
);

CKINVDCx5p33_ASAP7_75t_R g2466 ( 
.A(n_173),
.Y(n_2466)
);

CKINVDCx5p33_ASAP7_75t_R g2467 ( 
.A(n_1144),
.Y(n_2467)
);

CKINVDCx5p33_ASAP7_75t_R g2468 ( 
.A(n_1487),
.Y(n_2468)
);

CKINVDCx5p33_ASAP7_75t_R g2469 ( 
.A(n_1419),
.Y(n_2469)
);

CKINVDCx20_ASAP7_75t_R g2470 ( 
.A(n_1217),
.Y(n_2470)
);

CKINVDCx20_ASAP7_75t_R g2471 ( 
.A(n_947),
.Y(n_2471)
);

HB1xp67_ASAP7_75t_L g2472 ( 
.A(n_1004),
.Y(n_2472)
);

BUFx2_ASAP7_75t_SL g2473 ( 
.A(n_499),
.Y(n_2473)
);

CKINVDCx5p33_ASAP7_75t_R g2474 ( 
.A(n_1600),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_1070),
.Y(n_2475)
);

INVx2_ASAP7_75t_SL g2476 ( 
.A(n_418),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_480),
.Y(n_2477)
);

CKINVDCx5p33_ASAP7_75t_R g2478 ( 
.A(n_964),
.Y(n_2478)
);

BUFx6f_ASAP7_75t_L g2479 ( 
.A(n_1639),
.Y(n_2479)
);

CKINVDCx5p33_ASAP7_75t_R g2480 ( 
.A(n_252),
.Y(n_2480)
);

CKINVDCx5p33_ASAP7_75t_R g2481 ( 
.A(n_1425),
.Y(n_2481)
);

BUFx6f_ASAP7_75t_L g2482 ( 
.A(n_1687),
.Y(n_2482)
);

CKINVDCx5p33_ASAP7_75t_R g2483 ( 
.A(n_1218),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_1434),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_135),
.Y(n_2485)
);

CKINVDCx5p33_ASAP7_75t_R g2486 ( 
.A(n_405),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_699),
.Y(n_2487)
);

CKINVDCx5p33_ASAP7_75t_R g2488 ( 
.A(n_367),
.Y(n_2488)
);

CKINVDCx20_ASAP7_75t_R g2489 ( 
.A(n_1521),
.Y(n_2489)
);

CKINVDCx20_ASAP7_75t_R g2490 ( 
.A(n_1091),
.Y(n_2490)
);

CKINVDCx5p33_ASAP7_75t_R g2491 ( 
.A(n_1478),
.Y(n_2491)
);

INVx1_ASAP7_75t_SL g2492 ( 
.A(n_460),
.Y(n_2492)
);

CKINVDCx5p33_ASAP7_75t_R g2493 ( 
.A(n_1562),
.Y(n_2493)
);

CKINVDCx5p33_ASAP7_75t_R g2494 ( 
.A(n_1215),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_1012),
.Y(n_2495)
);

CKINVDCx5p33_ASAP7_75t_R g2496 ( 
.A(n_1497),
.Y(n_2496)
);

CKINVDCx20_ASAP7_75t_R g2497 ( 
.A(n_1532),
.Y(n_2497)
);

BUFx10_ASAP7_75t_L g2498 ( 
.A(n_809),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_556),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_1336),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_1538),
.Y(n_2501)
);

CKINVDCx20_ASAP7_75t_R g2502 ( 
.A(n_303),
.Y(n_2502)
);

CKINVDCx5p33_ASAP7_75t_R g2503 ( 
.A(n_555),
.Y(n_2503)
);

CKINVDCx5p33_ASAP7_75t_R g2504 ( 
.A(n_1220),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_776),
.Y(n_2505)
);

CKINVDCx5p33_ASAP7_75t_R g2506 ( 
.A(n_209),
.Y(n_2506)
);

CKINVDCx5p33_ASAP7_75t_R g2507 ( 
.A(n_1170),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_1594),
.Y(n_2508)
);

CKINVDCx5p33_ASAP7_75t_R g2509 ( 
.A(n_1611),
.Y(n_2509)
);

CKINVDCx5p33_ASAP7_75t_R g2510 ( 
.A(n_1648),
.Y(n_2510)
);

INVx1_ASAP7_75t_SL g2511 ( 
.A(n_860),
.Y(n_2511)
);

CKINVDCx5p33_ASAP7_75t_R g2512 ( 
.A(n_111),
.Y(n_2512)
);

CKINVDCx20_ASAP7_75t_R g2513 ( 
.A(n_106),
.Y(n_2513)
);

BUFx3_ASAP7_75t_L g2514 ( 
.A(n_489),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_1479),
.Y(n_2515)
);

INVx1_ASAP7_75t_SL g2516 ( 
.A(n_1252),
.Y(n_2516)
);

CKINVDCx5p33_ASAP7_75t_R g2517 ( 
.A(n_929),
.Y(n_2517)
);

CKINVDCx5p33_ASAP7_75t_R g2518 ( 
.A(n_794),
.Y(n_2518)
);

CKINVDCx20_ASAP7_75t_R g2519 ( 
.A(n_378),
.Y(n_2519)
);

CKINVDCx5p33_ASAP7_75t_R g2520 ( 
.A(n_783),
.Y(n_2520)
);

CKINVDCx5p33_ASAP7_75t_R g2521 ( 
.A(n_958),
.Y(n_2521)
);

CKINVDCx5p33_ASAP7_75t_R g2522 ( 
.A(n_341),
.Y(n_2522)
);

CKINVDCx20_ASAP7_75t_R g2523 ( 
.A(n_1642),
.Y(n_2523)
);

INVx2_ASAP7_75t_L g2524 ( 
.A(n_636),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_766),
.Y(n_2525)
);

CKINVDCx5p33_ASAP7_75t_R g2526 ( 
.A(n_1677),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_1181),
.Y(n_2527)
);

CKINVDCx5p33_ASAP7_75t_R g2528 ( 
.A(n_1250),
.Y(n_2528)
);

CKINVDCx5p33_ASAP7_75t_R g2529 ( 
.A(n_1514),
.Y(n_2529)
);

CKINVDCx5p33_ASAP7_75t_R g2530 ( 
.A(n_35),
.Y(n_2530)
);

INVx1_ASAP7_75t_SL g2531 ( 
.A(n_1215),
.Y(n_2531)
);

INVxp67_ASAP7_75t_L g2532 ( 
.A(n_971),
.Y(n_2532)
);

CKINVDCx5p33_ASAP7_75t_R g2533 ( 
.A(n_1184),
.Y(n_2533)
);

CKINVDCx20_ASAP7_75t_R g2534 ( 
.A(n_1619),
.Y(n_2534)
);

CKINVDCx5p33_ASAP7_75t_R g2535 ( 
.A(n_349),
.Y(n_2535)
);

CKINVDCx20_ASAP7_75t_R g2536 ( 
.A(n_995),
.Y(n_2536)
);

CKINVDCx5p33_ASAP7_75t_R g2537 ( 
.A(n_1265),
.Y(n_2537)
);

CKINVDCx5p33_ASAP7_75t_R g2538 ( 
.A(n_956),
.Y(n_2538)
);

CKINVDCx5p33_ASAP7_75t_R g2539 ( 
.A(n_1495),
.Y(n_2539)
);

BUFx3_ASAP7_75t_L g2540 ( 
.A(n_1263),
.Y(n_2540)
);

CKINVDCx5p33_ASAP7_75t_R g2541 ( 
.A(n_1603),
.Y(n_2541)
);

CKINVDCx5p33_ASAP7_75t_R g2542 ( 
.A(n_1659),
.Y(n_2542)
);

CKINVDCx5p33_ASAP7_75t_R g2543 ( 
.A(n_1067),
.Y(n_2543)
);

CKINVDCx5p33_ASAP7_75t_R g2544 ( 
.A(n_919),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_1649),
.Y(n_2545)
);

BUFx10_ASAP7_75t_L g2546 ( 
.A(n_1496),
.Y(n_2546)
);

CKINVDCx5p33_ASAP7_75t_R g2547 ( 
.A(n_1608),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_696),
.Y(n_2548)
);

CKINVDCx5p33_ASAP7_75t_R g2549 ( 
.A(n_1651),
.Y(n_2549)
);

CKINVDCx5p33_ASAP7_75t_R g2550 ( 
.A(n_1654),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_9),
.Y(n_2551)
);

INVx3_ASAP7_75t_L g2552 ( 
.A(n_1610),
.Y(n_2552)
);

CKINVDCx5p33_ASAP7_75t_R g2553 ( 
.A(n_248),
.Y(n_2553)
);

CKINVDCx5p33_ASAP7_75t_R g2554 ( 
.A(n_875),
.Y(n_2554)
);

BUFx6f_ASAP7_75t_L g2555 ( 
.A(n_1320),
.Y(n_2555)
);

INVx1_ASAP7_75t_SL g2556 ( 
.A(n_236),
.Y(n_2556)
);

CKINVDCx5p33_ASAP7_75t_R g2557 ( 
.A(n_1604),
.Y(n_2557)
);

CKINVDCx5p33_ASAP7_75t_R g2558 ( 
.A(n_904),
.Y(n_2558)
);

CKINVDCx5p33_ASAP7_75t_R g2559 ( 
.A(n_1442),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_1097),
.Y(n_2560)
);

CKINVDCx5p33_ASAP7_75t_R g2561 ( 
.A(n_1534),
.Y(n_2561)
);

CKINVDCx5p33_ASAP7_75t_R g2562 ( 
.A(n_744),
.Y(n_2562)
);

CKINVDCx5p33_ASAP7_75t_R g2563 ( 
.A(n_250),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_1517),
.Y(n_2564)
);

CKINVDCx5p33_ASAP7_75t_R g2565 ( 
.A(n_1172),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_1690),
.Y(n_2566)
);

CKINVDCx20_ASAP7_75t_R g2567 ( 
.A(n_1637),
.Y(n_2567)
);

CKINVDCx5p33_ASAP7_75t_R g2568 ( 
.A(n_1430),
.Y(n_2568)
);

CKINVDCx5p33_ASAP7_75t_R g2569 ( 
.A(n_836),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_1203),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_1176),
.Y(n_2571)
);

BUFx8_ASAP7_75t_SL g2572 ( 
.A(n_237),
.Y(n_2572)
);

INVxp33_ASAP7_75t_SL g2573 ( 
.A(n_1579),
.Y(n_2573)
);

CKINVDCx5p33_ASAP7_75t_R g2574 ( 
.A(n_1615),
.Y(n_2574)
);

CKINVDCx5p33_ASAP7_75t_R g2575 ( 
.A(n_765),
.Y(n_2575)
);

CKINVDCx5p33_ASAP7_75t_R g2576 ( 
.A(n_1261),
.Y(n_2576)
);

CKINVDCx5p33_ASAP7_75t_R g2577 ( 
.A(n_427),
.Y(n_2577)
);

CKINVDCx5p33_ASAP7_75t_R g2578 ( 
.A(n_798),
.Y(n_2578)
);

CKINVDCx5p33_ASAP7_75t_R g2579 ( 
.A(n_1593),
.Y(n_2579)
);

CKINVDCx5p33_ASAP7_75t_R g2580 ( 
.A(n_953),
.Y(n_2580)
);

CKINVDCx5p33_ASAP7_75t_R g2581 ( 
.A(n_799),
.Y(n_2581)
);

CKINVDCx5p33_ASAP7_75t_R g2582 ( 
.A(n_1093),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_388),
.Y(n_2583)
);

CKINVDCx5p33_ASAP7_75t_R g2584 ( 
.A(n_93),
.Y(n_2584)
);

INVx1_ASAP7_75t_SL g2585 ( 
.A(n_829),
.Y(n_2585)
);

INVx2_ASAP7_75t_L g2586 ( 
.A(n_717),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_1192),
.Y(n_2587)
);

CKINVDCx5p33_ASAP7_75t_R g2588 ( 
.A(n_1657),
.Y(n_2588)
);

CKINVDCx5p33_ASAP7_75t_R g2589 ( 
.A(n_1622),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_1584),
.Y(n_2590)
);

CKINVDCx5p33_ASAP7_75t_R g2591 ( 
.A(n_137),
.Y(n_2591)
);

CKINVDCx5p33_ASAP7_75t_R g2592 ( 
.A(n_1212),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_1364),
.Y(n_2593)
);

CKINVDCx16_ASAP7_75t_R g2594 ( 
.A(n_1586),
.Y(n_2594)
);

CKINVDCx20_ASAP7_75t_R g2595 ( 
.A(n_425),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_1076),
.Y(n_2596)
);

CKINVDCx5p33_ASAP7_75t_R g2597 ( 
.A(n_703),
.Y(n_2597)
);

CKINVDCx5p33_ASAP7_75t_R g2598 ( 
.A(n_954),
.Y(n_2598)
);

CKINVDCx5p33_ASAP7_75t_R g2599 ( 
.A(n_1465),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_272),
.Y(n_2600)
);

CKINVDCx5p33_ASAP7_75t_R g2601 ( 
.A(n_661),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_391),
.Y(n_2602)
);

BUFx8_ASAP7_75t_SL g2603 ( 
.A(n_1696),
.Y(n_2603)
);

INVx1_ASAP7_75t_SL g2604 ( 
.A(n_620),
.Y(n_2604)
);

CKINVDCx5p33_ASAP7_75t_R g2605 ( 
.A(n_1045),
.Y(n_2605)
);

CKINVDCx5p33_ASAP7_75t_R g2606 ( 
.A(n_1171),
.Y(n_2606)
);

CKINVDCx20_ASAP7_75t_R g2607 ( 
.A(n_510),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_1599),
.Y(n_2608)
);

CKINVDCx5p33_ASAP7_75t_R g2609 ( 
.A(n_16),
.Y(n_2609)
);

CKINVDCx5p33_ASAP7_75t_R g2610 ( 
.A(n_1505),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_1129),
.Y(n_2611)
);

CKINVDCx5p33_ASAP7_75t_R g2612 ( 
.A(n_322),
.Y(n_2612)
);

BUFx8_ASAP7_75t_SL g2613 ( 
.A(n_1582),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_48),
.Y(n_2614)
);

CKINVDCx5p33_ASAP7_75t_R g2615 ( 
.A(n_1653),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_986),
.Y(n_2616)
);

CKINVDCx5p33_ASAP7_75t_R g2617 ( 
.A(n_1441),
.Y(n_2617)
);

CKINVDCx20_ASAP7_75t_R g2618 ( 
.A(n_1433),
.Y(n_2618)
);

INVx2_ASAP7_75t_SL g2619 ( 
.A(n_1211),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_795),
.Y(n_2620)
);

CKINVDCx5p33_ASAP7_75t_R g2621 ( 
.A(n_715),
.Y(n_2621)
);

BUFx6f_ASAP7_75t_L g2622 ( 
.A(n_1470),
.Y(n_2622)
);

CKINVDCx5p33_ASAP7_75t_R g2623 ( 
.A(n_142),
.Y(n_2623)
);

BUFx3_ASAP7_75t_L g2624 ( 
.A(n_1412),
.Y(n_2624)
);

CKINVDCx5p33_ASAP7_75t_R g2625 ( 
.A(n_438),
.Y(n_2625)
);

BUFx10_ASAP7_75t_L g2626 ( 
.A(n_1501),
.Y(n_2626)
);

CKINVDCx5p33_ASAP7_75t_R g2627 ( 
.A(n_790),
.Y(n_2627)
);

BUFx6f_ASAP7_75t_L g2628 ( 
.A(n_805),
.Y(n_2628)
);

CKINVDCx5p33_ASAP7_75t_R g2629 ( 
.A(n_633),
.Y(n_2629)
);

CKINVDCx20_ASAP7_75t_R g2630 ( 
.A(n_114),
.Y(n_2630)
);

BUFx3_ASAP7_75t_L g2631 ( 
.A(n_185),
.Y(n_2631)
);

CKINVDCx5p33_ASAP7_75t_R g2632 ( 
.A(n_671),
.Y(n_2632)
);

INVxp33_ASAP7_75t_R g2633 ( 
.A(n_553),
.Y(n_2633)
);

CKINVDCx5p33_ASAP7_75t_R g2634 ( 
.A(n_859),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_1373),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_1101),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_1163),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_713),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_1046),
.Y(n_2639)
);

INVx1_ASAP7_75t_SL g2640 ( 
.A(n_1554),
.Y(n_2640)
);

INVx2_ASAP7_75t_L g2641 ( 
.A(n_1472),
.Y(n_2641)
);

INVx4_ASAP7_75t_R g2642 ( 
.A(n_1130),
.Y(n_2642)
);

BUFx3_ASAP7_75t_L g2643 ( 
.A(n_651),
.Y(n_2643)
);

CKINVDCx5p33_ASAP7_75t_R g2644 ( 
.A(n_973),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_404),
.Y(n_2645)
);

CKINVDCx5p33_ASAP7_75t_R g2646 ( 
.A(n_739),
.Y(n_2646)
);

CKINVDCx5p33_ASAP7_75t_R g2647 ( 
.A(n_329),
.Y(n_2647)
);

CKINVDCx5p33_ASAP7_75t_R g2648 ( 
.A(n_1043),
.Y(n_2648)
);

CKINVDCx5p33_ASAP7_75t_R g2649 ( 
.A(n_1022),
.Y(n_2649)
);

CKINVDCx5p33_ASAP7_75t_R g2650 ( 
.A(n_325),
.Y(n_2650)
);

CKINVDCx5p33_ASAP7_75t_R g2651 ( 
.A(n_251),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_899),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_1077),
.Y(n_2653)
);

CKINVDCx5p33_ASAP7_75t_R g2654 ( 
.A(n_1206),
.Y(n_2654)
);

CKINVDCx5p33_ASAP7_75t_R g2655 ( 
.A(n_342),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_1553),
.Y(n_2656)
);

CKINVDCx5p33_ASAP7_75t_R g2657 ( 
.A(n_27),
.Y(n_2657)
);

INVx2_ASAP7_75t_L g2658 ( 
.A(n_624),
.Y(n_2658)
);

CKINVDCx5p33_ASAP7_75t_R g2659 ( 
.A(n_1011),
.Y(n_2659)
);

CKINVDCx5p33_ASAP7_75t_R g2660 ( 
.A(n_1179),
.Y(n_2660)
);

CKINVDCx5p33_ASAP7_75t_R g2661 ( 
.A(n_610),
.Y(n_2661)
);

CKINVDCx5p33_ASAP7_75t_R g2662 ( 
.A(n_1587),
.Y(n_2662)
);

CKINVDCx14_ASAP7_75t_R g2663 ( 
.A(n_207),
.Y(n_2663)
);

CKINVDCx5p33_ASAP7_75t_R g2664 ( 
.A(n_1438),
.Y(n_2664)
);

CKINVDCx5p33_ASAP7_75t_R g2665 ( 
.A(n_861),
.Y(n_2665)
);

CKINVDCx5p33_ASAP7_75t_R g2666 ( 
.A(n_1424),
.Y(n_2666)
);

CKINVDCx5p33_ASAP7_75t_R g2667 ( 
.A(n_1123),
.Y(n_2667)
);

CKINVDCx5p33_ASAP7_75t_R g2668 ( 
.A(n_1061),
.Y(n_2668)
);

CKINVDCx5p33_ASAP7_75t_R g2669 ( 
.A(n_1617),
.Y(n_2669)
);

CKINVDCx20_ASAP7_75t_R g2670 ( 
.A(n_945),
.Y(n_2670)
);

CKINVDCx5p33_ASAP7_75t_R g2671 ( 
.A(n_1566),
.Y(n_2671)
);

CKINVDCx5p33_ASAP7_75t_R g2672 ( 
.A(n_1162),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_1301),
.Y(n_2673)
);

CKINVDCx5p33_ASAP7_75t_R g2674 ( 
.A(n_168),
.Y(n_2674)
);

CKINVDCx20_ASAP7_75t_R g2675 ( 
.A(n_180),
.Y(n_2675)
);

INVx2_ASAP7_75t_SL g2676 ( 
.A(n_313),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_1316),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_1227),
.Y(n_2678)
);

BUFx6f_ASAP7_75t_L g2679 ( 
.A(n_327),
.Y(n_2679)
);

CKINVDCx5p33_ASAP7_75t_R g2680 ( 
.A(n_1416),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_1203),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_420),
.Y(n_2682)
);

CKINVDCx5p33_ASAP7_75t_R g2683 ( 
.A(n_1030),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_258),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_955),
.Y(n_2685)
);

CKINVDCx5p33_ASAP7_75t_R g2686 ( 
.A(n_736),
.Y(n_2686)
);

CKINVDCx5p33_ASAP7_75t_R g2687 ( 
.A(n_17),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_1239),
.Y(n_2688)
);

CKINVDCx20_ASAP7_75t_R g2689 ( 
.A(n_439),
.Y(n_2689)
);

CKINVDCx5p33_ASAP7_75t_R g2690 ( 
.A(n_122),
.Y(n_2690)
);

CKINVDCx5p33_ASAP7_75t_R g2691 ( 
.A(n_1179),
.Y(n_2691)
);

BUFx10_ASAP7_75t_L g2692 ( 
.A(n_1375),
.Y(n_2692)
);

CKINVDCx5p33_ASAP7_75t_R g2693 ( 
.A(n_1141),
.Y(n_2693)
);

CKINVDCx5p33_ASAP7_75t_R g2694 ( 
.A(n_992),
.Y(n_2694)
);

CKINVDCx5p33_ASAP7_75t_R g2695 ( 
.A(n_84),
.Y(n_2695)
);

CKINVDCx5p33_ASAP7_75t_R g2696 ( 
.A(n_634),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_1444),
.Y(n_2697)
);

CKINVDCx5p33_ASAP7_75t_R g2698 ( 
.A(n_138),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_469),
.Y(n_2699)
);

CKINVDCx16_ASAP7_75t_R g2700 ( 
.A(n_121),
.Y(n_2700)
);

CKINVDCx5p33_ASAP7_75t_R g2701 ( 
.A(n_1680),
.Y(n_2701)
);

CKINVDCx5p33_ASAP7_75t_R g2702 ( 
.A(n_1576),
.Y(n_2702)
);

CKINVDCx20_ASAP7_75t_R g2703 ( 
.A(n_1109),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_880),
.Y(n_2704)
);

BUFx2_ASAP7_75t_L g2705 ( 
.A(n_1674),
.Y(n_2705)
);

CKINVDCx5p33_ASAP7_75t_R g2706 ( 
.A(n_584),
.Y(n_2706)
);

CKINVDCx16_ASAP7_75t_R g2707 ( 
.A(n_27),
.Y(n_2707)
);

BUFx10_ASAP7_75t_L g2708 ( 
.A(n_1211),
.Y(n_2708)
);

CKINVDCx5p33_ASAP7_75t_R g2709 ( 
.A(n_1533),
.Y(n_2709)
);

CKINVDCx5p33_ASAP7_75t_R g2710 ( 
.A(n_1634),
.Y(n_2710)
);

CKINVDCx5p33_ASAP7_75t_R g2711 ( 
.A(n_1431),
.Y(n_2711)
);

INVx1_ASAP7_75t_SL g2712 ( 
.A(n_1160),
.Y(n_2712)
);

CKINVDCx20_ASAP7_75t_R g2713 ( 
.A(n_906),
.Y(n_2713)
);

CKINVDCx5p33_ASAP7_75t_R g2714 ( 
.A(n_1308),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_683),
.Y(n_2715)
);

CKINVDCx5p33_ASAP7_75t_R g2716 ( 
.A(n_422),
.Y(n_2716)
);

INVxp67_ASAP7_75t_L g2717 ( 
.A(n_1544),
.Y(n_2717)
);

INVx2_ASAP7_75t_SL g2718 ( 
.A(n_1187),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_1577),
.Y(n_2719)
);

CKINVDCx5p33_ASAP7_75t_R g2720 ( 
.A(n_756),
.Y(n_2720)
);

CKINVDCx5p33_ASAP7_75t_R g2721 ( 
.A(n_473),
.Y(n_2721)
);

CKINVDCx5p33_ASAP7_75t_R g2722 ( 
.A(n_640),
.Y(n_2722)
);

CKINVDCx5p33_ASAP7_75t_R g2723 ( 
.A(n_65),
.Y(n_2723)
);

CKINVDCx5p33_ASAP7_75t_R g2724 ( 
.A(n_1277),
.Y(n_2724)
);

CKINVDCx5p33_ASAP7_75t_R g2725 ( 
.A(n_205),
.Y(n_2725)
);

CKINVDCx5p33_ASAP7_75t_R g2726 ( 
.A(n_1195),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_705),
.Y(n_2727)
);

CKINVDCx5p33_ASAP7_75t_R g2728 ( 
.A(n_1204),
.Y(n_2728)
);

CKINVDCx5p33_ASAP7_75t_R g2729 ( 
.A(n_1693),
.Y(n_2729)
);

BUFx6f_ASAP7_75t_L g2730 ( 
.A(n_1207),
.Y(n_2730)
);

INVx1_ASAP7_75t_SL g2731 ( 
.A(n_1530),
.Y(n_2731)
);

BUFx3_ASAP7_75t_L g2732 ( 
.A(n_968),
.Y(n_2732)
);

INVx2_ASAP7_75t_L g2733 ( 
.A(n_125),
.Y(n_2733)
);

CKINVDCx5p33_ASAP7_75t_R g2734 ( 
.A(n_350),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_1624),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_809),
.Y(n_2736)
);

CKINVDCx5p33_ASAP7_75t_R g2737 ( 
.A(n_134),
.Y(n_2737)
);

CKINVDCx5p33_ASAP7_75t_R g2738 ( 
.A(n_472),
.Y(n_2738)
);

CKINVDCx5p33_ASAP7_75t_R g2739 ( 
.A(n_1571),
.Y(n_2739)
);

CKINVDCx5p33_ASAP7_75t_R g2740 ( 
.A(n_1160),
.Y(n_2740)
);

BUFx3_ASAP7_75t_L g2741 ( 
.A(n_134),
.Y(n_2741)
);

CKINVDCx5p33_ASAP7_75t_R g2742 ( 
.A(n_1033),
.Y(n_2742)
);

CKINVDCx5p33_ASAP7_75t_R g2743 ( 
.A(n_1415),
.Y(n_2743)
);

CKINVDCx5p33_ASAP7_75t_R g2744 ( 
.A(n_478),
.Y(n_2744)
);

BUFx6f_ASAP7_75t_L g2745 ( 
.A(n_1221),
.Y(n_2745)
);

CKINVDCx5p33_ASAP7_75t_R g2746 ( 
.A(n_1443),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_1580),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_877),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_1543),
.Y(n_2749)
);

CKINVDCx5p33_ASAP7_75t_R g2750 ( 
.A(n_336),
.Y(n_2750)
);

INVx1_ASAP7_75t_SL g2751 ( 
.A(n_1173),
.Y(n_2751)
);

CKINVDCx5p33_ASAP7_75t_R g2752 ( 
.A(n_637),
.Y(n_2752)
);

CKINVDCx5p33_ASAP7_75t_R g2753 ( 
.A(n_1011),
.Y(n_2753)
);

CKINVDCx5p33_ASAP7_75t_R g2754 ( 
.A(n_1432),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_905),
.Y(n_2755)
);

BUFx3_ASAP7_75t_L g2756 ( 
.A(n_319),
.Y(n_2756)
);

CKINVDCx5p33_ASAP7_75t_R g2757 ( 
.A(n_377),
.Y(n_2757)
);

CKINVDCx5p33_ASAP7_75t_R g2758 ( 
.A(n_596),
.Y(n_2758)
);

CKINVDCx5p33_ASAP7_75t_R g2759 ( 
.A(n_43),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_162),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_621),
.Y(n_2761)
);

CKINVDCx5p33_ASAP7_75t_R g2762 ( 
.A(n_230),
.Y(n_2762)
);

CKINVDCx20_ASAP7_75t_R g2763 ( 
.A(n_1306),
.Y(n_2763)
);

CKINVDCx5p33_ASAP7_75t_R g2764 ( 
.A(n_205),
.Y(n_2764)
);

CKINVDCx5p33_ASAP7_75t_R g2765 ( 
.A(n_1145),
.Y(n_2765)
);

CKINVDCx5p33_ASAP7_75t_R g2766 ( 
.A(n_1447),
.Y(n_2766)
);

CKINVDCx5p33_ASAP7_75t_R g2767 ( 
.A(n_1511),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_461),
.Y(n_2768)
);

INVx1_ASAP7_75t_SL g2769 ( 
.A(n_1031),
.Y(n_2769)
);

CKINVDCx5p33_ASAP7_75t_R g2770 ( 
.A(n_768),
.Y(n_2770)
);

CKINVDCx5p33_ASAP7_75t_R g2771 ( 
.A(n_1310),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_1658),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_1695),
.Y(n_2773)
);

CKINVDCx5p33_ASAP7_75t_R g2774 ( 
.A(n_247),
.Y(n_2774)
);

CKINVDCx5p33_ASAP7_75t_R g2775 ( 
.A(n_1679),
.Y(n_2775)
);

CKINVDCx5p33_ASAP7_75t_R g2776 ( 
.A(n_1157),
.Y(n_2776)
);

CKINVDCx5p33_ASAP7_75t_R g2777 ( 
.A(n_171),
.Y(n_2777)
);

CKINVDCx5p33_ASAP7_75t_R g2778 ( 
.A(n_256),
.Y(n_2778)
);

CKINVDCx5p33_ASAP7_75t_R g2779 ( 
.A(n_1575),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_1184),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_878),
.Y(n_2781)
);

INVx1_ASAP7_75t_SL g2782 ( 
.A(n_354),
.Y(n_2782)
);

CKINVDCx5p33_ASAP7_75t_R g2783 ( 
.A(n_633),
.Y(n_2783)
);

CKINVDCx5p33_ASAP7_75t_R g2784 ( 
.A(n_372),
.Y(n_2784)
);

CKINVDCx20_ASAP7_75t_R g2785 ( 
.A(n_1130),
.Y(n_2785)
);

INVx2_ASAP7_75t_SL g2786 ( 
.A(n_1531),
.Y(n_2786)
);

BUFx2_ASAP7_75t_L g2787 ( 
.A(n_428),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2026),
.Y(n_2788)
);

INVxp67_ASAP7_75t_SL g2789 ( 
.A(n_2026),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_1884),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_1884),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_1884),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_1884),
.Y(n_2793)
);

CKINVDCx16_ASAP7_75t_R g2794 ( 
.A(n_1725),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_1884),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2439),
.Y(n_2796)
);

CKINVDCx20_ASAP7_75t_R g2797 ( 
.A(n_1760),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2439),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2439),
.Y(n_2799)
);

CKINVDCx20_ASAP7_75t_R g2800 ( 
.A(n_1864),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2439),
.Y(n_2801)
);

CKINVDCx14_ASAP7_75t_R g2802 ( 
.A(n_2663),
.Y(n_2802)
);

INVx2_ASAP7_75t_L g2803 ( 
.A(n_2439),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2464),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2464),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2464),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2464),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2464),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_1709),
.Y(n_2809)
);

CKINVDCx16_ASAP7_75t_R g2810 ( 
.A(n_1893),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_1713),
.Y(n_2811)
);

CKINVDCx16_ASAP7_75t_R g2812 ( 
.A(n_1962),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_1719),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_1723),
.Y(n_2814)
);

INVx2_ASAP7_75t_L g2815 ( 
.A(n_1752),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_1726),
.Y(n_2816)
);

INVxp67_ASAP7_75t_L g2817 ( 
.A(n_1956),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_1729),
.Y(n_2818)
);

CKINVDCx5p33_ASAP7_75t_R g2819 ( 
.A(n_2266),
.Y(n_2819)
);

INVxp33_ASAP7_75t_SL g2820 ( 
.A(n_2331),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_1752),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_1732),
.Y(n_2822)
);

INVxp67_ASAP7_75t_SL g2823 ( 
.A(n_1752),
.Y(n_2823)
);

INVx2_ASAP7_75t_L g2824 ( 
.A(n_1758),
.Y(n_2824)
);

CKINVDCx5p33_ASAP7_75t_R g2825 ( 
.A(n_2572),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_1736),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_1748),
.Y(n_2827)
);

INVxp67_ASAP7_75t_L g2828 ( 
.A(n_2083),
.Y(n_2828)
);

CKINVDCx20_ASAP7_75t_R g2829 ( 
.A(n_1738),
.Y(n_2829)
);

CKINVDCx20_ASAP7_75t_R g2830 ( 
.A(n_1929),
.Y(n_2830)
);

BUFx3_ASAP7_75t_L g2831 ( 
.A(n_2122),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_1753),
.Y(n_2832)
);

CKINVDCx16_ASAP7_75t_R g2833 ( 
.A(n_2101),
.Y(n_2833)
);

BUFx6f_ASAP7_75t_L g2834 ( 
.A(n_1952),
.Y(n_2834)
);

INVx2_ASAP7_75t_L g2835 ( 
.A(n_1758),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_1763),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_1766),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_1771),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_1773),
.Y(n_2839)
);

INVxp67_ASAP7_75t_L g2840 ( 
.A(n_2148),
.Y(n_2840)
);

CKINVDCx5p33_ASAP7_75t_R g2841 ( 
.A(n_2282),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_1778),
.Y(n_2842)
);

INVxp33_ASAP7_75t_L g2843 ( 
.A(n_2351),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_1813),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_1820),
.Y(n_2845)
);

INVx2_ASAP7_75t_L g2846 ( 
.A(n_1758),
.Y(n_2846)
);

CKINVDCx14_ASAP7_75t_R g2847 ( 
.A(n_1859),
.Y(n_2847)
);

INVx1_ASAP7_75t_SL g2848 ( 
.A(n_1779),
.Y(n_2848)
);

CKINVDCx5p33_ASAP7_75t_R g2849 ( 
.A(n_2603),
.Y(n_2849)
);

INVx1_ASAP7_75t_SL g2850 ( 
.A(n_1784),
.Y(n_2850)
);

CKINVDCx16_ASAP7_75t_R g2851 ( 
.A(n_2159),
.Y(n_2851)
);

INVxp67_ASAP7_75t_SL g2852 ( 
.A(n_1964),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_1823),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_1833),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_1837),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_1844),
.Y(n_2856)
);

CKINVDCx5p33_ASAP7_75t_R g2857 ( 
.A(n_2613),
.Y(n_2857)
);

BUFx3_ASAP7_75t_L g2858 ( 
.A(n_2144),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_1846),
.Y(n_2859)
);

CKINVDCx5p33_ASAP7_75t_R g2860 ( 
.A(n_2368),
.Y(n_2860)
);

CKINVDCx5p33_ASAP7_75t_R g2861 ( 
.A(n_2427),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_1851),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_1853),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_1964),
.Y(n_2864)
);

INVx1_ASAP7_75t_SL g2865 ( 
.A(n_1811),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_1857),
.Y(n_2866)
);

CKINVDCx16_ASAP7_75t_R g2867 ( 
.A(n_2700),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_1858),
.Y(n_2868)
);

BUFx2_ASAP7_75t_L g2869 ( 
.A(n_2392),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_1867),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_1870),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_1896),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_1902),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_1903),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_1914),
.Y(n_2875)
);

INVxp67_ASAP7_75t_SL g2876 ( 
.A(n_1964),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_1915),
.Y(n_2877)
);

INVxp33_ASAP7_75t_SL g2878 ( 
.A(n_2415),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_1918),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_1922),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_1923),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_1926),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_1932),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_1935),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_1936),
.Y(n_2885)
);

CKINVDCx14_ASAP7_75t_R g2886 ( 
.A(n_2453),
.Y(n_2886)
);

CKINVDCx5p33_ASAP7_75t_R g2887 ( 
.A(n_2707),
.Y(n_2887)
);

CKINVDCx20_ASAP7_75t_R g2888 ( 
.A(n_1994),
.Y(n_2888)
);

CKINVDCx5p33_ASAP7_75t_R g2889 ( 
.A(n_2006),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_1941),
.Y(n_2890)
);

INVxp67_ASAP7_75t_SL g2891 ( 
.A(n_1991),
.Y(n_2891)
);

CKINVDCx20_ASAP7_75t_R g2892 ( 
.A(n_2126),
.Y(n_2892)
);

CKINVDCx5p33_ASAP7_75t_R g2893 ( 
.A(n_2141),
.Y(n_2893)
);

CKINVDCx16_ASAP7_75t_R g2894 ( 
.A(n_1733),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_1945),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_1963),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_1966),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_1974),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_1981),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_1982),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_1995),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_1991),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2002),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2018),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2025),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_1991),
.Y(n_2906)
);

CKINVDCx20_ASAP7_75t_R g2907 ( 
.A(n_2219),
.Y(n_2907)
);

INVxp67_ASAP7_75t_SL g2908 ( 
.A(n_2036),
.Y(n_2908)
);

INVx2_ASAP7_75t_L g2909 ( 
.A(n_2036),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2060),
.Y(n_2910)
);

INVx2_ASAP7_75t_L g2911 ( 
.A(n_2036),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2065),
.Y(n_2912)
);

INVxp33_ASAP7_75t_L g2913 ( 
.A(n_2472),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2071),
.Y(n_2914)
);

CKINVDCx5p33_ASAP7_75t_R g2915 ( 
.A(n_2274),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2075),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2079),
.Y(n_2917)
);

INVxp67_ASAP7_75t_SL g2918 ( 
.A(n_2289),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2081),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2089),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2099),
.Y(n_2921)
);

CKINVDCx5p33_ASAP7_75t_R g2922 ( 
.A(n_2322),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2103),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2108),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2110),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2111),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2118),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2143),
.Y(n_2928)
);

INVxp33_ASAP7_75t_SL g2929 ( 
.A(n_2450),
.Y(n_2929)
);

CKINVDCx20_ASAP7_75t_R g2930 ( 
.A(n_2403),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2150),
.Y(n_2931)
);

INVx2_ASAP7_75t_L g2932 ( 
.A(n_2289),
.Y(n_2932)
);

NOR2xp67_ASAP7_75t_L g2933 ( 
.A(n_1742),
.B(n_0),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2157),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2168),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2178),
.Y(n_2936)
);

CKINVDCx5p33_ASAP7_75t_R g2937 ( 
.A(n_2489),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2187),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2188),
.Y(n_2939)
);

CKINVDCx5p33_ASAP7_75t_R g2940 ( 
.A(n_2497),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2190),
.Y(n_2941)
);

INVxp33_ASAP7_75t_L g2942 ( 
.A(n_2787),
.Y(n_2942)
);

INVxp33_ASAP7_75t_L g2943 ( 
.A(n_1737),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2193),
.Y(n_2944)
);

INVxp67_ASAP7_75t_L g2945 ( 
.A(n_1740),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2194),
.Y(n_2946)
);

CKINVDCx5p33_ASAP7_75t_R g2947 ( 
.A(n_2523),
.Y(n_2947)
);

HB1xp67_ASAP7_75t_L g2948 ( 
.A(n_1786),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2196),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2199),
.Y(n_2950)
);

INVxp67_ASAP7_75t_SL g2951 ( 
.A(n_2289),
.Y(n_2951)
);

INVx2_ASAP7_75t_L g2952 ( 
.A(n_2628),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2206),
.Y(n_2953)
);

CKINVDCx5p33_ASAP7_75t_R g2954 ( 
.A(n_2534),
.Y(n_2954)
);

INVxp67_ASAP7_75t_SL g2955 ( 
.A(n_2628),
.Y(n_2955)
);

INVxp67_ASAP7_75t_SL g2956 ( 
.A(n_2628),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2207),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2211),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2229),
.Y(n_2959)
);

CKINVDCx5p33_ASAP7_75t_R g2960 ( 
.A(n_2567),
.Y(n_2960)
);

NOR2xp33_ASAP7_75t_L g2961 ( 
.A(n_2105),
.B(n_0),
.Y(n_2961)
);

BUFx6f_ASAP7_75t_L g2962 ( 
.A(n_1952),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2230),
.Y(n_2963)
);

HB1xp67_ASAP7_75t_L g2964 ( 
.A(n_1799),
.Y(n_2964)
);

INVx1_ASAP7_75t_L g2965 ( 
.A(n_2233),
.Y(n_2965)
);

HB1xp67_ASAP7_75t_L g2966 ( 
.A(n_1826),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2237),
.Y(n_2967)
);

INVx4_ASAP7_75t_R g2968 ( 
.A(n_1720),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2241),
.Y(n_2969)
);

CKINVDCx16_ASAP7_75t_R g2970 ( 
.A(n_1933),
.Y(n_2970)
);

INVxp33_ASAP7_75t_SL g2971 ( 
.A(n_2399),
.Y(n_2971)
);

INVx2_ASAP7_75t_L g2972 ( 
.A(n_2679),
.Y(n_2972)
);

CKINVDCx5p33_ASAP7_75t_R g2973 ( 
.A(n_2618),
.Y(n_2973)
);

CKINVDCx20_ASAP7_75t_R g2974 ( 
.A(n_2763),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2243),
.Y(n_2975)
);

INVxp33_ASAP7_75t_L g2976 ( 
.A(n_1886),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2251),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2259),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2262),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2265),
.Y(n_2980)
);

INVx2_ASAP7_75t_L g2981 ( 
.A(n_2679),
.Y(n_2981)
);

INVxp67_ASAP7_75t_L g2982 ( 
.A(n_1855),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2300),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2316),
.Y(n_2984)
);

CKINVDCx20_ASAP7_75t_R g2985 ( 
.A(n_1815),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2319),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2325),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2334),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2343),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2348),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2352),
.Y(n_2991)
);

INVxp67_ASAP7_75t_L g2992 ( 
.A(n_1916),
.Y(n_2992)
);

INVx1_ASAP7_75t_SL g2993 ( 
.A(n_1831),
.Y(n_2993)
);

INVxp33_ASAP7_75t_L g2994 ( 
.A(n_1899),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2355),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2358),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2361),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2363),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2365),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2366),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2374),
.Y(n_3001)
);

INVxp67_ASAP7_75t_SL g3002 ( 
.A(n_2679),
.Y(n_3002)
);

BUFx2_ASAP7_75t_L g3003 ( 
.A(n_1951),
.Y(n_3003)
);

CKINVDCx16_ASAP7_75t_R g3004 ( 
.A(n_2594),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2386),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2390),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2391),
.Y(n_3007)
);

CKINVDCx20_ASAP7_75t_R g3008 ( 
.A(n_2785),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2402),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2404),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2414),
.Y(n_3011)
);

INVxp67_ASAP7_75t_SL g3012 ( 
.A(n_2730),
.Y(n_3012)
);

HB1xp67_ASAP7_75t_L g3013 ( 
.A(n_2057),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2417),
.Y(n_3014)
);

INVxp33_ASAP7_75t_SL g3015 ( 
.A(n_2473),
.Y(n_3015)
);

INVxp67_ASAP7_75t_SL g3016 ( 
.A(n_2730),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2431),
.Y(n_3017)
);

BUFx2_ASAP7_75t_L g3018 ( 
.A(n_2078),
.Y(n_3018)
);

CKINVDCx5p33_ASAP7_75t_R g3019 ( 
.A(n_1711),
.Y(n_3019)
);

CKINVDCx5p33_ASAP7_75t_R g3020 ( 
.A(n_1718),
.Y(n_3020)
);

INVx1_ASAP7_75t_SL g3021 ( 
.A(n_1850),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2432),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2433),
.Y(n_3023)
);

CKINVDCx5p33_ASAP7_75t_R g3024 ( 
.A(n_2774),
.Y(n_3024)
);

INVxp67_ASAP7_75t_SL g3025 ( 
.A(n_2730),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2446),
.Y(n_3026)
);

INVx3_ASAP7_75t_L g3027 ( 
.A(n_2183),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2451),
.Y(n_3028)
);

HB1xp67_ASAP7_75t_L g3029 ( 
.A(n_2514),
.Y(n_3029)
);

INVxp67_ASAP7_75t_SL g3030 ( 
.A(n_2745),
.Y(n_3030)
);

CKINVDCx5p33_ASAP7_75t_R g3031 ( 
.A(n_2783),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_2458),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_2460),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2477),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2485),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2487),
.Y(n_3036)
);

CKINVDCx5p33_ASAP7_75t_R g3037 ( 
.A(n_1724),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2499),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2505),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2525),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2527),
.Y(n_3041)
);

INVxp67_ASAP7_75t_L g3042 ( 
.A(n_2631),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2548),
.Y(n_3043)
);

CKINVDCx5p33_ASAP7_75t_R g3044 ( 
.A(n_2776),
.Y(n_3044)
);

CKINVDCx20_ASAP7_75t_R g3045 ( 
.A(n_1880),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2551),
.Y(n_3046)
);

NOR2xp67_ASAP7_75t_L g3047 ( 
.A(n_2044),
.B(n_1),
.Y(n_3047)
);

INVx2_ASAP7_75t_L g3048 ( 
.A(n_2834),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2789),
.B(n_2847),
.Y(n_3049)
);

BUFx2_ASAP7_75t_L g3050 ( 
.A(n_2860),
.Y(n_3050)
);

AND2x2_ASAP7_75t_L g3051 ( 
.A(n_2802),
.B(n_2705),
.Y(n_3051)
);

OAI22x1_ASAP7_75t_SL g3052 ( 
.A1(n_2985),
.A2(n_1912),
.B1(n_1928),
.B2(n_1890),
.Y(n_3052)
);

AND2x2_ASAP7_75t_L g3053 ( 
.A(n_2943),
.B(n_1728),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2823),
.Y(n_3054)
);

CKINVDCx16_ASAP7_75t_R g3055 ( 
.A(n_2794),
.Y(n_3055)
);

OAI22xp5_ASAP7_75t_L g3056 ( 
.A1(n_2817),
.A2(n_1992),
.B1(n_2017),
.B2(n_1944),
.Y(n_3056)
);

BUFx6f_ASAP7_75t_L g3057 ( 
.A(n_2834),
.Y(n_3057)
);

BUFx2_ASAP7_75t_L g3058 ( 
.A(n_2861),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2852),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2876),
.Y(n_3060)
);

BUFx2_ASAP7_75t_L g3061 ( 
.A(n_2887),
.Y(n_3061)
);

AND2x2_ASAP7_75t_L g3062 ( 
.A(n_2976),
.B(n_1728),
.Y(n_3062)
);

INVx2_ASAP7_75t_L g3063 ( 
.A(n_2834),
.Y(n_3063)
);

AOI22xp5_ASAP7_75t_L g3064 ( 
.A1(n_2929),
.A2(n_2113),
.B1(n_2186),
.B2(n_2109),
.Y(n_3064)
);

XNOR2x2_ASAP7_75t_L g3065 ( 
.A(n_2848),
.B(n_2633),
.Y(n_3065)
);

NOR2x1_ASAP7_75t_L g3066 ( 
.A(n_2831),
.B(n_2208),
.Y(n_3066)
);

BUFx8_ASAP7_75t_SL g3067 ( 
.A(n_3008),
.Y(n_3067)
);

AND2x2_ASAP7_75t_L g3068 ( 
.A(n_2994),
.B(n_1860),
.Y(n_3068)
);

BUFx2_ASAP7_75t_L g3069 ( 
.A(n_3019),
.Y(n_3069)
);

BUFx2_ASAP7_75t_L g3070 ( 
.A(n_3020),
.Y(n_3070)
);

HB1xp67_ASAP7_75t_L g3071 ( 
.A(n_2810),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_2891),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2886),
.B(n_2908),
.Y(n_3073)
);

INVx3_ASAP7_75t_L g3074 ( 
.A(n_3027),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2918),
.Y(n_3075)
);

AND2x4_ASAP7_75t_L g3076 ( 
.A(n_2858),
.B(n_2643),
.Y(n_3076)
);

INVx2_ASAP7_75t_L g3077 ( 
.A(n_2962),
.Y(n_3077)
);

BUFx2_ASAP7_75t_L g3078 ( 
.A(n_3024),
.Y(n_3078)
);

INVx4_ASAP7_75t_L g3079 ( 
.A(n_3031),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2951),
.Y(n_3080)
);

OAI21x1_ASAP7_75t_L g3081 ( 
.A1(n_2803),
.A2(n_2226),
.B(n_1791),
.Y(n_3081)
);

INVx2_ASAP7_75t_L g3082 ( 
.A(n_2962),
.Y(n_3082)
);

INVx2_ASAP7_75t_L g3083 ( 
.A(n_2962),
.Y(n_3083)
);

BUFx6f_ASAP7_75t_L g3084 ( 
.A(n_2815),
.Y(n_3084)
);

OAI21x1_ASAP7_75t_L g3085 ( 
.A1(n_2790),
.A2(n_2226),
.B(n_1791),
.Y(n_3085)
);

INVx2_ASAP7_75t_L g3086 ( 
.A(n_2821),
.Y(n_3086)
);

HB1xp67_ASAP7_75t_L g3087 ( 
.A(n_2812),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2955),
.Y(n_3088)
);

INVx5_ASAP7_75t_L g3089 ( 
.A(n_2833),
.Y(n_3089)
);

CKINVDCx5p33_ASAP7_75t_R g3090 ( 
.A(n_2889),
.Y(n_3090)
);

BUFx6f_ASAP7_75t_L g3091 ( 
.A(n_2824),
.Y(n_3091)
);

INVx2_ASAP7_75t_L g3092 ( 
.A(n_2835),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2956),
.Y(n_3093)
);

BUFx6f_ASAP7_75t_L g3094 ( 
.A(n_2846),
.Y(n_3094)
);

OA21x2_ASAP7_75t_L g3095 ( 
.A1(n_2791),
.A2(n_2793),
.B(n_2792),
.Y(n_3095)
);

INVx2_ASAP7_75t_L g3096 ( 
.A(n_2864),
.Y(n_3096)
);

OAI22xp5_ASAP7_75t_SL g3097 ( 
.A1(n_3045),
.A2(n_2249),
.B1(n_2250),
.B2(n_2209),
.Y(n_3097)
);

INVx2_ASAP7_75t_L g3098 ( 
.A(n_2902),
.Y(n_3098)
);

NOR2xp33_ASAP7_75t_L g3099 ( 
.A(n_2971),
.B(n_2299),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_3002),
.Y(n_3100)
);

OAI21x1_ASAP7_75t_L g3101 ( 
.A1(n_2795),
.A2(n_2552),
.B(n_1715),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_3012),
.Y(n_3102)
);

HB1xp67_ASAP7_75t_L g3103 ( 
.A(n_2851),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_3016),
.B(n_1714),
.Y(n_3104)
);

INVx3_ASAP7_75t_L g3105 ( 
.A(n_3027),
.Y(n_3105)
);

INVx6_ASAP7_75t_L g3106 ( 
.A(n_2867),
.Y(n_3106)
);

CKINVDCx20_ASAP7_75t_R g3107 ( 
.A(n_2829),
.Y(n_3107)
);

INVx5_ASAP7_75t_L g3108 ( 
.A(n_2869),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_3025),
.B(n_1721),
.Y(n_3109)
);

AND2x2_ASAP7_75t_L g3110 ( 
.A(n_2942),
.B(n_1860),
.Y(n_3110)
);

OAI21x1_ASAP7_75t_L g3111 ( 
.A1(n_2796),
.A2(n_2552),
.B(n_1761),
.Y(n_3111)
);

INVx2_ASAP7_75t_L g3112 ( 
.A(n_2906),
.Y(n_3112)
);

BUFx6f_ASAP7_75t_L g3113 ( 
.A(n_2909),
.Y(n_3113)
);

BUFx3_ASAP7_75t_L g3114 ( 
.A(n_3003),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_3030),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_L g3116 ( 
.A(n_2945),
.B(n_2982),
.Y(n_3116)
);

INVx2_ASAP7_75t_L g3117 ( 
.A(n_2911),
.Y(n_3117)
);

HB1xp67_ASAP7_75t_L g3118 ( 
.A(n_3037),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2788),
.Y(n_3119)
);

BUFx6f_ASAP7_75t_L g3120 ( 
.A(n_2932),
.Y(n_3120)
);

INVx2_ASAP7_75t_L g3121 ( 
.A(n_2952),
.Y(n_3121)
);

AND2x4_ASAP7_75t_L g3122 ( 
.A(n_2828),
.B(n_2732),
.Y(n_3122)
);

CKINVDCx16_ASAP7_75t_R g3123 ( 
.A(n_2894),
.Y(n_3123)
);

NOR2xp33_ASAP7_75t_L g3124 ( 
.A(n_3015),
.B(n_2573),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_2798),
.Y(n_3125)
);

HB1xp67_ASAP7_75t_L g3126 ( 
.A(n_3044),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_2799),
.Y(n_3127)
);

AND2x6_ASAP7_75t_L g3128 ( 
.A(n_2809),
.B(n_2741),
.Y(n_3128)
);

NOR2xp33_ASAP7_75t_SL g3129 ( 
.A(n_2841),
.B(n_2080),
.Y(n_3129)
);

AND2x6_ASAP7_75t_L g3130 ( 
.A(n_2811),
.B(n_2756),
.Y(n_3130)
);

INVx2_ASAP7_75t_L g3131 ( 
.A(n_2972),
.Y(n_3131)
);

HB1xp67_ASAP7_75t_L g3132 ( 
.A(n_2850),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2801),
.Y(n_3133)
);

BUFx6f_ASAP7_75t_L g3134 ( 
.A(n_2981),
.Y(n_3134)
);

BUFx6f_ASAP7_75t_L g3135 ( 
.A(n_3018),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2804),
.Y(n_3136)
);

HB1xp67_ASAP7_75t_L g3137 ( 
.A(n_2865),
.Y(n_3137)
);

BUFx6f_ASAP7_75t_L g3138 ( 
.A(n_2813),
.Y(n_3138)
);

BUFx3_ASAP7_75t_L g3139 ( 
.A(n_2805),
.Y(n_3139)
);

INVx4_ASAP7_75t_L g3140 ( 
.A(n_2849),
.Y(n_3140)
);

OA21x2_ASAP7_75t_L g3141 ( 
.A1(n_2806),
.A2(n_1769),
.B(n_1731),
.Y(n_3141)
);

HB1xp67_ASAP7_75t_L g3142 ( 
.A(n_2993),
.Y(n_3142)
);

BUFx6f_ASAP7_75t_L g3143 ( 
.A(n_2814),
.Y(n_3143)
);

BUFx6f_ASAP7_75t_L g3144 ( 
.A(n_2816),
.Y(n_3144)
);

NOR2x1_ASAP7_75t_L g3145 ( 
.A(n_2818),
.B(n_2349),
.Y(n_3145)
);

INVx2_ASAP7_75t_L g3146 ( 
.A(n_2807),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_2808),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2822),
.Y(n_3148)
);

BUFx6f_ASAP7_75t_L g3149 ( 
.A(n_2826),
.Y(n_3149)
);

AND2x4_ASAP7_75t_L g3150 ( 
.A(n_2840),
.B(n_1722),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_L g3151 ( 
.A(n_2992),
.B(n_1774),
.Y(n_3151)
);

INVx4_ASAP7_75t_L g3152 ( 
.A(n_2857),
.Y(n_3152)
);

INVx3_ASAP7_75t_L g3153 ( 
.A(n_2827),
.Y(n_3153)
);

AOI22xp5_ASAP7_75t_L g3154 ( 
.A1(n_2820),
.A2(n_2272),
.B1(n_2279),
.B2(n_2263),
.Y(n_3154)
);

BUFx6f_ASAP7_75t_L g3155 ( 
.A(n_2832),
.Y(n_3155)
);

BUFx2_ASAP7_75t_L g3156 ( 
.A(n_2819),
.Y(n_3156)
);

HB1xp67_ASAP7_75t_L g3157 ( 
.A(n_3021),
.Y(n_3157)
);

NAND2xp5_ASAP7_75t_L g3158 ( 
.A(n_3042),
.B(n_2836),
.Y(n_3158)
);

OAI21x1_ASAP7_75t_L g3159 ( 
.A1(n_2837),
.A2(n_1796),
.B(n_1793),
.Y(n_3159)
);

INVx3_ASAP7_75t_L g3160 ( 
.A(n_2838),
.Y(n_3160)
);

BUFx3_ASAP7_75t_L g3161 ( 
.A(n_2839),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2842),
.Y(n_3162)
);

INVxp67_ASAP7_75t_L g3163 ( 
.A(n_2948),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2844),
.Y(n_3164)
);

CKINVDCx5p33_ASAP7_75t_R g3165 ( 
.A(n_2893),
.Y(n_3165)
);

BUFx8_ASAP7_75t_L g3166 ( 
.A(n_2845),
.Y(n_3166)
);

AND2x4_ASAP7_75t_L g3167 ( 
.A(n_2964),
.B(n_1751),
.Y(n_3167)
);

BUFx2_ASAP7_75t_L g3168 ( 
.A(n_2825),
.Y(n_3168)
);

AND2x4_ASAP7_75t_L g3169 ( 
.A(n_2966),
.B(n_1939),
.Y(n_3169)
);

BUFx6f_ASAP7_75t_L g3170 ( 
.A(n_2853),
.Y(n_3170)
);

AOI22xp5_ASAP7_75t_SL g3171 ( 
.A1(n_2830),
.A2(n_2313),
.B1(n_2321),
.B2(n_2281),
.Y(n_3171)
);

INVx2_ASAP7_75t_L g3172 ( 
.A(n_2854),
.Y(n_3172)
);

INVx2_ASAP7_75t_L g3173 ( 
.A(n_2855),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_L g3174 ( 
.A(n_2856),
.B(n_1797),
.Y(n_3174)
);

INVx2_ASAP7_75t_L g3175 ( 
.A(n_2859),
.Y(n_3175)
);

INVx5_ASAP7_75t_L g3176 ( 
.A(n_2970),
.Y(n_3176)
);

INVx2_ASAP7_75t_L g3177 ( 
.A(n_2862),
.Y(n_3177)
);

OAI22x1_ASAP7_75t_R g3178 ( 
.A1(n_2888),
.A2(n_2328),
.B1(n_2339),
.B2(n_2326),
.Y(n_3178)
);

AND2x4_ASAP7_75t_L g3179 ( 
.A(n_3013),
.B(n_2171),
.Y(n_3179)
);

CKINVDCx16_ASAP7_75t_R g3180 ( 
.A(n_3004),
.Y(n_3180)
);

BUFx6f_ASAP7_75t_L g3181 ( 
.A(n_2863),
.Y(n_3181)
);

AND2x4_ASAP7_75t_L g3182 ( 
.A(n_3029),
.B(n_2217),
.Y(n_3182)
);

CKINVDCx5p33_ASAP7_75t_R g3183 ( 
.A(n_2915),
.Y(n_3183)
);

HB1xp67_ASAP7_75t_L g3184 ( 
.A(n_2922),
.Y(n_3184)
);

AND2x2_ASAP7_75t_L g3185 ( 
.A(n_2843),
.B(n_2080),
.Y(n_3185)
);

AND2x2_ASAP7_75t_L g3186 ( 
.A(n_2913),
.B(n_2104),
.Y(n_3186)
);

AND2x2_ASAP7_75t_L g3187 ( 
.A(n_2866),
.B(n_2104),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2868),
.Y(n_3188)
);

BUFx6f_ASAP7_75t_L g3189 ( 
.A(n_2870),
.Y(n_3189)
);

BUFx8_ASAP7_75t_L g3190 ( 
.A(n_2871),
.Y(n_3190)
);

INVx2_ASAP7_75t_L g3191 ( 
.A(n_2872),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_2873),
.Y(n_3192)
);

HB1xp67_ASAP7_75t_L g3193 ( 
.A(n_2937),
.Y(n_3193)
);

BUFx6f_ASAP7_75t_L g3194 ( 
.A(n_2874),
.Y(n_3194)
);

INVx2_ASAP7_75t_L g3195 ( 
.A(n_2875),
.Y(n_3195)
);

HB1xp67_ASAP7_75t_L g3196 ( 
.A(n_2940),
.Y(n_3196)
);

INVx2_ASAP7_75t_L g3197 ( 
.A(n_2877),
.Y(n_3197)
);

BUFx2_ASAP7_75t_L g3198 ( 
.A(n_2797),
.Y(n_3198)
);

INVx1_ASAP7_75t_SL g3199 ( 
.A(n_2947),
.Y(n_3199)
);

INVx2_ASAP7_75t_L g3200 ( 
.A(n_2879),
.Y(n_3200)
);

OAI21x1_ASAP7_75t_L g3201 ( 
.A1(n_2880),
.A2(n_1803),
.B(n_1798),
.Y(n_3201)
);

AND2x4_ASAP7_75t_L g3202 ( 
.A(n_2800),
.B(n_2881),
.Y(n_3202)
);

BUFx2_ASAP7_75t_L g3203 ( 
.A(n_2954),
.Y(n_3203)
);

INVx2_ASAP7_75t_L g3204 ( 
.A(n_2882),
.Y(n_3204)
);

OAI21x1_ASAP7_75t_L g3205 ( 
.A1(n_2883),
.A2(n_1827),
.B(n_1809),
.Y(n_3205)
);

BUFx2_ASAP7_75t_L g3206 ( 
.A(n_2960),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_2884),
.Y(n_3207)
);

INVxp33_ASAP7_75t_SL g3208 ( 
.A(n_2973),
.Y(n_3208)
);

BUFx6f_ASAP7_75t_L g3209 ( 
.A(n_2885),
.Y(n_3209)
);

INVx2_ASAP7_75t_L g3210 ( 
.A(n_2890),
.Y(n_3210)
);

BUFx6f_ASAP7_75t_L g3211 ( 
.A(n_2895),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_L g3212 ( 
.A(n_2896),
.B(n_1832),
.Y(n_3212)
);

INVx5_ASAP7_75t_L g3213 ( 
.A(n_2878),
.Y(n_3213)
);

OA21x2_ASAP7_75t_L g3214 ( 
.A1(n_2897),
.A2(n_1868),
.B(n_1838),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_2898),
.Y(n_3215)
);

NAND2xp5_ASAP7_75t_L g3216 ( 
.A(n_2899),
.B(n_2900),
.Y(n_3216)
);

BUFx8_ASAP7_75t_SL g3217 ( 
.A(n_2892),
.Y(n_3217)
);

INVx2_ASAP7_75t_L g3218 ( 
.A(n_2901),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_2903),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_2904),
.B(n_1874),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_2905),
.Y(n_3221)
);

INVx3_ASAP7_75t_L g3222 ( 
.A(n_2910),
.Y(n_3222)
);

HB1xp67_ASAP7_75t_L g3223 ( 
.A(n_2907),
.Y(n_3223)
);

AOI22xp5_ASAP7_75t_L g3224 ( 
.A1(n_2961),
.A2(n_2395),
.B1(n_2423),
.B2(n_2388),
.Y(n_3224)
);

BUFx12f_ASAP7_75t_L g3225 ( 
.A(n_2968),
.Y(n_3225)
);

NOR2xp33_ASAP7_75t_SL g3226 ( 
.A(n_2930),
.B(n_2454),
.Y(n_3226)
);

CKINVDCx5p33_ASAP7_75t_R g3227 ( 
.A(n_2974),
.Y(n_3227)
);

INVx2_ASAP7_75t_L g3228 ( 
.A(n_2912),
.Y(n_3228)
);

AND2x2_ASAP7_75t_L g3229 ( 
.A(n_2914),
.B(n_2454),
.Y(n_3229)
);

INVx2_ASAP7_75t_L g3230 ( 
.A(n_2916),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_2917),
.Y(n_3231)
);

INVx2_ASAP7_75t_L g3232 ( 
.A(n_2919),
.Y(n_3232)
);

BUFx6f_ASAP7_75t_L g3233 ( 
.A(n_2920),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_2921),
.Y(n_3234)
);

CKINVDCx5p33_ASAP7_75t_R g3235 ( 
.A(n_2923),
.Y(n_3235)
);

INVxp33_ASAP7_75t_SL g3236 ( 
.A(n_2933),
.Y(n_3236)
);

OAI22xp33_ASAP7_75t_SL g3237 ( 
.A1(n_2924),
.A2(n_1765),
.B1(n_1996),
.B2(n_1764),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_2925),
.Y(n_3238)
);

BUFx6f_ASAP7_75t_L g3239 ( 
.A(n_2926),
.Y(n_3239)
);

AND2x4_ASAP7_75t_L g3240 ( 
.A(n_2927),
.B(n_2240),
.Y(n_3240)
);

INVx3_ASAP7_75t_L g3241 ( 
.A(n_2928),
.Y(n_3241)
);

INVx3_ASAP7_75t_L g3242 ( 
.A(n_2931),
.Y(n_3242)
);

HB1xp67_ASAP7_75t_L g3243 ( 
.A(n_2934),
.Y(n_3243)
);

AND2x2_ASAP7_75t_L g3244 ( 
.A(n_2935),
.B(n_2546),
.Y(n_3244)
);

NAND2xp33_ASAP7_75t_L g3245 ( 
.A(n_2936),
.B(n_2745),
.Y(n_3245)
);

OAI22xp5_ASAP7_75t_L g3246 ( 
.A1(n_3047),
.A2(n_2461),
.B1(n_2470),
.B2(n_2442),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_2938),
.B(n_1875),
.Y(n_3247)
);

OA21x2_ASAP7_75t_L g3248 ( 
.A1(n_2939),
.A2(n_1894),
.B(n_1892),
.Y(n_3248)
);

INVx2_ASAP7_75t_L g3249 ( 
.A(n_2941),
.Y(n_3249)
);

BUFx6f_ASAP7_75t_L g3250 ( 
.A(n_2944),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_2946),
.Y(n_3251)
);

XOR2xp5_ASAP7_75t_L g3252 ( 
.A(n_2949),
.B(n_2471),
.Y(n_3252)
);

INVx2_ASAP7_75t_L g3253 ( 
.A(n_2950),
.Y(n_3253)
);

BUFx3_ASAP7_75t_L g3254 ( 
.A(n_2953),
.Y(n_3254)
);

BUFx3_ASAP7_75t_L g3255 ( 
.A(n_2957),
.Y(n_3255)
);

BUFx6f_ASAP7_75t_L g3256 ( 
.A(n_2958),
.Y(n_3256)
);

AOI22xp5_ASAP7_75t_SL g3257 ( 
.A1(n_2959),
.A2(n_2502),
.B1(n_2513),
.B2(n_2490),
.Y(n_3257)
);

INVx4_ASAP7_75t_L g3258 ( 
.A(n_2963),
.Y(n_3258)
);

INVx2_ASAP7_75t_L g3259 ( 
.A(n_2965),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_3119),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_L g3261 ( 
.A(n_3187),
.B(n_2967),
.Y(n_3261)
);

INVx2_ASAP7_75t_L g3262 ( 
.A(n_3084),
.Y(n_3262)
);

INVx3_ASAP7_75t_L g3263 ( 
.A(n_3135),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_3172),
.Y(n_3264)
);

INVx4_ASAP7_75t_L g3265 ( 
.A(n_3225),
.Y(n_3265)
);

INVx2_ASAP7_75t_L g3266 ( 
.A(n_3091),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_L g3267 ( 
.A(n_3229),
.B(n_2969),
.Y(n_3267)
);

INVx2_ASAP7_75t_L g3268 ( 
.A(n_3094),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_3173),
.Y(n_3269)
);

AND2x2_ASAP7_75t_L g3270 ( 
.A(n_3053),
.B(n_2975),
.Y(n_3270)
);

BUFx2_ASAP7_75t_L g3271 ( 
.A(n_3132),
.Y(n_3271)
);

OAI22xp5_ASAP7_75t_SL g3272 ( 
.A1(n_3097),
.A2(n_2536),
.B1(n_2595),
.B2(n_2519),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_3175),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_3177),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_L g3275 ( 
.A(n_3244),
.B(n_2977),
.Y(n_3275)
);

INVx2_ASAP7_75t_L g3276 ( 
.A(n_3113),
.Y(n_3276)
);

INVx1_ASAP7_75t_SL g3277 ( 
.A(n_3137),
.Y(n_3277)
);

INVx2_ASAP7_75t_L g3278 ( 
.A(n_3120),
.Y(n_3278)
);

INVx3_ASAP7_75t_L g3279 ( 
.A(n_3114),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_3191),
.Y(n_3280)
);

BUFx2_ASAP7_75t_L g3281 ( 
.A(n_3142),
.Y(n_3281)
);

HB1xp67_ASAP7_75t_L g3282 ( 
.A(n_3157),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_3195),
.Y(n_3283)
);

NOR2xp33_ASAP7_75t_L g3284 ( 
.A(n_3049),
.B(n_2978),
.Y(n_3284)
);

AND2x2_ASAP7_75t_L g3285 ( 
.A(n_3062),
.B(n_2979),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_3197),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_3200),
.Y(n_3287)
);

INVxp67_ASAP7_75t_L g3288 ( 
.A(n_3185),
.Y(n_3288)
);

INVx2_ASAP7_75t_L g3289 ( 
.A(n_3134),
.Y(n_3289)
);

BUFx6f_ASAP7_75t_L g3290 ( 
.A(n_3057),
.Y(n_3290)
);

BUFx6f_ASAP7_75t_L g3291 ( 
.A(n_3138),
.Y(n_3291)
);

INVx2_ASAP7_75t_L g3292 ( 
.A(n_3086),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_3204),
.Y(n_3293)
);

AND2x2_ASAP7_75t_L g3294 ( 
.A(n_3068),
.B(n_3186),
.Y(n_3294)
);

INVx2_ASAP7_75t_L g3295 ( 
.A(n_3092),
.Y(n_3295)
);

NOR2x1_ASAP7_75t_L g3296 ( 
.A(n_3140),
.B(n_2372),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_3210),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_3218),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_3228),
.Y(n_3299)
);

BUFx6f_ASAP7_75t_L g3300 ( 
.A(n_3143),
.Y(n_3300)
);

AND2x2_ASAP7_75t_L g3301 ( 
.A(n_3110),
.B(n_2980),
.Y(n_3301)
);

INVx2_ASAP7_75t_L g3302 ( 
.A(n_3096),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_3230),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_3232),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_3249),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_3125),
.B(n_2983),
.Y(n_3306)
);

INVx2_ASAP7_75t_L g3307 ( 
.A(n_3098),
.Y(n_3307)
);

OAI22xp5_ASAP7_75t_L g3308 ( 
.A1(n_3124),
.A2(n_2097),
.B1(n_2180),
.B2(n_2076),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_3253),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_3259),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_3144),
.Y(n_3311)
);

INVx1_ASAP7_75t_L g3312 ( 
.A(n_3149),
.Y(n_3312)
);

OAI22xp5_ASAP7_75t_SL g3313 ( 
.A1(n_3224),
.A2(n_2630),
.B1(n_2670),
.B2(n_2607),
.Y(n_3313)
);

INVx2_ASAP7_75t_L g3314 ( 
.A(n_3112),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_3155),
.Y(n_3315)
);

OAI22xp5_ASAP7_75t_L g3316 ( 
.A1(n_3099),
.A2(n_2532),
.B1(n_1734),
.B2(n_1977),
.Y(n_3316)
);

AND2x4_ASAP7_75t_L g3317 ( 
.A(n_3089),
.B(n_2984),
.Y(n_3317)
);

INVx2_ASAP7_75t_L g3318 ( 
.A(n_3117),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_3170),
.Y(n_3319)
);

AND2x4_ASAP7_75t_L g3320 ( 
.A(n_3176),
.B(n_2986),
.Y(n_3320)
);

NAND2x1_ASAP7_75t_L g3321 ( 
.A(n_3095),
.B(n_1901),
.Y(n_3321)
);

INVx2_ASAP7_75t_L g3322 ( 
.A(n_3121),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_3181),
.Y(n_3323)
);

HB1xp67_ASAP7_75t_L g3324 ( 
.A(n_3071),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_3189),
.Y(n_3325)
);

INVx2_ASAP7_75t_L g3326 ( 
.A(n_3131),
.Y(n_3326)
);

INVx3_ASAP7_75t_L g3327 ( 
.A(n_3194),
.Y(n_3327)
);

AND2x2_ASAP7_75t_L g3328 ( 
.A(n_3163),
.B(n_2987),
.Y(n_3328)
);

BUFx6f_ASAP7_75t_L g3329 ( 
.A(n_3209),
.Y(n_3329)
);

INVx2_ASAP7_75t_SL g3330 ( 
.A(n_3106),
.Y(n_3330)
);

AND2x2_ASAP7_75t_L g3331 ( 
.A(n_3069),
.B(n_2988),
.Y(n_3331)
);

BUFx12f_ASAP7_75t_L g3332 ( 
.A(n_3090),
.Y(n_3332)
);

BUFx12f_ASAP7_75t_L g3333 ( 
.A(n_3165),
.Y(n_3333)
);

BUFx2_ASAP7_75t_L g3334 ( 
.A(n_3087),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_3211),
.Y(n_3335)
);

INVx2_ASAP7_75t_L g3336 ( 
.A(n_3048),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_3233),
.Y(n_3337)
);

NOR2xp33_ASAP7_75t_L g3338 ( 
.A(n_3236),
.B(n_2989),
.Y(n_3338)
);

OAI22xp5_ASAP7_75t_L g3339 ( 
.A1(n_3235),
.A2(n_3079),
.B1(n_3243),
.B2(n_3078),
.Y(n_3339)
);

NAND2xp5_ASAP7_75t_L g3340 ( 
.A(n_3127),
.B(n_2990),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_L g3341 ( 
.A(n_3133),
.B(n_2991),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_3239),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_3250),
.Y(n_3343)
);

INVx2_ASAP7_75t_L g3344 ( 
.A(n_3063),
.Y(n_3344)
);

INVx2_ASAP7_75t_L g3345 ( 
.A(n_3077),
.Y(n_3345)
);

AND2x2_ASAP7_75t_L g3346 ( 
.A(n_3070),
.B(n_2995),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_3256),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_SL g3348 ( 
.A(n_3129),
.B(n_1730),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_3148),
.Y(n_3349)
);

INVx2_ASAP7_75t_L g3350 ( 
.A(n_3082),
.Y(n_3350)
);

BUFx2_ASAP7_75t_L g3351 ( 
.A(n_3103),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3162),
.Y(n_3352)
);

AND2x4_ASAP7_75t_L g3353 ( 
.A(n_3202),
.B(n_2996),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_3164),
.Y(n_3354)
);

AND2x2_ASAP7_75t_L g3355 ( 
.A(n_3050),
.B(n_2997),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_3188),
.Y(n_3356)
);

INVx2_ASAP7_75t_L g3357 ( 
.A(n_3083),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_3192),
.Y(n_3358)
);

NAND2xp33_ASAP7_75t_SL g3359 ( 
.A(n_3118),
.B(n_2675),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_3207),
.Y(n_3360)
);

AND2x4_ASAP7_75t_L g3361 ( 
.A(n_3076),
.B(n_2998),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3215),
.Y(n_3362)
);

INVx2_ASAP7_75t_L g3363 ( 
.A(n_3146),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_3219),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_3221),
.Y(n_3365)
);

INVx1_ASAP7_75t_L g3366 ( 
.A(n_3231),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_3234),
.Y(n_3367)
);

AND2x4_ASAP7_75t_L g3368 ( 
.A(n_3108),
.B(n_2999),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_3136),
.B(n_3000),
.Y(n_3369)
);

INVx2_ASAP7_75t_L g3370 ( 
.A(n_3139),
.Y(n_3370)
);

AND2x2_ASAP7_75t_L g3371 ( 
.A(n_3058),
.B(n_3001),
.Y(n_3371)
);

INVxp67_ASAP7_75t_L g3372 ( 
.A(n_3116),
.Y(n_3372)
);

BUFx2_ASAP7_75t_L g3373 ( 
.A(n_3183),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_3238),
.Y(n_3374)
);

AND2x4_ASAP7_75t_L g3375 ( 
.A(n_3061),
.B(n_3005),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_3251),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_3147),
.Y(n_3377)
);

INVx3_ASAP7_75t_L g3378 ( 
.A(n_3074),
.Y(n_3378)
);

INVx1_ASAP7_75t_L g3379 ( 
.A(n_3054),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_3059),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_3060),
.Y(n_3381)
);

HB1xp67_ASAP7_75t_L g3382 ( 
.A(n_3203),
.Y(n_3382)
);

INVx2_ASAP7_75t_L g3383 ( 
.A(n_3072),
.Y(n_3383)
);

INVx2_ASAP7_75t_L g3384 ( 
.A(n_3075),
.Y(n_3384)
);

AND2x2_ASAP7_75t_L g3385 ( 
.A(n_3122),
.B(n_3006),
.Y(n_3385)
);

AND2x2_ASAP7_75t_L g3386 ( 
.A(n_3051),
.B(n_3007),
.Y(n_3386)
);

INVx2_ASAP7_75t_L g3387 ( 
.A(n_3080),
.Y(n_3387)
);

INVx2_ASAP7_75t_L g3388 ( 
.A(n_3088),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_L g3389 ( 
.A(n_3093),
.B(n_3009),
.Y(n_3389)
);

INVx1_ASAP7_75t_L g3390 ( 
.A(n_3100),
.Y(n_3390)
);

INVx3_ASAP7_75t_L g3391 ( 
.A(n_3105),
.Y(n_3391)
);

AND2x2_ASAP7_75t_L g3392 ( 
.A(n_3126),
.B(n_3010),
.Y(n_3392)
);

INVx2_ASAP7_75t_L g3393 ( 
.A(n_3102),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_3115),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_3161),
.Y(n_3395)
);

BUFx6f_ASAP7_75t_L g3396 ( 
.A(n_3254),
.Y(n_3396)
);

INVx1_ASAP7_75t_L g3397 ( 
.A(n_3255),
.Y(n_3397)
);

BUFx2_ASAP7_75t_L g3398 ( 
.A(n_3206),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_3258),
.B(n_3011),
.Y(n_3399)
);

INVx2_ASAP7_75t_L g3400 ( 
.A(n_3153),
.Y(n_3400)
);

INVx3_ASAP7_75t_L g3401 ( 
.A(n_3160),
.Y(n_3401)
);

INVx2_ASAP7_75t_L g3402 ( 
.A(n_3222),
.Y(n_3402)
);

AND2x2_ASAP7_75t_L g3403 ( 
.A(n_3213),
.B(n_3014),
.Y(n_3403)
);

AND2x2_ASAP7_75t_L g3404 ( 
.A(n_3055),
.B(n_3017),
.Y(n_3404)
);

BUFx3_ASAP7_75t_L g3405 ( 
.A(n_3156),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3241),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_3242),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_3216),
.Y(n_3408)
);

INVx2_ASAP7_75t_L g3409 ( 
.A(n_3081),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3214),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_3248),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_3158),
.Y(n_3412)
);

AND2x4_ASAP7_75t_L g3413 ( 
.A(n_3167),
.B(n_3022),
.Y(n_3413)
);

BUFx6f_ASAP7_75t_L g3414 ( 
.A(n_3159),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_3104),
.Y(n_3415)
);

OAI21x1_ASAP7_75t_L g3416 ( 
.A1(n_3101),
.A2(n_1961),
.B(n_1960),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_3109),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_3174),
.Y(n_3418)
);

INVx2_ASAP7_75t_L g3419 ( 
.A(n_3141),
.Y(n_3419)
);

INVx2_ASAP7_75t_L g3420 ( 
.A(n_3201),
.Y(n_3420)
);

INVx2_ASAP7_75t_L g3421 ( 
.A(n_3205),
.Y(n_3421)
);

BUFx6f_ASAP7_75t_L g3422 ( 
.A(n_3168),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_3212),
.Y(n_3423)
);

HB1xp67_ASAP7_75t_L g3424 ( 
.A(n_3056),
.Y(n_3424)
);

INVx1_ASAP7_75t_L g3425 ( 
.A(n_3220),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3247),
.Y(n_3426)
);

AND2x4_ASAP7_75t_L g3427 ( 
.A(n_3169),
.B(n_3023),
.Y(n_3427)
);

INVx2_ASAP7_75t_L g3428 ( 
.A(n_3145),
.Y(n_3428)
);

INVx3_ASAP7_75t_L g3429 ( 
.A(n_3240),
.Y(n_3429)
);

NOR2xp33_ASAP7_75t_L g3430 ( 
.A(n_3073),
.B(n_3151),
.Y(n_3430)
);

INVx1_ASAP7_75t_L g3431 ( 
.A(n_3066),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_3085),
.Y(n_3432)
);

INVx2_ASAP7_75t_L g3433 ( 
.A(n_3111),
.Y(n_3433)
);

HB1xp67_ASAP7_75t_L g3434 ( 
.A(n_3199),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_L g3435 ( 
.A(n_3128),
.B(n_3026),
.Y(n_3435)
);

INVx2_ASAP7_75t_L g3436 ( 
.A(n_3179),
.Y(n_3436)
);

AND2x6_ASAP7_75t_L g3437 ( 
.A(n_3182),
.B(n_1970),
.Y(n_3437)
);

AND2x4_ASAP7_75t_L g3438 ( 
.A(n_3150),
.B(n_3028),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_3245),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3128),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_L g3441 ( 
.A(n_3130),
.B(n_3032),
.Y(n_3441)
);

CKINVDCx8_ASAP7_75t_R g3442 ( 
.A(n_3123),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_3130),
.Y(n_3443)
);

INVx1_ASAP7_75t_SL g3444 ( 
.A(n_3107),
.Y(n_3444)
);

INVx1_ASAP7_75t_L g3445 ( 
.A(n_3237),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_3166),
.Y(n_3446)
);

INVx1_ASAP7_75t_L g3447 ( 
.A(n_3190),
.Y(n_3447)
);

INVxp67_ASAP7_75t_L g3448 ( 
.A(n_3067),
.Y(n_3448)
);

INVx2_ASAP7_75t_L g3449 ( 
.A(n_3152),
.Y(n_3449)
);

INVxp67_ASAP7_75t_L g3450 ( 
.A(n_3223),
.Y(n_3450)
);

INVx1_ASAP7_75t_L g3451 ( 
.A(n_3184),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_3193),
.Y(n_3452)
);

BUFx6f_ASAP7_75t_L g3453 ( 
.A(n_3217),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_L g3454 ( 
.A(n_3180),
.B(n_3033),
.Y(n_3454)
);

INVx1_ASAP7_75t_L g3455 ( 
.A(n_3196),
.Y(n_3455)
);

INVx2_ASAP7_75t_L g3456 ( 
.A(n_3065),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_3246),
.Y(n_3457)
);

INVx3_ASAP7_75t_L g3458 ( 
.A(n_3227),
.Y(n_3458)
);

INVx3_ASAP7_75t_L g3459 ( 
.A(n_3198),
.Y(n_3459)
);

BUFx6f_ASAP7_75t_L g3460 ( 
.A(n_3208),
.Y(n_3460)
);

AND2x2_ASAP7_75t_L g3461 ( 
.A(n_3226),
.B(n_3034),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_3257),
.Y(n_3462)
);

INVx2_ASAP7_75t_L g3463 ( 
.A(n_3154),
.Y(n_3463)
);

INVxp67_ASAP7_75t_L g3464 ( 
.A(n_3064),
.Y(n_3464)
);

BUFx6f_ASAP7_75t_L g3465 ( 
.A(n_3178),
.Y(n_3465)
);

OA21x2_ASAP7_75t_L g3466 ( 
.A1(n_3171),
.A2(n_1997),
.B(n_1983),
.Y(n_3466)
);

INVx2_ASAP7_75t_L g3467 ( 
.A(n_3252),
.Y(n_3467)
);

INVx2_ASAP7_75t_L g3468 ( 
.A(n_3052),
.Y(n_3468)
);

INVx2_ASAP7_75t_L g3469 ( 
.A(n_3084),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_3119),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_3119),
.Y(n_3471)
);

BUFx6f_ASAP7_75t_L g3472 ( 
.A(n_3225),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3119),
.Y(n_3473)
);

XNOR2xp5_ASAP7_75t_L g3474 ( 
.A(n_3107),
.B(n_2689),
.Y(n_3474)
);

AND2x2_ASAP7_75t_L g3475 ( 
.A(n_3053),
.B(n_3035),
.Y(n_3475)
);

INVx2_ASAP7_75t_L g3476 ( 
.A(n_3084),
.Y(n_3476)
);

AND2x4_ASAP7_75t_L g3477 ( 
.A(n_3089),
.B(n_3036),
.Y(n_3477)
);

INVx2_ASAP7_75t_L g3478 ( 
.A(n_3084),
.Y(n_3478)
);

HB1xp67_ASAP7_75t_L g3479 ( 
.A(n_3132),
.Y(n_3479)
);

BUFx6f_ASAP7_75t_L g3480 ( 
.A(n_3225),
.Y(n_3480)
);

INVx2_ASAP7_75t_L g3481 ( 
.A(n_3084),
.Y(n_3481)
);

INVx3_ASAP7_75t_L g3482 ( 
.A(n_3135),
.Y(n_3482)
);

INVx1_ASAP7_75t_SL g3483 ( 
.A(n_3132),
.Y(n_3483)
);

INVx2_ASAP7_75t_L g3484 ( 
.A(n_3084),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_L g3485 ( 
.A(n_3187),
.B(n_3038),
.Y(n_3485)
);

INVx2_ASAP7_75t_L g3486 ( 
.A(n_3292),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3379),
.Y(n_3487)
);

OR2x2_ASAP7_75t_L g3488 ( 
.A(n_3277),
.B(n_2034),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_SL g3489 ( 
.A(n_3375),
.B(n_1739),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_SL g3490 ( 
.A(n_3294),
.B(n_1744),
.Y(n_3490)
);

INVx3_ASAP7_75t_L g3491 ( 
.A(n_3405),
.Y(n_3491)
);

INVx4_ASAP7_75t_SL g3492 ( 
.A(n_3453),
.Y(n_3492)
);

INVx1_ASAP7_75t_L g3493 ( 
.A(n_3380),
.Y(n_3493)
);

INVx2_ASAP7_75t_L g3494 ( 
.A(n_3295),
.Y(n_3494)
);

AOI22xp5_ASAP7_75t_L g3495 ( 
.A1(n_3430),
.A2(n_2072),
.B1(n_2717),
.B2(n_1971),
.Y(n_3495)
);

AND2x2_ASAP7_75t_L g3496 ( 
.A(n_3271),
.B(n_2703),
.Y(n_3496)
);

OR2x6_ASAP7_75t_L g3497 ( 
.A(n_3330),
.B(n_3039),
.Y(n_3497)
);

CKINVDCx5p33_ASAP7_75t_R g3498 ( 
.A(n_3332),
.Y(n_3498)
);

NOR2xp33_ASAP7_75t_L g3499 ( 
.A(n_3372),
.B(n_2107),
.Y(n_3499)
);

CKINVDCx6p67_ASAP7_75t_R g3500 ( 
.A(n_3333),
.Y(n_3500)
);

INVx2_ASAP7_75t_SL g3501 ( 
.A(n_3281),
.Y(n_3501)
);

AND2x2_ASAP7_75t_L g3502 ( 
.A(n_3483),
.B(n_2713),
.Y(n_3502)
);

INVx3_ASAP7_75t_L g3503 ( 
.A(n_3422),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3381),
.Y(n_3504)
);

INVx3_ASAP7_75t_L g3505 ( 
.A(n_3422),
.Y(n_3505)
);

INVx2_ASAP7_75t_L g3506 ( 
.A(n_3302),
.Y(n_3506)
);

INVx1_ASAP7_75t_SL g3507 ( 
.A(n_3444),
.Y(n_3507)
);

OAI22xp5_ASAP7_75t_L g3508 ( 
.A1(n_3408),
.A2(n_3423),
.B1(n_3425),
.B2(n_3418),
.Y(n_3508)
);

OR2x6_ASAP7_75t_L g3509 ( 
.A(n_3472),
.B(n_3040),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_L g3510 ( 
.A(n_3426),
.B(n_1825),
.Y(n_3510)
);

INVx2_ASAP7_75t_L g3511 ( 
.A(n_3307),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_L g3512 ( 
.A(n_3284),
.B(n_1839),
.Y(n_3512)
);

OAI22xp5_ASAP7_75t_L g3513 ( 
.A1(n_3412),
.A2(n_1747),
.B1(n_1754),
.B2(n_1746),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_L g3514 ( 
.A(n_3415),
.B(n_1975),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_SL g3515 ( 
.A(n_3339),
.B(n_1770),
.Y(n_3515)
);

NAND2xp5_ASAP7_75t_L g3516 ( 
.A(n_3417),
.B(n_3338),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_L g3517 ( 
.A(n_3270),
.B(n_2029),
.Y(n_3517)
);

NAND2xp5_ASAP7_75t_SL g3518 ( 
.A(n_3331),
.B(n_1772),
.Y(n_3518)
);

INVx5_ASAP7_75t_L g3519 ( 
.A(n_3472),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_SL g3520 ( 
.A(n_3346),
.B(n_1777),
.Y(n_3520)
);

INVxp67_ASAP7_75t_SL g3521 ( 
.A(n_3434),
.Y(n_3521)
);

INVx3_ASAP7_75t_L g3522 ( 
.A(n_3279),
.Y(n_3522)
);

NAND2xp5_ASAP7_75t_L g3523 ( 
.A(n_3285),
.B(n_2295),
.Y(n_3523)
);

OAI22xp5_ASAP7_75t_L g3524 ( 
.A1(n_3377),
.A2(n_1780),
.B1(n_1782),
.B2(n_1781),
.Y(n_3524)
);

INVx2_ASAP7_75t_L g3525 ( 
.A(n_3314),
.Y(n_3525)
);

AOI22xp33_ASAP7_75t_L g3526 ( 
.A1(n_3457),
.A2(n_3424),
.B1(n_3463),
.B2(n_3464),
.Y(n_3526)
);

BUFx6f_ASAP7_75t_L g3527 ( 
.A(n_3480),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_3475),
.B(n_2308),
.Y(n_3528)
);

AND2x2_ASAP7_75t_L g3529 ( 
.A(n_3355),
.B(n_3041),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_L g3530 ( 
.A(n_3301),
.B(n_2396),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_L g3531 ( 
.A(n_3261),
.B(n_2516),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_3390),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3394),
.Y(n_3533)
);

AND2x2_ASAP7_75t_L g3534 ( 
.A(n_3371),
.B(n_3043),
.Y(n_3534)
);

INVx2_ASAP7_75t_L g3535 ( 
.A(n_3318),
.Y(n_3535)
);

AOI22xp33_ASAP7_75t_L g3536 ( 
.A1(n_3383),
.A2(n_2260),
.B1(n_2353),
.B2(n_2340),
.Y(n_3536)
);

NAND2xp33_ASAP7_75t_SL g3537 ( 
.A(n_3460),
.B(n_3373),
.Y(n_3537)
);

BUFx3_ASAP7_75t_L g3538 ( 
.A(n_3453),
.Y(n_3538)
);

INVx2_ASAP7_75t_L g3539 ( 
.A(n_3322),
.Y(n_3539)
);

INVx6_ASAP7_75t_L g3540 ( 
.A(n_3480),
.Y(n_3540)
);

NOR2xp33_ASAP7_75t_L g3541 ( 
.A(n_3288),
.B(n_2380),
.Y(n_3541)
);

NOR3xp33_ASAP7_75t_L g3542 ( 
.A(n_3316),
.B(n_2445),
.C(n_2406),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_SL g3543 ( 
.A(n_3392),
.B(n_1785),
.Y(n_3543)
);

AOI22xp33_ASAP7_75t_L g3544 ( 
.A1(n_3384),
.A2(n_2511),
.B1(n_2531),
.B2(n_2492),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3387),
.Y(n_3545)
);

AOI22xp33_ASAP7_75t_L g3546 ( 
.A1(n_3388),
.A2(n_2585),
.B1(n_2604),
.B2(n_2556),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_SL g3547 ( 
.A(n_3267),
.B(n_1787),
.Y(n_3547)
);

INVx1_ASAP7_75t_L g3548 ( 
.A(n_3393),
.Y(n_3548)
);

OAI22xp5_ASAP7_75t_L g3549 ( 
.A1(n_3275),
.A2(n_1788),
.B1(n_1794),
.B2(n_1789),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_3485),
.B(n_2640),
.Y(n_3550)
);

BUFx10_ASAP7_75t_L g3551 ( 
.A(n_3460),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3349),
.Y(n_3552)
);

AND2x2_ASAP7_75t_L g3553 ( 
.A(n_3282),
.B(n_3046),
.Y(n_3553)
);

INVx2_ASAP7_75t_L g3554 ( 
.A(n_3326),
.Y(n_3554)
);

NOR2xp33_ASAP7_75t_L g3555 ( 
.A(n_3454),
.B(n_2712),
.Y(n_3555)
);

NAND2xp5_ASAP7_75t_SL g3556 ( 
.A(n_3396),
.B(n_1801),
.Y(n_3556)
);

INVx3_ASAP7_75t_L g3557 ( 
.A(n_3291),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_L g3558 ( 
.A(n_3386),
.B(n_2731),
.Y(n_3558)
);

INVx5_ASAP7_75t_L g3559 ( 
.A(n_3265),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3352),
.Y(n_3560)
);

INVx5_ASAP7_75t_L g3561 ( 
.A(n_3459),
.Y(n_3561)
);

BUFx6f_ASAP7_75t_SL g3562 ( 
.A(n_3446),
.Y(n_3562)
);

INVx5_ASAP7_75t_L g3563 ( 
.A(n_3334),
.Y(n_3563)
);

NOR3xp33_ASAP7_75t_L g3564 ( 
.A(n_3398),
.B(n_2769),
.C(n_2751),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3354),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_SL g3566 ( 
.A(n_3396),
.B(n_1802),
.Y(n_3566)
);

INVx2_ASAP7_75t_L g3567 ( 
.A(n_3363),
.Y(n_3567)
);

INVx1_ASAP7_75t_SL g3568 ( 
.A(n_3479),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3356),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_3358),
.Y(n_3570)
);

CKINVDCx14_ASAP7_75t_R g3571 ( 
.A(n_3474),
.Y(n_3571)
);

INVx2_ASAP7_75t_L g3572 ( 
.A(n_3264),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3360),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_3362),
.Y(n_3574)
);

INVxp33_ASAP7_75t_SL g3575 ( 
.A(n_3382),
.Y(n_3575)
);

AND2x2_ASAP7_75t_L g3576 ( 
.A(n_3328),
.B(n_1735),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3364),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3365),
.Y(n_3578)
);

AND2x2_ASAP7_75t_L g3579 ( 
.A(n_3404),
.B(n_1735),
.Y(n_3579)
);

BUFx10_ASAP7_75t_L g3580 ( 
.A(n_3317),
.Y(n_3580)
);

INVx1_ASAP7_75t_L g3581 ( 
.A(n_3366),
.Y(n_3581)
);

NOR2xp33_ASAP7_75t_L g3582 ( 
.A(n_3451),
.B(n_2782),
.Y(n_3582)
);

AND2x2_ASAP7_75t_L g3583 ( 
.A(n_3353),
.B(n_3461),
.Y(n_3583)
);

INVx2_ASAP7_75t_L g3584 ( 
.A(n_3269),
.Y(n_3584)
);

NOR2xp33_ASAP7_75t_L g3585 ( 
.A(n_3452),
.B(n_1808),
.Y(n_3585)
);

BUFx10_ASAP7_75t_L g3586 ( 
.A(n_3320),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_3367),
.Y(n_3587)
);

INVx1_ASAP7_75t_SL g3588 ( 
.A(n_3351),
.Y(n_3588)
);

INVx2_ASAP7_75t_L g3589 ( 
.A(n_3273),
.Y(n_3589)
);

INVx2_ASAP7_75t_L g3590 ( 
.A(n_3274),
.Y(n_3590)
);

NOR2xp33_ASAP7_75t_L g3591 ( 
.A(n_3455),
.B(n_3324),
.Y(n_3591)
);

INVx4_ASAP7_75t_L g3592 ( 
.A(n_3291),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_3374),
.Y(n_3593)
);

OR2x6_ASAP7_75t_L g3594 ( 
.A(n_3465),
.B(n_2253),
.Y(n_3594)
);

OR2x2_ASAP7_75t_L g3595 ( 
.A(n_3450),
.B(n_2290),
.Y(n_3595)
);

INVx1_ASAP7_75t_L g3596 ( 
.A(n_3376),
.Y(n_3596)
);

INVx4_ASAP7_75t_L g3597 ( 
.A(n_3300),
.Y(n_3597)
);

INVx6_ASAP7_75t_L g3598 ( 
.A(n_3465),
.Y(n_3598)
);

AOI22xp33_ASAP7_75t_L g3599 ( 
.A1(n_3260),
.A2(n_3470),
.B1(n_3473),
.B2(n_3471),
.Y(n_3599)
);

INVx5_ASAP7_75t_L g3600 ( 
.A(n_3458),
.Y(n_3600)
);

BUFx10_ASAP7_75t_L g3601 ( 
.A(n_3477),
.Y(n_3601)
);

NOR2xp33_ASAP7_75t_L g3602 ( 
.A(n_3370),
.B(n_1810),
.Y(n_3602)
);

BUFx10_ASAP7_75t_L g3603 ( 
.A(n_3368),
.Y(n_3603)
);

BUFx6f_ASAP7_75t_L g3604 ( 
.A(n_3300),
.Y(n_3604)
);

INVx4_ASAP7_75t_L g3605 ( 
.A(n_3329),
.Y(n_3605)
);

INVx2_ASAP7_75t_L g3606 ( 
.A(n_3280),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_3283),
.Y(n_3607)
);

INVx2_ASAP7_75t_L g3608 ( 
.A(n_3286),
.Y(n_3608)
);

INVx5_ASAP7_75t_L g3609 ( 
.A(n_3329),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3287),
.Y(n_3610)
);

OAI21xp5_ASAP7_75t_L g3611 ( 
.A1(n_3409),
.A2(n_2019),
.B(n_2016),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_SL g3612 ( 
.A(n_3401),
.B(n_1812),
.Y(n_3612)
);

NOR2xp33_ASAP7_75t_L g3613 ( 
.A(n_3378),
.B(n_3391),
.Y(n_3613)
);

BUFx8_ASAP7_75t_SL g3614 ( 
.A(n_3263),
.Y(n_3614)
);

INVx3_ASAP7_75t_L g3615 ( 
.A(n_3442),
.Y(n_3615)
);

BUFx2_ASAP7_75t_L g3616 ( 
.A(n_3359),
.Y(n_3616)
);

INVx2_ASAP7_75t_SL g3617 ( 
.A(n_3403),
.Y(n_3617)
);

INVx1_ASAP7_75t_L g3618 ( 
.A(n_3293),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_SL g3619 ( 
.A(n_3449),
.B(n_1814),
.Y(n_3619)
);

NAND2xp5_ASAP7_75t_L g3620 ( 
.A(n_3297),
.B(n_2324),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_SL g3621 ( 
.A(n_3435),
.B(n_1818),
.Y(n_3621)
);

NAND2xp5_ASAP7_75t_L g3622 ( 
.A(n_3298),
.B(n_2408),
.Y(n_3622)
);

NAND2xp5_ASAP7_75t_SL g3623 ( 
.A(n_3441),
.B(n_1819),
.Y(n_3623)
);

NOR2xp33_ASAP7_75t_L g3624 ( 
.A(n_3395),
.B(n_1822),
.Y(n_3624)
);

INVx1_ASAP7_75t_L g3625 ( 
.A(n_3299),
.Y(n_3625)
);

NAND2xp5_ASAP7_75t_L g3626 ( 
.A(n_3303),
.B(n_3304),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_L g3627 ( 
.A(n_3305),
.B(n_2476),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_SL g3628 ( 
.A(n_3361),
.B(n_1824),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_3309),
.Y(n_3629)
);

INVx5_ASAP7_75t_L g3630 ( 
.A(n_3482),
.Y(n_3630)
);

INVx1_ASAP7_75t_SL g3631 ( 
.A(n_3385),
.Y(n_3631)
);

INVx4_ASAP7_75t_L g3632 ( 
.A(n_3290),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_3310),
.B(n_2619),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_SL g3634 ( 
.A(n_3399),
.B(n_1828),
.Y(n_3634)
);

NOR2xp33_ASAP7_75t_L g3635 ( 
.A(n_3397),
.B(n_1829),
.Y(n_3635)
);

NOR2xp33_ASAP7_75t_SL g3636 ( 
.A(n_3448),
.B(n_2546),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_SL g3637 ( 
.A(n_3413),
.B(n_1834),
.Y(n_3637)
);

NOR2xp33_ASAP7_75t_L g3638 ( 
.A(n_3431),
.B(n_1840),
.Y(n_3638)
);

AND2x6_ASAP7_75t_L g3639 ( 
.A(n_3440),
.B(n_2560),
.Y(n_3639)
);

INVxp33_ASAP7_75t_SL g3640 ( 
.A(n_3308),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3306),
.Y(n_3641)
);

INVx1_ASAP7_75t_L g3642 ( 
.A(n_3340),
.Y(n_3642)
);

INVx4_ASAP7_75t_L g3643 ( 
.A(n_3290),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3341),
.Y(n_3644)
);

NOR2xp33_ASAP7_75t_L g3645 ( 
.A(n_3428),
.B(n_1841),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3369),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_L g3647 ( 
.A(n_3406),
.B(n_2676),
.Y(n_3647)
);

NAND2xp5_ASAP7_75t_SL g3648 ( 
.A(n_3427),
.B(n_1842),
.Y(n_3648)
);

BUFx3_ASAP7_75t_L g3649 ( 
.A(n_3327),
.Y(n_3649)
);

INVx2_ASAP7_75t_L g3650 ( 
.A(n_3400),
.Y(n_3650)
);

BUFx6f_ASAP7_75t_L g3651 ( 
.A(n_3262),
.Y(n_3651)
);

AOI22xp33_ASAP7_75t_L g3652 ( 
.A1(n_3313),
.A2(n_2718),
.B1(n_2692),
.B2(n_2626),
.Y(n_3652)
);

INVx1_ASAP7_75t_L g3653 ( 
.A(n_3402),
.Y(n_3653)
);

NOR2xp33_ASAP7_75t_L g3654 ( 
.A(n_3436),
.B(n_1845),
.Y(n_3654)
);

BUFx4f_ASAP7_75t_L g3655 ( 
.A(n_3447),
.Y(n_3655)
);

NOR2xp33_ASAP7_75t_SL g3656 ( 
.A(n_3272),
.B(n_2626),
.Y(n_3656)
);

BUFx4f_ASAP7_75t_L g3657 ( 
.A(n_3437),
.Y(n_3657)
);

OR2x6_ASAP7_75t_L g3658 ( 
.A(n_3468),
.B(n_2570),
.Y(n_3658)
);

INVx2_ASAP7_75t_SL g3659 ( 
.A(n_3438),
.Y(n_3659)
);

INVx2_ASAP7_75t_L g3660 ( 
.A(n_3336),
.Y(n_3660)
);

INVx1_ASAP7_75t_SL g3661 ( 
.A(n_3467),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_SL g3662 ( 
.A(n_3443),
.B(n_1849),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_SL g3663 ( 
.A(n_3296),
.B(n_1852),
.Y(n_3663)
);

NAND2xp5_ASAP7_75t_L g3664 ( 
.A(n_3407),
.B(n_2745),
.Y(n_3664)
);

BUFx10_ASAP7_75t_L g3665 ( 
.A(n_3437),
.Y(n_3665)
);

INVx4_ASAP7_75t_L g3666 ( 
.A(n_3429),
.Y(n_3666)
);

AND2x4_ASAP7_75t_L g3667 ( 
.A(n_3311),
.B(n_2571),
.Y(n_3667)
);

AND2x2_ASAP7_75t_L g3668 ( 
.A(n_3445),
.B(n_1806),
.Y(n_3668)
);

INVx2_ASAP7_75t_L g3669 ( 
.A(n_3344),
.Y(n_3669)
);

NAND2xp33_ASAP7_75t_R g3670 ( 
.A(n_3462),
.B(n_1856),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3389),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_SL g3672 ( 
.A(n_3348),
.B(n_3414),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_3345),
.Y(n_3673)
);

BUFx10_ASAP7_75t_L g3674 ( 
.A(n_3437),
.Y(n_3674)
);

INVx2_ASAP7_75t_L g3675 ( 
.A(n_3350),
.Y(n_3675)
);

INVx2_ASAP7_75t_L g3676 ( 
.A(n_3357),
.Y(n_3676)
);

INVx1_ASAP7_75t_L g3677 ( 
.A(n_3439),
.Y(n_3677)
);

NAND2x1p5_ASAP7_75t_L g3678 ( 
.A(n_3312),
.B(n_2587),
.Y(n_3678)
);

INVx2_ASAP7_75t_L g3679 ( 
.A(n_3419),
.Y(n_3679)
);

AND2x4_ASAP7_75t_L g3680 ( 
.A(n_3315),
.B(n_2596),
.Y(n_3680)
);

NAND2xp5_ASAP7_75t_SL g3681 ( 
.A(n_3414),
.B(n_1862),
.Y(n_3681)
);

INVx2_ASAP7_75t_L g3682 ( 
.A(n_3410),
.Y(n_3682)
);

INVx4_ASAP7_75t_L g3683 ( 
.A(n_3266),
.Y(n_3683)
);

NAND2xp5_ASAP7_75t_SL g3684 ( 
.A(n_3319),
.B(n_1863),
.Y(n_3684)
);

AOI22xp33_ASAP7_75t_L g3685 ( 
.A1(n_3411),
.A2(n_2692),
.B1(n_1919),
.B2(n_1947),
.Y(n_3685)
);

INVx5_ASAP7_75t_L g3686 ( 
.A(n_3268),
.Y(n_3686)
);

CKINVDCx20_ASAP7_75t_R g3687 ( 
.A(n_3466),
.Y(n_3687)
);

INVx2_ASAP7_75t_L g3688 ( 
.A(n_3276),
.Y(n_3688)
);

INVx5_ASAP7_75t_L g3689 ( 
.A(n_3278),
.Y(n_3689)
);

INVx2_ASAP7_75t_L g3690 ( 
.A(n_3289),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_3321),
.Y(n_3691)
);

BUFx10_ASAP7_75t_L g3692 ( 
.A(n_3323),
.Y(n_3692)
);

OAI22xp5_ASAP7_75t_L g3693 ( 
.A1(n_3432),
.A2(n_1876),
.B1(n_1879),
.B2(n_1871),
.Y(n_3693)
);

INVx5_ASAP7_75t_L g3694 ( 
.A(n_3469),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3476),
.Y(n_3695)
);

INVx3_ASAP7_75t_L g3696 ( 
.A(n_3478),
.Y(n_3696)
);

NAND2xp33_ASAP7_75t_L g3697 ( 
.A(n_3433),
.B(n_1887),
.Y(n_3697)
);

OR2x2_ASAP7_75t_L g3698 ( 
.A(n_3325),
.B(n_2600),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_3481),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3484),
.Y(n_3700)
);

BUFx6f_ASAP7_75t_L g3701 ( 
.A(n_3335),
.Y(n_3701)
);

INVx1_ASAP7_75t_L g3702 ( 
.A(n_3337),
.Y(n_3702)
);

INVx4_ASAP7_75t_L g3703 ( 
.A(n_3342),
.Y(n_3703)
);

INVx3_ASAP7_75t_L g3704 ( 
.A(n_3343),
.Y(n_3704)
);

NAND2xp5_ASAP7_75t_SL g3705 ( 
.A(n_3347),
.B(n_1888),
.Y(n_3705)
);

BUFx10_ASAP7_75t_L g3706 ( 
.A(n_3456),
.Y(n_3706)
);

AOI22xp5_ASAP7_75t_L g3707 ( 
.A1(n_3420),
.A2(n_2330),
.B1(n_2362),
.B2(n_2028),
.Y(n_3707)
);

INVx1_ASAP7_75t_L g3708 ( 
.A(n_3421),
.Y(n_3708)
);

INVx3_ASAP7_75t_L g3709 ( 
.A(n_3416),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_3379),
.Y(n_3710)
);

NOR2xp33_ASAP7_75t_L g3711 ( 
.A(n_3372),
.B(n_1891),
.Y(n_3711)
);

AND3x2_ASAP7_75t_L g3712 ( 
.A(n_3373),
.B(n_2001),
.C(n_1909),
.Y(n_3712)
);

AND2x2_ASAP7_75t_L g3713 ( 
.A(n_3271),
.B(n_1806),
.Y(n_3713)
);

INVx3_ASAP7_75t_L g3714 ( 
.A(n_3405),
.Y(n_3714)
);

INVx1_ASAP7_75t_L g3715 ( 
.A(n_3379),
.Y(n_3715)
);

AND2x2_ASAP7_75t_L g3716 ( 
.A(n_3271),
.B(n_1873),
.Y(n_3716)
);

INVx2_ASAP7_75t_L g3717 ( 
.A(n_3292),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3379),
.Y(n_3718)
);

INVx3_ASAP7_75t_L g3719 ( 
.A(n_3405),
.Y(n_3719)
);

AOI22xp33_ASAP7_75t_L g3720 ( 
.A1(n_3457),
.A2(n_2033),
.B1(n_2038),
.B2(n_2020),
.Y(n_3720)
);

AND2x2_ASAP7_75t_L g3721 ( 
.A(n_3271),
.B(n_1873),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_L g3722 ( 
.A(n_3430),
.B(n_1895),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_3379),
.Y(n_3723)
);

INVx3_ASAP7_75t_L g3724 ( 
.A(n_3405),
.Y(n_3724)
);

NAND2xp5_ASAP7_75t_L g3725 ( 
.A(n_3430),
.B(n_1897),
.Y(n_3725)
);

INVx4_ASAP7_75t_L g3726 ( 
.A(n_3472),
.Y(n_3726)
);

NOR2xp33_ASAP7_75t_L g3727 ( 
.A(n_3372),
.B(n_1898),
.Y(n_3727)
);

INVx3_ASAP7_75t_L g3728 ( 
.A(n_3405),
.Y(n_3728)
);

INVx1_ASAP7_75t_L g3729 ( 
.A(n_3379),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_L g3730 ( 
.A(n_3430),
.B(n_1907),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_L g3731 ( 
.A(n_3430),
.B(n_1910),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_3379),
.Y(n_3732)
);

BUFx3_ASAP7_75t_L g3733 ( 
.A(n_3332),
.Y(n_3733)
);

INVx2_ASAP7_75t_L g3734 ( 
.A(n_3292),
.Y(n_3734)
);

AOI22xp5_ASAP7_75t_L g3735 ( 
.A1(n_3430),
.A2(n_2786),
.B1(n_2434),
.B2(n_2041),
.Y(n_3735)
);

INVx2_ASAP7_75t_L g3736 ( 
.A(n_3292),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_L g3737 ( 
.A(n_3430),
.B(n_1913),
.Y(n_3737)
);

INVx6_ASAP7_75t_L g3738 ( 
.A(n_3453),
.Y(n_3738)
);

INVx4_ASAP7_75t_L g3739 ( 
.A(n_3472),
.Y(n_3739)
);

INVx3_ASAP7_75t_L g3740 ( 
.A(n_3405),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_L g3741 ( 
.A(n_3430),
.B(n_1917),
.Y(n_3741)
);

OR2x2_ASAP7_75t_L g3742 ( 
.A(n_3277),
.B(n_2602),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_SL g3743 ( 
.A(n_3375),
.B(n_1920),
.Y(n_3743)
);

NAND2xp5_ASAP7_75t_SL g3744 ( 
.A(n_3375),
.B(n_1924),
.Y(n_3744)
);

INVx3_ASAP7_75t_L g3745 ( 
.A(n_3405),
.Y(n_3745)
);

INVx3_ASAP7_75t_L g3746 ( 
.A(n_3405),
.Y(n_3746)
);

BUFx4f_ASAP7_75t_L g3747 ( 
.A(n_3453),
.Y(n_3747)
);

AND2x6_ASAP7_75t_L g3748 ( 
.A(n_3294),
.B(n_2611),
.Y(n_3748)
);

INVx2_ASAP7_75t_L g3749 ( 
.A(n_3292),
.Y(n_3749)
);

BUFx10_ASAP7_75t_L g3750 ( 
.A(n_3453),
.Y(n_3750)
);

AND2x4_ASAP7_75t_L g3751 ( 
.A(n_3330),
.B(n_2614),
.Y(n_3751)
);

AOI22xp33_ASAP7_75t_L g3752 ( 
.A1(n_3457),
.A2(n_2047),
.B1(n_2077),
.B2(n_2054),
.Y(n_3752)
);

INVx2_ASAP7_75t_L g3753 ( 
.A(n_3292),
.Y(n_3753)
);

INVx2_ASAP7_75t_L g3754 ( 
.A(n_3292),
.Y(n_3754)
);

BUFx10_ASAP7_75t_L g3755 ( 
.A(n_3453),
.Y(n_3755)
);

NAND2xp5_ASAP7_75t_L g3756 ( 
.A(n_3430),
.B(n_1927),
.Y(n_3756)
);

BUFx3_ASAP7_75t_L g3757 ( 
.A(n_3332),
.Y(n_3757)
);

OR2x6_ASAP7_75t_L g3758 ( 
.A(n_3330),
.B(n_2616),
.Y(n_3758)
);

NAND2xp33_ASAP7_75t_L g3759 ( 
.A(n_3449),
.B(n_1934),
.Y(n_3759)
);

AND3x2_ASAP7_75t_L g3760 ( 
.A(n_3373),
.B(n_2147),
.C(n_2124),
.Y(n_3760)
);

NAND2xp5_ASAP7_75t_L g3761 ( 
.A(n_3430),
.B(n_1938),
.Y(n_3761)
);

NAND2xp5_ASAP7_75t_L g3762 ( 
.A(n_3430),
.B(n_1943),
.Y(n_3762)
);

NOR2xp33_ASAP7_75t_L g3763 ( 
.A(n_3372),
.B(n_1946),
.Y(n_3763)
);

INVx4_ASAP7_75t_L g3764 ( 
.A(n_3472),
.Y(n_3764)
);

INVx5_ASAP7_75t_L g3765 ( 
.A(n_3472),
.Y(n_3765)
);

AND2x4_ASAP7_75t_L g3766 ( 
.A(n_3330),
.B(n_2620),
.Y(n_3766)
);

INVx2_ASAP7_75t_L g3767 ( 
.A(n_3292),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_3379),
.Y(n_3768)
);

INVx1_ASAP7_75t_SL g3769 ( 
.A(n_3277),
.Y(n_3769)
);

NAND2x1p5_ASAP7_75t_L g3770 ( 
.A(n_3265),
.B(n_2636),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_3379),
.Y(n_3771)
);

BUFx6f_ASAP7_75t_L g3772 ( 
.A(n_3472),
.Y(n_3772)
);

INVx2_ASAP7_75t_L g3773 ( 
.A(n_3292),
.Y(n_3773)
);

INVx1_ASAP7_75t_L g3774 ( 
.A(n_3379),
.Y(n_3774)
);

AND2x6_ASAP7_75t_L g3775 ( 
.A(n_3294),
.B(n_2637),
.Y(n_3775)
);

INVx4_ASAP7_75t_L g3776 ( 
.A(n_3472),
.Y(n_3776)
);

INVx2_ASAP7_75t_L g3777 ( 
.A(n_3292),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_L g3778 ( 
.A(n_3430),
.B(n_1949),
.Y(n_3778)
);

INVx2_ASAP7_75t_L g3779 ( 
.A(n_3292),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_SL g3780 ( 
.A(n_3375),
.B(n_1950),
.Y(n_3780)
);

BUFx6f_ASAP7_75t_L g3781 ( 
.A(n_3472),
.Y(n_3781)
);

BUFx6f_ASAP7_75t_L g3782 ( 
.A(n_3472),
.Y(n_3782)
);

AND2x4_ASAP7_75t_L g3783 ( 
.A(n_3330),
.B(n_2638),
.Y(n_3783)
);

INVx5_ASAP7_75t_L g3784 ( 
.A(n_3472),
.Y(n_3784)
);

NOR2xp33_ASAP7_75t_L g3785 ( 
.A(n_3372),
.B(n_1953),
.Y(n_3785)
);

NAND2xp33_ASAP7_75t_L g3786 ( 
.A(n_3516),
.B(n_1955),
.Y(n_3786)
);

AOI22xp33_ASAP7_75t_L g3787 ( 
.A1(n_3640),
.A2(n_2179),
.B1(n_2301),
.B2(n_1881),
.Y(n_3787)
);

INVx2_ASAP7_75t_L g3788 ( 
.A(n_3679),
.Y(n_3788)
);

NAND2xp5_ASAP7_75t_SL g3789 ( 
.A(n_3588),
.B(n_3508),
.Y(n_3789)
);

NAND2xp5_ASAP7_75t_SL g3790 ( 
.A(n_3575),
.B(n_1958),
.Y(n_3790)
);

NOR3xp33_ASAP7_75t_L g3791 ( 
.A(n_3722),
.B(n_2645),
.C(n_2639),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_L g3792 ( 
.A(n_3512),
.B(n_2652),
.Y(n_3792)
);

OAI22xp5_ASAP7_75t_L g3793 ( 
.A1(n_3725),
.A2(n_1967),
.B1(n_1968),
.B2(n_1965),
.Y(n_3793)
);

NAND2xp5_ASAP7_75t_SL g3794 ( 
.A(n_3657),
.B(n_1969),
.Y(n_3794)
);

NAND2xp5_ASAP7_75t_SL g3795 ( 
.A(n_3501),
.B(n_1972),
.Y(n_3795)
);

NOR2xp33_ASAP7_75t_L g3796 ( 
.A(n_3521),
.B(n_1973),
.Y(n_3796)
);

INVx5_ASAP7_75t_L g3797 ( 
.A(n_3665),
.Y(n_3797)
);

NAND2xp5_ASAP7_75t_L g3798 ( 
.A(n_3730),
.B(n_2653),
.Y(n_3798)
);

OAI21xp5_ASAP7_75t_L g3799 ( 
.A1(n_3611),
.A2(n_2048),
.B(n_2032),
.Y(n_3799)
);

INVx3_ASAP7_75t_L g3800 ( 
.A(n_3750),
.Y(n_3800)
);

BUFx3_ASAP7_75t_L g3801 ( 
.A(n_3738),
.Y(n_3801)
);

INVxp67_ASAP7_75t_L g3802 ( 
.A(n_3769),
.Y(n_3802)
);

CKINVDCx11_ASAP7_75t_R g3803 ( 
.A(n_3755),
.Y(n_3803)
);

OAI22xp5_ASAP7_75t_L g3804 ( 
.A1(n_3731),
.A2(n_1986),
.B1(n_1987),
.B2(n_1985),
.Y(n_3804)
);

NAND2xp5_ASAP7_75t_SL g3805 ( 
.A(n_3561),
.B(n_2000),
.Y(n_3805)
);

NOR2xp33_ASAP7_75t_L g3806 ( 
.A(n_3568),
.B(n_2003),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_3487),
.Y(n_3807)
);

NAND2xp5_ASAP7_75t_L g3808 ( 
.A(n_3737),
.B(n_2678),
.Y(n_3808)
);

NAND2xp5_ASAP7_75t_L g3809 ( 
.A(n_3741),
.B(n_2681),
.Y(n_3809)
);

INVx2_ASAP7_75t_L g3810 ( 
.A(n_3486),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_SL g3811 ( 
.A(n_3561),
.B(n_2004),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_L g3812 ( 
.A(n_3756),
.B(n_3761),
.Y(n_3812)
);

OR2x2_ASAP7_75t_L g3813 ( 
.A(n_3631),
.B(n_2682),
.Y(n_3813)
);

NOR2xp33_ASAP7_75t_SL g3814 ( 
.A(n_3498),
.B(n_1881),
.Y(n_3814)
);

INVx3_ASAP7_75t_L g3815 ( 
.A(n_3551),
.Y(n_3815)
);

NAND2xp5_ASAP7_75t_L g3816 ( 
.A(n_3762),
.B(n_2684),
.Y(n_3816)
);

NAND2xp5_ASAP7_75t_L g3817 ( 
.A(n_3778),
.B(n_2685),
.Y(n_3817)
);

O2A1O1Ixp5_ASAP7_75t_L g3818 ( 
.A1(n_3681),
.A2(n_3672),
.B(n_3634),
.C(n_3547),
.Y(n_3818)
);

NOR2xp67_ASAP7_75t_L g3819 ( 
.A(n_3519),
.B(n_2063),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_SL g3820 ( 
.A(n_3563),
.B(n_2005),
.Y(n_3820)
);

OAI21xp5_ASAP7_75t_L g3821 ( 
.A1(n_3708),
.A2(n_2091),
.B(n_2087),
.Y(n_3821)
);

NAND2xp5_ASAP7_75t_SL g3822 ( 
.A(n_3563),
.B(n_2007),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_SL g3823 ( 
.A(n_3600),
.B(n_2008),
.Y(n_3823)
);

INVx2_ASAP7_75t_L g3824 ( 
.A(n_3494),
.Y(n_3824)
);

INVxp33_ASAP7_75t_L g3825 ( 
.A(n_3502),
.Y(n_3825)
);

NAND2xp5_ASAP7_75t_L g3826 ( 
.A(n_3671),
.B(n_2699),
.Y(n_3826)
);

INVx2_ASAP7_75t_L g3827 ( 
.A(n_3506),
.Y(n_3827)
);

OAI22xp5_ASAP7_75t_L g3828 ( 
.A1(n_3495),
.A2(n_2012),
.B1(n_2021),
.B2(n_2011),
.Y(n_3828)
);

O2A1O1Ixp33_ASAP7_75t_L g3829 ( 
.A1(n_3711),
.A2(n_2715),
.B(n_2727),
.C(n_2704),
.Y(n_3829)
);

CKINVDCx5p33_ASAP7_75t_R g3830 ( 
.A(n_3500),
.Y(n_3830)
);

HB1xp67_ASAP7_75t_L g3831 ( 
.A(n_3507),
.Y(n_3831)
);

NAND2xp5_ASAP7_75t_L g3832 ( 
.A(n_3641),
.B(n_2736),
.Y(n_3832)
);

INVx1_ASAP7_75t_L g3833 ( 
.A(n_3493),
.Y(n_3833)
);

NOR2xp33_ASAP7_75t_L g3834 ( 
.A(n_3499),
.B(n_2023),
.Y(n_3834)
);

NAND2xp5_ASAP7_75t_L g3835 ( 
.A(n_3642),
.B(n_3644),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_L g3836 ( 
.A(n_3646),
.B(n_2748),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_3514),
.B(n_2755),
.Y(n_3837)
);

INVx2_ASAP7_75t_L g3838 ( 
.A(n_3511),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_3504),
.Y(n_3839)
);

AND2x2_ASAP7_75t_L g3840 ( 
.A(n_3583),
.B(n_2179),
.Y(n_3840)
);

INVx2_ASAP7_75t_L g3841 ( 
.A(n_3525),
.Y(n_3841)
);

OR2x2_ASAP7_75t_L g3842 ( 
.A(n_3488),
.B(n_2760),
.Y(n_3842)
);

NOR3xp33_ASAP7_75t_L g3843 ( 
.A(n_3591),
.B(n_3763),
.C(n_3727),
.Y(n_3843)
);

NAND2xp5_ASAP7_75t_L g3844 ( 
.A(n_3555),
.B(n_2761),
.Y(n_3844)
);

INVxp67_ASAP7_75t_SL g3845 ( 
.A(n_3491),
.Y(n_3845)
);

NAND2xp5_ASAP7_75t_L g3846 ( 
.A(n_3510),
.B(n_2768),
.Y(n_3846)
);

NOR2xp33_ASAP7_75t_L g3847 ( 
.A(n_3785),
.B(n_2027),
.Y(n_3847)
);

INVx2_ASAP7_75t_L g3848 ( 
.A(n_3535),
.Y(n_3848)
);

NAND2xp5_ASAP7_75t_L g3849 ( 
.A(n_3529),
.B(n_2780),
.Y(n_3849)
);

INVx1_ASAP7_75t_L g3850 ( 
.A(n_3532),
.Y(n_3850)
);

A2O1A1Ixp33_ASAP7_75t_L g3851 ( 
.A1(n_3735),
.A2(n_2119),
.B(n_2128),
.C(n_2116),
.Y(n_3851)
);

INVx2_ASAP7_75t_L g3852 ( 
.A(n_3539),
.Y(n_3852)
);

INVx2_ASAP7_75t_L g3853 ( 
.A(n_3554),
.Y(n_3853)
);

NAND2xp5_ASAP7_75t_SL g3854 ( 
.A(n_3600),
.B(n_2030),
.Y(n_3854)
);

INVx2_ASAP7_75t_L g3855 ( 
.A(n_3717),
.Y(n_3855)
);

AOI22xp33_ASAP7_75t_L g3856 ( 
.A1(n_3542),
.A2(n_2312),
.B1(n_2409),
.B2(n_2301),
.Y(n_3856)
);

NOR3xp33_ASAP7_75t_L g3857 ( 
.A(n_3714),
.B(n_2781),
.C(n_2037),
.Y(n_3857)
);

OR2x2_ASAP7_75t_L g3858 ( 
.A(n_3496),
.B(n_3742),
.Y(n_3858)
);

NAND2xp5_ASAP7_75t_L g3859 ( 
.A(n_3534),
.B(n_2031),
.Y(n_3859)
);

INVx1_ASAP7_75t_L g3860 ( 
.A(n_3533),
.Y(n_3860)
);

NAND2xp5_ASAP7_75t_L g3861 ( 
.A(n_3531),
.B(n_3550),
.Y(n_3861)
);

INVx2_ASAP7_75t_L g3862 ( 
.A(n_3734),
.Y(n_3862)
);

BUFx6f_ASAP7_75t_L g3863 ( 
.A(n_3527),
.Y(n_3863)
);

NAND2xp5_ASAP7_75t_L g3864 ( 
.A(n_3710),
.B(n_2039),
.Y(n_3864)
);

AND2x2_ASAP7_75t_L g3865 ( 
.A(n_3579),
.B(n_2312),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_L g3866 ( 
.A(n_3715),
.B(n_2040),
.Y(n_3866)
);

NAND2xp5_ASAP7_75t_L g3867 ( 
.A(n_3718),
.B(n_2042),
.Y(n_3867)
);

NAND2xp5_ASAP7_75t_L g3868 ( 
.A(n_3723),
.B(n_2045),
.Y(n_3868)
);

NOR2xp33_ASAP7_75t_L g3869 ( 
.A(n_3576),
.B(n_2046),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_L g3870 ( 
.A(n_3729),
.B(n_2049),
.Y(n_3870)
);

NOR2xp33_ASAP7_75t_SL g3871 ( 
.A(n_3747),
.B(n_2409),
.Y(n_3871)
);

NAND2xp5_ASAP7_75t_SL g3872 ( 
.A(n_3719),
.B(n_2050),
.Y(n_3872)
);

INVxp67_ASAP7_75t_L g3873 ( 
.A(n_3541),
.Y(n_3873)
);

INVx2_ASAP7_75t_L g3874 ( 
.A(n_3736),
.Y(n_3874)
);

AND2x6_ASAP7_75t_L g3875 ( 
.A(n_3691),
.B(n_2129),
.Y(n_3875)
);

INVx2_ASAP7_75t_L g3876 ( 
.A(n_3749),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3732),
.Y(n_3877)
);

AOI22xp5_ASAP7_75t_L g3878 ( 
.A1(n_3748),
.A2(n_2162),
.B1(n_2204),
.B2(n_2138),
.Y(n_3878)
);

NOR2xp33_ASAP7_75t_L g3879 ( 
.A(n_3724),
.B(n_2053),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_SL g3880 ( 
.A(n_3728),
.B(n_2055),
.Y(n_3880)
);

NOR3xp33_ASAP7_75t_L g3881 ( 
.A(n_3740),
.B(n_2064),
.C(n_2058),
.Y(n_3881)
);

NAND3xp33_ASAP7_75t_L g3882 ( 
.A(n_3582),
.B(n_2068),
.C(n_2067),
.Y(n_3882)
);

NOR2xp67_ASAP7_75t_L g3883 ( 
.A(n_3519),
.B(n_2210),
.Y(n_3883)
);

BUFx6f_ASAP7_75t_L g3884 ( 
.A(n_3527),
.Y(n_3884)
);

INVx2_ASAP7_75t_SL g3885 ( 
.A(n_3745),
.Y(n_3885)
);

NAND2xp5_ASAP7_75t_L g3886 ( 
.A(n_3768),
.B(n_2070),
.Y(n_3886)
);

NAND2xp5_ASAP7_75t_L g3887 ( 
.A(n_3771),
.B(n_2073),
.Y(n_3887)
);

NOR2xp33_ASAP7_75t_L g3888 ( 
.A(n_3746),
.B(n_2082),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_3774),
.Y(n_3889)
);

INVx2_ASAP7_75t_L g3890 ( 
.A(n_3753),
.Y(n_3890)
);

INVx2_ASAP7_75t_SL g3891 ( 
.A(n_3540),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_L g3892 ( 
.A(n_3526),
.B(n_2092),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_L g3893 ( 
.A(n_3517),
.B(n_2100),
.Y(n_3893)
);

BUFx3_ASAP7_75t_L g3894 ( 
.A(n_3538),
.Y(n_3894)
);

AOI21xp5_ASAP7_75t_L g3895 ( 
.A1(n_3709),
.A2(n_1712),
.B(n_1710),
.Y(n_3895)
);

INVx2_ASAP7_75t_L g3896 ( 
.A(n_3754),
.Y(n_3896)
);

NAND2xp5_ASAP7_75t_SL g3897 ( 
.A(n_3666),
.B(n_2106),
.Y(n_3897)
);

INVx1_ASAP7_75t_L g3898 ( 
.A(n_3552),
.Y(n_3898)
);

INVx2_ASAP7_75t_L g3899 ( 
.A(n_3767),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3560),
.Y(n_3900)
);

NAND2xp5_ASAP7_75t_SL g3901 ( 
.A(n_3674),
.B(n_2115),
.Y(n_3901)
);

INVx3_ASAP7_75t_L g3902 ( 
.A(n_3772),
.Y(n_3902)
);

INVx1_ASAP7_75t_L g3903 ( 
.A(n_3565),
.Y(n_3903)
);

INVx1_ASAP7_75t_L g3904 ( 
.A(n_3569),
.Y(n_3904)
);

INVx2_ASAP7_75t_SL g3905 ( 
.A(n_3609),
.Y(n_3905)
);

INVx1_ASAP7_75t_L g3906 ( 
.A(n_3570),
.Y(n_3906)
);

HB1xp67_ASAP7_75t_L g3907 ( 
.A(n_3659),
.Y(n_3907)
);

NAND2xp5_ASAP7_75t_L g3908 ( 
.A(n_3523),
.B(n_2117),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3573),
.Y(n_3909)
);

OAI22xp33_ASAP7_75t_L g3910 ( 
.A1(n_3656),
.A2(n_2123),
.B1(n_2125),
.B2(n_2120),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_L g3911 ( 
.A(n_3528),
.B(n_2127),
.Y(n_3911)
);

AO22x2_ASAP7_75t_L g3912 ( 
.A1(n_3661),
.A2(n_2174),
.B1(n_2214),
.B2(n_2153),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_3574),
.Y(n_3913)
);

INVx1_ASAP7_75t_L g3914 ( 
.A(n_3577),
.Y(n_3914)
);

NAND2xp5_ASAP7_75t_L g3915 ( 
.A(n_3530),
.B(n_2130),
.Y(n_3915)
);

INVx2_ASAP7_75t_L g3916 ( 
.A(n_3773),
.Y(n_3916)
);

NAND2xp33_ASAP7_75t_L g3917 ( 
.A(n_3578),
.B(n_2131),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3581),
.Y(n_3918)
);

NAND2xp5_ASAP7_75t_SL g3919 ( 
.A(n_3522),
.B(n_2133),
.Y(n_3919)
);

NAND2xp5_ASAP7_75t_SL g3920 ( 
.A(n_3503),
.B(n_2134),
.Y(n_3920)
);

NAND2xp33_ASAP7_75t_L g3921 ( 
.A(n_3587),
.B(n_3593),
.Y(n_3921)
);

BUFx8_ASAP7_75t_L g3922 ( 
.A(n_3562),
.Y(n_3922)
);

INVx2_ASAP7_75t_L g3923 ( 
.A(n_3777),
.Y(n_3923)
);

NAND2xp5_ASAP7_75t_SL g3924 ( 
.A(n_3505),
.B(n_2136),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3596),
.Y(n_3925)
);

BUFx3_ASAP7_75t_L g3926 ( 
.A(n_3784),
.Y(n_3926)
);

A2O1A1Ixp33_ASAP7_75t_L g3927 ( 
.A1(n_3638),
.A2(n_2224),
.B(n_2232),
.C(n_2212),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_L g3928 ( 
.A(n_3558),
.B(n_2137),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_3545),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_L g3930 ( 
.A(n_3599),
.B(n_2142),
.Y(n_3930)
);

INVxp33_ASAP7_75t_L g3931 ( 
.A(n_3713),
.Y(n_3931)
);

NAND3xp33_ASAP7_75t_L g3932 ( 
.A(n_3585),
.B(n_2146),
.C(n_2145),
.Y(n_3932)
);

NAND2xp5_ASAP7_75t_L g3933 ( 
.A(n_3548),
.B(n_2149),
.Y(n_3933)
);

AND2x2_ASAP7_75t_L g3934 ( 
.A(n_3553),
.B(n_2440),
.Y(n_3934)
);

NAND2xp5_ASAP7_75t_L g3935 ( 
.A(n_3677),
.B(n_2151),
.Y(n_3935)
);

INVx2_ASAP7_75t_L g3936 ( 
.A(n_3779),
.Y(n_3936)
);

OAI22xp5_ASAP7_75t_L g3937 ( 
.A1(n_3518),
.A2(n_2156),
.B1(n_2158),
.B2(n_2152),
.Y(n_3937)
);

INVx1_ASAP7_75t_L g3938 ( 
.A(n_3626),
.Y(n_3938)
);

NAND2xp5_ASAP7_75t_L g3939 ( 
.A(n_3607),
.B(n_3610),
.Y(n_3939)
);

BUFx2_ASAP7_75t_L g3940 ( 
.A(n_3497),
.Y(n_3940)
);

AND2x4_ASAP7_75t_L g3941 ( 
.A(n_3765),
.B(n_3784),
.Y(n_3941)
);

BUFx6f_ASAP7_75t_L g3942 ( 
.A(n_3772),
.Y(n_3942)
);

BUFx8_ASAP7_75t_L g3943 ( 
.A(n_3781),
.Y(n_3943)
);

NAND2xp5_ASAP7_75t_L g3944 ( 
.A(n_3618),
.B(n_2160),
.Y(n_3944)
);

INVx8_ASAP7_75t_L g3945 ( 
.A(n_3765),
.Y(n_3945)
);

OR2x2_ASAP7_75t_L g3946 ( 
.A(n_3716),
.B(n_2161),
.Y(n_3946)
);

INVx1_ASAP7_75t_L g3947 ( 
.A(n_3625),
.Y(n_3947)
);

INVx2_ASAP7_75t_L g3948 ( 
.A(n_3567),
.Y(n_3948)
);

NOR2xp33_ASAP7_75t_L g3949 ( 
.A(n_3616),
.B(n_2163),
.Y(n_3949)
);

INVx2_ASAP7_75t_L g3950 ( 
.A(n_3572),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_L g3951 ( 
.A(n_3629),
.B(n_2166),
.Y(n_3951)
);

INVx2_ASAP7_75t_L g3952 ( 
.A(n_3584),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_L g3953 ( 
.A(n_3639),
.B(n_2167),
.Y(n_3953)
);

INVx1_ASAP7_75t_L g3954 ( 
.A(n_3589),
.Y(n_3954)
);

BUFx3_ASAP7_75t_L g3955 ( 
.A(n_3781),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_3639),
.B(n_2169),
.Y(n_3956)
);

NOR2xp33_ASAP7_75t_L g3957 ( 
.A(n_3520),
.B(n_2172),
.Y(n_3957)
);

AOI22xp5_ASAP7_75t_L g3958 ( 
.A1(n_3748),
.A2(n_2256),
.B1(n_2268),
.B2(n_2247),
.Y(n_3958)
);

NOR2xp67_ASAP7_75t_L g3959 ( 
.A(n_3559),
.B(n_2270),
.Y(n_3959)
);

BUFx3_ASAP7_75t_L g3960 ( 
.A(n_3782),
.Y(n_3960)
);

INVxp67_ASAP7_75t_L g3961 ( 
.A(n_3721),
.Y(n_3961)
);

NAND3xp33_ASAP7_75t_L g3962 ( 
.A(n_3624),
.B(n_2181),
.C(n_2176),
.Y(n_3962)
);

O2A1O1Ixp5_ASAP7_75t_L g3963 ( 
.A1(n_3662),
.A2(n_2375),
.B(n_2416),
.C(n_2231),
.Y(n_3963)
);

NAND2xp5_ASAP7_75t_SL g3964 ( 
.A(n_3613),
.B(n_2182),
.Y(n_3964)
);

NAND2x1_ASAP7_75t_L g3965 ( 
.A(n_3650),
.B(n_1930),
.Y(n_3965)
);

NAND2xp5_ASAP7_75t_L g3966 ( 
.A(n_3590),
.B(n_2185),
.Y(n_3966)
);

NAND2xp33_ASAP7_75t_L g3967 ( 
.A(n_3537),
.B(n_2191),
.Y(n_3967)
);

NAND2xp33_ASAP7_75t_L g3968 ( 
.A(n_3775),
.B(n_2195),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_SL g3969 ( 
.A(n_3604),
.B(n_2197),
.Y(n_3969)
);

INVx2_ASAP7_75t_L g3970 ( 
.A(n_3606),
.Y(n_3970)
);

NAND2xp33_ASAP7_75t_L g3971 ( 
.A(n_3775),
.B(n_2198),
.Y(n_3971)
);

NOR2x1p5_ASAP7_75t_L g3972 ( 
.A(n_3733),
.B(n_2201),
.Y(n_3972)
);

NAND2xp5_ASAP7_75t_L g3973 ( 
.A(n_3608),
.B(n_2203),
.Y(n_3973)
);

INVx1_ASAP7_75t_L g3974 ( 
.A(n_3653),
.Y(n_3974)
);

INVx4_ASAP7_75t_L g3975 ( 
.A(n_3782),
.Y(n_3975)
);

NAND2xp5_ASAP7_75t_SL g3976 ( 
.A(n_3604),
.B(n_3636),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_SL g3977 ( 
.A(n_3707),
.B(n_2205),
.Y(n_3977)
);

INVx1_ASAP7_75t_L g3978 ( 
.A(n_3673),
.Y(n_3978)
);

NOR2xp67_ASAP7_75t_L g3979 ( 
.A(n_3559),
.B(n_2277),
.Y(n_3979)
);

OR2x6_ASAP7_75t_L g3980 ( 
.A(n_3598),
.B(n_2430),
.Y(n_3980)
);

AOI22xp5_ASAP7_75t_L g3981 ( 
.A1(n_3759),
.A2(n_2294),
.B1(n_2304),
.B2(n_2278),
.Y(n_3981)
);

BUFx10_ASAP7_75t_L g3982 ( 
.A(n_3654),
.Y(n_3982)
);

BUFx3_ASAP7_75t_L g3983 ( 
.A(n_3757),
.Y(n_3983)
);

INVx2_ASAP7_75t_SL g3984 ( 
.A(n_3609),
.Y(n_3984)
);

NAND2xp5_ASAP7_75t_L g3985 ( 
.A(n_3720),
.B(n_2213),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_L g3986 ( 
.A(n_3752),
.B(n_3668),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_3682),
.Y(n_3987)
);

NAND2xp5_ASAP7_75t_L g3988 ( 
.A(n_3685),
.B(n_2218),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_L g3989 ( 
.A(n_3635),
.B(n_2220),
.Y(n_3989)
);

INVx4_ASAP7_75t_L g3990 ( 
.A(n_3492),
.Y(n_3990)
);

INVx1_ASAP7_75t_L g3991 ( 
.A(n_3660),
.Y(n_3991)
);

INVx2_ASAP7_75t_L g3992 ( 
.A(n_3669),
.Y(n_3992)
);

NAND2xp5_ASAP7_75t_L g3993 ( 
.A(n_3645),
.B(n_2222),
.Y(n_3993)
);

INVx1_ASAP7_75t_L g3994 ( 
.A(n_3675),
.Y(n_3994)
);

AND2x6_ASAP7_75t_L g3995 ( 
.A(n_3615),
.B(n_2305),
.Y(n_3995)
);

INVxp67_ASAP7_75t_L g3996 ( 
.A(n_3602),
.Y(n_3996)
);

AND2x4_ASAP7_75t_L g3997 ( 
.A(n_3726),
.B(n_3739),
.Y(n_3997)
);

INVx2_ASAP7_75t_L g3998 ( 
.A(n_3676),
.Y(n_3998)
);

INVx1_ASAP7_75t_L g3999 ( 
.A(n_3620),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_SL g4000 ( 
.A(n_3704),
.B(n_2225),
.Y(n_4000)
);

NAND2xp5_ASAP7_75t_L g4001 ( 
.A(n_3549),
.B(n_2227),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_L g4002 ( 
.A(n_3617),
.B(n_2228),
.Y(n_4002)
);

NAND2xp5_ASAP7_75t_SL g4003 ( 
.A(n_3693),
.B(n_2234),
.Y(n_4003)
);

NAND2xp5_ASAP7_75t_L g4004 ( 
.A(n_3513),
.B(n_2235),
.Y(n_4004)
);

NAND2xp33_ASAP7_75t_L g4005 ( 
.A(n_3664),
.B(n_3647),
.Y(n_4005)
);

INVx4_ASAP7_75t_L g4006 ( 
.A(n_3764),
.Y(n_4006)
);

AND2x2_ASAP7_75t_L g4007 ( 
.A(n_3564),
.B(n_2440),
.Y(n_4007)
);

NAND2xp5_ASAP7_75t_SL g4008 ( 
.A(n_3701),
.B(n_2236),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_L g4009 ( 
.A(n_3751),
.B(n_2239),
.Y(n_4009)
);

NAND2xp5_ASAP7_75t_SL g4010 ( 
.A(n_3701),
.B(n_2242),
.Y(n_4010)
);

NAND2xp5_ASAP7_75t_L g4011 ( 
.A(n_3766),
.B(n_2244),
.Y(n_4011)
);

INVx2_ASAP7_75t_L g4012 ( 
.A(n_3688),
.Y(n_4012)
);

INVx1_ASAP7_75t_L g4013 ( 
.A(n_3622),
.Y(n_4013)
);

NAND2xp5_ASAP7_75t_SL g4014 ( 
.A(n_3783),
.B(n_2245),
.Y(n_4014)
);

NAND2xp5_ASAP7_75t_L g4015 ( 
.A(n_3621),
.B(n_2246),
.Y(n_4015)
);

NAND2xp5_ASAP7_75t_SL g4016 ( 
.A(n_3592),
.B(n_2258),
.Y(n_4016)
);

INVxp67_ASAP7_75t_SL g4017 ( 
.A(n_3557),
.Y(n_4017)
);

AOI22xp33_ASAP7_75t_L g4018 ( 
.A1(n_3652),
.A2(n_2708),
.B1(n_2498),
.B2(n_2441),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_L g4019 ( 
.A(n_3623),
.B(n_2261),
.Y(n_4019)
);

AOI22xp33_ASAP7_75t_L g4020 ( 
.A1(n_3536),
.A2(n_2708),
.B1(n_2498),
.B2(n_2449),
.Y(n_4020)
);

NAND2xp5_ASAP7_75t_SL g4021 ( 
.A(n_3597),
.B(n_2264),
.Y(n_4021)
);

NOR2xp33_ASAP7_75t_L g4022 ( 
.A(n_3543),
.B(n_3515),
.Y(n_4022)
);

NAND2xp5_ASAP7_75t_L g4023 ( 
.A(n_3544),
.B(n_2269),
.Y(n_4023)
);

NOR2xp67_ASAP7_75t_L g4024 ( 
.A(n_3776),
.B(n_2307),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3627),
.Y(n_4025)
);

INVx2_ASAP7_75t_SL g4026 ( 
.A(n_3580),
.Y(n_4026)
);

INVx1_ASAP7_75t_L g4027 ( 
.A(n_3633),
.Y(n_4027)
);

NAND2xp5_ASAP7_75t_L g4028 ( 
.A(n_3546),
.B(n_2271),
.Y(n_4028)
);

NAND2xp5_ASAP7_75t_L g4029 ( 
.A(n_3698),
.B(n_2273),
.Y(n_4029)
);

INVx1_ASAP7_75t_L g4030 ( 
.A(n_3702),
.Y(n_4030)
);

NOR2xp33_ASAP7_75t_L g4031 ( 
.A(n_3489),
.B(n_2275),
.Y(n_4031)
);

OR2x2_ASAP7_75t_L g4032 ( 
.A(n_3595),
.B(n_2280),
.Y(n_4032)
);

NOR2xp33_ASAP7_75t_SL g4033 ( 
.A(n_3655),
.B(n_3614),
.Y(n_4033)
);

INVx1_ASAP7_75t_L g4034 ( 
.A(n_3695),
.Y(n_4034)
);

INVx2_ASAP7_75t_L g4035 ( 
.A(n_3690),
.Y(n_4035)
);

NOR2xp33_ASAP7_75t_L g4036 ( 
.A(n_3743),
.B(n_2283),
.Y(n_4036)
);

NOR2xp33_ASAP7_75t_L g4037 ( 
.A(n_3744),
.B(n_2284),
.Y(n_4037)
);

INVx3_ASAP7_75t_L g4038 ( 
.A(n_3632),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_L g4039 ( 
.A(n_3619),
.B(n_2285),
.Y(n_4039)
);

NAND2xp5_ASAP7_75t_L g4040 ( 
.A(n_3663),
.B(n_2286),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_SL g4041 ( 
.A(n_3605),
.B(n_2287),
.Y(n_4041)
);

NAND2xp5_ASAP7_75t_SL g4042 ( 
.A(n_3586),
.B(n_2288),
.Y(n_4042)
);

NAND2xp5_ASAP7_75t_L g4043 ( 
.A(n_3490),
.B(n_2291),
.Y(n_4043)
);

NAND2xp5_ASAP7_75t_L g4044 ( 
.A(n_3699),
.B(n_3700),
.Y(n_4044)
);

NAND2xp5_ASAP7_75t_L g4045 ( 
.A(n_3524),
.B(n_2292),
.Y(n_4045)
);

OAI22xp5_ASAP7_75t_L g4046 ( 
.A1(n_3780),
.A2(n_2296),
.B1(n_2302),
.B2(n_2293),
.Y(n_4046)
);

AOI22xp33_ASAP7_75t_L g4047 ( 
.A1(n_3667),
.A2(n_3680),
.B1(n_3687),
.B2(n_3637),
.Y(n_4047)
);

NAND2xp5_ASAP7_75t_SL g4048 ( 
.A(n_3601),
.B(n_3630),
.Y(n_4048)
);

NAND2xp5_ASAP7_75t_L g4049 ( 
.A(n_3697),
.B(n_2303),
.Y(n_4049)
);

NAND2xp5_ASAP7_75t_L g4050 ( 
.A(n_3651),
.B(n_2306),
.Y(n_4050)
);

INVx2_ASAP7_75t_L g4051 ( 
.A(n_3696),
.Y(n_4051)
);

AOI22xp33_ASAP7_75t_L g4052 ( 
.A1(n_3648),
.A2(n_2475),
.B1(n_2495),
.B2(n_2438),
.Y(n_4052)
);

NOR2xp33_ASAP7_75t_L g4053 ( 
.A(n_3628),
.B(n_2309),
.Y(n_4053)
);

CKINVDCx5p33_ASAP7_75t_R g4054 ( 
.A(n_3571),
.Y(n_4054)
);

INVx1_ASAP7_75t_L g4055 ( 
.A(n_3651),
.Y(n_4055)
);

OR2x2_ASAP7_75t_L g4056 ( 
.A(n_3758),
.B(n_2310),
.Y(n_4056)
);

NOR3xp33_ASAP7_75t_L g4057 ( 
.A(n_3612),
.B(n_2315),
.C(n_2311),
.Y(n_4057)
);

NOR2xp33_ASAP7_75t_L g4058 ( 
.A(n_3703),
.B(n_2320),
.Y(n_4058)
);

BUFx6f_ASAP7_75t_SL g4059 ( 
.A(n_3509),
.Y(n_4059)
);

NOR2xp33_ASAP7_75t_L g4060 ( 
.A(n_3683),
.B(n_2323),
.Y(n_4060)
);

NAND2xp5_ASAP7_75t_L g4061 ( 
.A(n_3706),
.B(n_2333),
.Y(n_4061)
);

INVxp67_ASAP7_75t_L g4062 ( 
.A(n_3670),
.Y(n_4062)
);

NAND2xp5_ASAP7_75t_L g4063 ( 
.A(n_3684),
.B(n_2335),
.Y(n_4063)
);

NAND2xp5_ASAP7_75t_L g4064 ( 
.A(n_3705),
.B(n_2337),
.Y(n_4064)
);

NOR2xp33_ASAP7_75t_L g4065 ( 
.A(n_3556),
.B(n_3566),
.Y(n_4065)
);

NAND2xp5_ASAP7_75t_L g4066 ( 
.A(n_3678),
.B(n_2341),
.Y(n_4066)
);

NOR2x1p5_ASAP7_75t_L g4067 ( 
.A(n_3649),
.B(n_2342),
.Y(n_4067)
);

AOI22xp5_ASAP7_75t_L g4068 ( 
.A1(n_3643),
.A2(n_2318),
.B1(n_2336),
.B2(n_2314),
.Y(n_4068)
);

OAI22xp5_ASAP7_75t_SL g4069 ( 
.A1(n_3594),
.A2(n_2345),
.B1(n_2347),
.B2(n_2346),
.Y(n_4069)
);

INVx1_ASAP7_75t_L g4070 ( 
.A(n_3692),
.Y(n_4070)
);

INVx2_ASAP7_75t_L g4071 ( 
.A(n_3686),
.Y(n_4071)
);

INVx1_ASAP7_75t_L g4072 ( 
.A(n_3686),
.Y(n_4072)
);

INVx4_ASAP7_75t_L g4073 ( 
.A(n_3630),
.Y(n_4073)
);

OAI22xp33_ASAP7_75t_L g4074 ( 
.A1(n_3770),
.A2(n_3658),
.B1(n_3694),
.B2(n_3689),
.Y(n_4074)
);

NOR2xp67_ASAP7_75t_L g4075 ( 
.A(n_3689),
.B(n_2350),
.Y(n_4075)
);

NAND2xp5_ASAP7_75t_SL g4076 ( 
.A(n_3603),
.B(n_2354),
.Y(n_4076)
);

NOR2xp67_ASAP7_75t_L g4077 ( 
.A(n_3694),
.B(n_2367),
.Y(n_4077)
);

INVx2_ASAP7_75t_L g4078 ( 
.A(n_3712),
.Y(n_4078)
);

INVx3_ASAP7_75t_L g4079 ( 
.A(n_3760),
.Y(n_4079)
);

INVx1_ASAP7_75t_L g4080 ( 
.A(n_3487),
.Y(n_4080)
);

INVx2_ASAP7_75t_L g4081 ( 
.A(n_3679),
.Y(n_4081)
);

INVxp67_ASAP7_75t_L g4082 ( 
.A(n_3769),
.Y(n_4082)
);

INVx2_ASAP7_75t_L g4083 ( 
.A(n_3679),
.Y(n_4083)
);

INVx1_ASAP7_75t_L g4084 ( 
.A(n_3487),
.Y(n_4084)
);

OR2x2_ASAP7_75t_L g4085 ( 
.A(n_3588),
.B(n_2356),
.Y(n_4085)
);

INVx1_ASAP7_75t_L g4086 ( 
.A(n_3487),
.Y(n_4086)
);

NAND2xp5_ASAP7_75t_SL g4087 ( 
.A(n_3516),
.B(n_2357),
.Y(n_4087)
);

INVx1_ASAP7_75t_L g4088 ( 
.A(n_3487),
.Y(n_4088)
);

NAND2xp5_ASAP7_75t_L g4089 ( 
.A(n_3516),
.B(n_2359),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_L g4090 ( 
.A(n_3516),
.B(n_2364),
.Y(n_4090)
);

INVx3_ASAP7_75t_L g4091 ( 
.A(n_3750),
.Y(n_4091)
);

INVx2_ASAP7_75t_SL g4092 ( 
.A(n_3769),
.Y(n_4092)
);

NAND2xp5_ASAP7_75t_L g4093 ( 
.A(n_3516),
.B(n_2369),
.Y(n_4093)
);

AOI22xp5_ASAP7_75t_L g4094 ( 
.A1(n_3640),
.A2(n_2394),
.B1(n_2410),
.B2(n_2393),
.Y(n_4094)
);

OAI22xp5_ASAP7_75t_L g4095 ( 
.A1(n_3516),
.A2(n_2371),
.B1(n_2373),
.B2(n_2370),
.Y(n_4095)
);

AOI22xp5_ASAP7_75t_L g4096 ( 
.A1(n_3640),
.A2(n_2484),
.B1(n_2500),
.B2(n_2455),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_L g4097 ( 
.A(n_3516),
.B(n_2376),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_L g4098 ( 
.A(n_3516),
.B(n_2379),
.Y(n_4098)
);

AOI22xp5_ASAP7_75t_L g4099 ( 
.A1(n_3640),
.A2(n_2508),
.B1(n_2515),
.B2(n_2501),
.Y(n_4099)
);

BUFx3_ASAP7_75t_L g4100 ( 
.A(n_3738),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_3487),
.Y(n_4101)
);

INVx1_ASAP7_75t_L g4102 ( 
.A(n_3487),
.Y(n_4102)
);

NAND2xp5_ASAP7_75t_L g4103 ( 
.A(n_3516),
.B(n_2382),
.Y(n_4103)
);

NOR2xp33_ASAP7_75t_L g4104 ( 
.A(n_3640),
.B(n_2383),
.Y(n_4104)
);

INVx2_ASAP7_75t_L g4105 ( 
.A(n_3679),
.Y(n_4105)
);

INVx2_ASAP7_75t_L g4106 ( 
.A(n_3679),
.Y(n_4106)
);

AOI21xp5_ASAP7_75t_L g4107 ( 
.A1(n_3508),
.A2(n_1717),
.B(n_1716),
.Y(n_4107)
);

NAND2xp5_ASAP7_75t_L g4108 ( 
.A(n_3516),
.B(n_2387),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_L g4109 ( 
.A(n_3516),
.B(n_2389),
.Y(n_4109)
);

NOR3xp33_ASAP7_75t_L g4110 ( 
.A(n_3516),
.B(n_2398),
.C(n_2397),
.Y(n_4110)
);

INVx4_ASAP7_75t_L g4111 ( 
.A(n_3519),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_SL g4112 ( 
.A(n_3516),
.B(n_2400),
.Y(n_4112)
);

CKINVDCx5p33_ASAP7_75t_R g4113 ( 
.A(n_3498),
.Y(n_4113)
);

NOR2x1p5_ASAP7_75t_L g4114 ( 
.A(n_3500),
.B(n_2401),
.Y(n_4114)
);

NAND2xp5_ASAP7_75t_L g4115 ( 
.A(n_3516),
.B(n_2407),
.Y(n_4115)
);

NOR2xp33_ASAP7_75t_L g4116 ( 
.A(n_3640),
.B(n_2411),
.Y(n_4116)
);

INVx1_ASAP7_75t_SL g4117 ( 
.A(n_3769),
.Y(n_4117)
);

NAND2xp5_ASAP7_75t_L g4118 ( 
.A(n_3516),
.B(n_2412),
.Y(n_4118)
);

AOI22xp5_ASAP7_75t_L g4119 ( 
.A1(n_3640),
.A2(n_2564),
.B1(n_2566),
.B2(n_2545),
.Y(n_4119)
);

INVx2_ASAP7_75t_L g4120 ( 
.A(n_3679),
.Y(n_4120)
);

NAND2xp5_ASAP7_75t_L g4121 ( 
.A(n_3516),
.B(n_2413),
.Y(n_4121)
);

NAND2xp5_ASAP7_75t_SL g4122 ( 
.A(n_3516),
.B(n_2420),
.Y(n_4122)
);

NAND2xp5_ASAP7_75t_SL g4123 ( 
.A(n_3516),
.B(n_2422),
.Y(n_4123)
);

NAND2xp5_ASAP7_75t_SL g4124 ( 
.A(n_3516),
.B(n_2424),
.Y(n_4124)
);

NOR2xp33_ASAP7_75t_L g4125 ( 
.A(n_3640),
.B(n_2425),
.Y(n_4125)
);

NOR2xp33_ASAP7_75t_L g4126 ( 
.A(n_3640),
.B(n_2426),
.Y(n_4126)
);

NAND2xp5_ASAP7_75t_L g4127 ( 
.A(n_3516),
.B(n_2428),
.Y(n_4127)
);

NAND2xp5_ASAP7_75t_L g4128 ( 
.A(n_3516),
.B(n_2429),
.Y(n_4128)
);

AOI22xp33_ASAP7_75t_L g4129 ( 
.A1(n_3640),
.A2(n_2583),
.B1(n_2586),
.B2(n_2524),
.Y(n_4129)
);

INVx1_ASAP7_75t_L g4130 ( 
.A(n_3487),
.Y(n_4130)
);

OAI22xp5_ASAP7_75t_L g4131 ( 
.A1(n_3516),
.A2(n_2447),
.B1(n_2448),
.B2(n_2437),
.Y(n_4131)
);

NOR2xp33_ASAP7_75t_L g4132 ( 
.A(n_3640),
.B(n_2452),
.Y(n_4132)
);

INVx3_ASAP7_75t_L g4133 ( 
.A(n_3750),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_SL g4134 ( 
.A(n_3516),
.B(n_2456),
.Y(n_4134)
);

OAI22xp5_ASAP7_75t_L g4135 ( 
.A1(n_3516),
.A2(n_2459),
.B1(n_2463),
.B2(n_2457),
.Y(n_4135)
);

INVx4_ASAP7_75t_L g4136 ( 
.A(n_3519),
.Y(n_4136)
);

NAND2xp5_ASAP7_75t_SL g4137 ( 
.A(n_3516),
.B(n_2466),
.Y(n_4137)
);

NAND2xp5_ASAP7_75t_L g4138 ( 
.A(n_3516),
.B(n_2467),
.Y(n_4138)
);

AOI21xp5_ASAP7_75t_L g4139 ( 
.A1(n_3508),
.A2(n_1741),
.B(n_1727),
.Y(n_4139)
);

INVx1_ASAP7_75t_L g4140 ( 
.A(n_3487),
.Y(n_4140)
);

NAND2xp5_ASAP7_75t_L g4141 ( 
.A(n_3516),
.B(n_2478),
.Y(n_4141)
);

INVx2_ASAP7_75t_L g4142 ( 
.A(n_3679),
.Y(n_4142)
);

NAND2xp33_ASAP7_75t_L g4143 ( 
.A(n_3516),
.B(n_2480),
.Y(n_4143)
);

NOR2xp67_ASAP7_75t_L g4144 ( 
.A(n_3519),
.B(n_2593),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_3939),
.Y(n_4145)
);

INVx2_ASAP7_75t_L g4146 ( 
.A(n_3950),
.Y(n_4146)
);

INVx3_ASAP7_75t_L g4147 ( 
.A(n_3945),
.Y(n_4147)
);

BUFx3_ASAP7_75t_L g4148 ( 
.A(n_3945),
.Y(n_4148)
);

NOR2xp33_ASAP7_75t_L g4149 ( 
.A(n_4104),
.B(n_2483),
.Y(n_4149)
);

OR2x6_ASAP7_75t_L g4150 ( 
.A(n_3990),
.B(n_2658),
.Y(n_4150)
);

INVx2_ASAP7_75t_SL g4151 ( 
.A(n_3941),
.Y(n_4151)
);

INVx5_ASAP7_75t_L g4152 ( 
.A(n_4111),
.Y(n_4152)
);

INVx5_ASAP7_75t_L g4153 ( 
.A(n_4136),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_SL g4154 ( 
.A(n_3843),
.B(n_2486),
.Y(n_4154)
);

OR2x2_ASAP7_75t_L g4155 ( 
.A(n_3858),
.B(n_2488),
.Y(n_4155)
);

AOI22xp33_ASAP7_75t_L g4156 ( 
.A1(n_4116),
.A2(n_2503),
.B1(n_2504),
.B2(n_2494),
.Y(n_4156)
);

CKINVDCx5p33_ASAP7_75t_R g4157 ( 
.A(n_4113),
.Y(n_4157)
);

INVxp67_ASAP7_75t_L g4158 ( 
.A(n_3831),
.Y(n_4158)
);

NOR2xp33_ASAP7_75t_L g4159 ( 
.A(n_4125),
.B(n_2506),
.Y(n_4159)
);

AOI22xp5_ASAP7_75t_L g4160 ( 
.A1(n_4126),
.A2(n_2512),
.B1(n_2517),
.B2(n_2507),
.Y(n_4160)
);

BUFx6f_ASAP7_75t_L g4161 ( 
.A(n_3801),
.Y(n_4161)
);

AND2x2_ASAP7_75t_L g4162 ( 
.A(n_4132),
.B(n_2518),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_L g4163 ( 
.A(n_3873),
.B(n_2520),
.Y(n_4163)
);

AND2x2_ASAP7_75t_L g4164 ( 
.A(n_3934),
.B(n_2521),
.Y(n_4164)
);

AOI22xp33_ASAP7_75t_L g4165 ( 
.A1(n_3834),
.A2(n_2530),
.B1(n_2533),
.B2(n_2522),
.Y(n_4165)
);

AND2x4_ASAP7_75t_L g4166 ( 
.A(n_4100),
.B(n_2733),
.Y(n_4166)
);

CKINVDCx5p33_ASAP7_75t_R g4167 ( 
.A(n_3803),
.Y(n_4167)
);

AOI22xp5_ASAP7_75t_L g4168 ( 
.A1(n_3847),
.A2(n_2538),
.B1(n_2543),
.B2(n_2535),
.Y(n_4168)
);

INVx1_ASAP7_75t_L g4169 ( 
.A(n_3807),
.Y(n_4169)
);

NAND2xp5_ASAP7_75t_SL g4170 ( 
.A(n_3996),
.B(n_3982),
.Y(n_4170)
);

NAND2xp5_ASAP7_75t_L g4171 ( 
.A(n_3861),
.B(n_2544),
.Y(n_4171)
);

AND2x4_ASAP7_75t_L g4172 ( 
.A(n_3997),
.B(n_2608),
.Y(n_4172)
);

BUFx5_ASAP7_75t_L g4173 ( 
.A(n_3987),
.Y(n_4173)
);

OAI22xp5_ASAP7_75t_L g4174 ( 
.A1(n_3812),
.A2(n_2554),
.B1(n_2558),
.B2(n_2553),
.Y(n_4174)
);

AND2x4_ASAP7_75t_L g4175 ( 
.A(n_3800),
.B(n_2635),
.Y(n_4175)
);

NAND2xp5_ASAP7_75t_L g4176 ( 
.A(n_3835),
.B(n_2562),
.Y(n_4176)
);

AOI22x1_ASAP7_75t_L g4177 ( 
.A1(n_3895),
.A2(n_2565),
.B1(n_2569),
.B2(n_2563),
.Y(n_4177)
);

AND2x6_ASAP7_75t_L g4178 ( 
.A(n_3938),
.B(n_2656),
.Y(n_4178)
);

INVx1_ASAP7_75t_L g4179 ( 
.A(n_3833),
.Y(n_4179)
);

INVx1_ASAP7_75t_L g4180 ( 
.A(n_3839),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_3850),
.Y(n_4181)
);

INVx2_ASAP7_75t_L g4182 ( 
.A(n_3952),
.Y(n_4182)
);

AOI22xp33_ASAP7_75t_L g4183 ( 
.A1(n_3825),
.A2(n_2577),
.B1(n_2578),
.B2(n_2575),
.Y(n_4183)
);

INVx2_ASAP7_75t_L g4184 ( 
.A(n_3970),
.Y(n_4184)
);

NAND2xp5_ASAP7_75t_L g4185 ( 
.A(n_4089),
.B(n_2580),
.Y(n_4185)
);

INVx2_ASAP7_75t_L g4186 ( 
.A(n_3788),
.Y(n_4186)
);

BUFx6f_ASAP7_75t_L g4187 ( 
.A(n_3894),
.Y(n_4187)
);

INVx2_ASAP7_75t_SL g4188 ( 
.A(n_3943),
.Y(n_4188)
);

BUFx2_ASAP7_75t_L g4189 ( 
.A(n_3802),
.Y(n_4189)
);

INVx2_ASAP7_75t_L g4190 ( 
.A(n_4081),
.Y(n_4190)
);

CKINVDCx5p33_ASAP7_75t_R g4191 ( 
.A(n_3830),
.Y(n_4191)
);

INVx2_ASAP7_75t_L g4192 ( 
.A(n_4083),
.Y(n_4192)
);

CKINVDCx6p67_ASAP7_75t_R g4193 ( 
.A(n_4059),
.Y(n_4193)
);

INVxp67_ASAP7_75t_L g4194 ( 
.A(n_4092),
.Y(n_4194)
);

NOR3xp33_ASAP7_75t_SL g4195 ( 
.A(n_3897),
.B(n_2582),
.C(n_2581),
.Y(n_4195)
);

NAND2xp5_ASAP7_75t_SL g4196 ( 
.A(n_3863),
.B(n_2584),
.Y(n_4196)
);

NOR2xp33_ASAP7_75t_L g4197 ( 
.A(n_3931),
.B(n_2591),
.Y(n_4197)
);

BUFx3_ASAP7_75t_L g4198 ( 
.A(n_3926),
.Y(n_4198)
);

INVx4_ASAP7_75t_L g4199 ( 
.A(n_3863),
.Y(n_4199)
);

AND2x4_ASAP7_75t_L g4200 ( 
.A(n_4091),
.B(n_2673),
.Y(n_4200)
);

NOR2xp33_ASAP7_75t_L g4201 ( 
.A(n_3789),
.B(n_2592),
.Y(n_4201)
);

BUFx6f_ASAP7_75t_L g4202 ( 
.A(n_3884),
.Y(n_4202)
);

AOI22xp5_ASAP7_75t_L g4203 ( 
.A1(n_3806),
.A2(n_4094),
.B1(n_4099),
.B2(n_4096),
.Y(n_4203)
);

NOR2xp33_ASAP7_75t_R g4204 ( 
.A(n_4054),
.B(n_2597),
.Y(n_4204)
);

BUFx2_ASAP7_75t_L g4205 ( 
.A(n_4082),
.Y(n_4205)
);

NAND2xp5_ASAP7_75t_L g4206 ( 
.A(n_4090),
.B(n_2598),
.Y(n_4206)
);

INVx1_ASAP7_75t_L g4207 ( 
.A(n_3860),
.Y(n_4207)
);

AOI22xp5_ASAP7_75t_L g4208 ( 
.A1(n_4119),
.A2(n_3796),
.B1(n_3869),
.B2(n_3961),
.Y(n_4208)
);

INVx1_ASAP7_75t_L g4209 ( 
.A(n_3877),
.Y(n_4209)
);

BUFx6f_ASAP7_75t_L g4210 ( 
.A(n_3884),
.Y(n_4210)
);

NAND2xp5_ASAP7_75t_SL g4211 ( 
.A(n_3942),
.B(n_2601),
.Y(n_4211)
);

NAND2xp5_ASAP7_75t_L g4212 ( 
.A(n_4093),
.B(n_2605),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_L g4213 ( 
.A(n_4097),
.B(n_2606),
.Y(n_4213)
);

NAND2xp5_ASAP7_75t_SL g4214 ( 
.A(n_3942),
.B(n_2609),
.Y(n_4214)
);

BUFx6f_ASAP7_75t_L g4215 ( 
.A(n_3955),
.Y(n_4215)
);

INVx1_ASAP7_75t_L g4216 ( 
.A(n_3889),
.Y(n_4216)
);

OR2x4_ASAP7_75t_L g4217 ( 
.A(n_4032),
.B(n_1998),
.Y(n_4217)
);

AO22x1_ASAP7_75t_L g4218 ( 
.A1(n_3995),
.A2(n_2621),
.B1(n_2623),
.B2(n_2612),
.Y(n_4218)
);

AOI22xp5_ASAP7_75t_L g4219 ( 
.A1(n_3865),
.A2(n_2627),
.B1(n_2629),
.B2(n_2625),
.Y(n_4219)
);

INVx3_ASAP7_75t_L g4220 ( 
.A(n_3983),
.Y(n_4220)
);

NOR2xp33_ASAP7_75t_L g4221 ( 
.A(n_3949),
.B(n_2632),
.Y(n_4221)
);

NAND2xp5_ASAP7_75t_L g4222 ( 
.A(n_4098),
.B(n_2634),
.Y(n_4222)
);

NOR3xp33_ASAP7_75t_SL g4223 ( 
.A(n_4087),
.B(n_2646),
.C(n_2644),
.Y(n_4223)
);

INVx1_ASAP7_75t_L g4224 ( 
.A(n_3898),
.Y(n_4224)
);

AOI22xp33_ASAP7_75t_L g4225 ( 
.A1(n_4047),
.A2(n_2648),
.B1(n_2649),
.B2(n_2647),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_3900),
.Y(n_4226)
);

NOR2xp33_ASAP7_75t_R g4227 ( 
.A(n_4033),
.B(n_2650),
.Y(n_4227)
);

INVx5_ASAP7_75t_L g4228 ( 
.A(n_3980),
.Y(n_4228)
);

OR2x6_ASAP7_75t_L g4229 ( 
.A(n_3980),
.B(n_2405),
.Y(n_4229)
);

CKINVDCx5p33_ASAP7_75t_R g4230 ( 
.A(n_3922),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_3903),
.Y(n_4231)
);

NOR2x1_ASAP7_75t_R g4232 ( 
.A(n_4006),
.B(n_2651),
.Y(n_4232)
);

INVx1_ASAP7_75t_L g4233 ( 
.A(n_3904),
.Y(n_4233)
);

OAI22xp5_ASAP7_75t_SL g4234 ( 
.A1(n_4069),
.A2(n_2654),
.B1(n_2657),
.B2(n_2655),
.Y(n_4234)
);

INVx2_ASAP7_75t_L g4235 ( 
.A(n_4105),
.Y(n_4235)
);

INVx2_ASAP7_75t_SL g4236 ( 
.A(n_3960),
.Y(n_4236)
);

BUFx12f_ASAP7_75t_L g4237 ( 
.A(n_3891),
.Y(n_4237)
);

INVx1_ASAP7_75t_L g4238 ( 
.A(n_3906),
.Y(n_4238)
);

INVx5_ASAP7_75t_L g4239 ( 
.A(n_4133),
.Y(n_4239)
);

INVx2_ASAP7_75t_L g4240 ( 
.A(n_4106),
.Y(n_4240)
);

NAND2xp5_ASAP7_75t_L g4241 ( 
.A(n_4103),
.B(n_2659),
.Y(n_4241)
);

BUFx2_ASAP7_75t_L g4242 ( 
.A(n_4117),
.Y(n_4242)
);

AND2x2_ASAP7_75t_SL g4243 ( 
.A(n_3871),
.B(n_2677),
.Y(n_4243)
);

INVx2_ASAP7_75t_L g4244 ( 
.A(n_4120),
.Y(n_4244)
);

NAND2xp5_ASAP7_75t_L g4245 ( 
.A(n_4108),
.B(n_2660),
.Y(n_4245)
);

INVx1_ASAP7_75t_L g4246 ( 
.A(n_3909),
.Y(n_4246)
);

HB1xp67_ASAP7_75t_L g4247 ( 
.A(n_3940),
.Y(n_4247)
);

NAND2xp5_ASAP7_75t_L g4248 ( 
.A(n_4109),
.B(n_2661),
.Y(n_4248)
);

INVxp67_ASAP7_75t_SL g4249 ( 
.A(n_3921),
.Y(n_4249)
);

AOI21xp5_ASAP7_75t_L g4250 ( 
.A1(n_4005),
.A2(n_2697),
.B(n_2688),
.Y(n_4250)
);

OR2x2_ASAP7_75t_L g4251 ( 
.A(n_4085),
.B(n_2665),
.Y(n_4251)
);

BUFx4f_ASAP7_75t_L g4252 ( 
.A(n_3815),
.Y(n_4252)
);

INVx3_ASAP7_75t_L g4253 ( 
.A(n_3975),
.Y(n_4253)
);

NAND2xp5_ASAP7_75t_L g4254 ( 
.A(n_4115),
.B(n_2667),
.Y(n_4254)
);

AOI22xp33_ASAP7_75t_L g4255 ( 
.A1(n_4062),
.A2(n_2672),
.B1(n_2674),
.B2(n_2668),
.Y(n_4255)
);

INVx5_ASAP7_75t_L g4256 ( 
.A(n_3995),
.Y(n_4256)
);

AOI21xp5_ASAP7_75t_L g4257 ( 
.A1(n_3786),
.A2(n_2735),
.B(n_2719),
.Y(n_4257)
);

NAND2xp5_ASAP7_75t_L g4258 ( 
.A(n_4118),
.B(n_2683),
.Y(n_4258)
);

AOI22xp5_ASAP7_75t_L g4259 ( 
.A1(n_3791),
.A2(n_2687),
.B1(n_2690),
.B2(n_2686),
.Y(n_4259)
);

NAND2xp5_ASAP7_75t_L g4260 ( 
.A(n_4121),
.B(n_2691),
.Y(n_4260)
);

AOI22xp5_ASAP7_75t_L g4261 ( 
.A1(n_3910),
.A2(n_2694),
.B1(n_2695),
.B2(n_2693),
.Y(n_4261)
);

NAND2xp5_ASAP7_75t_SL g4262 ( 
.A(n_4074),
.B(n_2696),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_3913),
.Y(n_4263)
);

INVx2_ASAP7_75t_L g4264 ( 
.A(n_4142),
.Y(n_4264)
);

NAND2xp5_ASAP7_75t_L g4265 ( 
.A(n_4127),
.B(n_2698),
.Y(n_4265)
);

INVx3_ASAP7_75t_L g4266 ( 
.A(n_4073),
.Y(n_4266)
);

AND2x4_ASAP7_75t_L g4267 ( 
.A(n_3797),
.B(n_2747),
.Y(n_4267)
);

BUFx6f_ASAP7_75t_SL g4268 ( 
.A(n_4026),
.Y(n_4268)
);

NAND2xp5_ASAP7_75t_SL g4269 ( 
.A(n_3797),
.B(n_3885),
.Y(n_4269)
);

NAND2xp5_ASAP7_75t_L g4270 ( 
.A(n_4128),
.B(n_2706),
.Y(n_4270)
);

OR2x6_ASAP7_75t_L g4271 ( 
.A(n_3905),
.B(n_2540),
.Y(n_4271)
);

NAND2xp5_ASAP7_75t_SL g4272 ( 
.A(n_3797),
.B(n_2716),
.Y(n_4272)
);

NAND2xp5_ASAP7_75t_L g4273 ( 
.A(n_4138),
.B(n_2720),
.Y(n_4273)
);

NAND2xp5_ASAP7_75t_L g4274 ( 
.A(n_4141),
.B(n_3844),
.Y(n_4274)
);

AND2x2_ASAP7_75t_L g4275 ( 
.A(n_3840),
.B(n_2721),
.Y(n_4275)
);

INVx2_ASAP7_75t_L g4276 ( 
.A(n_3954),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_3914),
.Y(n_4277)
);

NAND2xp5_ASAP7_75t_L g4278 ( 
.A(n_3792),
.B(n_2722),
.Y(n_4278)
);

INVx5_ASAP7_75t_L g4279 ( 
.A(n_3995),
.Y(n_4279)
);

AND3x2_ASAP7_75t_SL g4280 ( 
.A(n_4078),
.B(n_2642),
.C(n_1807),
.Y(n_4280)
);

NAND2xp5_ASAP7_75t_L g4281 ( 
.A(n_3798),
.B(n_2723),
.Y(n_4281)
);

NAND2xp5_ASAP7_75t_L g4282 ( 
.A(n_3808),
.B(n_2725),
.Y(n_4282)
);

INVx1_ASAP7_75t_L g4283 ( 
.A(n_3918),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_3925),
.Y(n_4284)
);

AND2x4_ASAP7_75t_L g4285 ( 
.A(n_3902),
.B(n_2749),
.Y(n_4285)
);

AOI22xp33_ASAP7_75t_L g4286 ( 
.A1(n_3799),
.A2(n_2726),
.B1(n_2734),
.B2(n_2728),
.Y(n_4286)
);

AOI22xp5_ASAP7_75t_L g4287 ( 
.A1(n_3917),
.A2(n_2738),
.B1(n_2740),
.B2(n_2737),
.Y(n_4287)
);

NAND2xp5_ASAP7_75t_SL g4288 ( 
.A(n_4058),
.B(n_2742),
.Y(n_4288)
);

BUFx6f_ASAP7_75t_L g4289 ( 
.A(n_3984),
.Y(n_4289)
);

INVx1_ASAP7_75t_L g4290 ( 
.A(n_4080),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_4084),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_4086),
.Y(n_4292)
);

INVx5_ASAP7_75t_L g4293 ( 
.A(n_3875),
.Y(n_4293)
);

INVx1_ASAP7_75t_L g4294 ( 
.A(n_4088),
.Y(n_4294)
);

AOI22xp5_ASAP7_75t_L g4295 ( 
.A1(n_3968),
.A2(n_2750),
.B1(n_2752),
.B2(n_2744),
.Y(n_4295)
);

CKINVDCx11_ASAP7_75t_R g4296 ( 
.A(n_4071),
.Y(n_4296)
);

BUFx12f_ASAP7_75t_L g4297 ( 
.A(n_4114),
.Y(n_4297)
);

HB1xp67_ASAP7_75t_L g4298 ( 
.A(n_3907),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_4101),
.Y(n_4299)
);

NOR2xp33_ASAP7_75t_R g4300 ( 
.A(n_3814),
.B(n_3967),
.Y(n_4300)
);

BUFx6f_ASAP7_75t_L g4301 ( 
.A(n_4038),
.Y(n_4301)
);

INVx1_ASAP7_75t_L g4302 ( 
.A(n_4102),
.Y(n_4302)
);

INVx1_ASAP7_75t_L g4303 ( 
.A(n_4130),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_4140),
.Y(n_4304)
);

OAI21xp5_ASAP7_75t_L g4305 ( 
.A1(n_3818),
.A2(n_2773),
.B(n_2772),
.Y(n_4305)
);

NAND3xp33_ASAP7_75t_SL g4306 ( 
.A(n_3829),
.B(n_2757),
.C(n_2753),
.Y(n_4306)
);

BUFx6f_ASAP7_75t_L g4307 ( 
.A(n_4048),
.Y(n_4307)
);

NAND2xp5_ASAP7_75t_L g4308 ( 
.A(n_3809),
.B(n_2758),
.Y(n_4308)
);

INVx2_ASAP7_75t_SL g4309 ( 
.A(n_4067),
.Y(n_4309)
);

INVx1_ASAP7_75t_L g4310 ( 
.A(n_3947),
.Y(n_4310)
);

INVxp67_ASAP7_75t_L g4311 ( 
.A(n_3813),
.Y(n_4311)
);

NOR3xp33_ASAP7_75t_SL g4312 ( 
.A(n_4112),
.B(n_2762),
.C(n_2759),
.Y(n_4312)
);

NAND2xp5_ASAP7_75t_SL g4313 ( 
.A(n_4110),
.B(n_2764),
.Y(n_4313)
);

CKINVDCx5p33_ASAP7_75t_R g4314 ( 
.A(n_3972),
.Y(n_4314)
);

NAND2xp5_ASAP7_75t_L g4315 ( 
.A(n_3816),
.B(n_2765),
.Y(n_4315)
);

NAND3xp33_ASAP7_75t_SL g4316 ( 
.A(n_3989),
.B(n_2777),
.C(n_2770),
.Y(n_4316)
);

NAND2xp5_ASAP7_75t_SL g4317 ( 
.A(n_4022),
.B(n_2778),
.Y(n_4317)
);

AOI22x1_ASAP7_75t_L g4318 ( 
.A1(n_3999),
.A2(n_2784),
.B1(n_1816),
.B2(n_1905),
.Y(n_4318)
);

INVx2_ASAP7_75t_SL g4319 ( 
.A(n_4070),
.Y(n_4319)
);

AND2x2_ASAP7_75t_SL g4320 ( 
.A(n_3971),
.B(n_1776),
.Y(n_4320)
);

NAND2xp5_ASAP7_75t_L g4321 ( 
.A(n_3817),
.B(n_1),
.Y(n_4321)
);

INVx1_ASAP7_75t_L g4322 ( 
.A(n_4030),
.Y(n_4322)
);

INVx2_ASAP7_75t_L g4323 ( 
.A(n_3974),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_3929),
.Y(n_4324)
);

AND2x6_ASAP7_75t_L g4325 ( 
.A(n_4013),
.B(n_1931),
.Y(n_4325)
);

AOI22xp5_ASAP7_75t_L g4326 ( 
.A1(n_4143),
.A2(n_1745),
.B1(n_1749),
.B2(n_1743),
.Y(n_4326)
);

INVx1_ASAP7_75t_L g4327 ( 
.A(n_3978),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_4034),
.Y(n_4328)
);

NOR2xp33_ASAP7_75t_L g4329 ( 
.A(n_3993),
.B(n_1750),
.Y(n_4329)
);

INVx2_ASAP7_75t_L g4330 ( 
.A(n_3810),
.Y(n_4330)
);

NAND2xp5_ASAP7_75t_L g4331 ( 
.A(n_3986),
.B(n_2),
.Y(n_4331)
);

AOI21xp5_ASAP7_75t_L g4332 ( 
.A1(n_4122),
.A2(n_2267),
.B(n_2009),
.Y(n_4332)
);

INVx2_ASAP7_75t_SL g4333 ( 
.A(n_3976),
.Y(n_4333)
);

CKINVDCx5p33_ASAP7_75t_R g4334 ( 
.A(n_4079),
.Y(n_4334)
);

INVx2_ASAP7_75t_SL g4335 ( 
.A(n_4055),
.Y(n_4335)
);

AND2x2_ASAP7_75t_L g4336 ( 
.A(n_3842),
.B(n_2),
.Y(n_4336)
);

INVx2_ASAP7_75t_L g4337 ( 
.A(n_3824),
.Y(n_4337)
);

AOI21xp5_ASAP7_75t_L g4338 ( 
.A1(n_4123),
.A2(n_2641),
.B(n_2590),
.Y(n_4338)
);

AOI21xp5_ASAP7_75t_L g4339 ( 
.A1(n_4124),
.A2(n_1756),
.B(n_1755),
.Y(n_4339)
);

NAND2xp5_ASAP7_75t_L g4340 ( 
.A(n_3837),
.B(n_3),
.Y(n_4340)
);

BUFx6f_ASAP7_75t_L g4341 ( 
.A(n_4072),
.Y(n_4341)
);

NAND2xp5_ASAP7_75t_SL g4342 ( 
.A(n_3879),
.B(n_1757),
.Y(n_4342)
);

NAND2xp5_ASAP7_75t_L g4343 ( 
.A(n_3846),
.B(n_3),
.Y(n_4343)
);

INVx1_ASAP7_75t_L g4344 ( 
.A(n_3991),
.Y(n_4344)
);

NAND2xp5_ASAP7_75t_L g4345 ( 
.A(n_3849),
.B(n_4),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_3994),
.Y(n_4346)
);

INVx2_ASAP7_75t_L g4347 ( 
.A(n_3827),
.Y(n_4347)
);

NAND2xp5_ASAP7_75t_L g4348 ( 
.A(n_3859),
.B(n_4),
.Y(n_4348)
);

NOR2x1p5_ASAP7_75t_L g4349 ( 
.A(n_3845),
.B(n_2624),
.Y(n_4349)
);

CKINVDCx5p33_ASAP7_75t_R g4350 ( 
.A(n_3790),
.Y(n_4350)
);

NAND2xp5_ASAP7_75t_SL g4351 ( 
.A(n_3888),
.B(n_1759),
.Y(n_4351)
);

BUFx2_ASAP7_75t_L g4352 ( 
.A(n_3875),
.Y(n_4352)
);

NAND2xp5_ASAP7_75t_L g4353 ( 
.A(n_3893),
.B(n_5),
.Y(n_4353)
);

NAND2xp5_ASAP7_75t_SL g4354 ( 
.A(n_4060),
.B(n_1762),
.Y(n_4354)
);

INVx1_ASAP7_75t_L g4355 ( 
.A(n_4044),
.Y(n_4355)
);

NAND2xp5_ASAP7_75t_L g4356 ( 
.A(n_3908),
.B(n_5),
.Y(n_4356)
);

INVx3_ASAP7_75t_L g4357 ( 
.A(n_4051),
.Y(n_4357)
);

NOR2xp33_ASAP7_75t_L g4358 ( 
.A(n_4025),
.B(n_1767),
.Y(n_4358)
);

NAND2xp5_ASAP7_75t_L g4359 ( 
.A(n_3911),
.B(n_6),
.Y(n_4359)
);

NOR2x1p5_ASAP7_75t_L g4360 ( 
.A(n_3946),
.B(n_1768),
.Y(n_4360)
);

NAND2xp5_ASAP7_75t_L g4361 ( 
.A(n_3915),
.B(n_6),
.Y(n_4361)
);

NOR2xp33_ASAP7_75t_L g4362 ( 
.A(n_4027),
.B(n_3882),
.Y(n_4362)
);

NAND2xp5_ASAP7_75t_L g4363 ( 
.A(n_3928),
.B(n_7),
.Y(n_4363)
);

AOI22xp5_ASAP7_75t_L g4364 ( 
.A1(n_4031),
.A2(n_4036),
.B1(n_4037),
.B2(n_3787),
.Y(n_4364)
);

INVx4_ASAP7_75t_L g4365 ( 
.A(n_3875),
.Y(n_4365)
);

NOR2xp33_ASAP7_75t_SL g4366 ( 
.A(n_3959),
.B(n_1775),
.Y(n_4366)
);

AND2x4_ASAP7_75t_L g4367 ( 
.A(n_4017),
.B(n_4024),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_3838),
.Y(n_4368)
);

NOR2xp33_ASAP7_75t_L g4369 ( 
.A(n_4134),
.B(n_4137),
.Y(n_4369)
);

INVx3_ASAP7_75t_L g4370 ( 
.A(n_3965),
.Y(n_4370)
);

NOR3xp33_ASAP7_75t_SL g4371 ( 
.A(n_4095),
.B(n_1790),
.C(n_1783),
.Y(n_4371)
);

NAND2xp5_ASAP7_75t_SL g4372 ( 
.A(n_3878),
.B(n_1792),
.Y(n_4372)
);

INVx1_ASAP7_75t_L g4373 ( 
.A(n_3841),
.Y(n_4373)
);

NAND2xp5_ASAP7_75t_SL g4374 ( 
.A(n_3958),
.B(n_1795),
.Y(n_4374)
);

NAND2xp5_ASAP7_75t_L g4375 ( 
.A(n_3826),
.B(n_7),
.Y(n_4375)
);

NAND2xp5_ASAP7_75t_L g4376 ( 
.A(n_3832),
.B(n_8),
.Y(n_4376)
);

INVx1_ASAP7_75t_L g4377 ( 
.A(n_3848),
.Y(n_4377)
);

NAND2xp5_ASAP7_75t_L g4378 ( 
.A(n_3836),
.B(n_8),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_3852),
.Y(n_4379)
);

INVx1_ASAP7_75t_SL g4380 ( 
.A(n_4050),
.Y(n_4380)
);

INVx1_ASAP7_75t_L g4381 ( 
.A(n_3853),
.Y(n_4381)
);

AND3x1_ASAP7_75t_L g4382 ( 
.A(n_3881),
.B(n_9),
.C(n_10),
.Y(n_4382)
);

INVx2_ASAP7_75t_L g4383 ( 
.A(n_3855),
.Y(n_4383)
);

INVx1_ASAP7_75t_L g4384 ( 
.A(n_3862),
.Y(n_4384)
);

AOI22xp33_ASAP7_75t_L g4385 ( 
.A1(n_3892),
.A2(n_3828),
.B1(n_4129),
.B2(n_4028),
.Y(n_4385)
);

BUFx6f_ASAP7_75t_L g4386 ( 
.A(n_3874),
.Y(n_4386)
);

HB1xp67_ASAP7_75t_L g4387 ( 
.A(n_4012),
.Y(n_4387)
);

AOI21xp5_ASAP7_75t_L g4388 ( 
.A1(n_3964),
.A2(n_1804),
.B(n_1800),
.Y(n_4388)
);

AND2x2_ASAP7_75t_L g4389 ( 
.A(n_4007),
.B(n_10),
.Y(n_4389)
);

CKINVDCx5p33_ASAP7_75t_R g4390 ( 
.A(n_4065),
.Y(n_4390)
);

INVx2_ASAP7_75t_L g4391 ( 
.A(n_3876),
.Y(n_4391)
);

NOR3xp33_ASAP7_75t_SL g4392 ( 
.A(n_4131),
.B(n_1817),
.C(n_1805),
.Y(n_4392)
);

INVx1_ASAP7_75t_L g4393 ( 
.A(n_3890),
.Y(n_4393)
);

AND2x4_ASAP7_75t_L g4394 ( 
.A(n_3819),
.B(n_11),
.Y(n_4394)
);

INVx5_ASAP7_75t_L g4395 ( 
.A(n_4035),
.Y(n_4395)
);

BUFx4f_ASAP7_75t_L g4396 ( 
.A(n_4056),
.Y(n_4396)
);

BUFx6f_ASAP7_75t_L g4397 ( 
.A(n_3896),
.Y(n_4397)
);

NAND2xp5_ASAP7_75t_L g4398 ( 
.A(n_4135),
.B(n_11),
.Y(n_4398)
);

INVx1_ASAP7_75t_L g4399 ( 
.A(n_3899),
.Y(n_4399)
);

OAI22xp5_ASAP7_75t_L g4400 ( 
.A1(n_4004),
.A2(n_1830),
.B1(n_1835),
.B2(n_1821),
.Y(n_4400)
);

AOI22xp5_ASAP7_75t_L g4401 ( 
.A1(n_3957),
.A2(n_1843),
.B1(n_1847),
.B2(n_1836),
.Y(n_4401)
);

AND3x1_ASAP7_75t_L g4402 ( 
.A(n_4057),
.B(n_12),
.C(n_13),
.Y(n_4402)
);

NAND2xp5_ASAP7_75t_SL g4403 ( 
.A(n_3981),
.B(n_1848),
.Y(n_4403)
);

NAND2xp5_ASAP7_75t_SL g4404 ( 
.A(n_3932),
.B(n_1854),
.Y(n_4404)
);

INVx2_ASAP7_75t_L g4405 ( 
.A(n_3916),
.Y(n_4405)
);

NAND2xp5_ASAP7_75t_L g4406 ( 
.A(n_4029),
.B(n_12),
.Y(n_4406)
);

BUFx4f_ASAP7_75t_L g4407 ( 
.A(n_3923),
.Y(n_4407)
);

AO21x1_ASAP7_75t_L g4408 ( 
.A1(n_3821),
.A2(n_2085),
.B(n_1878),
.Y(n_4408)
);

NAND2xp5_ASAP7_75t_L g4409 ( 
.A(n_3864),
.B(n_13),
.Y(n_4409)
);

NOR2xp33_ASAP7_75t_L g4410 ( 
.A(n_4014),
.B(n_1861),
.Y(n_4410)
);

INVx1_ASAP7_75t_L g4411 ( 
.A(n_3936),
.Y(n_4411)
);

CKINVDCx5p33_ASAP7_75t_R g4412 ( 
.A(n_3820),
.Y(n_4412)
);

AOI22xp5_ASAP7_75t_L g4413 ( 
.A1(n_3793),
.A2(n_1866),
.B1(n_1869),
.B2(n_1865),
.Y(n_4413)
);

INVx1_ASAP7_75t_L g4414 ( 
.A(n_3948),
.Y(n_4414)
);

BUFx2_ASAP7_75t_L g4415 ( 
.A(n_4061),
.Y(n_4415)
);

INVx1_ASAP7_75t_L g4416 ( 
.A(n_3992),
.Y(n_4416)
);

NAND2xp5_ASAP7_75t_L g4417 ( 
.A(n_3866),
.B(n_14),
.Y(n_4417)
);

NAND2xp33_ASAP7_75t_L g4418 ( 
.A(n_3962),
.B(n_1878),
.Y(n_4418)
);

AND2x2_ASAP7_75t_L g4419 ( 
.A(n_3912),
.B(n_15),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_3998),
.Y(n_4420)
);

AOI22xp5_ASAP7_75t_L g4421 ( 
.A1(n_3804),
.A2(n_1877),
.B1(n_1882),
.B2(n_1872),
.Y(n_4421)
);

OAI22xp33_ASAP7_75t_L g4422 ( 
.A1(n_4045),
.A2(n_1885),
.B1(n_1889),
.B2(n_1883),
.Y(n_4422)
);

NOR3xp33_ASAP7_75t_SL g4423 ( 
.A(n_3823),
.B(n_1904),
.C(n_1900),
.Y(n_4423)
);

NAND2x1p5_ASAP7_75t_L g4424 ( 
.A(n_3979),
.B(n_3883),
.Y(n_4424)
);

CKINVDCx20_ASAP7_75t_R g4425 ( 
.A(n_3822),
.Y(n_4425)
);

AND3x1_ASAP7_75t_SL g4426 ( 
.A(n_4018),
.B(n_15),
.C(n_16),
.Y(n_4426)
);

AND3x2_ASAP7_75t_SL g4427 ( 
.A(n_3912),
.B(n_18),
.C(n_19),
.Y(n_4427)
);

AOI22xp5_ASAP7_75t_L g4428 ( 
.A1(n_4053),
.A2(n_1906),
.B1(n_1911),
.B2(n_1908),
.Y(n_4428)
);

INVx1_ASAP7_75t_L g4429 ( 
.A(n_3966),
.Y(n_4429)
);

BUFx2_ASAP7_75t_L g4430 ( 
.A(n_3953),
.Y(n_4430)
);

INVx1_ASAP7_75t_L g4431 ( 
.A(n_3973),
.Y(n_4431)
);

AND3x1_ASAP7_75t_SL g4432 ( 
.A(n_4046),
.B(n_18),
.C(n_20),
.Y(n_4432)
);

CKINVDCx5p33_ASAP7_75t_R g4433 ( 
.A(n_3854),
.Y(n_4433)
);

INVx2_ASAP7_75t_L g4434 ( 
.A(n_3933),
.Y(n_4434)
);

BUFx8_ASAP7_75t_L g4435 ( 
.A(n_4144),
.Y(n_4435)
);

CKINVDCx20_ASAP7_75t_R g4436 ( 
.A(n_3805),
.Y(n_4436)
);

INVx2_ASAP7_75t_L g4437 ( 
.A(n_3935),
.Y(n_4437)
);

AOI22xp33_ASAP7_75t_L g4438 ( 
.A1(n_4023),
.A2(n_1952),
.B1(n_2102),
.B2(n_2022),
.Y(n_4438)
);

INVx1_ASAP7_75t_L g4439 ( 
.A(n_4323),
.Y(n_4439)
);

NAND2xp5_ASAP7_75t_L g4440 ( 
.A(n_4145),
.B(n_4020),
.Y(n_4440)
);

NOR2xp33_ASAP7_75t_L g4441 ( 
.A(n_4390),
.B(n_3956),
.Y(n_4441)
);

NAND2xp5_ASAP7_75t_L g4442 ( 
.A(n_4311),
.B(n_4009),
.Y(n_4442)
);

BUFx6f_ASAP7_75t_L g4443 ( 
.A(n_4161),
.Y(n_4443)
);

INVx2_ASAP7_75t_L g4444 ( 
.A(n_4276),
.Y(n_4444)
);

NOR2xp33_ASAP7_75t_L g4445 ( 
.A(n_4149),
.B(n_3795),
.Y(n_4445)
);

CKINVDCx14_ASAP7_75t_R g4446 ( 
.A(n_4204),
.Y(n_4446)
);

INVx3_ASAP7_75t_L g4447 ( 
.A(n_4161),
.Y(n_4447)
);

INVx1_ASAP7_75t_L g4448 ( 
.A(n_4169),
.Y(n_4448)
);

NAND2xp5_ASAP7_75t_L g4449 ( 
.A(n_4274),
.B(n_4011),
.Y(n_4449)
);

AND3x2_ASAP7_75t_SL g4450 ( 
.A(n_4427),
.B(n_3856),
.C(n_3857),
.Y(n_4450)
);

NAND2xp5_ASAP7_75t_SL g4451 ( 
.A(n_4203),
.B(n_4075),
.Y(n_4451)
);

NOR2xp67_ASAP7_75t_L g4452 ( 
.A(n_4228),
.B(n_3794),
.Y(n_4452)
);

NAND2xp5_ASAP7_75t_SL g4453 ( 
.A(n_4208),
.B(n_4077),
.Y(n_4453)
);

NAND2xp5_ASAP7_75t_L g4454 ( 
.A(n_4159),
.B(n_4355),
.Y(n_4454)
);

NOR2xp33_ASAP7_75t_L g4455 ( 
.A(n_4364),
.B(n_4003),
.Y(n_4455)
);

INVx4_ASAP7_75t_L g4456 ( 
.A(n_4157),
.Y(n_4456)
);

OAI21xp33_ASAP7_75t_L g4457 ( 
.A1(n_4221),
.A2(n_4001),
.B(n_3927),
.Y(n_4457)
);

INVxp67_ASAP7_75t_L g4458 ( 
.A(n_4189),
.Y(n_4458)
);

BUFx6f_ASAP7_75t_L g4459 ( 
.A(n_4148),
.Y(n_4459)
);

NOR2xp33_ASAP7_75t_L g4460 ( 
.A(n_4162),
.B(n_4066),
.Y(n_4460)
);

O2A1O1Ixp33_ASAP7_75t_L g4461 ( 
.A1(n_4406),
.A2(n_3977),
.B(n_3851),
.C(n_4049),
.Y(n_4461)
);

NAND2xp5_ASAP7_75t_SL g4462 ( 
.A(n_4243),
.B(n_4068),
.Y(n_4462)
);

INVx2_ASAP7_75t_SL g4463 ( 
.A(n_4252),
.Y(n_4463)
);

INVx1_ASAP7_75t_L g4464 ( 
.A(n_4179),
.Y(n_4464)
);

INVx1_ASAP7_75t_L g4465 ( 
.A(n_4180),
.Y(n_4465)
);

NAND2xp5_ASAP7_75t_L g4466 ( 
.A(n_4380),
.B(n_4242),
.Y(n_4466)
);

INVx2_ASAP7_75t_L g4467 ( 
.A(n_4146),
.Y(n_4467)
);

INVx3_ASAP7_75t_L g4468 ( 
.A(n_4187),
.Y(n_4468)
);

BUFx2_ASAP7_75t_L g4469 ( 
.A(n_4205),
.Y(n_4469)
);

INVx1_ASAP7_75t_L g4470 ( 
.A(n_4181),
.Y(n_4470)
);

CKINVDCx6p67_ASAP7_75t_R g4471 ( 
.A(n_4228),
.Y(n_4471)
);

AOI22xp5_ASAP7_75t_L g4472 ( 
.A1(n_4178),
.A2(n_4008),
.B1(n_4010),
.B2(n_3937),
.Y(n_4472)
);

BUFx3_ASAP7_75t_L g4473 ( 
.A(n_4187),
.Y(n_4473)
);

INVx1_ASAP7_75t_L g4474 ( 
.A(n_4207),
.Y(n_4474)
);

BUFx4f_ASAP7_75t_L g4475 ( 
.A(n_4193),
.Y(n_4475)
);

NAND2xp5_ASAP7_75t_L g4476 ( 
.A(n_4164),
.B(n_3867),
.Y(n_4476)
);

CKINVDCx5p33_ASAP7_75t_R g4477 ( 
.A(n_4230),
.Y(n_4477)
);

NAND2xp5_ASAP7_75t_L g4478 ( 
.A(n_4437),
.B(n_3868),
.Y(n_4478)
);

INVx1_ASAP7_75t_SL g4479 ( 
.A(n_4247),
.Y(n_4479)
);

INVx1_ASAP7_75t_L g4480 ( 
.A(n_4209),
.Y(n_4480)
);

INVx1_ASAP7_75t_L g4481 ( 
.A(n_4216),
.Y(n_4481)
);

BUFx6f_ASAP7_75t_L g4482 ( 
.A(n_4215),
.Y(n_4482)
);

AND2x4_ASAP7_75t_L g4483 ( 
.A(n_4198),
.B(n_3811),
.Y(n_4483)
);

BUFx4f_ASAP7_75t_L g4484 ( 
.A(n_4297),
.Y(n_4484)
);

INVx2_ASAP7_75t_L g4485 ( 
.A(n_4182),
.Y(n_4485)
);

NAND2xp5_ASAP7_75t_L g4486 ( 
.A(n_4178),
.B(n_3870),
.Y(n_4486)
);

AND2x4_ASAP7_75t_L g4487 ( 
.A(n_4151),
.B(n_4042),
.Y(n_4487)
);

AND2x2_ASAP7_75t_L g4488 ( 
.A(n_4336),
.B(n_3886),
.Y(n_4488)
);

NAND2xp5_ASAP7_75t_L g4489 ( 
.A(n_4178),
.B(n_3887),
.Y(n_4489)
);

O2A1O1Ixp33_ASAP7_75t_L g4490 ( 
.A1(n_4398),
.A2(n_4043),
.B(n_4039),
.C(n_4000),
.Y(n_4490)
);

A2O1A1Ixp33_ASAP7_75t_L g4491 ( 
.A1(n_4329),
.A2(n_4107),
.B(n_4139),
.C(n_3963),
.Y(n_4491)
);

AND2x4_ASAP7_75t_L g4492 ( 
.A(n_4220),
.B(n_4076),
.Y(n_4492)
);

BUFx3_ASAP7_75t_L g4493 ( 
.A(n_4237),
.Y(n_4493)
);

AND2x2_ASAP7_75t_L g4494 ( 
.A(n_4275),
.B(n_4002),
.Y(n_4494)
);

AND2x2_ASAP7_75t_L g4495 ( 
.A(n_4419),
.B(n_4396),
.Y(n_4495)
);

NAND2xp5_ASAP7_75t_L g4496 ( 
.A(n_4171),
.B(n_3930),
.Y(n_4496)
);

INVx2_ASAP7_75t_L g4497 ( 
.A(n_4184),
.Y(n_4497)
);

INVx2_ASAP7_75t_L g4498 ( 
.A(n_4186),
.Y(n_4498)
);

NAND2xp5_ASAP7_75t_L g4499 ( 
.A(n_4158),
.B(n_3944),
.Y(n_4499)
);

INVx2_ASAP7_75t_L g4500 ( 
.A(n_4190),
.Y(n_4500)
);

NAND2xp5_ASAP7_75t_SL g4501 ( 
.A(n_4293),
.B(n_3951),
.Y(n_4501)
);

NAND2xp5_ASAP7_75t_L g4502 ( 
.A(n_4429),
.B(n_3988),
.Y(n_4502)
);

INVx1_ASAP7_75t_SL g4503 ( 
.A(n_4215),
.Y(n_4503)
);

OR2x2_ASAP7_75t_L g4504 ( 
.A(n_4155),
.B(n_3985),
.Y(n_4504)
);

NOR2xp33_ASAP7_75t_L g4505 ( 
.A(n_4170),
.B(n_4040),
.Y(n_4505)
);

BUFx2_ASAP7_75t_L g4506 ( 
.A(n_4202),
.Y(n_4506)
);

HB1xp67_ASAP7_75t_L g4507 ( 
.A(n_4298),
.Y(n_4507)
);

AOI22xp33_ASAP7_75t_L g4508 ( 
.A1(n_4320),
.A2(n_4052),
.B1(n_4019),
.B2(n_4015),
.Y(n_4508)
);

CKINVDCx16_ASAP7_75t_R g4509 ( 
.A(n_4300),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_4224),
.Y(n_4510)
);

INVx4_ASAP7_75t_L g4511 ( 
.A(n_4152),
.Y(n_4511)
);

AND2x2_ASAP7_75t_L g4512 ( 
.A(n_4389),
.B(n_4063),
.Y(n_4512)
);

INVx1_ASAP7_75t_L g4513 ( 
.A(n_4226),
.Y(n_4513)
);

BUFx3_ASAP7_75t_L g4514 ( 
.A(n_4202),
.Y(n_4514)
);

INVx2_ASAP7_75t_L g4515 ( 
.A(n_4192),
.Y(n_4515)
);

OAI22xp5_ASAP7_75t_L g4516 ( 
.A1(n_4249),
.A2(n_3880),
.B1(n_3872),
.B2(n_4064),
.Y(n_4516)
);

NAND2xp5_ASAP7_75t_L g4517 ( 
.A(n_4431),
.B(n_3901),
.Y(n_4517)
);

INVx1_ASAP7_75t_L g4518 ( 
.A(n_4231),
.Y(n_4518)
);

NAND2xp5_ASAP7_75t_L g4519 ( 
.A(n_4434),
.B(n_4016),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_L g4520 ( 
.A(n_4362),
.B(n_4021),
.Y(n_4520)
);

AND2x4_ASAP7_75t_L g4521 ( 
.A(n_4239),
.B(n_3969),
.Y(n_4521)
);

INVxp67_ASAP7_75t_L g4522 ( 
.A(n_4210),
.Y(n_4522)
);

INVx2_ASAP7_75t_L g4523 ( 
.A(n_4235),
.Y(n_4523)
);

INVx3_ASAP7_75t_L g4524 ( 
.A(n_4210),
.Y(n_4524)
);

NAND2xp5_ASAP7_75t_L g4525 ( 
.A(n_4194),
.B(n_4041),
.Y(n_4525)
);

NAND2xp5_ASAP7_75t_L g4526 ( 
.A(n_4358),
.B(n_4233),
.Y(n_4526)
);

INVx2_ASAP7_75t_L g4527 ( 
.A(n_4240),
.Y(n_4527)
);

BUFx6f_ASAP7_75t_L g4528 ( 
.A(n_4407),
.Y(n_4528)
);

INVx1_ASAP7_75t_L g4529 ( 
.A(n_4238),
.Y(n_4529)
);

NAND2xp5_ASAP7_75t_L g4530 ( 
.A(n_4246),
.B(n_3920),
.Y(n_4530)
);

AO22x1_ASAP7_75t_L g4531 ( 
.A1(n_4256),
.A2(n_4279),
.B1(n_4293),
.B2(n_4325),
.Y(n_4531)
);

AOI21xp5_ASAP7_75t_L g4532 ( 
.A1(n_4342),
.A2(n_3919),
.B(n_3924),
.Y(n_4532)
);

BUFx2_ASAP7_75t_L g4533 ( 
.A(n_4236),
.Y(n_4533)
);

CKINVDCx5p33_ASAP7_75t_R g4534 ( 
.A(n_4167),
.Y(n_4534)
);

INVx1_ASAP7_75t_SL g4535 ( 
.A(n_4296),
.Y(n_4535)
);

NAND2xp5_ASAP7_75t_L g4536 ( 
.A(n_4263),
.B(n_20),
.Y(n_4536)
);

BUFx6f_ASAP7_75t_L g4537 ( 
.A(n_4152),
.Y(n_4537)
);

INVx3_ASAP7_75t_L g4538 ( 
.A(n_4199),
.Y(n_4538)
);

NAND2xp5_ASAP7_75t_L g4539 ( 
.A(n_4277),
.B(n_21),
.Y(n_4539)
);

NAND2xp5_ASAP7_75t_L g4540 ( 
.A(n_4283),
.B(n_4284),
.Y(n_4540)
);

AOI22x1_ASAP7_75t_L g4541 ( 
.A1(n_4257),
.A2(n_1925),
.B1(n_1937),
.B2(n_1921),
.Y(n_4541)
);

AND2x2_ASAP7_75t_L g4542 ( 
.A(n_4251),
.B(n_21),
.Y(n_4542)
);

INVx3_ASAP7_75t_L g4543 ( 
.A(n_4153),
.Y(n_4543)
);

NAND2xp5_ASAP7_75t_L g4544 ( 
.A(n_4290),
.B(n_22),
.Y(n_4544)
);

OAI22xp5_ASAP7_75t_L g4545 ( 
.A1(n_4286),
.A2(n_1942),
.B1(n_1948),
.B2(n_1940),
.Y(n_4545)
);

NAND2xp5_ASAP7_75t_L g4546 ( 
.A(n_4291),
.B(n_22),
.Y(n_4546)
);

INVx1_ASAP7_75t_L g4547 ( 
.A(n_4292),
.Y(n_4547)
);

BUFx2_ASAP7_75t_L g4548 ( 
.A(n_4425),
.Y(n_4548)
);

NAND2xp5_ASAP7_75t_L g4549 ( 
.A(n_4294),
.B(n_23),
.Y(n_4549)
);

AOI22xp5_ASAP7_75t_L g4550 ( 
.A1(n_4201),
.A2(n_1954),
.B1(n_1959),
.B2(n_1957),
.Y(n_4550)
);

HB1xp67_ASAP7_75t_SL g4551 ( 
.A(n_4191),
.Y(n_4551)
);

INVx2_ASAP7_75t_L g4552 ( 
.A(n_4244),
.Y(n_4552)
);

AND2x4_ASAP7_75t_L g4553 ( 
.A(n_4239),
.B(n_1231),
.Y(n_4553)
);

INVx3_ASAP7_75t_L g4554 ( 
.A(n_4153),
.Y(n_4554)
);

BUFx2_ASAP7_75t_L g4555 ( 
.A(n_4350),
.Y(n_4555)
);

HB1xp67_ASAP7_75t_L g4556 ( 
.A(n_4334),
.Y(n_4556)
);

HB1xp67_ASAP7_75t_L g4557 ( 
.A(n_4299),
.Y(n_4557)
);

INVxp33_ASAP7_75t_SL g4558 ( 
.A(n_4232),
.Y(n_4558)
);

NAND2xp5_ASAP7_75t_L g4559 ( 
.A(n_4302),
.B(n_23),
.Y(n_4559)
);

INVx2_ASAP7_75t_L g4560 ( 
.A(n_4264),
.Y(n_4560)
);

BUFx2_ASAP7_75t_L g4561 ( 
.A(n_4412),
.Y(n_4561)
);

NOR2xp33_ASAP7_75t_L g4562 ( 
.A(n_4288),
.B(n_1976),
.Y(n_4562)
);

NAND2xp5_ASAP7_75t_L g4563 ( 
.A(n_4303),
.B(n_24),
.Y(n_4563)
);

INVx1_ASAP7_75t_L g4564 ( 
.A(n_4304),
.Y(n_4564)
);

INVx1_ASAP7_75t_SL g4565 ( 
.A(n_4430),
.Y(n_4565)
);

INVx1_ASAP7_75t_L g4566 ( 
.A(n_4310),
.Y(n_4566)
);

NOR2xp33_ASAP7_75t_L g4567 ( 
.A(n_4415),
.B(n_1978),
.Y(n_4567)
);

INVx1_ASAP7_75t_L g4568 ( 
.A(n_4322),
.Y(n_4568)
);

NAND2xp5_ASAP7_75t_L g4569 ( 
.A(n_4176),
.B(n_24),
.Y(n_4569)
);

BUFx2_ASAP7_75t_L g4570 ( 
.A(n_4436),
.Y(n_4570)
);

NAND2xp5_ASAP7_75t_L g4571 ( 
.A(n_4281),
.B(n_25),
.Y(n_4571)
);

BUFx3_ASAP7_75t_L g4572 ( 
.A(n_4147),
.Y(n_4572)
);

NAND2xp5_ASAP7_75t_L g4573 ( 
.A(n_4282),
.B(n_4308),
.Y(n_4573)
);

INVx1_ASAP7_75t_L g4574 ( 
.A(n_4324),
.Y(n_4574)
);

AND2x2_ASAP7_75t_L g4575 ( 
.A(n_4160),
.B(n_25),
.Y(n_4575)
);

INVx2_ASAP7_75t_SL g4576 ( 
.A(n_4289),
.Y(n_4576)
);

AND2x2_ASAP7_75t_L g4577 ( 
.A(n_4156),
.B(n_26),
.Y(n_4577)
);

INVx3_ASAP7_75t_L g4578 ( 
.A(n_4289),
.Y(n_4578)
);

INVx1_ASAP7_75t_L g4579 ( 
.A(n_4327),
.Y(n_4579)
);

BUFx6f_ASAP7_75t_L g4580 ( 
.A(n_4301),
.Y(n_4580)
);

INVx1_ASAP7_75t_L g4581 ( 
.A(n_4328),
.Y(n_4581)
);

INVx2_ASAP7_75t_L g4582 ( 
.A(n_4330),
.Y(n_4582)
);

NOR2xp33_ASAP7_75t_L g4583 ( 
.A(n_4316),
.B(n_1979),
.Y(n_4583)
);

BUFx3_ASAP7_75t_L g4584 ( 
.A(n_4307),
.Y(n_4584)
);

HB1xp67_ASAP7_75t_L g4585 ( 
.A(n_4172),
.Y(n_4585)
);

INVx1_ASAP7_75t_L g4586 ( 
.A(n_4344),
.Y(n_4586)
);

INVx3_ASAP7_75t_L g4587 ( 
.A(n_4301),
.Y(n_4587)
);

BUFx6f_ASAP7_75t_L g4588 ( 
.A(n_4307),
.Y(n_4588)
);

NAND2xp5_ASAP7_75t_SL g4589 ( 
.A(n_4256),
.B(n_1980),
.Y(n_4589)
);

AND2x2_ASAP7_75t_L g4590 ( 
.A(n_4197),
.B(n_4261),
.Y(n_4590)
);

INVx1_ASAP7_75t_L g4591 ( 
.A(n_4346),
.Y(n_4591)
);

NAND2xp5_ASAP7_75t_L g4592 ( 
.A(n_4315),
.B(n_26),
.Y(n_4592)
);

OAI22xp5_ASAP7_75t_L g4593 ( 
.A1(n_4165),
.A2(n_1988),
.B1(n_1989),
.B2(n_1984),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_4387),
.Y(n_4594)
);

INVx2_ASAP7_75t_L g4595 ( 
.A(n_4337),
.Y(n_4595)
);

AOI22xp33_ASAP7_75t_L g4596 ( 
.A1(n_4385),
.A2(n_4325),
.B1(n_4306),
.B2(n_4225),
.Y(n_4596)
);

INVx4_ASAP7_75t_L g4597 ( 
.A(n_4268),
.Y(n_4597)
);

CKINVDCx5p33_ASAP7_75t_R g4598 ( 
.A(n_4314),
.Y(n_4598)
);

NOR2xp33_ASAP7_75t_R g4599 ( 
.A(n_4188),
.B(n_1990),
.Y(n_4599)
);

BUFx3_ASAP7_75t_L g4600 ( 
.A(n_4341),
.Y(n_4600)
);

AND2x2_ASAP7_75t_L g4601 ( 
.A(n_4285),
.B(n_28),
.Y(n_4601)
);

AOI221xp5_ASAP7_75t_L g4602 ( 
.A1(n_4234),
.A2(n_2010),
.B1(n_2013),
.B2(n_1999),
.C(n_1993),
.Y(n_4602)
);

AND2x4_ASAP7_75t_L g4603 ( 
.A(n_4279),
.B(n_1232),
.Y(n_4603)
);

INVx3_ASAP7_75t_L g4604 ( 
.A(n_4253),
.Y(n_4604)
);

NAND2xp5_ASAP7_75t_L g4605 ( 
.A(n_4278),
.B(n_28),
.Y(n_4605)
);

BUFx2_ASAP7_75t_L g4606 ( 
.A(n_4433),
.Y(n_4606)
);

INVx3_ASAP7_75t_L g4607 ( 
.A(n_4367),
.Y(n_4607)
);

AND2x2_ASAP7_75t_L g4608 ( 
.A(n_4219),
.B(n_29),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_4368),
.Y(n_4609)
);

NAND2xp5_ASAP7_75t_L g4610 ( 
.A(n_4325),
.B(n_29),
.Y(n_4610)
);

NAND2xp5_ASAP7_75t_L g4611 ( 
.A(n_4345),
.B(n_30),
.Y(n_4611)
);

INVx1_ASAP7_75t_L g4612 ( 
.A(n_4373),
.Y(n_4612)
);

OR2x2_ASAP7_75t_L g4613 ( 
.A(n_4229),
.B(n_31),
.Y(n_4613)
);

BUFx3_ASAP7_75t_L g4614 ( 
.A(n_4341),
.Y(n_4614)
);

INVx4_ASAP7_75t_L g4615 ( 
.A(n_4150),
.Y(n_4615)
);

INVx1_ASAP7_75t_L g4616 ( 
.A(n_4377),
.Y(n_4616)
);

INVx2_ASAP7_75t_SL g4617 ( 
.A(n_4395),
.Y(n_4617)
);

AND2x2_ASAP7_75t_L g4618 ( 
.A(n_4360),
.B(n_31),
.Y(n_4618)
);

AOI22xp5_ASAP7_75t_L g4619 ( 
.A1(n_4168),
.A2(n_2014),
.B1(n_2024),
.B2(n_2015),
.Y(n_4619)
);

INVx2_ASAP7_75t_L g4620 ( 
.A(n_4347),
.Y(n_4620)
);

AOI22xp5_ASAP7_75t_L g4621 ( 
.A1(n_4366),
.A2(n_2035),
.B1(n_2051),
.B2(n_2043),
.Y(n_4621)
);

NAND2xp5_ASAP7_75t_SL g4622 ( 
.A(n_4173),
.B(n_2052),
.Y(n_4622)
);

AND2x4_ASAP7_75t_L g4623 ( 
.A(n_4309),
.B(n_1233),
.Y(n_4623)
);

AND2x2_ASAP7_75t_L g4624 ( 
.A(n_4166),
.B(n_32),
.Y(n_4624)
);

NAND2xp5_ASAP7_75t_L g4625 ( 
.A(n_4352),
.B(n_32),
.Y(n_4625)
);

NOR2xp33_ASAP7_75t_L g4626 ( 
.A(n_4154),
.B(n_2056),
.Y(n_4626)
);

OAI221xp5_ASAP7_75t_L g4627 ( 
.A1(n_4259),
.A2(n_2061),
.B1(n_2066),
.B2(n_2062),
.C(n_2059),
.Y(n_4627)
);

CKINVDCx20_ASAP7_75t_R g4628 ( 
.A(n_4227),
.Y(n_4628)
);

NAND2xp5_ASAP7_75t_SL g4629 ( 
.A(n_4173),
.B(n_4365),
.Y(n_4629)
);

AOI22xp33_ASAP7_75t_L g4630 ( 
.A1(n_4383),
.A2(n_2022),
.B1(n_2479),
.B2(n_2102),
.Y(n_4630)
);

INVx2_ASAP7_75t_L g4631 ( 
.A(n_4391),
.Y(n_4631)
);

AOI22xp5_ASAP7_75t_L g4632 ( 
.A1(n_4402),
.A2(n_2069),
.B1(n_2084),
.B2(n_2074),
.Y(n_4632)
);

CKINVDCx5p33_ASAP7_75t_R g4633 ( 
.A(n_4435),
.Y(n_4633)
);

BUFx6f_ASAP7_75t_L g4634 ( 
.A(n_4386),
.Y(n_4634)
);

A2O1A1Ixp33_ASAP7_75t_L g4635 ( 
.A1(n_4321),
.A2(n_2088),
.B(n_2090),
.C(n_2086),
.Y(n_4635)
);

NAND2xp5_ASAP7_75t_L g4636 ( 
.A(n_4163),
.B(n_33),
.Y(n_4636)
);

A2O1A1Ixp33_ASAP7_75t_L g4637 ( 
.A1(n_4353),
.A2(n_2094),
.B(n_2095),
.C(n_2093),
.Y(n_4637)
);

INVx1_ASAP7_75t_L g4638 ( 
.A(n_4379),
.Y(n_4638)
);

INVx3_ASAP7_75t_SL g4639 ( 
.A(n_4150),
.Y(n_4639)
);

AOI22xp5_ASAP7_75t_L g4640 ( 
.A1(n_4426),
.A2(n_2098),
.B1(n_2112),
.B2(n_2096),
.Y(n_4640)
);

AND2x2_ASAP7_75t_L g4641 ( 
.A(n_4175),
.B(n_33),
.Y(n_4641)
);

NAND2xp5_ASAP7_75t_SL g4642 ( 
.A(n_4173),
.B(n_2114),
.Y(n_4642)
);

INVx1_ASAP7_75t_L g4643 ( 
.A(n_4381),
.Y(n_4643)
);

NAND2xp5_ASAP7_75t_L g4644 ( 
.A(n_4340),
.B(n_34),
.Y(n_4644)
);

NAND2xp5_ASAP7_75t_L g4645 ( 
.A(n_4343),
.B(n_35),
.Y(n_4645)
);

CKINVDCx5p33_ASAP7_75t_R g4646 ( 
.A(n_4319),
.Y(n_4646)
);

INVx1_ASAP7_75t_L g4647 ( 
.A(n_4384),
.Y(n_4647)
);

OR2x6_ASAP7_75t_L g4648 ( 
.A(n_4229),
.B(n_2022),
.Y(n_4648)
);

INVx3_ASAP7_75t_L g4649 ( 
.A(n_4266),
.Y(n_4649)
);

BUFx6f_ASAP7_75t_L g4650 ( 
.A(n_4386),
.Y(n_4650)
);

INVx2_ASAP7_75t_L g4651 ( 
.A(n_4405),
.Y(n_4651)
);

CKINVDCx5p33_ASAP7_75t_R g4652 ( 
.A(n_4223),
.Y(n_4652)
);

INVx2_ASAP7_75t_L g4653 ( 
.A(n_4393),
.Y(n_4653)
);

HB1xp67_ASAP7_75t_L g4654 ( 
.A(n_4357),
.Y(n_4654)
);

INVx1_ASAP7_75t_L g4655 ( 
.A(n_4399),
.Y(n_4655)
);

AND2x2_ASAP7_75t_L g4656 ( 
.A(n_4200),
.B(n_36),
.Y(n_4656)
);

AND3x1_ASAP7_75t_SL g4657 ( 
.A(n_4349),
.B(n_37),
.C(n_38),
.Y(n_4657)
);

A2O1A1Ixp33_ASAP7_75t_L g4658 ( 
.A1(n_4356),
.A2(n_4361),
.B(n_4363),
.C(n_4359),
.Y(n_4658)
);

BUFx6f_ASAP7_75t_L g4659 ( 
.A(n_4397),
.Y(n_4659)
);

INVx2_ASAP7_75t_L g4660 ( 
.A(n_4411),
.Y(n_4660)
);

INVx1_ASAP7_75t_L g4661 ( 
.A(n_4414),
.Y(n_4661)
);

CKINVDCx5p33_ASAP7_75t_R g4662 ( 
.A(n_4312),
.Y(n_4662)
);

NAND2xp5_ASAP7_75t_SL g4663 ( 
.A(n_4395),
.B(n_2121),
.Y(n_4663)
);

BUFx3_ASAP7_75t_L g4664 ( 
.A(n_4217),
.Y(n_4664)
);

NAND2xp5_ASAP7_75t_L g4665 ( 
.A(n_4375),
.B(n_37),
.Y(n_4665)
);

BUFx12f_ASAP7_75t_L g4666 ( 
.A(n_4271),
.Y(n_4666)
);

BUFx2_ASAP7_75t_L g4667 ( 
.A(n_4267),
.Y(n_4667)
);

AOI221xp5_ASAP7_75t_SL g4668 ( 
.A1(n_4174),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.C(n_41),
.Y(n_4668)
);

INVx2_ASAP7_75t_SL g4669 ( 
.A(n_4397),
.Y(n_4669)
);

INVx2_ASAP7_75t_SL g4670 ( 
.A(n_4333),
.Y(n_4670)
);

NAND2xp5_ASAP7_75t_L g4671 ( 
.A(n_4376),
.B(n_39),
.Y(n_4671)
);

INVxp67_ASAP7_75t_L g4672 ( 
.A(n_4335),
.Y(n_4672)
);

INVx2_ASAP7_75t_L g4673 ( 
.A(n_4416),
.Y(n_4673)
);

INVx2_ASAP7_75t_L g4674 ( 
.A(n_4420),
.Y(n_4674)
);

INVx1_ASAP7_75t_SL g4675 ( 
.A(n_4271),
.Y(n_4675)
);

AOI22xp33_ASAP7_75t_L g4676 ( 
.A1(n_4318),
.A2(n_2479),
.B1(n_2482),
.B2(n_2102),
.Y(n_4676)
);

CKINVDCx5p33_ASAP7_75t_R g4677 ( 
.A(n_4195),
.Y(n_4677)
);

NOR2xp33_ASAP7_75t_L g4678 ( 
.A(n_4317),
.B(n_2132),
.Y(n_4678)
);

AND2x2_ASAP7_75t_L g4679 ( 
.A(n_4394),
.B(n_41),
.Y(n_4679)
);

BUFx12f_ASAP7_75t_L g4680 ( 
.A(n_4424),
.Y(n_4680)
);

NOR2xp33_ASAP7_75t_L g4681 ( 
.A(n_4354),
.B(n_2135),
.Y(n_4681)
);

AND2x2_ASAP7_75t_L g4682 ( 
.A(n_4287),
.B(n_42),
.Y(n_4682)
);

NOR2xp33_ASAP7_75t_L g4683 ( 
.A(n_4369),
.B(n_2139),
.Y(n_4683)
);

NAND2xp5_ASAP7_75t_L g4684 ( 
.A(n_4378),
.B(n_42),
.Y(n_4684)
);

NAND2xp5_ASAP7_75t_L g4685 ( 
.A(n_4185),
.B(n_4206),
.Y(n_4685)
);

AND2x4_ASAP7_75t_SL g4686 ( 
.A(n_4423),
.B(n_2479),
.Y(n_4686)
);

AND2x2_ASAP7_75t_SL g4687 ( 
.A(n_4382),
.B(n_2482),
.Y(n_4687)
);

BUFx2_ASAP7_75t_L g4688 ( 
.A(n_4370),
.Y(n_4688)
);

INVx4_ASAP7_75t_L g4689 ( 
.A(n_4218),
.Y(n_4689)
);

BUFx3_ASAP7_75t_L g4690 ( 
.A(n_4348),
.Y(n_4690)
);

NAND2xp5_ASAP7_75t_L g4691 ( 
.A(n_4212),
.B(n_44),
.Y(n_4691)
);

BUFx6f_ASAP7_75t_L g4692 ( 
.A(n_4269),
.Y(n_4692)
);

BUFx3_ASAP7_75t_L g4693 ( 
.A(n_4409),
.Y(n_4693)
);

INVx3_ASAP7_75t_SL g4694 ( 
.A(n_4196),
.Y(n_4694)
);

OAI22xp5_ASAP7_75t_SL g4695 ( 
.A1(n_4410),
.A2(n_2154),
.B1(n_2155),
.B2(n_2140),
.Y(n_4695)
);

NAND2xp5_ASAP7_75t_L g4696 ( 
.A(n_4213),
.B(n_46),
.Y(n_4696)
);

NAND2xp5_ASAP7_75t_L g4697 ( 
.A(n_4222),
.B(n_46),
.Y(n_4697)
);

INVx4_ASAP7_75t_L g4698 ( 
.A(n_4432),
.Y(n_4698)
);

NAND2xp5_ASAP7_75t_L g4699 ( 
.A(n_4241),
.B(n_47),
.Y(n_4699)
);

INVx2_ASAP7_75t_L g4700 ( 
.A(n_4331),
.Y(n_4700)
);

INVx2_ASAP7_75t_L g4701 ( 
.A(n_4417),
.Y(n_4701)
);

NAND2xp5_ASAP7_75t_L g4702 ( 
.A(n_4245),
.B(n_47),
.Y(n_4702)
);

INVx2_ASAP7_75t_L g4703 ( 
.A(n_4177),
.Y(n_4703)
);

NAND2xp5_ASAP7_75t_L g4704 ( 
.A(n_4248),
.B(n_4254),
.Y(n_4704)
);

OAI22xp5_ASAP7_75t_L g4705 ( 
.A1(n_4258),
.A2(n_2165),
.B1(n_2170),
.B2(n_2164),
.Y(n_4705)
);

AND2x2_ASAP7_75t_SL g4706 ( 
.A(n_4418),
.B(n_2482),
.Y(n_4706)
);

CKINVDCx5p33_ASAP7_75t_R g4707 ( 
.A(n_4371),
.Y(n_4707)
);

BUFx6f_ASAP7_75t_L g4708 ( 
.A(n_4272),
.Y(n_4708)
);

AND2x2_ASAP7_75t_SL g4709 ( 
.A(n_4438),
.B(n_2555),
.Y(n_4709)
);

NAND2xp5_ASAP7_75t_L g4710 ( 
.A(n_4260),
.B(n_48),
.Y(n_4710)
);

INVx1_ASAP7_75t_L g4711 ( 
.A(n_4305),
.Y(n_4711)
);

NAND2xp5_ASAP7_75t_L g4712 ( 
.A(n_4265),
.B(n_4270),
.Y(n_4712)
);

INVx1_ASAP7_75t_L g4713 ( 
.A(n_4250),
.Y(n_4713)
);

INVx2_ASAP7_75t_SL g4714 ( 
.A(n_4211),
.Y(n_4714)
);

INVx1_ASAP7_75t_L g4715 ( 
.A(n_4273),
.Y(n_4715)
);

INVx2_ASAP7_75t_L g4716 ( 
.A(n_4404),
.Y(n_4716)
);

NOR2xp33_ASAP7_75t_L g4717 ( 
.A(n_4262),
.B(n_2173),
.Y(n_4717)
);

OR2x6_ASAP7_75t_L g4718 ( 
.A(n_4214),
.B(n_2555),
.Y(n_4718)
);

INVx2_ASAP7_75t_L g4719 ( 
.A(n_4403),
.Y(n_4719)
);

NAND2xp5_ASAP7_75t_L g4720 ( 
.A(n_4428),
.B(n_49),
.Y(n_4720)
);

BUFx2_ASAP7_75t_L g4721 ( 
.A(n_4392),
.Y(n_4721)
);

INVx1_ASAP7_75t_L g4722 ( 
.A(n_4332),
.Y(n_4722)
);

BUFx6f_ASAP7_75t_L g4723 ( 
.A(n_4313),
.Y(n_4723)
);

NOR2xp33_ASAP7_75t_L g4724 ( 
.A(n_4351),
.B(n_2175),
.Y(n_4724)
);

AOI22xp5_ASAP7_75t_L g4725 ( 
.A1(n_4401),
.A2(n_2189),
.B1(n_2192),
.B2(n_2177),
.Y(n_4725)
);

INVx1_ASAP7_75t_L g4726 ( 
.A(n_4338),
.Y(n_4726)
);

AND2x4_ASAP7_75t_L g4727 ( 
.A(n_4372),
.B(n_1234),
.Y(n_4727)
);

AND2x6_ASAP7_75t_L g4728 ( 
.A(n_4280),
.B(n_2555),
.Y(n_4728)
);

CKINVDCx6p67_ASAP7_75t_R g4729 ( 
.A(n_4374),
.Y(n_4729)
);

AND2x4_ASAP7_75t_L g4730 ( 
.A(n_4183),
.B(n_4255),
.Y(n_4730)
);

AND2x2_ASAP7_75t_L g4731 ( 
.A(n_4295),
.B(n_49),
.Y(n_4731)
);

BUFx2_ASAP7_75t_L g4732 ( 
.A(n_4326),
.Y(n_4732)
);

OR2x2_ASAP7_75t_SL g4733 ( 
.A(n_4422),
.B(n_2622),
.Y(n_4733)
);

AND2x4_ASAP7_75t_L g4734 ( 
.A(n_4339),
.B(n_1235),
.Y(n_4734)
);

HB1xp67_ASAP7_75t_L g4735 ( 
.A(n_4400),
.Y(n_4735)
);

AOI22xp5_ASAP7_75t_L g4736 ( 
.A1(n_4413),
.A2(n_2202),
.B1(n_2215),
.B2(n_2200),
.Y(n_4736)
);

BUFx2_ASAP7_75t_L g4737 ( 
.A(n_4421),
.Y(n_4737)
);

HB1xp67_ASAP7_75t_L g4738 ( 
.A(n_4408),
.Y(n_4738)
);

NAND3xp33_ASAP7_75t_L g4739 ( 
.A(n_4455),
.B(n_4388),
.C(n_2221),
.Y(n_4739)
);

BUFx6f_ASAP7_75t_L g4740 ( 
.A(n_4528),
.Y(n_4740)
);

OR2x2_ASAP7_75t_L g4741 ( 
.A(n_4557),
.B(n_50),
.Y(n_4741)
);

INVx1_ASAP7_75t_SL g4742 ( 
.A(n_4555),
.Y(n_4742)
);

OAI21x1_ASAP7_75t_L g4743 ( 
.A1(n_4722),
.A2(n_2085),
.B(n_1878),
.Y(n_4743)
);

NAND2x1p5_ASAP7_75t_L g4744 ( 
.A(n_4528),
.B(n_2622),
.Y(n_4744)
);

NAND2xp5_ASAP7_75t_L g4745 ( 
.A(n_4454),
.B(n_50),
.Y(n_4745)
);

OAI21x1_ASAP7_75t_SL g4746 ( 
.A1(n_4486),
.A2(n_51),
.B(n_52),
.Y(n_4746)
);

AND2x4_ASAP7_75t_L g4747 ( 
.A(n_4473),
.B(n_51),
.Y(n_4747)
);

NAND2xp5_ASAP7_75t_SL g4748 ( 
.A(n_4526),
.B(n_4489),
.Y(n_4748)
);

HB1xp67_ASAP7_75t_L g4749 ( 
.A(n_4507),
.Y(n_4749)
);

OAI21x1_ASAP7_75t_L g4750 ( 
.A1(n_4726),
.A2(n_2085),
.B(n_1878),
.Y(n_4750)
);

BUFx3_ASAP7_75t_L g4751 ( 
.A(n_4443),
.Y(n_4751)
);

OAI21xp5_ASAP7_75t_L g4752 ( 
.A1(n_4457),
.A2(n_2223),
.B(n_2216),
.Y(n_4752)
);

OAI21x1_ASAP7_75t_L g4753 ( 
.A1(n_4713),
.A2(n_2085),
.B(n_1878),
.Y(n_4753)
);

NOR2xp67_ASAP7_75t_L g4754 ( 
.A(n_4456),
.B(n_1236),
.Y(n_4754)
);

INVx1_ASAP7_75t_SL g4755 ( 
.A(n_4561),
.Y(n_4755)
);

INVx3_ASAP7_75t_L g4756 ( 
.A(n_4482),
.Y(n_4756)
);

AOI21xp5_ASAP7_75t_L g4757 ( 
.A1(n_4658),
.A2(n_2622),
.B(n_2248),
.Y(n_4757)
);

AO31x2_ASAP7_75t_L g4758 ( 
.A1(n_4711),
.A2(n_2184),
.A3(n_2085),
.B(n_1241),
.Y(n_4758)
);

OAI21x1_ASAP7_75t_L g4759 ( 
.A1(n_4738),
.A2(n_2184),
.B(n_1242),
.Y(n_4759)
);

INVx2_ASAP7_75t_L g4760 ( 
.A(n_4444),
.Y(n_4760)
);

BUFx3_ASAP7_75t_L g4761 ( 
.A(n_4443),
.Y(n_4761)
);

NAND2xp5_ASAP7_75t_L g4762 ( 
.A(n_4449),
.B(n_52),
.Y(n_4762)
);

OAI21x1_ASAP7_75t_L g4763 ( 
.A1(n_4629),
.A2(n_4700),
.B(n_4703),
.Y(n_4763)
);

OAI21xp5_ASAP7_75t_L g4764 ( 
.A1(n_4445),
.A2(n_2252),
.B(n_2238),
.Y(n_4764)
);

AOI21xp5_ASAP7_75t_L g4765 ( 
.A1(n_4706),
.A2(n_2255),
.B(n_2254),
.Y(n_4765)
);

CKINVDCx5p33_ASAP7_75t_R g4766 ( 
.A(n_4477),
.Y(n_4766)
);

INVx3_ASAP7_75t_L g4767 ( 
.A(n_4482),
.Y(n_4767)
);

NAND2x1p5_ASAP7_75t_L g4768 ( 
.A(n_4484),
.B(n_4463),
.Y(n_4768)
);

NAND2x1p5_ASAP7_75t_L g4769 ( 
.A(n_4475),
.B(n_1238),
.Y(n_4769)
);

OAI21xp5_ASAP7_75t_L g4770 ( 
.A1(n_4683),
.A2(n_2276),
.B(n_2257),
.Y(n_4770)
);

OAI21x1_ASAP7_75t_L g4771 ( 
.A1(n_4586),
.A2(n_2184),
.B(n_1248),
.Y(n_4771)
);

INVx2_ASAP7_75t_SL g4772 ( 
.A(n_4459),
.Y(n_4772)
);

INVx3_ASAP7_75t_L g4773 ( 
.A(n_4680),
.Y(n_4773)
);

OAI21x1_ASAP7_75t_L g4774 ( 
.A1(n_4591),
.A2(n_2184),
.B(n_1249),
.Y(n_4774)
);

AO31x2_ASAP7_75t_L g4775 ( 
.A1(n_4491),
.A2(n_2184),
.A3(n_1253),
.B(n_1255),
.Y(n_4775)
);

AOI21xp5_ASAP7_75t_L g4776 ( 
.A1(n_4451),
.A2(n_4704),
.B(n_4685),
.Y(n_4776)
);

BUFx8_ASAP7_75t_L g4777 ( 
.A(n_4606),
.Y(n_4777)
);

NAND2xp5_ASAP7_75t_SL g4778 ( 
.A(n_4687),
.B(n_2297),
.Y(n_4778)
);

AOI21xp5_ASAP7_75t_L g4779 ( 
.A1(n_4712),
.A2(n_2317),
.B(n_2298),
.Y(n_4779)
);

OAI21xp5_ASAP7_75t_L g4780 ( 
.A1(n_4460),
.A2(n_4590),
.B(n_4573),
.Y(n_4780)
);

NAND2xp5_ASAP7_75t_SL g4781 ( 
.A(n_4737),
.B(n_2327),
.Y(n_4781)
);

OAI21x1_ASAP7_75t_L g4782 ( 
.A1(n_4540),
.A2(n_4464),
.B(n_4448),
.Y(n_4782)
);

OAI21x1_ASAP7_75t_L g4783 ( 
.A1(n_4465),
.A2(n_1256),
.B(n_1243),
.Y(n_4783)
);

AOI21x1_ASAP7_75t_L g4784 ( 
.A1(n_4453),
.A2(n_2332),
.B(n_2329),
.Y(n_4784)
);

INVx2_ASAP7_75t_SL g4785 ( 
.A(n_4459),
.Y(n_4785)
);

NOR2xp33_ASAP7_75t_L g4786 ( 
.A(n_4441),
.B(n_53),
.Y(n_4786)
);

AOI21xp5_ASAP7_75t_L g4787 ( 
.A1(n_4622),
.A2(n_2344),
.B(n_2338),
.Y(n_4787)
);

AOI21xp5_ASAP7_75t_L g4788 ( 
.A1(n_4642),
.A2(n_2377),
.B(n_2360),
.Y(n_4788)
);

NAND2xp5_ASAP7_75t_L g4789 ( 
.A(n_4715),
.B(n_53),
.Y(n_4789)
);

CKINVDCx20_ASAP7_75t_R g4790 ( 
.A(n_4628),
.Y(n_4790)
);

OAI21xp5_ASAP7_75t_L g4791 ( 
.A1(n_4735),
.A2(n_2381),
.B(n_2378),
.Y(n_4791)
);

NOR2x1_ASAP7_75t_SL g4792 ( 
.A(n_4648),
.B(n_54),
.Y(n_4792)
);

INVx1_ASAP7_75t_L g4793 ( 
.A(n_4439),
.Y(n_4793)
);

NAND2x1p5_ASAP7_75t_L g4794 ( 
.A(n_4537),
.B(n_4514),
.Y(n_4794)
);

AOI21xp5_ASAP7_75t_L g4795 ( 
.A1(n_4496),
.A2(n_2385),
.B(n_2384),
.Y(n_4795)
);

INVx2_ASAP7_75t_L g4796 ( 
.A(n_4653),
.Y(n_4796)
);

OAI21xp33_ASAP7_75t_L g4797 ( 
.A1(n_4720),
.A2(n_2419),
.B(n_2418),
.Y(n_4797)
);

INVx1_ASAP7_75t_L g4798 ( 
.A(n_4470),
.Y(n_4798)
);

NAND2xp5_ASAP7_75t_SL g4799 ( 
.A(n_4689),
.B(n_2421),
.Y(n_4799)
);

AO31x2_ASAP7_75t_L g4800 ( 
.A1(n_4701),
.A2(n_1260),
.A3(n_1266),
.B(n_1258),
.Y(n_4800)
);

A2O1A1Ixp33_ASAP7_75t_L g4801 ( 
.A1(n_4490),
.A2(n_2436),
.B(n_2443),
.C(n_2435),
.Y(n_4801)
);

INVx1_ASAP7_75t_L g4802 ( 
.A(n_4474),
.Y(n_4802)
);

AOI21xp5_ASAP7_75t_L g4803 ( 
.A1(n_4461),
.A2(n_2462),
.B(n_2444),
.Y(n_4803)
);

AOI21xp5_ASAP7_75t_L g4804 ( 
.A1(n_4516),
.A2(n_2468),
.B(n_2465),
.Y(n_4804)
);

OAI21x1_ASAP7_75t_L g4805 ( 
.A1(n_4480),
.A2(n_1269),
.B(n_1267),
.Y(n_4805)
);

AO21x1_ASAP7_75t_L g4806 ( 
.A1(n_4462),
.A2(n_54),
.B(n_55),
.Y(n_4806)
);

O2A1O1Ixp5_ASAP7_75t_L g4807 ( 
.A1(n_4698),
.A2(n_59),
.B(n_57),
.C(n_58),
.Y(n_4807)
);

OAI21x1_ASAP7_75t_L g4808 ( 
.A1(n_4481),
.A2(n_1272),
.B(n_1270),
.Y(n_4808)
);

AO31x2_ASAP7_75t_L g4809 ( 
.A1(n_4609),
.A2(n_1274),
.A3(n_1275),
.B(n_1273),
.Y(n_4809)
);

BUFx3_ASAP7_75t_L g4810 ( 
.A(n_4447),
.Y(n_4810)
);

AOI22xp5_ASAP7_75t_L g4811 ( 
.A1(n_4732),
.A2(n_2474),
.B1(n_2481),
.B2(n_2469),
.Y(n_4811)
);

NAND2xp5_ASAP7_75t_L g4812 ( 
.A(n_4478),
.B(n_59),
.Y(n_4812)
);

BUFx6f_ASAP7_75t_L g4813 ( 
.A(n_4537),
.Y(n_4813)
);

OAI21x1_ASAP7_75t_L g4814 ( 
.A1(n_4510),
.A2(n_1282),
.B(n_1279),
.Y(n_4814)
);

OAI21xp5_ASAP7_75t_L g4815 ( 
.A1(n_4520),
.A2(n_2493),
.B(n_2491),
.Y(n_4815)
);

AO21x1_ASAP7_75t_L g4816 ( 
.A1(n_4610),
.A2(n_60),
.B(n_61),
.Y(n_4816)
);

AND2x2_ASAP7_75t_L g4817 ( 
.A(n_4542),
.B(n_60),
.Y(n_4817)
);

BUFx12f_ASAP7_75t_L g4818 ( 
.A(n_4633),
.Y(n_4818)
);

NAND2xp5_ASAP7_75t_L g4819 ( 
.A(n_4458),
.B(n_61),
.Y(n_4819)
);

OAI21x1_ASAP7_75t_L g4820 ( 
.A1(n_4513),
.A2(n_4529),
.B(n_4518),
.Y(n_4820)
);

AOI21xp5_ASAP7_75t_L g4821 ( 
.A1(n_4665),
.A2(n_2509),
.B(n_2496),
.Y(n_4821)
);

NAND2xp5_ASAP7_75t_L g4822 ( 
.A(n_4488),
.B(n_62),
.Y(n_4822)
);

AND2x2_ASAP7_75t_L g4823 ( 
.A(n_4494),
.B(n_62),
.Y(n_4823)
);

OR2x2_ASAP7_75t_L g4824 ( 
.A(n_4594),
.B(n_63),
.Y(n_4824)
);

OAI21x1_ASAP7_75t_L g4825 ( 
.A1(n_4547),
.A2(n_1285),
.B(n_1284),
.Y(n_4825)
);

HB1xp67_ASAP7_75t_L g4826 ( 
.A(n_4469),
.Y(n_4826)
);

INVx2_ASAP7_75t_L g4827 ( 
.A(n_4660),
.Y(n_4827)
);

NAND2xp5_ASAP7_75t_SL g4828 ( 
.A(n_4690),
.B(n_4693),
.Y(n_4828)
);

OAI21x1_ASAP7_75t_L g4829 ( 
.A1(n_4564),
.A2(n_1287),
.B(n_1286),
.Y(n_4829)
);

OAI21x1_ASAP7_75t_L g4830 ( 
.A1(n_4566),
.A2(n_1289),
.B(n_1288),
.Y(n_4830)
);

INVxp67_ASAP7_75t_SL g4831 ( 
.A(n_4466),
.Y(n_4831)
);

AOI21xp5_ASAP7_75t_L g4832 ( 
.A1(n_4671),
.A2(n_2526),
.B(n_2510),
.Y(n_4832)
);

BUFx2_ASAP7_75t_L g4833 ( 
.A(n_4646),
.Y(n_4833)
);

CKINVDCx20_ASAP7_75t_R g4834 ( 
.A(n_4446),
.Y(n_4834)
);

OA22x2_ASAP7_75t_L g4835 ( 
.A1(n_4472),
.A2(n_2529),
.B1(n_2537),
.B2(n_2528),
.Y(n_4835)
);

BUFx4_ASAP7_75t_SL g4836 ( 
.A(n_4534),
.Y(n_4836)
);

A2O1A1Ixp33_ASAP7_75t_L g4837 ( 
.A1(n_4596),
.A2(n_2541),
.B(n_2542),
.C(n_2539),
.Y(n_4837)
);

AND2x2_ASAP7_75t_L g4838 ( 
.A(n_4679),
.B(n_63),
.Y(n_4838)
);

OAI21x1_ASAP7_75t_L g4839 ( 
.A1(n_4568),
.A2(n_1292),
.B(n_1290),
.Y(n_4839)
);

NAND2xp5_ASAP7_75t_L g4840 ( 
.A(n_4479),
.B(n_64),
.Y(n_4840)
);

INVxp67_ASAP7_75t_SL g4841 ( 
.A(n_4574),
.Y(n_4841)
);

A2O1A1Ixp33_ASAP7_75t_L g4842 ( 
.A1(n_4691),
.A2(n_2549),
.B(n_2550),
.C(n_2547),
.Y(n_4842)
);

AND2x6_ASAP7_75t_SL g4843 ( 
.A(n_4483),
.B(n_64),
.Y(n_4843)
);

NOR2xp33_ASAP7_75t_L g4844 ( 
.A(n_4558),
.B(n_4721),
.Y(n_4844)
);

AND2x2_ASAP7_75t_L g4845 ( 
.A(n_4512),
.B(n_4601),
.Y(n_4845)
);

OAI21x1_ASAP7_75t_L g4846 ( 
.A1(n_4579),
.A2(n_1295),
.B(n_1293),
.Y(n_4846)
);

INVx2_ASAP7_75t_L g4847 ( 
.A(n_4673),
.Y(n_4847)
);

AOI221x1_ASAP7_75t_L g4848 ( 
.A1(n_4644),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.C(n_68),
.Y(n_4848)
);

AOI21xp5_ASAP7_75t_SL g4849 ( 
.A1(n_4501),
.A2(n_2559),
.B(n_2557),
.Y(n_4849)
);

AND2x2_ASAP7_75t_L g4850 ( 
.A(n_4641),
.B(n_66),
.Y(n_4850)
);

A2O1A1Ixp33_ASAP7_75t_L g4851 ( 
.A1(n_4696),
.A2(n_2568),
.B(n_2574),
.C(n_2561),
.Y(n_4851)
);

OAI21x1_ASAP7_75t_L g4852 ( 
.A1(n_4581),
.A2(n_4616),
.B(n_4612),
.Y(n_4852)
);

OA21x2_ASAP7_75t_L g4853 ( 
.A1(n_4668),
.A2(n_2579),
.B(n_2576),
.Y(n_4853)
);

INVx1_ASAP7_75t_L g4854 ( 
.A(n_4638),
.Y(n_4854)
);

AOI21xp5_ASAP7_75t_L g4855 ( 
.A1(n_4684),
.A2(n_2589),
.B(n_2588),
.Y(n_4855)
);

OAI22xp5_ASAP7_75t_L g4856 ( 
.A1(n_4640),
.A2(n_2610),
.B1(n_2615),
.B2(n_2599),
.Y(n_4856)
);

AOI21xp5_ASAP7_75t_L g4857 ( 
.A1(n_4645),
.A2(n_2662),
.B(n_2617),
.Y(n_4857)
);

AND2x2_ASAP7_75t_L g4858 ( 
.A(n_4656),
.B(n_67),
.Y(n_4858)
);

AOI21xp5_ASAP7_75t_L g4859 ( 
.A1(n_4611),
.A2(n_2666),
.B(n_2664),
.Y(n_4859)
);

AND2x2_ASAP7_75t_L g4860 ( 
.A(n_4608),
.B(n_68),
.Y(n_4860)
);

OAI22xp5_ASAP7_75t_L g4861 ( 
.A1(n_4697),
.A2(n_2671),
.B1(n_2680),
.B2(n_2669),
.Y(n_4861)
);

BUFx3_ASAP7_75t_L g4862 ( 
.A(n_4468),
.Y(n_4862)
);

OAI21x1_ASAP7_75t_L g4863 ( 
.A1(n_4643),
.A2(n_1299),
.B(n_1298),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4647),
.Y(n_4864)
);

OAI21xp5_ASAP7_75t_L g4865 ( 
.A1(n_4550),
.A2(n_2702),
.B(n_2701),
.Y(n_4865)
);

OAI22xp5_ASAP7_75t_L g4866 ( 
.A1(n_4699),
.A2(n_2710),
.B1(n_2711),
.B2(n_2709),
.Y(n_4866)
);

AOI21xp5_ASAP7_75t_L g4867 ( 
.A1(n_4532),
.A2(n_2724),
.B(n_2714),
.Y(n_4867)
);

A2O1A1Ixp33_ASAP7_75t_L g4868 ( 
.A1(n_4702),
.A2(n_2739),
.B(n_2743),
.C(n_2729),
.Y(n_4868)
);

OAI22xp5_ASAP7_75t_L g4869 ( 
.A1(n_4710),
.A2(n_2754),
.B1(n_2766),
.B2(n_2746),
.Y(n_4869)
);

NAND2xp5_ASAP7_75t_L g4870 ( 
.A(n_4565),
.B(n_69),
.Y(n_4870)
);

OAI21x1_ASAP7_75t_L g4871 ( 
.A1(n_4655),
.A2(n_1302),
.B(n_1300),
.Y(n_4871)
);

A2O1A1Ixp33_ASAP7_75t_L g4872 ( 
.A1(n_4571),
.A2(n_4592),
.B(n_4605),
.C(n_4583),
.Y(n_4872)
);

NAND2xp5_ASAP7_75t_L g4873 ( 
.A(n_4502),
.B(n_69),
.Y(n_4873)
);

CKINVDCx20_ASAP7_75t_R g4874 ( 
.A(n_4509),
.Y(n_4874)
);

AND2x2_ASAP7_75t_L g4875 ( 
.A(n_4624),
.B(n_4575),
.Y(n_4875)
);

BUFx2_ASAP7_75t_L g4876 ( 
.A(n_4506),
.Y(n_4876)
);

INVxp67_ASAP7_75t_L g4877 ( 
.A(n_4654),
.Y(n_4877)
);

OAI21x1_ASAP7_75t_L g4878 ( 
.A1(n_4661),
.A2(n_1305),
.B(n_1303),
.Y(n_4878)
);

AOI221x1_ASAP7_75t_L g4879 ( 
.A1(n_4440),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.C(n_73),
.Y(n_4879)
);

OAI21xp33_ASAP7_75t_L g4880 ( 
.A1(n_4569),
.A2(n_2771),
.B(n_2767),
.Y(n_4880)
);

NAND2xp5_ASAP7_75t_L g4881 ( 
.A(n_4476),
.B(n_70),
.Y(n_4881)
);

OAI21x1_ASAP7_75t_L g4882 ( 
.A1(n_4716),
.A2(n_1315),
.B(n_1313),
.Y(n_4882)
);

INVx1_ASAP7_75t_L g4883 ( 
.A(n_4674),
.Y(n_4883)
);

AND2x4_ASAP7_75t_L g4884 ( 
.A(n_4503),
.B(n_71),
.Y(n_4884)
);

INVx1_ASAP7_75t_L g4885 ( 
.A(n_4467),
.Y(n_4885)
);

NAND2xp5_ASAP7_75t_L g4886 ( 
.A(n_4499),
.B(n_72),
.Y(n_4886)
);

OAI21x1_ASAP7_75t_L g4887 ( 
.A1(n_4676),
.A2(n_4539),
.B(n_4536),
.Y(n_4887)
);

NOR2xp33_ASAP7_75t_L g4888 ( 
.A(n_4707),
.B(n_73),
.Y(n_4888)
);

A2O1A1Ixp33_ASAP7_75t_L g4889 ( 
.A1(n_4724),
.A2(n_2779),
.B(n_2775),
.C(n_76),
.Y(n_4889)
);

NAND2xp5_ASAP7_75t_L g4890 ( 
.A(n_4607),
.B(n_74),
.Y(n_4890)
);

AOI22xp5_ASAP7_75t_L g4891 ( 
.A1(n_4730),
.A2(n_77),
.B1(n_74),
.B2(n_75),
.Y(n_4891)
);

OAI21x1_ASAP7_75t_SL g4892 ( 
.A1(n_4544),
.A2(n_75),
.B(n_77),
.Y(n_4892)
);

AOI21xp5_ASAP7_75t_L g4893 ( 
.A1(n_4709),
.A2(n_78),
.B(n_79),
.Y(n_4893)
);

HB1xp67_ASAP7_75t_L g4894 ( 
.A(n_4672),
.Y(n_4894)
);

AO31x2_ASAP7_75t_L g4895 ( 
.A1(n_4485),
.A2(n_1318),
.A3(n_1319),
.B(n_1317),
.Y(n_4895)
);

INVx1_ASAP7_75t_L g4896 ( 
.A(n_4497),
.Y(n_4896)
);

NAND2xp5_ASAP7_75t_L g4897 ( 
.A(n_4442),
.B(n_78),
.Y(n_4897)
);

OAI21x1_ASAP7_75t_L g4898 ( 
.A1(n_4546),
.A2(n_1323),
.B(n_1322),
.Y(n_4898)
);

BUFx10_ASAP7_75t_L g4899 ( 
.A(n_4598),
.Y(n_4899)
);

AOI21xp5_ASAP7_75t_L g4900 ( 
.A1(n_4531),
.A2(n_79),
.B(n_80),
.Y(n_4900)
);

OAI21xp5_ASAP7_75t_L g4901 ( 
.A1(n_4562),
.A2(n_80),
.B(n_82),
.Y(n_4901)
);

OAI21x1_ASAP7_75t_L g4902 ( 
.A1(n_4549),
.A2(n_1325),
.B(n_1324),
.Y(n_4902)
);

AOI211x1_ASAP7_75t_L g4903 ( 
.A1(n_4682),
.A2(n_84),
.B(n_82),
.C(n_83),
.Y(n_4903)
);

OAI21x1_ASAP7_75t_L g4904 ( 
.A1(n_4559),
.A2(n_1329),
.B(n_1328),
.Y(n_4904)
);

AOI21xp5_ASAP7_75t_L g4905 ( 
.A1(n_4505),
.A2(n_83),
.B(n_85),
.Y(n_4905)
);

BUFx12f_ASAP7_75t_L g4906 ( 
.A(n_4666),
.Y(n_4906)
);

AO31x2_ASAP7_75t_L g4907 ( 
.A1(n_4498),
.A2(n_1332),
.A3(n_1338),
.B(n_1331),
.Y(n_4907)
);

AOI21xp5_ASAP7_75t_L g4908 ( 
.A1(n_4636),
.A2(n_85),
.B(n_86),
.Y(n_4908)
);

OAI21x1_ASAP7_75t_L g4909 ( 
.A1(n_4563),
.A2(n_1341),
.B(n_1340),
.Y(n_4909)
);

INVx3_ASAP7_75t_L g4910 ( 
.A(n_4580),
.Y(n_4910)
);

NOR2xp33_ASAP7_75t_L g4911 ( 
.A(n_4556),
.B(n_86),
.Y(n_4911)
);

NAND2xp5_ASAP7_75t_L g4912 ( 
.A(n_4585),
.B(n_87),
.Y(n_4912)
);

AOI21x1_ASAP7_75t_SL g4913 ( 
.A1(n_4731),
.A2(n_87),
.B(n_88),
.Y(n_4913)
);

NAND2x1p5_ASAP7_75t_L g4914 ( 
.A(n_4580),
.B(n_1344),
.Y(n_4914)
);

OAI21x1_ASAP7_75t_SL g4915 ( 
.A1(n_4625),
.A2(n_88),
.B(n_89),
.Y(n_4915)
);

NAND2xp5_ASAP7_75t_L g4916 ( 
.A(n_4504),
.B(n_90),
.Y(n_4916)
);

OAI21x1_ASAP7_75t_L g4917 ( 
.A1(n_4719),
.A2(n_1350),
.B(n_1345),
.Y(n_4917)
);

AOI21xp5_ASAP7_75t_L g4918 ( 
.A1(n_4530),
.A2(n_90),
.B(n_91),
.Y(n_4918)
);

OAI21x1_ASAP7_75t_L g4919 ( 
.A1(n_4630),
.A2(n_1353),
.B(n_1351),
.Y(n_4919)
);

AO31x2_ASAP7_75t_L g4920 ( 
.A1(n_4500),
.A2(n_4515),
.A3(n_4527),
.B(n_4523),
.Y(n_4920)
);

NAND2xp5_ASAP7_75t_L g4921 ( 
.A(n_4670),
.B(n_91),
.Y(n_4921)
);

A2O1A1Ixp33_ASAP7_75t_L g4922 ( 
.A1(n_4681),
.A2(n_94),
.B(n_92),
.C(n_93),
.Y(n_4922)
);

NAND2xp5_ASAP7_75t_L g4923 ( 
.A(n_4667),
.B(n_92),
.Y(n_4923)
);

NAND2xp5_ASAP7_75t_L g4924 ( 
.A(n_4495),
.B(n_94),
.Y(n_4924)
);

OAI21x1_ASAP7_75t_L g4925 ( 
.A1(n_4552),
.A2(n_1355),
.B(n_1354),
.Y(n_4925)
);

AND2x2_ASAP7_75t_L g4926 ( 
.A(n_4577),
.B(n_95),
.Y(n_4926)
);

AO31x2_ASAP7_75t_L g4927 ( 
.A1(n_4560),
.A2(n_1357),
.A3(n_1359),
.B(n_1356),
.Y(n_4927)
);

AOI22xp5_ASAP7_75t_L g4928 ( 
.A1(n_4677),
.A2(n_99),
.B1(n_96),
.B2(n_98),
.Y(n_4928)
);

OAI21x1_ASAP7_75t_L g4929 ( 
.A1(n_4582),
.A2(n_4620),
.B(n_4595),
.Y(n_4929)
);

BUFx6f_ASAP7_75t_L g4930 ( 
.A(n_4471),
.Y(n_4930)
);

OAI21x1_ASAP7_75t_L g4931 ( 
.A1(n_4631),
.A2(n_1361),
.B(n_1360),
.Y(n_4931)
);

NAND2xp5_ASAP7_75t_L g4932 ( 
.A(n_4675),
.B(n_96),
.Y(n_4932)
);

NAND2xp5_ASAP7_75t_L g4933 ( 
.A(n_4533),
.B(n_98),
.Y(n_4933)
);

AOI21xp5_ASAP7_75t_L g4934 ( 
.A1(n_4637),
.A2(n_99),
.B(n_100),
.Y(n_4934)
);

OAI21x1_ASAP7_75t_L g4935 ( 
.A1(n_4651),
.A2(n_1363),
.B(n_1362),
.Y(n_4935)
);

AO31x2_ASAP7_75t_L g4936 ( 
.A1(n_4635),
.A2(n_1366),
.A3(n_1367),
.B(n_1365),
.Y(n_4936)
);

AO31x2_ASAP7_75t_L g4937 ( 
.A1(n_4688),
.A2(n_1369),
.A3(n_1371),
.B(n_1368),
.Y(n_4937)
);

NAND2xp5_ASAP7_75t_L g4938 ( 
.A(n_4517),
.B(n_100),
.Y(n_4938)
);

OAI21x1_ASAP7_75t_L g4939 ( 
.A1(n_4589),
.A2(n_1376),
.B(n_1372),
.Y(n_4939)
);

NAND2xp5_ASAP7_75t_L g4940 ( 
.A(n_4669),
.B(n_101),
.Y(n_4940)
);

OA22x2_ASAP7_75t_L g4941 ( 
.A1(n_4648),
.A2(n_103),
.B1(n_101),
.B2(n_102),
.Y(n_4941)
);

BUFx6f_ASAP7_75t_L g4942 ( 
.A(n_4588),
.Y(n_4942)
);

NAND2xp33_ASAP7_75t_L g4943 ( 
.A(n_4652),
.B(n_102),
.Y(n_4943)
);

OAI22xp5_ASAP7_75t_L g4944 ( 
.A1(n_4632),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.Y(n_4944)
);

AO31x2_ASAP7_75t_L g4945 ( 
.A1(n_4705),
.A2(n_1378),
.A3(n_1379),
.B(n_1377),
.Y(n_4945)
);

NAND2xp5_ASAP7_75t_L g4946 ( 
.A(n_4634),
.B(n_105),
.Y(n_4946)
);

INVxp67_ASAP7_75t_L g4947 ( 
.A(n_4548),
.Y(n_4947)
);

BUFx2_ASAP7_75t_SL g4948 ( 
.A(n_4452),
.Y(n_4948)
);

NAND2xp5_ASAP7_75t_L g4949 ( 
.A(n_4634),
.B(n_106),
.Y(n_4949)
);

OAI21x1_ASAP7_75t_L g4950 ( 
.A1(n_4663),
.A2(n_1382),
.B(n_1381),
.Y(n_4950)
);

NAND2xp5_ASAP7_75t_L g4951 ( 
.A(n_4650),
.B(n_107),
.Y(n_4951)
);

A2O1A1Ixp33_ASAP7_75t_L g4952 ( 
.A1(n_4678),
.A2(n_109),
.B(n_107),
.C(n_108),
.Y(n_4952)
);

NAND3xp33_ASAP7_75t_L g4953 ( 
.A(n_4508),
.B(n_108),
.C(n_110),
.Y(n_4953)
);

NAND2xp5_ASAP7_75t_L g4954 ( 
.A(n_4650),
.B(n_110),
.Y(n_4954)
);

OAI21x1_ASAP7_75t_L g4955 ( 
.A1(n_4519),
.A2(n_4554),
.B(n_4543),
.Y(n_4955)
);

OAI21x1_ASAP7_75t_L g4956 ( 
.A1(n_4541),
.A2(n_1384),
.B(n_1383),
.Y(n_4956)
);

AOI31xp67_ASAP7_75t_L g4957 ( 
.A1(n_4727),
.A2(n_1388),
.A3(n_1390),
.B(n_1385),
.Y(n_4957)
);

OAI21x1_ASAP7_75t_L g4958 ( 
.A1(n_4524),
.A2(n_1392),
.B(n_1391),
.Y(n_4958)
);

OAI21xp5_ASAP7_75t_L g4959 ( 
.A1(n_4627),
.A2(n_111),
.B(n_112),
.Y(n_4959)
);

INVx5_ASAP7_75t_L g4960 ( 
.A(n_4588),
.Y(n_4960)
);

BUFx3_ASAP7_75t_L g4961 ( 
.A(n_4584),
.Y(n_4961)
);

NAND2xp5_ASAP7_75t_L g4962 ( 
.A(n_4659),
.B(n_112),
.Y(n_4962)
);

OAI21xp5_ASAP7_75t_L g4963 ( 
.A1(n_4736),
.A2(n_113),
.B(n_114),
.Y(n_4963)
);

AO21x2_ASAP7_75t_L g4964 ( 
.A1(n_4621),
.A2(n_1395),
.B(n_1394),
.Y(n_4964)
);

AOI21xp5_ASAP7_75t_SL g4965 ( 
.A1(n_4603),
.A2(n_113),
.B(n_116),
.Y(n_4965)
);

AOI21x1_ASAP7_75t_L g4966 ( 
.A1(n_4718),
.A2(n_1397),
.B(n_1396),
.Y(n_4966)
);

AOI221x1_ASAP7_75t_L g4967 ( 
.A1(n_4618),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.C(n_120),
.Y(n_4967)
);

INVx4_ASAP7_75t_L g4968 ( 
.A(n_4597),
.Y(n_4968)
);

OAI22x1_ASAP7_75t_L g4969 ( 
.A1(n_4639),
.A2(n_120),
.B1(n_117),
.B2(n_119),
.Y(n_4969)
);

INVx1_ASAP7_75t_L g4970 ( 
.A(n_4659),
.Y(n_4970)
);

O2A1O1Ixp33_ASAP7_75t_L g4971 ( 
.A1(n_4626),
.A2(n_124),
.B(n_121),
.C(n_123),
.Y(n_4971)
);

AOI21xp5_ASAP7_75t_L g4972 ( 
.A1(n_4734),
.A2(n_4718),
.B(n_4525),
.Y(n_4972)
);

NAND2xp5_ASAP7_75t_L g4973 ( 
.A(n_4831),
.B(n_4600),
.Y(n_4973)
);

NAND2xp5_ASAP7_75t_SL g4974 ( 
.A(n_4776),
.B(n_4692),
.Y(n_4974)
);

INVx1_ASAP7_75t_L g4975 ( 
.A(n_4841),
.Y(n_4975)
);

AND2x2_ASAP7_75t_L g4976 ( 
.A(n_4845),
.B(n_4570),
.Y(n_4976)
);

AOI21xp5_ASAP7_75t_L g4977 ( 
.A1(n_4872),
.A2(n_4686),
.B(n_4695),
.Y(n_4977)
);

AOI21xp5_ASAP7_75t_L g4978 ( 
.A1(n_4752),
.A2(n_4553),
.B(n_4717),
.Y(n_4978)
);

NAND2xp5_ASAP7_75t_L g4979 ( 
.A(n_4749),
.B(n_4614),
.Y(n_4979)
);

AND2x2_ASAP7_75t_L g4980 ( 
.A(n_4875),
.B(n_4613),
.Y(n_4980)
);

O2A1O1Ixp33_ASAP7_75t_L g4981 ( 
.A1(n_4901),
.A2(n_4714),
.B(n_4593),
.C(n_4694),
.Y(n_4981)
);

OAI22xp5_ASAP7_75t_L g4982 ( 
.A1(n_4786),
.A2(n_4733),
.B1(n_4662),
.B2(n_4729),
.Y(n_4982)
);

AOI222xp33_ASAP7_75t_L g4983 ( 
.A1(n_4943),
.A2(n_4728),
.B1(n_4450),
.B2(n_4602),
.C1(n_4623),
.C2(n_4567),
.Y(n_4983)
);

AND2x4_ASAP7_75t_L g4984 ( 
.A(n_4876),
.B(n_4493),
.Y(n_4984)
);

INVx1_ASAP7_75t_L g4985 ( 
.A(n_4798),
.Y(n_4985)
);

INVx2_ASAP7_75t_L g4986 ( 
.A(n_4796),
.Y(n_4986)
);

INVx1_ASAP7_75t_L g4987 ( 
.A(n_4802),
.Y(n_4987)
);

NAND2xp5_ASAP7_75t_L g4988 ( 
.A(n_4780),
.B(n_4692),
.Y(n_4988)
);

AO21x2_ASAP7_75t_L g4989 ( 
.A1(n_4753),
.A2(n_4599),
.B(n_4725),
.Y(n_4989)
);

BUFx3_ASAP7_75t_L g4990 ( 
.A(n_4961),
.Y(n_4990)
);

BUFx3_ASAP7_75t_L g4991 ( 
.A(n_4790),
.Y(n_4991)
);

AOI21xp5_ASAP7_75t_L g4992 ( 
.A1(n_4801),
.A2(n_4723),
.B(n_4545),
.Y(n_4992)
);

AND2x2_ASAP7_75t_L g4993 ( 
.A(n_4826),
.B(n_4522),
.Y(n_4993)
);

INVx1_ASAP7_75t_L g4994 ( 
.A(n_4820),
.Y(n_4994)
);

NAND2xp5_ASAP7_75t_L g4995 ( 
.A(n_4748),
.B(n_4877),
.Y(n_4995)
);

OR2x2_ASAP7_75t_L g4996 ( 
.A(n_4854),
.B(n_4535),
.Y(n_4996)
);

AOI21xp5_ASAP7_75t_L g4997 ( 
.A1(n_4757),
.A2(n_4723),
.B(n_4617),
.Y(n_4997)
);

NAND2xp5_ASAP7_75t_L g4998 ( 
.A(n_4894),
.B(n_4576),
.Y(n_4998)
);

O2A1O1Ixp33_ASAP7_75t_L g4999 ( 
.A1(n_4889),
.A2(n_4521),
.B(n_4492),
.C(n_4578),
.Y(n_4999)
);

INVx3_ASAP7_75t_SL g5000 ( 
.A(n_4766),
.Y(n_5000)
);

A2O1A1Ixp33_ASAP7_75t_L g5001 ( 
.A1(n_4959),
.A2(n_4619),
.B(n_4708),
.C(n_4487),
.Y(n_5001)
);

AND2x4_ASAP7_75t_L g5002 ( 
.A(n_4742),
.B(n_4615),
.Y(n_5002)
);

INVx2_ASAP7_75t_L g5003 ( 
.A(n_4827),
.Y(n_5003)
);

INVx2_ASAP7_75t_L g5004 ( 
.A(n_4847),
.Y(n_5004)
);

INVx2_ASAP7_75t_L g5005 ( 
.A(n_4760),
.Y(n_5005)
);

INVx1_ASAP7_75t_L g5006 ( 
.A(n_4864),
.Y(n_5006)
);

NAND2xp5_ASAP7_75t_SL g5007 ( 
.A(n_4972),
.B(n_4708),
.Y(n_5007)
);

INVx1_ASAP7_75t_L g5008 ( 
.A(n_4852),
.Y(n_5008)
);

BUFx2_ASAP7_75t_L g5009 ( 
.A(n_4777),
.Y(n_5009)
);

OR2x2_ASAP7_75t_L g5010 ( 
.A(n_4741),
.B(n_4587),
.Y(n_5010)
);

NAND2xp5_ASAP7_75t_L g5011 ( 
.A(n_4782),
.B(n_4728),
.Y(n_5011)
);

NOR2x1_ASAP7_75t_SL g5012 ( 
.A(n_4828),
.B(n_4511),
.Y(n_5012)
);

INVx2_ASAP7_75t_L g5013 ( 
.A(n_4883),
.Y(n_5013)
);

NOR2xp67_ASAP7_75t_L g5014 ( 
.A(n_4960),
.B(n_4649),
.Y(n_5014)
);

AND2x2_ASAP7_75t_L g5015 ( 
.A(n_4823),
.B(n_4604),
.Y(n_5015)
);

NAND2xp5_ASAP7_75t_L g5016 ( 
.A(n_4755),
.B(n_4728),
.Y(n_5016)
);

INVx2_ASAP7_75t_L g5017 ( 
.A(n_4885),
.Y(n_5017)
);

INVx3_ASAP7_75t_L g5018 ( 
.A(n_4813),
.Y(n_5018)
);

NAND2xp5_ASAP7_75t_L g5019 ( 
.A(n_4926),
.B(n_4538),
.Y(n_5019)
);

OR2x6_ASAP7_75t_L g5020 ( 
.A(n_4948),
.B(n_4664),
.Y(n_5020)
);

BUFx2_ASAP7_75t_L g5021 ( 
.A(n_4947),
.Y(n_5021)
);

OAI21x1_ASAP7_75t_SL g5022 ( 
.A1(n_4963),
.A2(n_4657),
.B(n_4551),
.Y(n_5022)
);

INVx3_ASAP7_75t_SL g5023 ( 
.A(n_4834),
.Y(n_5023)
);

OR2x6_ASAP7_75t_L g5024 ( 
.A(n_4965),
.B(n_4572),
.Y(n_5024)
);

INVx2_ASAP7_75t_SL g5025 ( 
.A(n_4960),
.Y(n_5025)
);

OR2x2_ASAP7_75t_L g5026 ( 
.A(n_4824),
.B(n_123),
.Y(n_5026)
);

NAND2xp5_ASAP7_75t_L g5027 ( 
.A(n_4762),
.B(n_124),
.Y(n_5027)
);

AOI21xp5_ASAP7_75t_SL g5028 ( 
.A1(n_4837),
.A2(n_125),
.B(n_126),
.Y(n_5028)
);

CKINVDCx5p33_ASAP7_75t_R g5029 ( 
.A(n_4836),
.Y(n_5029)
);

OAI21xp33_ASAP7_75t_L g5030 ( 
.A1(n_4922),
.A2(n_4952),
.B(n_4891),
.Y(n_5030)
);

BUFx6f_ASAP7_75t_SL g5031 ( 
.A(n_4899),
.Y(n_5031)
);

AND2x4_ASAP7_75t_L g5032 ( 
.A(n_4751),
.B(n_1399),
.Y(n_5032)
);

BUFx3_ASAP7_75t_L g5033 ( 
.A(n_4761),
.Y(n_5033)
);

O2A1O1Ixp5_ASAP7_75t_SL g5034 ( 
.A1(n_4970),
.A2(n_129),
.B(n_127),
.C(n_128),
.Y(n_5034)
);

AND2x2_ASAP7_75t_L g5035 ( 
.A(n_4860),
.B(n_127),
.Y(n_5035)
);

AOI21xp5_ASAP7_75t_L g5036 ( 
.A1(n_4791),
.A2(n_129),
.B(n_130),
.Y(n_5036)
);

CKINVDCx8_ASAP7_75t_R g5037 ( 
.A(n_4843),
.Y(n_5037)
);

INVx1_ASAP7_75t_SL g5038 ( 
.A(n_4833),
.Y(n_5038)
);

INVxp67_ASAP7_75t_L g5039 ( 
.A(n_4942),
.Y(n_5039)
);

NAND2xp5_ASAP7_75t_L g5040 ( 
.A(n_4873),
.B(n_130),
.Y(n_5040)
);

A2O1A1Ixp33_ASAP7_75t_SL g5041 ( 
.A1(n_4911),
.A2(n_133),
.B(n_131),
.C(n_132),
.Y(n_5041)
);

NOR2xp33_ASAP7_75t_L g5042 ( 
.A(n_4874),
.B(n_131),
.Y(n_5042)
);

NOR2xp33_ASAP7_75t_L g5043 ( 
.A(n_4844),
.B(n_132),
.Y(n_5043)
);

INVx1_ASAP7_75t_L g5044 ( 
.A(n_4793),
.Y(n_5044)
);

AND2x4_ASAP7_75t_L g5045 ( 
.A(n_4810),
.B(n_1401),
.Y(n_5045)
);

OR2x6_ASAP7_75t_L g5046 ( 
.A(n_4769),
.B(n_1402),
.Y(n_5046)
);

HB1xp67_ASAP7_75t_L g5047 ( 
.A(n_4955),
.Y(n_5047)
);

INVx1_ASAP7_75t_L g5048 ( 
.A(n_4896),
.Y(n_5048)
);

HB1xp67_ASAP7_75t_L g5049 ( 
.A(n_4763),
.Y(n_5049)
);

INVx2_ASAP7_75t_SL g5050 ( 
.A(n_4942),
.Y(n_5050)
);

HB1xp67_ASAP7_75t_L g5051 ( 
.A(n_4775),
.Y(n_5051)
);

NAND2xp5_ASAP7_75t_L g5052 ( 
.A(n_4745),
.B(n_133),
.Y(n_5052)
);

INVx3_ASAP7_75t_SL g5053 ( 
.A(n_4740),
.Y(n_5053)
);

INVx1_ASAP7_75t_L g5054 ( 
.A(n_4920),
.Y(n_5054)
);

AND2x4_ASAP7_75t_L g5055 ( 
.A(n_4862),
.B(n_1405),
.Y(n_5055)
);

INVx1_ASAP7_75t_L g5056 ( 
.A(n_4920),
.Y(n_5056)
);

INVx2_ASAP7_75t_L g5057 ( 
.A(n_4929),
.Y(n_5057)
);

AOI22xp33_ASAP7_75t_L g5058 ( 
.A1(n_4835),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_5058)
);

INVx1_ASAP7_75t_L g5059 ( 
.A(n_4789),
.Y(n_5059)
);

INVxp67_ASAP7_75t_L g5060 ( 
.A(n_4910),
.Y(n_5060)
);

INVx2_ASAP7_75t_L g5061 ( 
.A(n_4758),
.Y(n_5061)
);

NAND2xp5_ASAP7_75t_L g5062 ( 
.A(n_4812),
.B(n_136),
.Y(n_5062)
);

NAND2xp5_ASAP7_75t_L g5063 ( 
.A(n_4886),
.B(n_138),
.Y(n_5063)
);

NAND2x1p5_ASAP7_75t_L g5064 ( 
.A(n_4740),
.B(n_1406),
.Y(n_5064)
);

OAI21xp5_ASAP7_75t_L g5065 ( 
.A1(n_4953),
.A2(n_4764),
.B(n_4905),
.Y(n_5065)
);

NAND2xp5_ASAP7_75t_L g5066 ( 
.A(n_4881),
.B(n_139),
.Y(n_5066)
);

INVx1_ASAP7_75t_L g5067 ( 
.A(n_4938),
.Y(n_5067)
);

NOR2xp33_ASAP7_75t_L g5068 ( 
.A(n_4888),
.B(n_139),
.Y(n_5068)
);

OR2x6_ASAP7_75t_L g5069 ( 
.A(n_4744),
.B(n_4930),
.Y(n_5069)
);

NAND2x1p5_ASAP7_75t_L g5070 ( 
.A(n_4813),
.B(n_1407),
.Y(n_5070)
);

AOI22xp33_ASAP7_75t_SL g5071 ( 
.A1(n_4941),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.Y(n_5071)
);

AOI22xp33_ASAP7_75t_L g5072 ( 
.A1(n_4806),
.A2(n_143),
.B1(n_140),
.B2(n_141),
.Y(n_5072)
);

NOR2xp33_ASAP7_75t_L g5073 ( 
.A(n_4756),
.B(n_4767),
.Y(n_5073)
);

AND2x2_ASAP7_75t_L g5074 ( 
.A(n_4817),
.B(n_143),
.Y(n_5074)
);

NOR2xp33_ASAP7_75t_L g5075 ( 
.A(n_4768),
.B(n_144),
.Y(n_5075)
);

OR2x2_ASAP7_75t_L g5076 ( 
.A(n_4822),
.B(n_145),
.Y(n_5076)
);

NAND2xp5_ASAP7_75t_L g5077 ( 
.A(n_4897),
.B(n_145),
.Y(n_5077)
);

INVx1_ASAP7_75t_L g5078 ( 
.A(n_4840),
.Y(n_5078)
);

AOI21xp5_ASAP7_75t_L g5079 ( 
.A1(n_4803),
.A2(n_146),
.B(n_147),
.Y(n_5079)
);

CKINVDCx6p67_ASAP7_75t_R g5080 ( 
.A(n_4818),
.Y(n_5080)
);

INVx2_ASAP7_75t_SL g5081 ( 
.A(n_4794),
.Y(n_5081)
);

A2O1A1Ixp33_ASAP7_75t_L g5082 ( 
.A1(n_4971),
.A2(n_149),
.B(n_147),
.C(n_148),
.Y(n_5082)
);

NAND2xp5_ASAP7_75t_L g5083 ( 
.A(n_4916),
.B(n_148),
.Y(n_5083)
);

INVx1_ASAP7_75t_L g5084 ( 
.A(n_4758),
.Y(n_5084)
);

OR2x2_ASAP7_75t_L g5085 ( 
.A(n_4924),
.B(n_149),
.Y(n_5085)
);

A2O1A1Ixp33_ASAP7_75t_L g5086 ( 
.A1(n_4880),
.A2(n_152),
.B(n_150),
.C(n_151),
.Y(n_5086)
);

INVx1_ASAP7_75t_L g5087 ( 
.A(n_4870),
.Y(n_5087)
);

AOI21x1_ASAP7_75t_SL g5088 ( 
.A1(n_4819),
.A2(n_150),
.B(n_152),
.Y(n_5088)
);

INVx4_ASAP7_75t_L g5089 ( 
.A(n_4930),
.Y(n_5089)
);

OR2x2_ASAP7_75t_L g5090 ( 
.A(n_4912),
.B(n_155),
.Y(n_5090)
);

INVx1_ASAP7_75t_L g5091 ( 
.A(n_4746),
.Y(n_5091)
);

BUFx4_ASAP7_75t_SL g5092 ( 
.A(n_4739),
.Y(n_5092)
);

OR2x2_ASAP7_75t_L g5093 ( 
.A(n_4923),
.B(n_156),
.Y(n_5093)
);

HB1xp67_ASAP7_75t_L g5094 ( 
.A(n_4775),
.Y(n_5094)
);

AND2x2_ASAP7_75t_L g5095 ( 
.A(n_4850),
.B(n_156),
.Y(n_5095)
);

BUFx3_ASAP7_75t_L g5096 ( 
.A(n_4906),
.Y(n_5096)
);

BUFx3_ASAP7_75t_L g5097 ( 
.A(n_4772),
.Y(n_5097)
);

AND2x2_ASAP7_75t_L g5098 ( 
.A(n_4858),
.B(n_157),
.Y(n_5098)
);

INVx1_ASAP7_75t_L g5099 ( 
.A(n_4940),
.Y(n_5099)
);

BUFx5_ASAP7_75t_L g5100 ( 
.A(n_4759),
.Y(n_5100)
);

BUFx3_ASAP7_75t_L g5101 ( 
.A(n_4785),
.Y(n_5101)
);

CKINVDCx5p33_ASAP7_75t_R g5102 ( 
.A(n_4968),
.Y(n_5102)
);

NAND2xp5_ASAP7_75t_L g5103 ( 
.A(n_4903),
.B(n_158),
.Y(n_5103)
);

NAND2xp5_ASAP7_75t_L g5104 ( 
.A(n_4838),
.B(n_158),
.Y(n_5104)
);

INVx2_ASAP7_75t_SL g5105 ( 
.A(n_4773),
.Y(n_5105)
);

AOI21xp5_ASAP7_75t_L g5106 ( 
.A1(n_4964),
.A2(n_162),
.B(n_160),
.Y(n_5106)
);

BUFx12f_ASAP7_75t_L g5107 ( 
.A(n_4747),
.Y(n_5107)
);

AOI22xp5_ASAP7_75t_L g5108 ( 
.A1(n_4778),
.A2(n_164),
.B1(n_159),
.B2(n_163),
.Y(n_5108)
);

INVx1_ASAP7_75t_L g5109 ( 
.A(n_4816),
.Y(n_5109)
);

AND2x4_ASAP7_75t_L g5110 ( 
.A(n_4884),
.B(n_1408),
.Y(n_5110)
);

INVx1_ASAP7_75t_L g5111 ( 
.A(n_4933),
.Y(n_5111)
);

AOI21xp33_ASAP7_75t_SL g5112 ( 
.A1(n_4928),
.A2(n_4969),
.B(n_4944),
.Y(n_5112)
);

AOI21xp5_ASAP7_75t_L g5113 ( 
.A1(n_4887),
.A2(n_164),
.B(n_163),
.Y(n_5113)
);

INVx1_ASAP7_75t_L g5114 ( 
.A(n_4921),
.Y(n_5114)
);

INVx1_ASAP7_75t_SL g5115 ( 
.A(n_4781),
.Y(n_5115)
);

OAI22xp5_ASAP7_75t_L g5116 ( 
.A1(n_4811),
.A2(n_166),
.B1(n_159),
.B2(n_165),
.Y(n_5116)
);

OAI22xp5_ASAP7_75t_L g5117 ( 
.A1(n_4815),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.Y(n_5117)
);

NAND2x1p5_ASAP7_75t_L g5118 ( 
.A(n_4799),
.B(n_1409),
.Y(n_5118)
);

NAND2xp5_ASAP7_75t_L g5119 ( 
.A(n_4890),
.B(n_169),
.Y(n_5119)
);

NAND2xp5_ASAP7_75t_L g5120 ( 
.A(n_4967),
.B(n_169),
.Y(n_5120)
);

CKINVDCx11_ASAP7_75t_R g5121 ( 
.A(n_4856),
.Y(n_5121)
);

INVx1_ASAP7_75t_L g5122 ( 
.A(n_4946),
.Y(n_5122)
);

NAND3xp33_ASAP7_75t_L g5123 ( 
.A(n_4848),
.B(n_170),
.C(n_171),
.Y(n_5123)
);

AND2x2_ASAP7_75t_L g5124 ( 
.A(n_4949),
.B(n_170),
.Y(n_5124)
);

NAND2xp5_ASAP7_75t_L g5125 ( 
.A(n_4951),
.B(n_172),
.Y(n_5125)
);

AOI222xp33_ASAP7_75t_L g5126 ( 
.A1(n_4797),
.A2(n_174),
.B1(n_176),
.B2(n_172),
.C1(n_173),
.C2(n_175),
.Y(n_5126)
);

OR2x2_ASAP7_75t_L g5127 ( 
.A(n_4932),
.B(n_174),
.Y(n_5127)
);

BUFx6f_ASAP7_75t_L g5128 ( 
.A(n_4954),
.Y(n_5128)
);

OR2x6_ASAP7_75t_L g5129 ( 
.A(n_4914),
.B(n_1410),
.Y(n_5129)
);

INVx2_ASAP7_75t_L g5130 ( 
.A(n_4937),
.Y(n_5130)
);

NAND2xp5_ASAP7_75t_L g5131 ( 
.A(n_4962),
.B(n_176),
.Y(n_5131)
);

A2O1A1Ixp33_ASAP7_75t_SL g5132 ( 
.A1(n_4908),
.A2(n_179),
.B(n_177),
.C(n_178),
.Y(n_5132)
);

AND2x2_ASAP7_75t_L g5133 ( 
.A(n_4792),
.B(n_177),
.Y(n_5133)
);

NOR2xp33_ASAP7_75t_L g5134 ( 
.A(n_4770),
.B(n_180),
.Y(n_5134)
);

AOI22xp33_ASAP7_75t_L g5135 ( 
.A1(n_4893),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.Y(n_5135)
);

HB1xp67_ASAP7_75t_SL g5136 ( 
.A(n_4861),
.Y(n_5136)
);

OAI22xp5_ASAP7_75t_L g5137 ( 
.A1(n_5136),
.A2(n_4918),
.B1(n_4934),
.B2(n_4900),
.Y(n_5137)
);

BUFx6f_ASAP7_75t_L g5138 ( 
.A(n_4990),
.Y(n_5138)
);

OR2x2_ASAP7_75t_L g5139 ( 
.A(n_4975),
.B(n_4937),
.Y(n_5139)
);

NAND2xp5_ASAP7_75t_L g5140 ( 
.A(n_4995),
.B(n_4879),
.Y(n_5140)
);

NAND2xp5_ASAP7_75t_L g5141 ( 
.A(n_5059),
.B(n_4915),
.Y(n_5141)
);

NAND2xp5_ASAP7_75t_L g5142 ( 
.A(n_5067),
.B(n_4754),
.Y(n_5142)
);

HB1xp67_ASAP7_75t_L g5143 ( 
.A(n_5021),
.Y(n_5143)
);

BUFx3_ASAP7_75t_L g5144 ( 
.A(n_4991),
.Y(n_5144)
);

INVx1_ASAP7_75t_L g5145 ( 
.A(n_4985),
.Y(n_5145)
);

AND2x2_ASAP7_75t_L g5146 ( 
.A(n_4980),
.B(n_4945),
.Y(n_5146)
);

A2O1A1Ixp33_ASAP7_75t_SL g5147 ( 
.A1(n_5134),
.A2(n_4779),
.B(n_4832),
.C(n_4821),
.Y(n_5147)
);

OAI22xp5_ASAP7_75t_L g5148 ( 
.A1(n_5071),
.A2(n_4851),
.B1(n_4868),
.B2(n_4842),
.Y(n_5148)
);

AND2x4_ASAP7_75t_L g5149 ( 
.A(n_4993),
.B(n_4984),
.Y(n_5149)
);

AND2x2_ASAP7_75t_L g5150 ( 
.A(n_4976),
.B(n_4945),
.Y(n_5150)
);

AND2x4_ASAP7_75t_L g5151 ( 
.A(n_5038),
.B(n_4966),
.Y(n_5151)
);

A2O1A1Ixp33_ASAP7_75t_L g5152 ( 
.A1(n_4977),
.A2(n_4807),
.B(n_4804),
.C(n_4795),
.Y(n_5152)
);

AND2x4_ASAP7_75t_L g5153 ( 
.A(n_5033),
.B(n_4800),
.Y(n_5153)
);

A2O1A1Ixp33_ASAP7_75t_L g5154 ( 
.A1(n_4978),
.A2(n_4865),
.B(n_4765),
.C(n_4857),
.Y(n_5154)
);

NAND2xp5_ASAP7_75t_L g5155 ( 
.A(n_4987),
.B(n_4892),
.Y(n_5155)
);

A2O1A1Ixp33_ASAP7_75t_L g5156 ( 
.A1(n_5030),
.A2(n_4859),
.B(n_4855),
.C(n_4867),
.Y(n_5156)
);

AND2x2_ASAP7_75t_L g5157 ( 
.A(n_5015),
.B(n_4936),
.Y(n_5157)
);

AND2x2_ASAP7_75t_L g5158 ( 
.A(n_4979),
.B(n_4936),
.Y(n_5158)
);

NAND2xp5_ASAP7_75t_L g5159 ( 
.A(n_5006),
.B(n_4853),
.Y(n_5159)
);

NOR2xp33_ASAP7_75t_L g5160 ( 
.A(n_5000),
.B(n_181),
.Y(n_5160)
);

NAND2xp5_ASAP7_75t_L g5161 ( 
.A(n_5044),
.B(n_183),
.Y(n_5161)
);

A2O1A1Ixp33_ASAP7_75t_L g5162 ( 
.A1(n_5112),
.A2(n_4869),
.B(n_4866),
.C(n_4774),
.Y(n_5162)
);

INVx1_ASAP7_75t_SL g5163 ( 
.A(n_5053),
.Y(n_5163)
);

AOI22xp5_ASAP7_75t_L g5164 ( 
.A1(n_4982),
.A2(n_4902),
.B1(n_4904),
.B2(n_4898),
.Y(n_5164)
);

AND2x2_ASAP7_75t_L g5165 ( 
.A(n_5002),
.B(n_4771),
.Y(n_5165)
);

NOR2xp67_ASAP7_75t_L g5166 ( 
.A(n_5025),
.B(n_4784),
.Y(n_5166)
);

AND2x4_ASAP7_75t_L g5167 ( 
.A(n_4973),
.B(n_4800),
.Y(n_5167)
);

AND2x2_ASAP7_75t_L g5168 ( 
.A(n_5097),
.B(n_4958),
.Y(n_5168)
);

INVx2_ASAP7_75t_L g5169 ( 
.A(n_5013),
.Y(n_5169)
);

INVxp67_ASAP7_75t_L g5170 ( 
.A(n_4998),
.Y(n_5170)
);

NOR2xp33_ASAP7_75t_L g5171 ( 
.A(n_5023),
.B(n_184),
.Y(n_5171)
);

O2A1O1Ixp33_ASAP7_75t_L g5172 ( 
.A1(n_5082),
.A2(n_4788),
.B(n_4787),
.C(n_4913),
.Y(n_5172)
);

NAND2xp5_ASAP7_75t_L g5173 ( 
.A(n_5111),
.B(n_184),
.Y(n_5173)
);

NAND2xp5_ASAP7_75t_SL g5174 ( 
.A(n_4983),
.B(n_5016),
.Y(n_5174)
);

NOR2xp33_ASAP7_75t_SL g5175 ( 
.A(n_5089),
.B(n_4849),
.Y(n_5175)
);

OR2x6_ASAP7_75t_L g5176 ( 
.A(n_5020),
.B(n_4957),
.Y(n_5176)
);

AOI22xp5_ASAP7_75t_L g5177 ( 
.A1(n_5068),
.A2(n_4909),
.B1(n_4950),
.B2(n_4805),
.Y(n_5177)
);

AND2x4_ASAP7_75t_L g5178 ( 
.A(n_5101),
.B(n_4809),
.Y(n_5178)
);

INVx1_ASAP7_75t_SL g5179 ( 
.A(n_5107),
.Y(n_5179)
);

AO22x2_ASAP7_75t_L g5180 ( 
.A1(n_5054),
.A2(n_4809),
.B1(n_4907),
.B2(n_4895),
.Y(n_5180)
);

O2A1O1Ixp5_ASAP7_75t_L g5181 ( 
.A1(n_5036),
.A2(n_4939),
.B(n_194),
.C(n_202),
.Y(n_5181)
);

NAND2xp5_ASAP7_75t_L g5182 ( 
.A(n_5114),
.B(n_185),
.Y(n_5182)
);

AND2x2_ASAP7_75t_L g5183 ( 
.A(n_4996),
.B(n_4783),
.Y(n_5183)
);

NAND2xp5_ASAP7_75t_L g5184 ( 
.A(n_5099),
.B(n_186),
.Y(n_5184)
);

INVxp67_ASAP7_75t_L g5185 ( 
.A(n_5128),
.Y(n_5185)
);

INVx1_ASAP7_75t_L g5186 ( 
.A(n_5048),
.Y(n_5186)
);

INVx1_ASAP7_75t_L g5187 ( 
.A(n_5017),
.Y(n_5187)
);

INVx1_ASAP7_75t_L g5188 ( 
.A(n_4986),
.Y(n_5188)
);

NAND2xp5_ASAP7_75t_L g5189 ( 
.A(n_5087),
.B(n_186),
.Y(n_5189)
);

OR2x6_ASAP7_75t_SL g5190 ( 
.A(n_5029),
.B(n_4895),
.Y(n_5190)
);

INVx2_ASAP7_75t_L g5191 ( 
.A(n_5003),
.Y(n_5191)
);

OR2x2_ASAP7_75t_L g5192 ( 
.A(n_5078),
.B(n_5010),
.Y(n_5192)
);

AND2x2_ASAP7_75t_L g5193 ( 
.A(n_5019),
.B(n_4808),
.Y(n_5193)
);

CKINVDCx9p33_ASAP7_75t_R g5194 ( 
.A(n_5009),
.Y(n_5194)
);

INVx1_ASAP7_75t_L g5195 ( 
.A(n_5004),
.Y(n_5195)
);

INVx3_ASAP7_75t_L g5196 ( 
.A(n_5018),
.Y(n_5196)
);

INVxp67_ASAP7_75t_L g5197 ( 
.A(n_5128),
.Y(n_5197)
);

NOR2xp33_ASAP7_75t_SL g5198 ( 
.A(n_5037),
.B(n_4907),
.Y(n_5198)
);

O2A1O1Ixp33_ASAP7_75t_L g5199 ( 
.A1(n_5041),
.A2(n_189),
.B(n_187),
.C(n_188),
.Y(n_5199)
);

O2A1O1Ixp33_ASAP7_75t_L g5200 ( 
.A1(n_5065),
.A2(n_191),
.B(n_188),
.C(n_189),
.Y(n_5200)
);

INVx1_ASAP7_75t_L g5201 ( 
.A(n_5005),
.Y(n_5201)
);

AND2x4_ASAP7_75t_L g5202 ( 
.A(n_5020),
.B(n_4927),
.Y(n_5202)
);

INVxp67_ASAP7_75t_L g5203 ( 
.A(n_5122),
.Y(n_5203)
);

INVx1_ASAP7_75t_L g5204 ( 
.A(n_4994),
.Y(n_5204)
);

AND2x2_ASAP7_75t_L g5205 ( 
.A(n_5035),
.B(n_5074),
.Y(n_5205)
);

AND2x4_ASAP7_75t_L g5206 ( 
.A(n_5069),
.B(n_4927),
.Y(n_5206)
);

BUFx3_ASAP7_75t_L g5207 ( 
.A(n_5096),
.Y(n_5207)
);

OAI22xp5_ASAP7_75t_L g5208 ( 
.A1(n_5135),
.A2(n_5123),
.B1(n_5058),
.B2(n_5120),
.Y(n_5208)
);

AND2x4_ASAP7_75t_L g5209 ( 
.A(n_5069),
.B(n_4743),
.Y(n_5209)
);

O2A1O1Ixp33_ASAP7_75t_L g5210 ( 
.A1(n_5086),
.A2(n_193),
.B(n_191),
.C(n_192),
.Y(n_5210)
);

OR2x2_ASAP7_75t_L g5211 ( 
.A(n_4988),
.B(n_4750),
.Y(n_5211)
);

OR2x2_ASAP7_75t_L g5212 ( 
.A(n_5026),
.B(n_193),
.Y(n_5212)
);

A2O1A1Ixp33_ASAP7_75t_L g5213 ( 
.A1(n_4981),
.A2(n_4825),
.B(n_4830),
.C(n_4829),
.Y(n_5213)
);

OAI21x1_ASAP7_75t_SL g5214 ( 
.A1(n_5022),
.A2(n_5012),
.B(n_5091),
.Y(n_5214)
);

INVx1_ASAP7_75t_L g5215 ( 
.A(n_5008),
.Y(n_5215)
);

NAND2xp5_ASAP7_75t_L g5216 ( 
.A(n_5109),
.B(n_195),
.Y(n_5216)
);

AND2x2_ASAP7_75t_L g5217 ( 
.A(n_5095),
.B(n_4814),
.Y(n_5217)
);

NAND2x1p5_ASAP7_75t_L g5218 ( 
.A(n_5014),
.B(n_4839),
.Y(n_5218)
);

NOR2xp33_ASAP7_75t_L g5219 ( 
.A(n_5043),
.B(n_196),
.Y(n_5219)
);

AOI21xp5_ASAP7_75t_L g5220 ( 
.A1(n_5051),
.A2(n_4956),
.B(n_4871),
.Y(n_5220)
);

AND2x2_ASAP7_75t_L g5221 ( 
.A(n_5098),
.B(n_4846),
.Y(n_5221)
);

NAND2xp5_ASAP7_75t_L g5222 ( 
.A(n_5062),
.B(n_197),
.Y(n_5222)
);

NAND2xp5_ASAP7_75t_L g5223 ( 
.A(n_5040),
.B(n_197),
.Y(n_5223)
);

O2A1O1Ixp33_ASAP7_75t_SL g5224 ( 
.A1(n_5052),
.A2(n_200),
.B(n_198),
.C(n_199),
.Y(n_5224)
);

HB1xp67_ASAP7_75t_L g5225 ( 
.A(n_5047),
.Y(n_5225)
);

OA22x2_ASAP7_75t_L g5226 ( 
.A1(n_5007),
.A2(n_4878),
.B1(n_4863),
.B2(n_4882),
.Y(n_5226)
);

INVx1_ASAP7_75t_L g5227 ( 
.A(n_5084),
.Y(n_5227)
);

INVx2_ASAP7_75t_L g5228 ( 
.A(n_5056),
.Y(n_5228)
);

AOI21xp5_ASAP7_75t_L g5229 ( 
.A1(n_5094),
.A2(n_4919),
.B(n_4917),
.Y(n_5229)
);

INVx2_ASAP7_75t_L g5230 ( 
.A(n_5057),
.Y(n_5230)
);

INVx1_ASAP7_75t_L g5231 ( 
.A(n_5011),
.Y(n_5231)
);

HB1xp67_ASAP7_75t_L g5232 ( 
.A(n_5049),
.Y(n_5232)
);

NAND2xp5_ASAP7_75t_L g5233 ( 
.A(n_5027),
.B(n_201),
.Y(n_5233)
);

AOI21xp5_ASAP7_75t_SL g5234 ( 
.A1(n_5129),
.A2(n_4931),
.B(n_4925),
.Y(n_5234)
);

A2O1A1Ixp33_ASAP7_75t_L g5235 ( 
.A1(n_4992),
.A2(n_4935),
.B(n_203),
.C(n_201),
.Y(n_5235)
);

O2A1O1Ixp33_ASAP7_75t_L g5236 ( 
.A1(n_5116),
.A2(n_204),
.B(n_202),
.C(n_203),
.Y(n_5236)
);

INVx1_ASAP7_75t_L g5237 ( 
.A(n_5061),
.Y(n_5237)
);

INVx2_ASAP7_75t_L g5238 ( 
.A(n_5130),
.Y(n_5238)
);

OR2x2_ASAP7_75t_L g5239 ( 
.A(n_5076),
.B(n_5085),
.Y(n_5239)
);

BUFx2_ASAP7_75t_SL g5240 ( 
.A(n_5031),
.Y(n_5240)
);

CKINVDCx20_ASAP7_75t_R g5241 ( 
.A(n_5080),
.Y(n_5241)
);

INVx2_ASAP7_75t_L g5242 ( 
.A(n_5100),
.Y(n_5242)
);

AOI21xp5_ASAP7_75t_L g5243 ( 
.A1(n_4974),
.A2(n_204),
.B(n_206),
.Y(n_5243)
);

INVx1_ASAP7_75t_L g5244 ( 
.A(n_5103),
.Y(n_5244)
);

NOR2xp67_ASAP7_75t_L g5245 ( 
.A(n_5105),
.B(n_206),
.Y(n_5245)
);

AOI21xp5_ASAP7_75t_L g5246 ( 
.A1(n_5106),
.A2(n_207),
.B(n_208),
.Y(n_5246)
);

INVx1_ASAP7_75t_L g5247 ( 
.A(n_5060),
.Y(n_5247)
);

BUFx3_ASAP7_75t_L g5248 ( 
.A(n_5102),
.Y(n_5248)
);

INVx2_ASAP7_75t_L g5249 ( 
.A(n_5100),
.Y(n_5249)
);

AND2x2_ASAP7_75t_L g5250 ( 
.A(n_5039),
.B(n_208),
.Y(n_5250)
);

NAND2xp5_ASAP7_75t_L g5251 ( 
.A(n_5063),
.B(n_210),
.Y(n_5251)
);

INVx2_ASAP7_75t_L g5252 ( 
.A(n_5100),
.Y(n_5252)
);

AND2x2_ASAP7_75t_L g5253 ( 
.A(n_5124),
.B(n_211),
.Y(n_5253)
);

AOI21xp5_ASAP7_75t_L g5254 ( 
.A1(n_5113),
.A2(n_211),
.B(n_212),
.Y(n_5254)
);

AND2x4_ASAP7_75t_L g5255 ( 
.A(n_5081),
.B(n_5050),
.Y(n_5255)
);

NAND2xp5_ASAP7_75t_L g5256 ( 
.A(n_5077),
.B(n_212),
.Y(n_5256)
);

OA21x2_ASAP7_75t_L g5257 ( 
.A1(n_4997),
.A2(n_213),
.B(n_215),
.Y(n_5257)
);

AND2x2_ASAP7_75t_L g5258 ( 
.A(n_5042),
.B(n_216),
.Y(n_5258)
);

BUFx3_ASAP7_75t_L g5259 ( 
.A(n_5073),
.Y(n_5259)
);

NAND2xp5_ASAP7_75t_L g5260 ( 
.A(n_5066),
.B(n_216),
.Y(n_5260)
);

INVx1_ASAP7_75t_L g5261 ( 
.A(n_5125),
.Y(n_5261)
);

AND2x2_ASAP7_75t_L g5262 ( 
.A(n_5093),
.B(n_217),
.Y(n_5262)
);

AND2x2_ASAP7_75t_L g5263 ( 
.A(n_5104),
.B(n_5090),
.Y(n_5263)
);

O2A1O1Ixp33_ASAP7_75t_L g5264 ( 
.A1(n_5117),
.A2(n_219),
.B(n_217),
.C(n_218),
.Y(n_5264)
);

A2O1A1Ixp33_ASAP7_75t_L g5265 ( 
.A1(n_5001),
.A2(n_221),
.B(n_219),
.C(n_220),
.Y(n_5265)
);

A2O1A1Ixp33_ASAP7_75t_L g5266 ( 
.A1(n_5079),
.A2(n_223),
.B(n_221),
.C(n_222),
.Y(n_5266)
);

INVx1_ASAP7_75t_L g5267 ( 
.A(n_5131),
.Y(n_5267)
);

OR2x2_ASAP7_75t_L g5268 ( 
.A(n_5127),
.B(n_222),
.Y(n_5268)
);

NOR2xp67_ASAP7_75t_L g5269 ( 
.A(n_5119),
.B(n_224),
.Y(n_5269)
);

NOR2xp33_ASAP7_75t_L g5270 ( 
.A(n_5121),
.B(n_224),
.Y(n_5270)
);

NOR2xp67_ASAP7_75t_L g5271 ( 
.A(n_5083),
.B(n_225),
.Y(n_5271)
);

NAND2xp5_ASAP7_75t_L g5272 ( 
.A(n_5115),
.B(n_225),
.Y(n_5272)
);

OAI22xp5_ASAP7_75t_L g5273 ( 
.A1(n_5072),
.A2(n_229),
.B1(n_226),
.B2(n_227),
.Y(n_5273)
);

AND2x2_ASAP7_75t_L g5274 ( 
.A(n_5133),
.B(n_226),
.Y(n_5274)
);

NAND2xp5_ASAP7_75t_L g5275 ( 
.A(n_5075),
.B(n_227),
.Y(n_5275)
);

AND2x2_ASAP7_75t_L g5276 ( 
.A(n_5024),
.B(n_5045),
.Y(n_5276)
);

BUFx5_ASAP7_75t_L g5277 ( 
.A(n_5100),
.Y(n_5277)
);

INVx2_ASAP7_75t_L g5278 ( 
.A(n_4989),
.Y(n_5278)
);

INVx1_ASAP7_75t_L g5279 ( 
.A(n_4999),
.Y(n_5279)
);

INVx2_ASAP7_75t_L g5280 ( 
.A(n_5129),
.Y(n_5280)
);

INVx3_ASAP7_75t_L g5281 ( 
.A(n_5055),
.Y(n_5281)
);

INVx1_ASAP7_75t_SL g5282 ( 
.A(n_5092),
.Y(n_5282)
);

HB1xp67_ASAP7_75t_L g5283 ( 
.A(n_5024),
.Y(n_5283)
);

AOI21xp5_ASAP7_75t_L g5284 ( 
.A1(n_5028),
.A2(n_229),
.B(n_230),
.Y(n_5284)
);

INVx3_ASAP7_75t_L g5285 ( 
.A(n_5138),
.Y(n_5285)
);

BUFx2_ASAP7_75t_L g5286 ( 
.A(n_5143),
.Y(n_5286)
);

BUFx6f_ASAP7_75t_L g5287 ( 
.A(n_5138),
.Y(n_5287)
);

INVx1_ASAP7_75t_L g5288 ( 
.A(n_5145),
.Y(n_5288)
);

INVx1_ASAP7_75t_L g5289 ( 
.A(n_5186),
.Y(n_5289)
);

OAI22xp5_ASAP7_75t_L g5290 ( 
.A1(n_5162),
.A2(n_5046),
.B1(n_5108),
.B2(n_5118),
.Y(n_5290)
);

NAND2xp5_ASAP7_75t_L g5291 ( 
.A(n_5203),
.B(n_5132),
.Y(n_5291)
);

INVx2_ASAP7_75t_L g5292 ( 
.A(n_5169),
.Y(n_5292)
);

OA21x2_ASAP7_75t_L g5293 ( 
.A1(n_5231),
.A2(n_5110),
.B(n_5032),
.Y(n_5293)
);

INVx2_ASAP7_75t_L g5294 ( 
.A(n_5191),
.Y(n_5294)
);

INVx1_ASAP7_75t_L g5295 ( 
.A(n_5187),
.Y(n_5295)
);

HB1xp67_ASAP7_75t_L g5296 ( 
.A(n_5225),
.Y(n_5296)
);

HB1xp67_ASAP7_75t_L g5297 ( 
.A(n_5232),
.Y(n_5297)
);

INVx2_ASAP7_75t_L g5298 ( 
.A(n_5188),
.Y(n_5298)
);

INVx2_ASAP7_75t_L g5299 ( 
.A(n_5195),
.Y(n_5299)
);

HB1xp67_ASAP7_75t_L g5300 ( 
.A(n_5170),
.Y(n_5300)
);

INVx2_ASAP7_75t_L g5301 ( 
.A(n_5201),
.Y(n_5301)
);

INVx2_ASAP7_75t_L g5302 ( 
.A(n_5192),
.Y(n_5302)
);

NAND2xp5_ASAP7_75t_L g5303 ( 
.A(n_5261),
.B(n_5126),
.Y(n_5303)
);

INVx2_ASAP7_75t_L g5304 ( 
.A(n_5228),
.Y(n_5304)
);

AND2x2_ASAP7_75t_L g5305 ( 
.A(n_5149),
.B(n_5046),
.Y(n_5305)
);

OAI21x1_ASAP7_75t_L g5306 ( 
.A1(n_5220),
.A2(n_5088),
.B(n_5034),
.Y(n_5306)
);

INVx1_ASAP7_75t_L g5307 ( 
.A(n_5227),
.Y(n_5307)
);

INVx1_ASAP7_75t_L g5308 ( 
.A(n_5204),
.Y(n_5308)
);

OAI221xp5_ASAP7_75t_L g5309 ( 
.A1(n_5265),
.A2(n_5064),
.B1(n_5070),
.B2(n_233),
.C(n_231),
.Y(n_5309)
);

INVx1_ASAP7_75t_L g5310 ( 
.A(n_5215),
.Y(n_5310)
);

INVx1_ASAP7_75t_SL g5311 ( 
.A(n_5194),
.Y(n_5311)
);

AOI21xp5_ASAP7_75t_L g5312 ( 
.A1(n_5213),
.A2(n_232),
.B(n_233),
.Y(n_5312)
);

INVx1_ASAP7_75t_L g5313 ( 
.A(n_5139),
.Y(n_5313)
);

INVx2_ASAP7_75t_L g5314 ( 
.A(n_5238),
.Y(n_5314)
);

OR2x2_ASAP7_75t_L g5315 ( 
.A(n_5239),
.B(n_232),
.Y(n_5315)
);

INVx2_ASAP7_75t_L g5316 ( 
.A(n_5230),
.Y(n_5316)
);

INVx1_ASAP7_75t_L g5317 ( 
.A(n_5155),
.Y(n_5317)
);

INVx1_ASAP7_75t_L g5318 ( 
.A(n_5247),
.Y(n_5318)
);

INVx2_ASAP7_75t_L g5319 ( 
.A(n_5237),
.Y(n_5319)
);

NAND2xp5_ASAP7_75t_SL g5320 ( 
.A(n_5259),
.B(n_234),
.Y(n_5320)
);

INVx1_ASAP7_75t_L g5321 ( 
.A(n_5159),
.Y(n_5321)
);

AND2x2_ASAP7_75t_L g5322 ( 
.A(n_5150),
.B(n_234),
.Y(n_5322)
);

INVx1_ASAP7_75t_L g5323 ( 
.A(n_5141),
.Y(n_5323)
);

INVx1_ASAP7_75t_L g5324 ( 
.A(n_5161),
.Y(n_5324)
);

INVxp33_ASAP7_75t_L g5325 ( 
.A(n_5270),
.Y(n_5325)
);

INVx1_ASAP7_75t_L g5326 ( 
.A(n_5167),
.Y(n_5326)
);

INVx2_ASAP7_75t_L g5327 ( 
.A(n_5278),
.Y(n_5327)
);

AND2x2_ASAP7_75t_L g5328 ( 
.A(n_5205),
.B(n_235),
.Y(n_5328)
);

AND2x2_ASAP7_75t_L g5329 ( 
.A(n_5263),
.B(n_235),
.Y(n_5329)
);

INVx3_ASAP7_75t_L g5330 ( 
.A(n_5255),
.Y(n_5330)
);

INVx2_ASAP7_75t_L g5331 ( 
.A(n_5211),
.Y(n_5331)
);

INVx2_ASAP7_75t_L g5332 ( 
.A(n_5146),
.Y(n_5332)
);

NAND2xp5_ASAP7_75t_L g5333 ( 
.A(n_5267),
.B(n_236),
.Y(n_5333)
);

INVx2_ASAP7_75t_L g5334 ( 
.A(n_5157),
.Y(n_5334)
);

INVx1_ASAP7_75t_L g5335 ( 
.A(n_5158),
.Y(n_5335)
);

OAI21x1_ASAP7_75t_L g5336 ( 
.A1(n_5229),
.A2(n_237),
.B(n_238),
.Y(n_5336)
);

INVx2_ASAP7_75t_L g5337 ( 
.A(n_5183),
.Y(n_5337)
);

INVx1_ASAP7_75t_L g5338 ( 
.A(n_5244),
.Y(n_5338)
);

INVx3_ASAP7_75t_L g5339 ( 
.A(n_5196),
.Y(n_5339)
);

INVx1_ASAP7_75t_L g5340 ( 
.A(n_5193),
.Y(n_5340)
);

OAI21x1_ASAP7_75t_L g5341 ( 
.A1(n_5226),
.A2(n_238),
.B(n_239),
.Y(n_5341)
);

INVx1_ASAP7_75t_L g5342 ( 
.A(n_5216),
.Y(n_5342)
);

AO21x1_ASAP7_75t_SL g5343 ( 
.A1(n_5140),
.A2(n_241),
.B(n_242),
.Y(n_5343)
);

INVx1_ASAP7_75t_L g5344 ( 
.A(n_5142),
.Y(n_5344)
);

INVx1_ASAP7_75t_L g5345 ( 
.A(n_5283),
.Y(n_5345)
);

BUFx3_ASAP7_75t_L g5346 ( 
.A(n_5207),
.Y(n_5346)
);

AND2x4_ASAP7_75t_L g5347 ( 
.A(n_5153),
.B(n_241),
.Y(n_5347)
);

INVx6_ASAP7_75t_L g5348 ( 
.A(n_5144),
.Y(n_5348)
);

BUFx4f_ASAP7_75t_L g5349 ( 
.A(n_5281),
.Y(n_5349)
);

OA21x2_ASAP7_75t_L g5350 ( 
.A1(n_5174),
.A2(n_242),
.B(n_243),
.Y(n_5350)
);

INVx2_ASAP7_75t_L g5351 ( 
.A(n_5178),
.Y(n_5351)
);

OR2x6_ASAP7_75t_L g5352 ( 
.A(n_5240),
.B(n_244),
.Y(n_5352)
);

AND2x2_ASAP7_75t_L g5353 ( 
.A(n_5163),
.B(n_245),
.Y(n_5353)
);

INVx1_ASAP7_75t_L g5354 ( 
.A(n_5189),
.Y(n_5354)
);

BUFx3_ASAP7_75t_L g5355 ( 
.A(n_5248),
.Y(n_5355)
);

BUFx3_ASAP7_75t_L g5356 ( 
.A(n_5241),
.Y(n_5356)
);

INVx1_ASAP7_75t_L g5357 ( 
.A(n_5182),
.Y(n_5357)
);

INVx2_ASAP7_75t_L g5358 ( 
.A(n_5242),
.Y(n_5358)
);

INVx2_ASAP7_75t_L g5359 ( 
.A(n_5249),
.Y(n_5359)
);

CKINVDCx14_ASAP7_75t_R g5360 ( 
.A(n_5258),
.Y(n_5360)
);

INVx2_ASAP7_75t_L g5361 ( 
.A(n_5252),
.Y(n_5361)
);

INVx1_ASAP7_75t_L g5362 ( 
.A(n_5184),
.Y(n_5362)
);

BUFx6f_ASAP7_75t_L g5363 ( 
.A(n_5276),
.Y(n_5363)
);

INVx1_ASAP7_75t_L g5364 ( 
.A(n_5173),
.Y(n_5364)
);

O2A1O1Ixp33_ASAP7_75t_L g5365 ( 
.A1(n_5224),
.A2(n_247),
.B(n_245),
.C(n_246),
.Y(n_5365)
);

INVxp67_ASAP7_75t_R g5366 ( 
.A(n_5262),
.Y(n_5366)
);

INVxp67_ASAP7_75t_L g5367 ( 
.A(n_5160),
.Y(n_5367)
);

INVx1_ASAP7_75t_L g5368 ( 
.A(n_5180),
.Y(n_5368)
);

BUFx2_ASAP7_75t_L g5369 ( 
.A(n_5168),
.Y(n_5369)
);

INVx2_ASAP7_75t_L g5370 ( 
.A(n_5180),
.Y(n_5370)
);

INVx2_ASAP7_75t_L g5371 ( 
.A(n_5280),
.Y(n_5371)
);

INVx3_ASAP7_75t_L g5372 ( 
.A(n_5202),
.Y(n_5372)
);

INVx1_ASAP7_75t_L g5373 ( 
.A(n_5165),
.Y(n_5373)
);

INVx2_ASAP7_75t_SL g5374 ( 
.A(n_5179),
.Y(n_5374)
);

INVx1_ASAP7_75t_L g5375 ( 
.A(n_5185),
.Y(n_5375)
);

BUFx3_ASAP7_75t_L g5376 ( 
.A(n_5282),
.Y(n_5376)
);

INVx1_ASAP7_75t_L g5377 ( 
.A(n_5197),
.Y(n_5377)
);

AO21x2_ASAP7_75t_L g5378 ( 
.A1(n_5166),
.A2(n_246),
.B(n_248),
.Y(n_5378)
);

OAI21x1_ASAP7_75t_L g5379 ( 
.A1(n_5218),
.A2(n_249),
.B(n_251),
.Y(n_5379)
);

BUFx3_ASAP7_75t_L g5380 ( 
.A(n_5250),
.Y(n_5380)
);

BUFx5_ASAP7_75t_L g5381 ( 
.A(n_5279),
.Y(n_5381)
);

BUFx6f_ASAP7_75t_L g5382 ( 
.A(n_5209),
.Y(n_5382)
);

INVx2_ASAP7_75t_L g5383 ( 
.A(n_5206),
.Y(n_5383)
);

AOI21x1_ASAP7_75t_L g5384 ( 
.A1(n_5176),
.A2(n_249),
.B(n_252),
.Y(n_5384)
);

INVx2_ASAP7_75t_L g5385 ( 
.A(n_5277),
.Y(n_5385)
);

NAND2xp5_ASAP7_75t_L g5386 ( 
.A(n_5217),
.B(n_253),
.Y(n_5386)
);

INVx2_ASAP7_75t_L g5387 ( 
.A(n_5277),
.Y(n_5387)
);

INVx1_ASAP7_75t_L g5388 ( 
.A(n_5221),
.Y(n_5388)
);

HB1xp67_ASAP7_75t_L g5389 ( 
.A(n_5176),
.Y(n_5389)
);

AND2x2_ASAP7_75t_L g5390 ( 
.A(n_5253),
.B(n_253),
.Y(n_5390)
);

INVx1_ASAP7_75t_L g5391 ( 
.A(n_5151),
.Y(n_5391)
);

INVx1_ASAP7_75t_L g5392 ( 
.A(n_5190),
.Y(n_5392)
);

AOI22xp33_ASAP7_75t_L g5393 ( 
.A1(n_5208),
.A2(n_256),
.B1(n_254),
.B2(n_255),
.Y(n_5393)
);

INVx1_ASAP7_75t_L g5394 ( 
.A(n_5272),
.Y(n_5394)
);

OR2x6_ASAP7_75t_L g5395 ( 
.A(n_5234),
.B(n_254),
.Y(n_5395)
);

INVx1_ASAP7_75t_L g5396 ( 
.A(n_5257),
.Y(n_5396)
);

AO21x2_ASAP7_75t_L g5397 ( 
.A1(n_5164),
.A2(n_255),
.B(n_257),
.Y(n_5397)
);

INVx2_ASAP7_75t_L g5398 ( 
.A(n_5277),
.Y(n_5398)
);

AOI21xp5_ASAP7_75t_L g5399 ( 
.A1(n_5137),
.A2(n_257),
.B(n_258),
.Y(n_5399)
);

OAI21xp5_ASAP7_75t_L g5400 ( 
.A1(n_5284),
.A2(n_259),
.B(n_260),
.Y(n_5400)
);

INVx1_ASAP7_75t_L g5401 ( 
.A(n_5214),
.Y(n_5401)
);

HB1xp67_ASAP7_75t_L g5402 ( 
.A(n_5245),
.Y(n_5402)
);

INVx2_ASAP7_75t_L g5403 ( 
.A(n_5277),
.Y(n_5403)
);

NAND2xp5_ASAP7_75t_L g5404 ( 
.A(n_5219),
.B(n_5269),
.Y(n_5404)
);

INVx2_ASAP7_75t_L g5405 ( 
.A(n_5268),
.Y(n_5405)
);

INVx2_ASAP7_75t_L g5406 ( 
.A(n_5212),
.Y(n_5406)
);

INVx2_ASAP7_75t_L g5407 ( 
.A(n_5274),
.Y(n_5407)
);

AND2x2_ASAP7_75t_L g5408 ( 
.A(n_5171),
.B(n_259),
.Y(n_5408)
);

INVx1_ASAP7_75t_L g5409 ( 
.A(n_5222),
.Y(n_5409)
);

AND2x2_ASAP7_75t_L g5410 ( 
.A(n_5271),
.B(n_5275),
.Y(n_5410)
);

HB1xp67_ASAP7_75t_L g5411 ( 
.A(n_5223),
.Y(n_5411)
);

BUFx2_ASAP7_75t_L g5412 ( 
.A(n_5177),
.Y(n_5412)
);

AND2x2_ASAP7_75t_L g5413 ( 
.A(n_5233),
.B(n_260),
.Y(n_5413)
);

INVx1_ASAP7_75t_L g5414 ( 
.A(n_5251),
.Y(n_5414)
);

INVx2_ASAP7_75t_L g5415 ( 
.A(n_5256),
.Y(n_5415)
);

INVx2_ASAP7_75t_L g5416 ( 
.A(n_5260),
.Y(n_5416)
);

INVx2_ASAP7_75t_L g5417 ( 
.A(n_5181),
.Y(n_5417)
);

OAI22xp5_ASAP7_75t_L g5418 ( 
.A1(n_5154),
.A2(n_263),
.B1(n_261),
.B2(n_262),
.Y(n_5418)
);

BUFx2_ASAP7_75t_SL g5419 ( 
.A(n_5243),
.Y(n_5419)
);

NOR2x1_ASAP7_75t_SL g5420 ( 
.A(n_5148),
.B(n_261),
.Y(n_5420)
);

BUFx6f_ASAP7_75t_L g5421 ( 
.A(n_5175),
.Y(n_5421)
);

INVx1_ASAP7_75t_L g5422 ( 
.A(n_5198),
.Y(n_5422)
);

INVx1_ASAP7_75t_L g5423 ( 
.A(n_5200),
.Y(n_5423)
);

INVx2_ASAP7_75t_L g5424 ( 
.A(n_5273),
.Y(n_5424)
);

AOI221x1_ASAP7_75t_L g5425 ( 
.A1(n_5246),
.A2(n_266),
.B1(n_263),
.B2(n_265),
.C(n_267),
.Y(n_5425)
);

INVx2_ASAP7_75t_L g5426 ( 
.A(n_5235),
.Y(n_5426)
);

OR2x2_ASAP7_75t_L g5427 ( 
.A(n_5266),
.B(n_265),
.Y(n_5427)
);

BUFx2_ASAP7_75t_L g5428 ( 
.A(n_5152),
.Y(n_5428)
);

OAI22xp5_ASAP7_75t_L g5429 ( 
.A1(n_5156),
.A2(n_270),
.B1(n_268),
.B2(n_269),
.Y(n_5429)
);

INVx1_ASAP7_75t_L g5430 ( 
.A(n_5199),
.Y(n_5430)
);

INVx1_ASAP7_75t_L g5431 ( 
.A(n_5210),
.Y(n_5431)
);

BUFx3_ASAP7_75t_L g5432 ( 
.A(n_5147),
.Y(n_5432)
);

INVx2_ASAP7_75t_L g5433 ( 
.A(n_5254),
.Y(n_5433)
);

AO31x2_ASAP7_75t_L g5434 ( 
.A1(n_5264),
.A2(n_278),
.A3(n_287),
.B(n_268),
.Y(n_5434)
);

OAI22xp33_ASAP7_75t_SL g5435 ( 
.A1(n_5236),
.A2(n_272),
.B1(n_269),
.B2(n_270),
.Y(n_5435)
);

INVx2_ASAP7_75t_L g5436 ( 
.A(n_5172),
.Y(n_5436)
);

AND2x2_ASAP7_75t_L g5437 ( 
.A(n_5143),
.B(n_273),
.Y(n_5437)
);

INVx1_ASAP7_75t_L g5438 ( 
.A(n_5145),
.Y(n_5438)
);

AND2x2_ASAP7_75t_L g5439 ( 
.A(n_5143),
.B(n_274),
.Y(n_5439)
);

AOI221xp5_ASAP7_75t_L g5440 ( 
.A1(n_5200),
.A2(n_277),
.B1(n_274),
.B2(n_276),
.C(n_278),
.Y(n_5440)
);

INVx1_ASAP7_75t_L g5441 ( 
.A(n_5145),
.Y(n_5441)
);

INVx3_ASAP7_75t_L g5442 ( 
.A(n_5138),
.Y(n_5442)
);

INVx2_ASAP7_75t_L g5443 ( 
.A(n_5169),
.Y(n_5443)
);

NAND2xp5_ASAP7_75t_L g5444 ( 
.A(n_5203),
.B(n_276),
.Y(n_5444)
);

INVx1_ASAP7_75t_L g5445 ( 
.A(n_5145),
.Y(n_5445)
);

INVx1_ASAP7_75t_L g5446 ( 
.A(n_5145),
.Y(n_5446)
);

INVx3_ASAP7_75t_L g5447 ( 
.A(n_5138),
.Y(n_5447)
);

INVx1_ASAP7_75t_L g5448 ( 
.A(n_5307),
.Y(n_5448)
);

BUFx3_ASAP7_75t_L g5449 ( 
.A(n_5356),
.Y(n_5449)
);

BUFx2_ASAP7_75t_L g5450 ( 
.A(n_5286),
.Y(n_5450)
);

BUFx3_ASAP7_75t_L g5451 ( 
.A(n_5376),
.Y(n_5451)
);

OR2x2_ASAP7_75t_L g5452 ( 
.A(n_5300),
.B(n_277),
.Y(n_5452)
);

INVx1_ASAP7_75t_L g5453 ( 
.A(n_5308),
.Y(n_5453)
);

AND2x2_ASAP7_75t_L g5454 ( 
.A(n_5369),
.B(n_279),
.Y(n_5454)
);

AND2x2_ASAP7_75t_L g5455 ( 
.A(n_5388),
.B(n_279),
.Y(n_5455)
);

INVx1_ASAP7_75t_L g5456 ( 
.A(n_5310),
.Y(n_5456)
);

AND2x2_ASAP7_75t_L g5457 ( 
.A(n_5373),
.B(n_280),
.Y(n_5457)
);

AO31x2_ASAP7_75t_L g5458 ( 
.A1(n_5412),
.A2(n_283),
.A3(n_280),
.B(n_282),
.Y(n_5458)
);

AND2x2_ASAP7_75t_L g5459 ( 
.A(n_5330),
.B(n_284),
.Y(n_5459)
);

INVx1_ASAP7_75t_L g5460 ( 
.A(n_5338),
.Y(n_5460)
);

OR2x2_ASAP7_75t_L g5461 ( 
.A(n_5302),
.B(n_284),
.Y(n_5461)
);

INVx2_ASAP7_75t_L g5462 ( 
.A(n_5358),
.Y(n_5462)
);

AND2x2_ASAP7_75t_L g5463 ( 
.A(n_5337),
.B(n_285),
.Y(n_5463)
);

AND2x4_ASAP7_75t_L g5464 ( 
.A(n_5363),
.B(n_285),
.Y(n_5464)
);

INVx1_ASAP7_75t_L g5465 ( 
.A(n_5288),
.Y(n_5465)
);

AND2x2_ASAP7_75t_L g5466 ( 
.A(n_5340),
.B(n_286),
.Y(n_5466)
);

INVx2_ASAP7_75t_L g5467 ( 
.A(n_5359),
.Y(n_5467)
);

AND2x2_ASAP7_75t_L g5468 ( 
.A(n_5296),
.B(n_288),
.Y(n_5468)
);

INVx2_ASAP7_75t_SL g5469 ( 
.A(n_5348),
.Y(n_5469)
);

BUFx2_ASAP7_75t_L g5470 ( 
.A(n_5297),
.Y(n_5470)
);

AND2x2_ASAP7_75t_L g5471 ( 
.A(n_5366),
.B(n_288),
.Y(n_5471)
);

INVx2_ASAP7_75t_SL g5472 ( 
.A(n_5346),
.Y(n_5472)
);

AND2x4_ASAP7_75t_L g5473 ( 
.A(n_5363),
.B(n_5339),
.Y(n_5473)
);

INVx3_ASAP7_75t_L g5474 ( 
.A(n_5287),
.Y(n_5474)
);

HB1xp67_ASAP7_75t_L g5475 ( 
.A(n_5321),
.Y(n_5475)
);

INVx2_ASAP7_75t_L g5476 ( 
.A(n_5361),
.Y(n_5476)
);

INVx2_ASAP7_75t_L g5477 ( 
.A(n_5391),
.Y(n_5477)
);

INVx1_ASAP7_75t_L g5478 ( 
.A(n_5289),
.Y(n_5478)
);

INVx5_ASAP7_75t_L g5479 ( 
.A(n_5352),
.Y(n_5479)
);

INVx1_ASAP7_75t_L g5480 ( 
.A(n_5438),
.Y(n_5480)
);

AND2x2_ASAP7_75t_L g5481 ( 
.A(n_5345),
.B(n_289),
.Y(n_5481)
);

INVx1_ASAP7_75t_L g5482 ( 
.A(n_5441),
.Y(n_5482)
);

AND2x4_ASAP7_75t_L g5483 ( 
.A(n_5382),
.B(n_5372),
.Y(n_5483)
);

INVx1_ASAP7_75t_L g5484 ( 
.A(n_5445),
.Y(n_5484)
);

INVx1_ASAP7_75t_L g5485 ( 
.A(n_5446),
.Y(n_5485)
);

OR2x2_ASAP7_75t_L g5486 ( 
.A(n_5335),
.B(n_290),
.Y(n_5486)
);

BUFx6f_ASAP7_75t_L g5487 ( 
.A(n_5287),
.Y(n_5487)
);

INVx1_ASAP7_75t_L g5488 ( 
.A(n_5368),
.Y(n_5488)
);

AND2x4_ASAP7_75t_L g5489 ( 
.A(n_5382),
.B(n_291),
.Y(n_5489)
);

NAND2xp5_ASAP7_75t_L g5490 ( 
.A(n_5323),
.B(n_291),
.Y(n_5490)
);

AND2x2_ASAP7_75t_L g5491 ( 
.A(n_5392),
.B(n_292),
.Y(n_5491)
);

INVx1_ASAP7_75t_L g5492 ( 
.A(n_5295),
.Y(n_5492)
);

OR2x2_ASAP7_75t_L g5493 ( 
.A(n_5331),
.B(n_293),
.Y(n_5493)
);

BUFx3_ASAP7_75t_L g5494 ( 
.A(n_5355),
.Y(n_5494)
);

INVx1_ASAP7_75t_L g5495 ( 
.A(n_5313),
.Y(n_5495)
);

AND2x2_ASAP7_75t_L g5496 ( 
.A(n_5311),
.B(n_293),
.Y(n_5496)
);

AND2x2_ASAP7_75t_L g5497 ( 
.A(n_5317),
.B(n_295),
.Y(n_5497)
);

AND2x2_ASAP7_75t_L g5498 ( 
.A(n_5380),
.B(n_295),
.Y(n_5498)
);

INVx1_ASAP7_75t_L g5499 ( 
.A(n_5318),
.Y(n_5499)
);

AOI22xp33_ASAP7_75t_L g5500 ( 
.A1(n_5428),
.A2(n_298),
.B1(n_296),
.B2(n_297),
.Y(n_5500)
);

NAND2xp5_ASAP7_75t_L g5501 ( 
.A(n_5344),
.B(n_296),
.Y(n_5501)
);

INVx1_ASAP7_75t_L g5502 ( 
.A(n_5370),
.Y(n_5502)
);

INVx3_ASAP7_75t_L g5503 ( 
.A(n_5285),
.Y(n_5503)
);

INVx2_ASAP7_75t_L g5504 ( 
.A(n_5304),
.Y(n_5504)
);

NAND2xp5_ASAP7_75t_L g5505 ( 
.A(n_5324),
.B(n_298),
.Y(n_5505)
);

BUFx3_ASAP7_75t_L g5506 ( 
.A(n_5374),
.Y(n_5506)
);

INVxp67_ASAP7_75t_L g5507 ( 
.A(n_5343),
.Y(n_5507)
);

AOI22xp33_ASAP7_75t_L g5508 ( 
.A1(n_5426),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.Y(n_5508)
);

INVx1_ASAP7_75t_L g5509 ( 
.A(n_5342),
.Y(n_5509)
);

AND2x4_ASAP7_75t_L g5510 ( 
.A(n_5351),
.B(n_299),
.Y(n_5510)
);

AND2x4_ASAP7_75t_L g5511 ( 
.A(n_5375),
.B(n_300),
.Y(n_5511)
);

OR2x2_ASAP7_75t_L g5512 ( 
.A(n_5334),
.B(n_301),
.Y(n_5512)
);

INVx2_ASAP7_75t_L g5513 ( 
.A(n_5319),
.Y(n_5513)
);

OAI22xp5_ASAP7_75t_L g5514 ( 
.A1(n_5395),
.A2(n_305),
.B1(n_302),
.B2(n_304),
.Y(n_5514)
);

OR2x2_ASAP7_75t_L g5515 ( 
.A(n_5406),
.B(n_302),
.Y(n_5515)
);

NAND2xp5_ASAP7_75t_L g5516 ( 
.A(n_5354),
.B(n_305),
.Y(n_5516)
);

AND2x4_ASAP7_75t_L g5517 ( 
.A(n_5377),
.B(n_307),
.Y(n_5517)
);

INVx1_ASAP7_75t_L g5518 ( 
.A(n_5298),
.Y(n_5518)
);

AOI22xp33_ASAP7_75t_L g5519 ( 
.A1(n_5423),
.A2(n_309),
.B1(n_307),
.B2(n_308),
.Y(n_5519)
);

NAND2xp5_ASAP7_75t_L g5520 ( 
.A(n_5357),
.B(n_308),
.Y(n_5520)
);

INVx1_ASAP7_75t_L g5521 ( 
.A(n_5299),
.Y(n_5521)
);

HB1xp67_ASAP7_75t_L g5522 ( 
.A(n_5411),
.Y(n_5522)
);

INVx2_ASAP7_75t_L g5523 ( 
.A(n_5314),
.Y(n_5523)
);

NAND2xp5_ASAP7_75t_L g5524 ( 
.A(n_5362),
.B(n_309),
.Y(n_5524)
);

INVx2_ASAP7_75t_L g5525 ( 
.A(n_5327),
.Y(n_5525)
);

AND2x2_ASAP7_75t_L g5526 ( 
.A(n_5360),
.B(n_310),
.Y(n_5526)
);

HB1xp67_ASAP7_75t_L g5527 ( 
.A(n_5389),
.Y(n_5527)
);

HB1xp67_ASAP7_75t_L g5528 ( 
.A(n_5364),
.Y(n_5528)
);

AND2x2_ASAP7_75t_L g5529 ( 
.A(n_5305),
.B(n_310),
.Y(n_5529)
);

BUFx2_ASAP7_75t_L g5530 ( 
.A(n_5442),
.Y(n_5530)
);

AND2x2_ASAP7_75t_L g5531 ( 
.A(n_5407),
.B(n_311),
.Y(n_5531)
);

AND2x2_ASAP7_75t_L g5532 ( 
.A(n_5447),
.B(n_311),
.Y(n_5532)
);

AND2x2_ASAP7_75t_L g5533 ( 
.A(n_5349),
.B(n_312),
.Y(n_5533)
);

INVx1_ASAP7_75t_L g5534 ( 
.A(n_5301),
.Y(n_5534)
);

INVx1_ASAP7_75t_L g5535 ( 
.A(n_5396),
.Y(n_5535)
);

INVx2_ASAP7_75t_L g5536 ( 
.A(n_5326),
.Y(n_5536)
);

OR2x2_ASAP7_75t_L g5537 ( 
.A(n_5405),
.B(n_312),
.Y(n_5537)
);

AND2x2_ASAP7_75t_L g5538 ( 
.A(n_5367),
.B(n_313),
.Y(n_5538)
);

NOR2xp33_ASAP7_75t_L g5539 ( 
.A(n_5325),
.B(n_315),
.Y(n_5539)
);

INVx1_ASAP7_75t_L g5540 ( 
.A(n_5292),
.Y(n_5540)
);

AND2x2_ASAP7_75t_L g5541 ( 
.A(n_5332),
.B(n_315),
.Y(n_5541)
);

NOR2x1p5_ASAP7_75t_L g5542 ( 
.A(n_5404),
.B(n_316),
.Y(n_5542)
);

INVx2_ASAP7_75t_L g5543 ( 
.A(n_5316),
.Y(n_5543)
);

NAND2xp5_ASAP7_75t_L g5544 ( 
.A(n_5409),
.B(n_316),
.Y(n_5544)
);

INVx3_ASAP7_75t_L g5545 ( 
.A(n_5347),
.Y(n_5545)
);

AND2x2_ASAP7_75t_L g5546 ( 
.A(n_5383),
.B(n_317),
.Y(n_5546)
);

AND2x2_ASAP7_75t_L g5547 ( 
.A(n_5414),
.B(n_317),
.Y(n_5547)
);

INVx3_ASAP7_75t_SL g5548 ( 
.A(n_5352),
.Y(n_5548)
);

BUFx6f_ASAP7_75t_L g5549 ( 
.A(n_5421),
.Y(n_5549)
);

INVx1_ASAP7_75t_L g5550 ( 
.A(n_5443),
.Y(n_5550)
);

OR2x2_ASAP7_75t_L g5551 ( 
.A(n_5315),
.B(n_318),
.Y(n_5551)
);

INVx1_ASAP7_75t_L g5552 ( 
.A(n_5394),
.Y(n_5552)
);

INVx1_ASAP7_75t_L g5553 ( 
.A(n_5371),
.Y(n_5553)
);

NAND2xp5_ASAP7_75t_L g5554 ( 
.A(n_5381),
.B(n_318),
.Y(n_5554)
);

OAI22xp5_ASAP7_75t_L g5555 ( 
.A1(n_5395),
.A2(n_321),
.B1(n_319),
.B2(n_320),
.Y(n_5555)
);

AND2x2_ASAP7_75t_L g5556 ( 
.A(n_5401),
.B(n_320),
.Y(n_5556)
);

INVx1_ASAP7_75t_L g5557 ( 
.A(n_5294),
.Y(n_5557)
);

BUFx3_ASAP7_75t_L g5558 ( 
.A(n_5353),
.Y(n_5558)
);

INVx1_ASAP7_75t_L g5559 ( 
.A(n_5415),
.Y(n_5559)
);

INVx2_ASAP7_75t_L g5560 ( 
.A(n_5381),
.Y(n_5560)
);

AND2x2_ASAP7_75t_L g5561 ( 
.A(n_5322),
.B(n_321),
.Y(n_5561)
);

AOI22xp5_ASAP7_75t_L g5562 ( 
.A1(n_5290),
.A2(n_326),
.B1(n_324),
.B2(n_325),
.Y(n_5562)
);

OR2x2_ASAP7_75t_L g5563 ( 
.A(n_5416),
.B(n_324),
.Y(n_5563)
);

AND2x2_ASAP7_75t_L g5564 ( 
.A(n_5437),
.B(n_326),
.Y(n_5564)
);

INVx1_ASAP7_75t_L g5565 ( 
.A(n_5291),
.Y(n_5565)
);

INVx1_ASAP7_75t_L g5566 ( 
.A(n_5381),
.Y(n_5566)
);

OR2x6_ASAP7_75t_L g5567 ( 
.A(n_5421),
.B(n_327),
.Y(n_5567)
);

INVx1_ASAP7_75t_L g5568 ( 
.A(n_5444),
.Y(n_5568)
);

AND2x2_ASAP7_75t_L g5569 ( 
.A(n_5439),
.B(n_328),
.Y(n_5569)
);

INVxp67_ASAP7_75t_SL g5570 ( 
.A(n_5386),
.Y(n_5570)
);

INVx2_ASAP7_75t_L g5571 ( 
.A(n_5422),
.Y(n_5571)
);

INVx2_ASAP7_75t_L g5572 ( 
.A(n_5293),
.Y(n_5572)
);

INVx4_ASAP7_75t_L g5573 ( 
.A(n_5408),
.Y(n_5573)
);

INVx1_ASAP7_75t_L g5574 ( 
.A(n_5333),
.Y(n_5574)
);

OR2x2_ASAP7_75t_L g5575 ( 
.A(n_5303),
.B(n_328),
.Y(n_5575)
);

INVx1_ASAP7_75t_L g5576 ( 
.A(n_5385),
.Y(n_5576)
);

INVx3_ASAP7_75t_L g5577 ( 
.A(n_5410),
.Y(n_5577)
);

INVx1_ASAP7_75t_L g5578 ( 
.A(n_5387),
.Y(n_5578)
);

BUFx2_ASAP7_75t_L g5579 ( 
.A(n_5398),
.Y(n_5579)
);

OA21x2_ASAP7_75t_L g5580 ( 
.A1(n_5306),
.A2(n_329),
.B(n_330),
.Y(n_5580)
);

AOI22xp33_ASAP7_75t_L g5581 ( 
.A1(n_5431),
.A2(n_333),
.B1(n_330),
.B2(n_332),
.Y(n_5581)
);

OR2x2_ASAP7_75t_L g5582 ( 
.A(n_5403),
.B(n_332),
.Y(n_5582)
);

INVx1_ASAP7_75t_L g5583 ( 
.A(n_5336),
.Y(n_5583)
);

NAND2xp5_ASAP7_75t_L g5584 ( 
.A(n_5436),
.B(n_333),
.Y(n_5584)
);

AND2x2_ASAP7_75t_L g5585 ( 
.A(n_5328),
.B(n_334),
.Y(n_5585)
);

INVx1_ASAP7_75t_L g5586 ( 
.A(n_5397),
.Y(n_5586)
);

OAI222xp33_ASAP7_75t_L g5587 ( 
.A1(n_5312),
.A2(n_337),
.B1(n_339),
.B2(n_334),
.C1(n_335),
.C2(n_338),
.Y(n_5587)
);

INVx2_ASAP7_75t_L g5588 ( 
.A(n_5341),
.Y(n_5588)
);

OR2x2_ASAP7_75t_L g5589 ( 
.A(n_5329),
.B(n_335),
.Y(n_5589)
);

INVxp67_ASAP7_75t_L g5590 ( 
.A(n_5402),
.Y(n_5590)
);

AND2x2_ASAP7_75t_L g5591 ( 
.A(n_5390),
.B(n_339),
.Y(n_5591)
);

INVx1_ASAP7_75t_L g5592 ( 
.A(n_5417),
.Y(n_5592)
);

AO21x2_ASAP7_75t_L g5593 ( 
.A1(n_5384),
.A2(n_340),
.B(n_341),
.Y(n_5593)
);

AOI22xp33_ASAP7_75t_L g5594 ( 
.A1(n_5430),
.A2(n_343),
.B1(n_340),
.B2(n_342),
.Y(n_5594)
);

INVx2_ASAP7_75t_L g5595 ( 
.A(n_5378),
.Y(n_5595)
);

INVxp67_ASAP7_75t_SL g5596 ( 
.A(n_5432),
.Y(n_5596)
);

NAND2xp5_ASAP7_75t_L g5597 ( 
.A(n_5433),
.B(n_344),
.Y(n_5597)
);

HB1xp67_ASAP7_75t_L g5598 ( 
.A(n_5424),
.Y(n_5598)
);

CKINVDCx5p33_ASAP7_75t_R g5599 ( 
.A(n_5413),
.Y(n_5599)
);

INVx1_ASAP7_75t_L g5600 ( 
.A(n_5350),
.Y(n_5600)
);

INVx1_ASAP7_75t_L g5601 ( 
.A(n_5434),
.Y(n_5601)
);

INVx1_ASAP7_75t_L g5602 ( 
.A(n_5434),
.Y(n_5602)
);

AND2x2_ASAP7_75t_L g5603 ( 
.A(n_5420),
.B(n_344),
.Y(n_5603)
);

INVx1_ASAP7_75t_SL g5604 ( 
.A(n_5320),
.Y(n_5604)
);

INVx2_ASAP7_75t_L g5605 ( 
.A(n_5379),
.Y(n_5605)
);

NAND2xp5_ASAP7_75t_L g5606 ( 
.A(n_5399),
.B(n_345),
.Y(n_5606)
);

HB1xp67_ASAP7_75t_L g5607 ( 
.A(n_5418),
.Y(n_5607)
);

INVx1_ASAP7_75t_L g5608 ( 
.A(n_5427),
.Y(n_5608)
);

AO31x2_ASAP7_75t_L g5609 ( 
.A1(n_5429),
.A2(n_347),
.A3(n_345),
.B(n_346),
.Y(n_5609)
);

BUFx2_ASAP7_75t_SL g5610 ( 
.A(n_5419),
.Y(n_5610)
);

AOI222xp33_ASAP7_75t_L g5611 ( 
.A1(n_5440),
.A2(n_349),
.B1(n_352),
.B2(n_347),
.C1(n_348),
.C2(n_351),
.Y(n_5611)
);

AOI22xp33_ASAP7_75t_L g5612 ( 
.A1(n_5309),
.A2(n_353),
.B1(n_351),
.B2(n_352),
.Y(n_5612)
);

INVx2_ASAP7_75t_L g5613 ( 
.A(n_5400),
.Y(n_5613)
);

HB1xp67_ASAP7_75t_L g5614 ( 
.A(n_5435),
.Y(n_5614)
);

OAI22xp5_ASAP7_75t_L g5615 ( 
.A1(n_5393),
.A2(n_357),
.B1(n_355),
.B2(n_356),
.Y(n_5615)
);

INVx1_ASAP7_75t_L g5616 ( 
.A(n_5365),
.Y(n_5616)
);

AOI22xp33_ASAP7_75t_L g5617 ( 
.A1(n_5425),
.A2(n_357),
.B1(n_355),
.B2(n_356),
.Y(n_5617)
);

INVx2_ASAP7_75t_L g5618 ( 
.A(n_5358),
.Y(n_5618)
);

INVx2_ASAP7_75t_L g5619 ( 
.A(n_5358),
.Y(n_5619)
);

BUFx2_ASAP7_75t_L g5620 ( 
.A(n_5286),
.Y(n_5620)
);

NAND2xp5_ASAP7_75t_L g5621 ( 
.A(n_5323),
.B(n_358),
.Y(n_5621)
);

INVx2_ASAP7_75t_R g5622 ( 
.A(n_5396),
.Y(n_5622)
);

AOI22xp33_ASAP7_75t_L g5623 ( 
.A1(n_5428),
.A2(n_362),
.B1(n_359),
.B2(n_360),
.Y(n_5623)
);

OR2x2_ASAP7_75t_L g5624 ( 
.A(n_5300),
.B(n_359),
.Y(n_5624)
);

AND2x2_ASAP7_75t_L g5625 ( 
.A(n_5369),
.B(n_360),
.Y(n_5625)
);

INVx2_ASAP7_75t_L g5626 ( 
.A(n_5358),
.Y(n_5626)
);

AND2x2_ASAP7_75t_L g5627 ( 
.A(n_5369),
.B(n_362),
.Y(n_5627)
);

AOI22xp5_ASAP7_75t_L g5628 ( 
.A1(n_5428),
.A2(n_366),
.B1(n_363),
.B2(n_364),
.Y(n_5628)
);

AO21x2_ASAP7_75t_L g5629 ( 
.A1(n_5392),
.A2(n_363),
.B(n_364),
.Y(n_5629)
);

INVxp67_ASAP7_75t_SL g5630 ( 
.A(n_5596),
.Y(n_5630)
);

INVx2_ASAP7_75t_L g5631 ( 
.A(n_5572),
.Y(n_5631)
);

OR2x2_ASAP7_75t_L g5632 ( 
.A(n_5565),
.B(n_366),
.Y(n_5632)
);

AND2x2_ASAP7_75t_L g5633 ( 
.A(n_5577),
.B(n_368),
.Y(n_5633)
);

INVx2_ASAP7_75t_L g5634 ( 
.A(n_5571),
.Y(n_5634)
);

INVx2_ASAP7_75t_L g5635 ( 
.A(n_5462),
.Y(n_5635)
);

INVx1_ASAP7_75t_L g5636 ( 
.A(n_5528),
.Y(n_5636)
);

AND2x4_ASAP7_75t_L g5637 ( 
.A(n_5450),
.B(n_369),
.Y(n_5637)
);

AND2x4_ASAP7_75t_L g5638 ( 
.A(n_5620),
.B(n_370),
.Y(n_5638)
);

AND2x2_ASAP7_75t_L g5639 ( 
.A(n_5530),
.B(n_370),
.Y(n_5639)
);

HB1xp67_ASAP7_75t_L g5640 ( 
.A(n_5592),
.Y(n_5640)
);

INVx1_ASAP7_75t_L g5641 ( 
.A(n_5488),
.Y(n_5641)
);

AND2x2_ASAP7_75t_L g5642 ( 
.A(n_5473),
.B(n_371),
.Y(n_5642)
);

BUFx2_ASAP7_75t_L g5643 ( 
.A(n_5451),
.Y(n_5643)
);

INVx2_ASAP7_75t_L g5644 ( 
.A(n_5467),
.Y(n_5644)
);

INVxp67_ASAP7_75t_L g5645 ( 
.A(n_5470),
.Y(n_5645)
);

NOR2xp33_ASAP7_75t_R g5646 ( 
.A(n_5548),
.B(n_5599),
.Y(n_5646)
);

INVx1_ASAP7_75t_L g5647 ( 
.A(n_5475),
.Y(n_5647)
);

HB1xp67_ASAP7_75t_L g5648 ( 
.A(n_5522),
.Y(n_5648)
);

INVx2_ASAP7_75t_SL g5649 ( 
.A(n_5479),
.Y(n_5649)
);

INVx1_ASAP7_75t_L g5650 ( 
.A(n_5535),
.Y(n_5650)
);

AND2x2_ASAP7_75t_L g5651 ( 
.A(n_5503),
.B(n_371),
.Y(n_5651)
);

INVxp67_ASAP7_75t_SL g5652 ( 
.A(n_5598),
.Y(n_5652)
);

INVx1_ASAP7_75t_L g5653 ( 
.A(n_5495),
.Y(n_5653)
);

AO31x2_ASAP7_75t_L g5654 ( 
.A1(n_5586),
.A2(n_381),
.A3(n_389),
.B(n_373),
.Y(n_5654)
);

INVx2_ASAP7_75t_L g5655 ( 
.A(n_5476),
.Y(n_5655)
);

INVx3_ASAP7_75t_L g5656 ( 
.A(n_5506),
.Y(n_5656)
);

HB1xp67_ASAP7_75t_L g5657 ( 
.A(n_5527),
.Y(n_5657)
);

AND2x2_ASAP7_75t_L g5658 ( 
.A(n_5590),
.B(n_373),
.Y(n_5658)
);

AND2x2_ASAP7_75t_L g5659 ( 
.A(n_5573),
.B(n_374),
.Y(n_5659)
);

INVx2_ASAP7_75t_L g5660 ( 
.A(n_5618),
.Y(n_5660)
);

HB1xp67_ASAP7_75t_L g5661 ( 
.A(n_5583),
.Y(n_5661)
);

INVx1_ASAP7_75t_L g5662 ( 
.A(n_5552),
.Y(n_5662)
);

INVx1_ASAP7_75t_L g5663 ( 
.A(n_5448),
.Y(n_5663)
);

NOR2x1_ASAP7_75t_L g5664 ( 
.A(n_5494),
.B(n_375),
.Y(n_5664)
);

INVx2_ASAP7_75t_SL g5665 ( 
.A(n_5479),
.Y(n_5665)
);

NAND2xp33_ASAP7_75t_L g5666 ( 
.A(n_5607),
.B(n_375),
.Y(n_5666)
);

INVx1_ASAP7_75t_L g5667 ( 
.A(n_5453),
.Y(n_5667)
);

AND2x2_ASAP7_75t_L g5668 ( 
.A(n_5610),
.B(n_376),
.Y(n_5668)
);

AND2x2_ASAP7_75t_L g5669 ( 
.A(n_5568),
.B(n_377),
.Y(n_5669)
);

AND2x4_ASAP7_75t_L g5670 ( 
.A(n_5472),
.B(n_378),
.Y(n_5670)
);

INVx2_ASAP7_75t_L g5671 ( 
.A(n_5619),
.Y(n_5671)
);

OR2x2_ASAP7_75t_L g5672 ( 
.A(n_5570),
.B(n_379),
.Y(n_5672)
);

INVx1_ASAP7_75t_L g5673 ( 
.A(n_5456),
.Y(n_5673)
);

INVx1_ASAP7_75t_SL g5674 ( 
.A(n_5558),
.Y(n_5674)
);

AND2x2_ASAP7_75t_L g5675 ( 
.A(n_5545),
.B(n_5474),
.Y(n_5675)
);

BUFx2_ASAP7_75t_L g5676 ( 
.A(n_5449),
.Y(n_5676)
);

OR2x2_ASAP7_75t_L g5677 ( 
.A(n_5509),
.B(n_379),
.Y(n_5677)
);

AND2x4_ASAP7_75t_L g5678 ( 
.A(n_5483),
.B(n_380),
.Y(n_5678)
);

AND2x2_ASAP7_75t_L g5679 ( 
.A(n_5579),
.B(n_380),
.Y(n_5679)
);

INVx1_ASAP7_75t_L g5680 ( 
.A(n_5465),
.Y(n_5680)
);

BUFx2_ASAP7_75t_L g5681 ( 
.A(n_5507),
.Y(n_5681)
);

INVx1_ASAP7_75t_L g5682 ( 
.A(n_5478),
.Y(n_5682)
);

INVx1_ASAP7_75t_L g5683 ( 
.A(n_5480),
.Y(n_5683)
);

INVx2_ASAP7_75t_R g5684 ( 
.A(n_5601),
.Y(n_5684)
);

INVxp67_ASAP7_75t_L g5685 ( 
.A(n_5608),
.Y(n_5685)
);

INVx1_ASAP7_75t_L g5686 ( 
.A(n_5482),
.Y(n_5686)
);

INVx1_ASAP7_75t_L g5687 ( 
.A(n_5484),
.Y(n_5687)
);

AND2x2_ASAP7_75t_L g5688 ( 
.A(n_5454),
.B(n_381),
.Y(n_5688)
);

AND2x2_ASAP7_75t_L g5689 ( 
.A(n_5625),
.B(n_382),
.Y(n_5689)
);

AOI222xp33_ASAP7_75t_L g5690 ( 
.A1(n_5616),
.A2(n_385),
.B1(n_387),
.B2(n_383),
.C1(n_384),
.C2(n_386),
.Y(n_5690)
);

INVx5_ASAP7_75t_L g5691 ( 
.A(n_5567),
.Y(n_5691)
);

INVx2_ASAP7_75t_L g5692 ( 
.A(n_5626),
.Y(n_5692)
);

INVx1_ASAP7_75t_L g5693 ( 
.A(n_5485),
.Y(n_5693)
);

INVx1_ASAP7_75t_L g5694 ( 
.A(n_5492),
.Y(n_5694)
);

AND2x2_ASAP7_75t_L g5695 ( 
.A(n_5627),
.B(n_383),
.Y(n_5695)
);

INVx2_ASAP7_75t_L g5696 ( 
.A(n_5605),
.Y(n_5696)
);

OR2x2_ASAP7_75t_L g5697 ( 
.A(n_5574),
.B(n_385),
.Y(n_5697)
);

INVx2_ASAP7_75t_L g5698 ( 
.A(n_5595),
.Y(n_5698)
);

INVx2_ASAP7_75t_L g5699 ( 
.A(n_5525),
.Y(n_5699)
);

INVx2_ASAP7_75t_L g5700 ( 
.A(n_5477),
.Y(n_5700)
);

INVx2_ASAP7_75t_L g5701 ( 
.A(n_5576),
.Y(n_5701)
);

OR2x2_ASAP7_75t_L g5702 ( 
.A(n_5499),
.B(n_386),
.Y(n_5702)
);

NAND2xp5_ASAP7_75t_L g5703 ( 
.A(n_5497),
.B(n_387),
.Y(n_5703)
);

INVx1_ASAP7_75t_L g5704 ( 
.A(n_5460),
.Y(n_5704)
);

HB1xp67_ASAP7_75t_L g5705 ( 
.A(n_5600),
.Y(n_5705)
);

AND2x2_ASAP7_75t_L g5706 ( 
.A(n_5466),
.B(n_388),
.Y(n_5706)
);

INVx2_ASAP7_75t_L g5707 ( 
.A(n_5578),
.Y(n_5707)
);

HB1xp67_ASAP7_75t_L g5708 ( 
.A(n_5588),
.Y(n_5708)
);

INVx1_ASAP7_75t_L g5709 ( 
.A(n_5518),
.Y(n_5709)
);

AND2x2_ASAP7_75t_L g5710 ( 
.A(n_5622),
.B(n_389),
.Y(n_5710)
);

NAND2xp5_ASAP7_75t_L g5711 ( 
.A(n_5468),
.B(n_5490),
.Y(n_5711)
);

INVx1_ASAP7_75t_L g5712 ( 
.A(n_5521),
.Y(n_5712)
);

INVx2_ASAP7_75t_SL g5713 ( 
.A(n_5469),
.Y(n_5713)
);

NAND2xp5_ASAP7_75t_L g5714 ( 
.A(n_5621),
.B(n_390),
.Y(n_5714)
);

OR2x2_ASAP7_75t_L g5715 ( 
.A(n_5486),
.B(n_390),
.Y(n_5715)
);

HB1xp67_ASAP7_75t_L g5716 ( 
.A(n_5452),
.Y(n_5716)
);

HB1xp67_ASAP7_75t_L g5717 ( 
.A(n_5624),
.Y(n_5717)
);

BUFx6f_ASAP7_75t_L g5718 ( 
.A(n_5487),
.Y(n_5718)
);

NAND2xp5_ASAP7_75t_L g5719 ( 
.A(n_5501),
.B(n_391),
.Y(n_5719)
);

INVx1_ASAP7_75t_L g5720 ( 
.A(n_5534),
.Y(n_5720)
);

INVx2_ASAP7_75t_L g5721 ( 
.A(n_5513),
.Y(n_5721)
);

INVx2_ASAP7_75t_L g5722 ( 
.A(n_5502),
.Y(n_5722)
);

NAND2xp5_ASAP7_75t_L g5723 ( 
.A(n_5602),
.B(n_5613),
.Y(n_5723)
);

INVx1_ASAP7_75t_L g5724 ( 
.A(n_5559),
.Y(n_5724)
);

INVx1_ASAP7_75t_L g5725 ( 
.A(n_5536),
.Y(n_5725)
);

INVx2_ASAP7_75t_L g5726 ( 
.A(n_5504),
.Y(n_5726)
);

AND2x2_ASAP7_75t_L g5727 ( 
.A(n_5457),
.B(n_392),
.Y(n_5727)
);

AND2x4_ASAP7_75t_L g5728 ( 
.A(n_5463),
.B(n_392),
.Y(n_5728)
);

BUFx4f_ASAP7_75t_L g5729 ( 
.A(n_5567),
.Y(n_5729)
);

OAI211xp5_ASAP7_75t_L g5730 ( 
.A1(n_5614),
.A2(n_395),
.B(n_393),
.C(n_394),
.Y(n_5730)
);

AND2x2_ASAP7_75t_L g5731 ( 
.A(n_5455),
.B(n_395),
.Y(n_5731)
);

OR2x2_ASAP7_75t_L g5732 ( 
.A(n_5493),
.B(n_5512),
.Y(n_5732)
);

AND2x2_ASAP7_75t_L g5733 ( 
.A(n_5487),
.B(n_396),
.Y(n_5733)
);

INVx2_ASAP7_75t_L g5734 ( 
.A(n_5523),
.Y(n_5734)
);

BUFx2_ASAP7_75t_L g5735 ( 
.A(n_5526),
.Y(n_5735)
);

INVx2_ASAP7_75t_L g5736 ( 
.A(n_5543),
.Y(n_5736)
);

OR2x2_ASAP7_75t_L g5737 ( 
.A(n_5461),
.B(n_396),
.Y(n_5737)
);

INVx1_ASAP7_75t_L g5738 ( 
.A(n_5515),
.Y(n_5738)
);

INVx1_ASAP7_75t_L g5739 ( 
.A(n_5537),
.Y(n_5739)
);

INVx2_ASAP7_75t_L g5740 ( 
.A(n_5540),
.Y(n_5740)
);

BUFx2_ASAP7_75t_L g5741 ( 
.A(n_5511),
.Y(n_5741)
);

HB1xp67_ASAP7_75t_L g5742 ( 
.A(n_5597),
.Y(n_5742)
);

AND2x4_ASAP7_75t_L g5743 ( 
.A(n_5541),
.B(n_5464),
.Y(n_5743)
);

AND2x2_ASAP7_75t_L g5744 ( 
.A(n_5560),
.B(n_397),
.Y(n_5744)
);

AND2x4_ASAP7_75t_L g5745 ( 
.A(n_5582),
.B(n_398),
.Y(n_5745)
);

INVx2_ASAP7_75t_L g5746 ( 
.A(n_5550),
.Y(n_5746)
);

INVx2_ASAP7_75t_L g5747 ( 
.A(n_5557),
.Y(n_5747)
);

NAND2xp5_ASAP7_75t_L g5748 ( 
.A(n_5547),
.B(n_399),
.Y(n_5748)
);

INVx2_ASAP7_75t_L g5749 ( 
.A(n_5553),
.Y(n_5749)
);

INVx2_ASAP7_75t_SL g5750 ( 
.A(n_5498),
.Y(n_5750)
);

INVx2_ASAP7_75t_L g5751 ( 
.A(n_5566),
.Y(n_5751)
);

OR2x2_ASAP7_75t_L g5752 ( 
.A(n_5575),
.B(n_399),
.Y(n_5752)
);

AND2x4_ASAP7_75t_L g5753 ( 
.A(n_5546),
.B(n_400),
.Y(n_5753)
);

INVx1_ASAP7_75t_L g5754 ( 
.A(n_5563),
.Y(n_5754)
);

INVx2_ASAP7_75t_L g5755 ( 
.A(n_5510),
.Y(n_5755)
);

NAND2xp5_ASAP7_75t_L g5756 ( 
.A(n_5584),
.B(n_5604),
.Y(n_5756)
);

INVx2_ASAP7_75t_L g5757 ( 
.A(n_5554),
.Y(n_5757)
);

BUFx2_ASAP7_75t_L g5758 ( 
.A(n_5517),
.Y(n_5758)
);

INVx2_ASAP7_75t_L g5759 ( 
.A(n_5491),
.Y(n_5759)
);

OR2x2_ASAP7_75t_L g5760 ( 
.A(n_5551),
.B(n_5589),
.Y(n_5760)
);

AND2x2_ASAP7_75t_L g5761 ( 
.A(n_5481),
.B(n_400),
.Y(n_5761)
);

INVx2_ASAP7_75t_L g5762 ( 
.A(n_5458),
.Y(n_5762)
);

OR2x2_ASAP7_75t_L g5763 ( 
.A(n_5544),
.B(n_402),
.Y(n_5763)
);

INVxp67_ASAP7_75t_L g5764 ( 
.A(n_5629),
.Y(n_5764)
);

BUFx3_ASAP7_75t_L g5765 ( 
.A(n_5591),
.Y(n_5765)
);

AND2x4_ASAP7_75t_L g5766 ( 
.A(n_5459),
.B(n_402),
.Y(n_5766)
);

INVx1_ASAP7_75t_L g5767 ( 
.A(n_5505),
.Y(n_5767)
);

NAND2xp5_ASAP7_75t_L g5768 ( 
.A(n_5516),
.B(n_403),
.Y(n_5768)
);

AND2x2_ASAP7_75t_L g5769 ( 
.A(n_5556),
.B(n_5471),
.Y(n_5769)
);

INVx1_ASAP7_75t_L g5770 ( 
.A(n_5520),
.Y(n_5770)
);

INVx1_ASAP7_75t_L g5771 ( 
.A(n_5524),
.Y(n_5771)
);

AO22x2_ASAP7_75t_L g5772 ( 
.A1(n_5514),
.A2(n_405),
.B1(n_403),
.B2(n_404),
.Y(n_5772)
);

AOI22xp33_ASAP7_75t_SL g5773 ( 
.A1(n_5555),
.A2(n_414),
.B1(n_423),
.B2(n_406),
.Y(n_5773)
);

HB1xp67_ASAP7_75t_L g5774 ( 
.A(n_5580),
.Y(n_5774)
);

AND2x2_ASAP7_75t_L g5775 ( 
.A(n_5564),
.B(n_5569),
.Y(n_5775)
);

AND2x2_ASAP7_75t_L g5776 ( 
.A(n_5585),
.B(n_406),
.Y(n_5776)
);

NAND2xp5_ASAP7_75t_L g5777 ( 
.A(n_5531),
.B(n_407),
.Y(n_5777)
);

AO21x2_ASAP7_75t_L g5778 ( 
.A1(n_5496),
.A2(n_408),
.B(n_409),
.Y(n_5778)
);

BUFx3_ASAP7_75t_L g5779 ( 
.A(n_5529),
.Y(n_5779)
);

INVx1_ASAP7_75t_L g5780 ( 
.A(n_5458),
.Y(n_5780)
);

BUFx3_ASAP7_75t_L g5781 ( 
.A(n_5489),
.Y(n_5781)
);

AND2x2_ASAP7_75t_L g5782 ( 
.A(n_5561),
.B(n_409),
.Y(n_5782)
);

AND2x2_ASAP7_75t_L g5783 ( 
.A(n_5538),
.B(n_410),
.Y(n_5783)
);

AND2x4_ASAP7_75t_L g5784 ( 
.A(n_5549),
.B(n_410),
.Y(n_5784)
);

NOR4xp25_ASAP7_75t_SL g5785 ( 
.A(n_5542),
.B(n_5549),
.C(n_5593),
.D(n_5562),
.Y(n_5785)
);

NAND2xp5_ASAP7_75t_L g5786 ( 
.A(n_5539),
.B(n_411),
.Y(n_5786)
);

AND2x2_ASAP7_75t_L g5787 ( 
.A(n_5533),
.B(n_412),
.Y(n_5787)
);

AND2x2_ASAP7_75t_L g5788 ( 
.A(n_5532),
.B(n_412),
.Y(n_5788)
);

HB1xp67_ASAP7_75t_L g5789 ( 
.A(n_5609),
.Y(n_5789)
);

AND2x2_ASAP7_75t_L g5790 ( 
.A(n_5603),
.B(n_413),
.Y(n_5790)
);

NAND2xp5_ASAP7_75t_L g5791 ( 
.A(n_5606),
.B(n_414),
.Y(n_5791)
);

INVx1_ASAP7_75t_L g5792 ( 
.A(n_5609),
.Y(n_5792)
);

INVx1_ASAP7_75t_L g5793 ( 
.A(n_5628),
.Y(n_5793)
);

BUFx2_ASAP7_75t_L g5794 ( 
.A(n_5615),
.Y(n_5794)
);

AND2x2_ASAP7_75t_L g5795 ( 
.A(n_5519),
.B(n_415),
.Y(n_5795)
);

OR2x2_ASAP7_75t_L g5796 ( 
.A(n_5594),
.B(n_415),
.Y(n_5796)
);

INVx2_ASAP7_75t_L g5797 ( 
.A(n_5587),
.Y(n_5797)
);

AOI22xp33_ASAP7_75t_SL g5798 ( 
.A1(n_5612),
.A2(n_426),
.B1(n_435),
.B2(n_416),
.Y(n_5798)
);

BUFx2_ASAP7_75t_L g5799 ( 
.A(n_5611),
.Y(n_5799)
);

HB1xp67_ASAP7_75t_L g5800 ( 
.A(n_5508),
.Y(n_5800)
);

INVx2_ASAP7_75t_L g5801 ( 
.A(n_5581),
.Y(n_5801)
);

INVx1_ASAP7_75t_L g5802 ( 
.A(n_5617),
.Y(n_5802)
);

AND2x2_ASAP7_75t_L g5803 ( 
.A(n_5500),
.B(n_416),
.Y(n_5803)
);

BUFx3_ASAP7_75t_L g5804 ( 
.A(n_5623),
.Y(n_5804)
);

INVx1_ASAP7_75t_L g5805 ( 
.A(n_5528),
.Y(n_5805)
);

BUFx2_ASAP7_75t_L g5806 ( 
.A(n_5451),
.Y(n_5806)
);

INVx1_ASAP7_75t_L g5807 ( 
.A(n_5528),
.Y(n_5807)
);

AOI21xp5_ASAP7_75t_L g5808 ( 
.A1(n_5596),
.A2(n_417),
.B(n_418),
.Y(n_5808)
);

INVx2_ASAP7_75t_L g5809 ( 
.A(n_5572),
.Y(n_5809)
);

AND2x2_ASAP7_75t_L g5810 ( 
.A(n_5577),
.B(n_417),
.Y(n_5810)
);

AND2x2_ASAP7_75t_L g5811 ( 
.A(n_5577),
.B(n_419),
.Y(n_5811)
);

AND2x2_ASAP7_75t_L g5812 ( 
.A(n_5577),
.B(n_419),
.Y(n_5812)
);

NAND2xp5_ASAP7_75t_L g5813 ( 
.A(n_5565),
.B(n_421),
.Y(n_5813)
);

INVx2_ASAP7_75t_L g5814 ( 
.A(n_5572),
.Y(n_5814)
);

INVx1_ASAP7_75t_L g5815 ( 
.A(n_5528),
.Y(n_5815)
);

INVxp67_ASAP7_75t_L g5816 ( 
.A(n_5596),
.Y(n_5816)
);

INVx2_ASAP7_75t_L g5817 ( 
.A(n_5572),
.Y(n_5817)
);

INVx2_ASAP7_75t_L g5818 ( 
.A(n_5572),
.Y(n_5818)
);

NAND2xp5_ASAP7_75t_L g5819 ( 
.A(n_5565),
.B(n_421),
.Y(n_5819)
);

AND2x2_ASAP7_75t_L g5820 ( 
.A(n_5577),
.B(n_422),
.Y(n_5820)
);

OR2x2_ASAP7_75t_L g5821 ( 
.A(n_5565),
.B(n_424),
.Y(n_5821)
);

AND2x2_ASAP7_75t_L g5822 ( 
.A(n_5577),
.B(n_424),
.Y(n_5822)
);

AND2x2_ASAP7_75t_L g5823 ( 
.A(n_5577),
.B(n_425),
.Y(n_5823)
);

OR2x2_ASAP7_75t_L g5824 ( 
.A(n_5565),
.B(n_426),
.Y(n_5824)
);

INVx2_ASAP7_75t_L g5825 ( 
.A(n_5572),
.Y(n_5825)
);

INVx2_ASAP7_75t_L g5826 ( 
.A(n_5572),
.Y(n_5826)
);

INVx1_ASAP7_75t_L g5827 ( 
.A(n_5528),
.Y(n_5827)
);

INVx2_ASAP7_75t_L g5828 ( 
.A(n_5572),
.Y(n_5828)
);

HB1xp67_ASAP7_75t_L g5829 ( 
.A(n_5592),
.Y(n_5829)
);

AND2x2_ASAP7_75t_L g5830 ( 
.A(n_5577),
.B(n_428),
.Y(n_5830)
);

INVx2_ASAP7_75t_L g5831 ( 
.A(n_5572),
.Y(n_5831)
);

INVx2_ASAP7_75t_L g5832 ( 
.A(n_5572),
.Y(n_5832)
);

INVx2_ASAP7_75t_L g5833 ( 
.A(n_5572),
.Y(n_5833)
);

INVx1_ASAP7_75t_L g5834 ( 
.A(n_5663),
.Y(n_5834)
);

INVx1_ASAP7_75t_L g5835 ( 
.A(n_5667),
.Y(n_5835)
);

INVx1_ASAP7_75t_L g5836 ( 
.A(n_5673),
.Y(n_5836)
);

AND2x2_ASAP7_75t_L g5837 ( 
.A(n_5681),
.B(n_429),
.Y(n_5837)
);

INVx2_ASAP7_75t_L g5838 ( 
.A(n_5654),
.Y(n_5838)
);

NAND2xp5_ASAP7_75t_L g5839 ( 
.A(n_5742),
.B(n_430),
.Y(n_5839)
);

NOR2xp33_ASAP7_75t_L g5840 ( 
.A(n_5676),
.B(n_431),
.Y(n_5840)
);

AND2x2_ASAP7_75t_L g5841 ( 
.A(n_5630),
.B(n_431),
.Y(n_5841)
);

AND2x2_ASAP7_75t_L g5842 ( 
.A(n_5816),
.B(n_432),
.Y(n_5842)
);

NAND2xp5_ASAP7_75t_L g5843 ( 
.A(n_5685),
.B(n_432),
.Y(n_5843)
);

AND2x2_ASAP7_75t_L g5844 ( 
.A(n_5741),
.B(n_433),
.Y(n_5844)
);

BUFx8_ASAP7_75t_L g5845 ( 
.A(n_5776),
.Y(n_5845)
);

INVx2_ASAP7_75t_L g5846 ( 
.A(n_5654),
.Y(n_5846)
);

AND2x4_ASAP7_75t_L g5847 ( 
.A(n_5649),
.B(n_433),
.Y(n_5847)
);

AND2x4_ASAP7_75t_L g5848 ( 
.A(n_5665),
.B(n_5643),
.Y(n_5848)
);

AND2x2_ASAP7_75t_L g5849 ( 
.A(n_5758),
.B(n_434),
.Y(n_5849)
);

INVx3_ASAP7_75t_L g5850 ( 
.A(n_5656),
.Y(n_5850)
);

NAND2xp5_ASAP7_75t_L g5851 ( 
.A(n_5652),
.B(n_434),
.Y(n_5851)
);

NOR2xp33_ASAP7_75t_L g5852 ( 
.A(n_5806),
.B(n_435),
.Y(n_5852)
);

AND2x4_ASAP7_75t_L g5853 ( 
.A(n_5735),
.B(n_436),
.Y(n_5853)
);

INVx2_ASAP7_75t_L g5854 ( 
.A(n_5631),
.Y(n_5854)
);

AND2x4_ASAP7_75t_L g5855 ( 
.A(n_5713),
.B(n_436),
.Y(n_5855)
);

OR2x2_ASAP7_75t_L g5856 ( 
.A(n_5648),
.B(n_438),
.Y(n_5856)
);

INVx1_ASAP7_75t_SL g5857 ( 
.A(n_5646),
.Y(n_5857)
);

AND2x2_ASAP7_75t_L g5858 ( 
.A(n_5775),
.B(n_439),
.Y(n_5858)
);

AND2x2_ASAP7_75t_L g5859 ( 
.A(n_5675),
.B(n_440),
.Y(n_5859)
);

AND2x4_ASAP7_75t_SL g5860 ( 
.A(n_5678),
.B(n_440),
.Y(n_5860)
);

AND2x2_ASAP7_75t_L g5861 ( 
.A(n_5716),
.B(n_442),
.Y(n_5861)
);

BUFx6f_ASAP7_75t_L g5862 ( 
.A(n_5729),
.Y(n_5862)
);

INVx2_ASAP7_75t_L g5863 ( 
.A(n_5809),
.Y(n_5863)
);

NOR2xp67_ASAP7_75t_L g5864 ( 
.A(n_5764),
.B(n_442),
.Y(n_5864)
);

INVx1_ASAP7_75t_L g5865 ( 
.A(n_5680),
.Y(n_5865)
);

BUFx3_ASAP7_75t_L g5866 ( 
.A(n_5753),
.Y(n_5866)
);

AND2x2_ASAP7_75t_L g5867 ( 
.A(n_5717),
.B(n_443),
.Y(n_5867)
);

INVx1_ASAP7_75t_L g5868 ( 
.A(n_5682),
.Y(n_5868)
);

AND2x2_ASAP7_75t_L g5869 ( 
.A(n_5769),
.B(n_5765),
.Y(n_5869)
);

AND2x4_ASAP7_75t_L g5870 ( 
.A(n_5779),
.B(n_445),
.Y(n_5870)
);

OR2x2_ASAP7_75t_L g5871 ( 
.A(n_5657),
.B(n_446),
.Y(n_5871)
);

INVx1_ASAP7_75t_L g5872 ( 
.A(n_5683),
.Y(n_5872)
);

INVx2_ASAP7_75t_L g5873 ( 
.A(n_5814),
.Y(n_5873)
);

INVx1_ASAP7_75t_L g5874 ( 
.A(n_5686),
.Y(n_5874)
);

AND2x2_ASAP7_75t_L g5875 ( 
.A(n_5674),
.B(n_447),
.Y(n_5875)
);

INVx2_ASAP7_75t_L g5876 ( 
.A(n_5817),
.Y(n_5876)
);

INVx1_ASAP7_75t_L g5877 ( 
.A(n_5687),
.Y(n_5877)
);

INVx2_ASAP7_75t_L g5878 ( 
.A(n_5818),
.Y(n_5878)
);

INVx1_ASAP7_75t_L g5879 ( 
.A(n_5693),
.Y(n_5879)
);

INVx1_ASAP7_75t_L g5880 ( 
.A(n_5694),
.Y(n_5880)
);

NAND3xp33_ASAP7_75t_L g5881 ( 
.A(n_5666),
.B(n_5774),
.C(n_5799),
.Y(n_5881)
);

INVx1_ASAP7_75t_L g5882 ( 
.A(n_5704),
.Y(n_5882)
);

INVx1_ASAP7_75t_L g5883 ( 
.A(n_5641),
.Y(n_5883)
);

INVx1_ASAP7_75t_L g5884 ( 
.A(n_5662),
.Y(n_5884)
);

AND2x2_ASAP7_75t_L g5885 ( 
.A(n_5645),
.B(n_448),
.Y(n_5885)
);

NAND2xp5_ASAP7_75t_L g5886 ( 
.A(n_5767),
.B(n_5770),
.Y(n_5886)
);

AND2x4_ASAP7_75t_L g5887 ( 
.A(n_5750),
.B(n_448),
.Y(n_5887)
);

AND2x2_ASAP7_75t_L g5888 ( 
.A(n_5757),
.B(n_449),
.Y(n_5888)
);

INVx2_ASAP7_75t_L g5889 ( 
.A(n_5825),
.Y(n_5889)
);

NAND2xp5_ASAP7_75t_L g5890 ( 
.A(n_5771),
.B(n_449),
.Y(n_5890)
);

AND2x2_ASAP7_75t_L g5891 ( 
.A(n_5636),
.B(n_450),
.Y(n_5891)
);

AND2x2_ASAP7_75t_L g5892 ( 
.A(n_5647),
.B(n_451),
.Y(n_5892)
);

AND2x2_ASAP7_75t_L g5893 ( 
.A(n_5805),
.B(n_451),
.Y(n_5893)
);

AOI22xp33_ASAP7_75t_L g5894 ( 
.A1(n_5797),
.A2(n_454),
.B1(n_452),
.B2(n_453),
.Y(n_5894)
);

INVx1_ASAP7_75t_L g5895 ( 
.A(n_5653),
.Y(n_5895)
);

INVx1_ASAP7_75t_L g5896 ( 
.A(n_5789),
.Y(n_5896)
);

INVx2_ASAP7_75t_L g5897 ( 
.A(n_5826),
.Y(n_5897)
);

INVx2_ASAP7_75t_L g5898 ( 
.A(n_5828),
.Y(n_5898)
);

AND2x2_ASAP7_75t_L g5899 ( 
.A(n_5807),
.B(n_452),
.Y(n_5899)
);

INVx2_ASAP7_75t_L g5900 ( 
.A(n_5831),
.Y(n_5900)
);

AND2x2_ASAP7_75t_L g5901 ( 
.A(n_5815),
.B(n_453),
.Y(n_5901)
);

INVx1_ASAP7_75t_L g5902 ( 
.A(n_5792),
.Y(n_5902)
);

INVxp67_ASAP7_75t_SL g5903 ( 
.A(n_5640),
.Y(n_5903)
);

INVx1_ASAP7_75t_L g5904 ( 
.A(n_5650),
.Y(n_5904)
);

NOR2x1_ASAP7_75t_R g5905 ( 
.A(n_5691),
.B(n_454),
.Y(n_5905)
);

INVx2_ASAP7_75t_L g5906 ( 
.A(n_5832),
.Y(n_5906)
);

INVx2_ASAP7_75t_L g5907 ( 
.A(n_5833),
.Y(n_5907)
);

OR2x2_ASAP7_75t_L g5908 ( 
.A(n_5760),
.B(n_455),
.Y(n_5908)
);

A2O1A1Ixp33_ASAP7_75t_L g5909 ( 
.A1(n_5730),
.A2(n_457),
.B(n_455),
.C(n_456),
.Y(n_5909)
);

OR2x6_ASAP7_75t_L g5910 ( 
.A(n_5659),
.B(n_456),
.Y(n_5910)
);

INVx1_ASAP7_75t_L g5911 ( 
.A(n_5723),
.Y(n_5911)
);

INVx3_ASAP7_75t_L g5912 ( 
.A(n_5718),
.Y(n_5912)
);

BUFx3_ASAP7_75t_L g5913 ( 
.A(n_5728),
.Y(n_5913)
);

INVx1_ASAP7_75t_L g5914 ( 
.A(n_5709),
.Y(n_5914)
);

OR2x2_ASAP7_75t_L g5915 ( 
.A(n_5827),
.B(n_457),
.Y(n_5915)
);

AND2x2_ASAP7_75t_L g5916 ( 
.A(n_5705),
.B(n_458),
.Y(n_5916)
);

OR2x2_ASAP7_75t_L g5917 ( 
.A(n_5829),
.B(n_458),
.Y(n_5917)
);

INVx1_ASAP7_75t_L g5918 ( 
.A(n_5712),
.Y(n_5918)
);

NAND2xp5_ASAP7_75t_L g5919 ( 
.A(n_5813),
.B(n_459),
.Y(n_5919)
);

AND2x4_ASAP7_75t_L g5920 ( 
.A(n_5759),
.B(n_459),
.Y(n_5920)
);

INVx2_ASAP7_75t_L g5921 ( 
.A(n_5634),
.Y(n_5921)
);

INVx3_ASAP7_75t_L g5922 ( 
.A(n_5718),
.Y(n_5922)
);

INVx2_ASAP7_75t_L g5923 ( 
.A(n_5762),
.Y(n_5923)
);

AND2x2_ASAP7_75t_L g5924 ( 
.A(n_5633),
.B(n_460),
.Y(n_5924)
);

AOI22xp33_ASAP7_75t_L g5925 ( 
.A1(n_5802),
.A2(n_464),
.B1(n_461),
.B2(n_463),
.Y(n_5925)
);

INVx2_ASAP7_75t_L g5926 ( 
.A(n_5696),
.Y(n_5926)
);

BUFx6f_ASAP7_75t_L g5927 ( 
.A(n_5784),
.Y(n_5927)
);

INVxp67_ASAP7_75t_L g5928 ( 
.A(n_5800),
.Y(n_5928)
);

INVx4_ASAP7_75t_L g5929 ( 
.A(n_5670),
.Y(n_5929)
);

AND2x2_ASAP7_75t_L g5930 ( 
.A(n_5810),
.B(n_5811),
.Y(n_5930)
);

INVx1_ASAP7_75t_L g5931 ( 
.A(n_5720),
.Y(n_5931)
);

NAND2xp5_ASAP7_75t_L g5932 ( 
.A(n_5819),
.B(n_464),
.Y(n_5932)
);

INVx1_ASAP7_75t_L g5933 ( 
.A(n_5724),
.Y(n_5933)
);

AND2x2_ASAP7_75t_L g5934 ( 
.A(n_5812),
.B(n_465),
.Y(n_5934)
);

AND2x2_ASAP7_75t_L g5935 ( 
.A(n_5820),
.B(n_465),
.Y(n_5935)
);

AND2x2_ASAP7_75t_L g5936 ( 
.A(n_5822),
.B(n_466),
.Y(n_5936)
);

INVx2_ASAP7_75t_L g5937 ( 
.A(n_5698),
.Y(n_5937)
);

INVx2_ASAP7_75t_L g5938 ( 
.A(n_5700),
.Y(n_5938)
);

INVx2_ASAP7_75t_SL g5939 ( 
.A(n_5637),
.Y(n_5939)
);

AND2x2_ASAP7_75t_SL g5940 ( 
.A(n_5794),
.B(n_466),
.Y(n_5940)
);

INVxp67_ASAP7_75t_SL g5941 ( 
.A(n_5708),
.Y(n_5941)
);

AND2x2_ASAP7_75t_L g5942 ( 
.A(n_5823),
.B(n_467),
.Y(n_5942)
);

INVxp67_ASAP7_75t_L g5943 ( 
.A(n_5664),
.Y(n_5943)
);

AND2x2_ASAP7_75t_L g5944 ( 
.A(n_5830),
.B(n_467),
.Y(n_5944)
);

NAND2xp5_ASAP7_75t_L g5945 ( 
.A(n_5672),
.B(n_468),
.Y(n_5945)
);

INVx1_ASAP7_75t_L g5946 ( 
.A(n_5780),
.Y(n_5946)
);

OR2x2_ASAP7_75t_L g5947 ( 
.A(n_5756),
.B(n_468),
.Y(n_5947)
);

AND2x2_ASAP7_75t_L g5948 ( 
.A(n_5638),
.B(n_469),
.Y(n_5948)
);

INVx2_ASAP7_75t_L g5949 ( 
.A(n_5722),
.Y(n_5949)
);

INVx2_ASAP7_75t_L g5950 ( 
.A(n_5751),
.Y(n_5950)
);

AND2x2_ASAP7_75t_L g5951 ( 
.A(n_5679),
.B(n_470),
.Y(n_5951)
);

INVx1_ASAP7_75t_L g5952 ( 
.A(n_5661),
.Y(n_5952)
);

OR2x2_ASAP7_75t_L g5953 ( 
.A(n_5677),
.B(n_471),
.Y(n_5953)
);

AND2x2_ASAP7_75t_L g5954 ( 
.A(n_5711),
.B(n_471),
.Y(n_5954)
);

AND2x4_ASAP7_75t_SL g5955 ( 
.A(n_5668),
.B(n_472),
.Y(n_5955)
);

INVx2_ASAP7_75t_L g5956 ( 
.A(n_5701),
.Y(n_5956)
);

AND2x4_ASAP7_75t_L g5957 ( 
.A(n_5743),
.B(n_5639),
.Y(n_5957)
);

HB1xp67_ASAP7_75t_L g5958 ( 
.A(n_5702),
.Y(n_5958)
);

INVx1_ASAP7_75t_L g5959 ( 
.A(n_5725),
.Y(n_5959)
);

NAND2xp5_ASAP7_75t_L g5960 ( 
.A(n_5669),
.B(n_473),
.Y(n_5960)
);

INVx2_ASAP7_75t_L g5961 ( 
.A(n_5707),
.Y(n_5961)
);

BUFx3_ASAP7_75t_L g5962 ( 
.A(n_5781),
.Y(n_5962)
);

INVx1_ASAP7_75t_L g5963 ( 
.A(n_5738),
.Y(n_5963)
);

OR2x2_ASAP7_75t_L g5964 ( 
.A(n_5632),
.B(n_474),
.Y(n_5964)
);

INVx1_ASAP7_75t_L g5965 ( 
.A(n_5739),
.Y(n_5965)
);

NOR2x1p5_ASAP7_75t_L g5966 ( 
.A(n_5786),
.B(n_475),
.Y(n_5966)
);

AND2x2_ASAP7_75t_L g5967 ( 
.A(n_5710),
.B(n_476),
.Y(n_5967)
);

AND2x4_ASAP7_75t_L g5968 ( 
.A(n_5745),
.B(n_477),
.Y(n_5968)
);

AND2x2_ASAP7_75t_L g5969 ( 
.A(n_5744),
.B(n_478),
.Y(n_5969)
);

INVx1_ASAP7_75t_L g5970 ( 
.A(n_5754),
.Y(n_5970)
);

NOR2xp33_ASAP7_75t_L g5971 ( 
.A(n_5763),
.B(n_479),
.Y(n_5971)
);

AND2x2_ASAP7_75t_L g5972 ( 
.A(n_5658),
.B(n_479),
.Y(n_5972)
);

INVx1_ASAP7_75t_L g5973 ( 
.A(n_5740),
.Y(n_5973)
);

AND2x2_ASAP7_75t_L g5974 ( 
.A(n_5642),
.B(n_480),
.Y(n_5974)
);

NAND2xp5_ASAP7_75t_L g5975 ( 
.A(n_5821),
.B(n_5824),
.Y(n_5975)
);

AND2x2_ASAP7_75t_L g5976 ( 
.A(n_5651),
.B(n_481),
.Y(n_5976)
);

INVx1_ASAP7_75t_L g5977 ( 
.A(n_5746),
.Y(n_5977)
);

INVx1_ASAP7_75t_L g5978 ( 
.A(n_5747),
.Y(n_5978)
);

INVx1_ASAP7_75t_L g5979 ( 
.A(n_5749),
.Y(n_5979)
);

AND2x4_ASAP7_75t_L g5980 ( 
.A(n_5766),
.B(n_482),
.Y(n_5980)
);

AND2x2_ASAP7_75t_L g5981 ( 
.A(n_5790),
.B(n_5783),
.Y(n_5981)
);

AND2x4_ASAP7_75t_L g5982 ( 
.A(n_5691),
.B(n_482),
.Y(n_5982)
);

INVx2_ASAP7_75t_L g5983 ( 
.A(n_5635),
.Y(n_5983)
);

NOR2xp67_ASAP7_75t_L g5984 ( 
.A(n_5752),
.B(n_483),
.Y(n_5984)
);

AND2x2_ASAP7_75t_L g5985 ( 
.A(n_5688),
.B(n_484),
.Y(n_5985)
);

AND2x2_ASAP7_75t_L g5986 ( 
.A(n_5689),
.B(n_485),
.Y(n_5986)
);

INVx1_ASAP7_75t_L g5987 ( 
.A(n_5697),
.Y(n_5987)
);

AND2x2_ASAP7_75t_L g5988 ( 
.A(n_5695),
.B(n_486),
.Y(n_5988)
);

AND2x2_ASAP7_75t_L g5989 ( 
.A(n_5684),
.B(n_486),
.Y(n_5989)
);

INVx1_ASAP7_75t_L g5990 ( 
.A(n_5732),
.Y(n_5990)
);

INVx1_ASAP7_75t_L g5991 ( 
.A(n_5793),
.Y(n_5991)
);

INVx1_ASAP7_75t_L g5992 ( 
.A(n_5721),
.Y(n_5992)
);

AND2x2_ASAP7_75t_L g5993 ( 
.A(n_5761),
.B(n_487),
.Y(n_5993)
);

NOR2xp33_ASAP7_75t_R g5994 ( 
.A(n_5791),
.B(n_488),
.Y(n_5994)
);

AND2x2_ASAP7_75t_L g5995 ( 
.A(n_5706),
.B(n_488),
.Y(n_5995)
);

INVxp67_ASAP7_75t_L g5996 ( 
.A(n_5778),
.Y(n_5996)
);

HB1xp67_ASAP7_75t_L g5997 ( 
.A(n_5715),
.Y(n_5997)
);

NAND2xp5_ASAP7_75t_SL g5998 ( 
.A(n_5755),
.B(n_490),
.Y(n_5998)
);

INVx1_ASAP7_75t_L g5999 ( 
.A(n_5737),
.Y(n_5999)
);

INVx1_ASAP7_75t_L g6000 ( 
.A(n_5801),
.Y(n_6000)
);

INVx2_ASAP7_75t_L g6001 ( 
.A(n_5644),
.Y(n_6001)
);

NAND2xp5_ASAP7_75t_L g6002 ( 
.A(n_5714),
.B(n_490),
.Y(n_6002)
);

NAND2xp5_ASAP7_75t_L g6003 ( 
.A(n_5719),
.B(n_491),
.Y(n_6003)
);

INVx1_ASAP7_75t_L g6004 ( 
.A(n_5655),
.Y(n_6004)
);

INVx2_ASAP7_75t_L g6005 ( 
.A(n_5660),
.Y(n_6005)
);

INVxp33_ASAP7_75t_L g6006 ( 
.A(n_5787),
.Y(n_6006)
);

INVx2_ASAP7_75t_L g6007 ( 
.A(n_5671),
.Y(n_6007)
);

INVx1_ASAP7_75t_L g6008 ( 
.A(n_5692),
.Y(n_6008)
);

AND2x2_ASAP7_75t_L g6009 ( 
.A(n_5727),
.B(n_492),
.Y(n_6009)
);

INVx3_ASAP7_75t_L g6010 ( 
.A(n_5788),
.Y(n_6010)
);

NOR2x1_ASAP7_75t_L g6011 ( 
.A(n_5703),
.B(n_5748),
.Y(n_6011)
);

NAND2xp5_ASAP7_75t_L g6012 ( 
.A(n_5768),
.B(n_492),
.Y(n_6012)
);

OR2x2_ASAP7_75t_L g6013 ( 
.A(n_5777),
.B(n_493),
.Y(n_6013)
);

INVx2_ASAP7_75t_L g6014 ( 
.A(n_5699),
.Y(n_6014)
);

AOI22xp33_ASAP7_75t_L g6015 ( 
.A1(n_5804),
.A2(n_495),
.B1(n_493),
.B2(n_494),
.Y(n_6015)
);

OR2x2_ASAP7_75t_L g6016 ( 
.A(n_5726),
.B(n_494),
.Y(n_6016)
);

INVx2_ASAP7_75t_L g6017 ( 
.A(n_5734),
.Y(n_6017)
);

INVx1_ASAP7_75t_L g6018 ( 
.A(n_5736),
.Y(n_6018)
);

INVx1_ASAP7_75t_L g6019 ( 
.A(n_5772),
.Y(n_6019)
);

HB1xp67_ASAP7_75t_L g6020 ( 
.A(n_5731),
.Y(n_6020)
);

INVx2_ASAP7_75t_L g6021 ( 
.A(n_5733),
.Y(n_6021)
);

INVx2_ASAP7_75t_L g6022 ( 
.A(n_5782),
.Y(n_6022)
);

INVx1_ASAP7_75t_L g6023 ( 
.A(n_5772),
.Y(n_6023)
);

AND2x2_ASAP7_75t_L g6024 ( 
.A(n_5785),
.B(n_495),
.Y(n_6024)
);

INVx2_ASAP7_75t_L g6025 ( 
.A(n_5796),
.Y(n_6025)
);

NOR2xp67_ASAP7_75t_L g6026 ( 
.A(n_5808),
.B(n_496),
.Y(n_6026)
);

BUFx2_ASAP7_75t_L g6027 ( 
.A(n_5795),
.Y(n_6027)
);

AND2x2_ASAP7_75t_L g6028 ( 
.A(n_5690),
.B(n_497),
.Y(n_6028)
);

INVx1_ASAP7_75t_L g6029 ( 
.A(n_5803),
.Y(n_6029)
);

AND2x4_ASAP7_75t_SL g6030 ( 
.A(n_5773),
.B(n_497),
.Y(n_6030)
);

INVx1_ASAP7_75t_L g6031 ( 
.A(n_5798),
.Y(n_6031)
);

INVx2_ASAP7_75t_L g6032 ( 
.A(n_5654),
.Y(n_6032)
);

OR2x2_ASAP7_75t_L g6033 ( 
.A(n_5685),
.B(n_498),
.Y(n_6033)
);

INVx2_ASAP7_75t_SL g6034 ( 
.A(n_5646),
.Y(n_6034)
);

OR2x2_ASAP7_75t_L g6035 ( 
.A(n_5685),
.B(n_499),
.Y(n_6035)
);

AND2x2_ASAP7_75t_L g6036 ( 
.A(n_5681),
.B(n_500),
.Y(n_6036)
);

NAND2xp5_ASAP7_75t_L g6037 ( 
.A(n_5742),
.B(n_501),
.Y(n_6037)
);

INVx1_ASAP7_75t_L g6038 ( 
.A(n_5663),
.Y(n_6038)
);

INVx2_ASAP7_75t_SL g6039 ( 
.A(n_5646),
.Y(n_6039)
);

AND2x2_ASAP7_75t_L g6040 ( 
.A(n_5681),
.B(n_501),
.Y(n_6040)
);

INVx1_ASAP7_75t_L g6041 ( 
.A(n_5663),
.Y(n_6041)
);

AND2x2_ASAP7_75t_L g6042 ( 
.A(n_5681),
.B(n_502),
.Y(n_6042)
);

INVx2_ASAP7_75t_L g6043 ( 
.A(n_5654),
.Y(n_6043)
);

INVx1_ASAP7_75t_L g6044 ( 
.A(n_5663),
.Y(n_6044)
);

OR2x2_ASAP7_75t_L g6045 ( 
.A(n_5685),
.B(n_502),
.Y(n_6045)
);

OR2x6_ASAP7_75t_L g6046 ( 
.A(n_5649),
.B(n_503),
.Y(n_6046)
);

INVx1_ASAP7_75t_L g6047 ( 
.A(n_5663),
.Y(n_6047)
);

INVx2_ASAP7_75t_L g6048 ( 
.A(n_5654),
.Y(n_6048)
);

INVx2_ASAP7_75t_SL g6049 ( 
.A(n_5646),
.Y(n_6049)
);

INVx2_ASAP7_75t_L g6050 ( 
.A(n_5654),
.Y(n_6050)
);

INVx1_ASAP7_75t_L g6051 ( 
.A(n_5663),
.Y(n_6051)
);

INVx2_ASAP7_75t_L g6052 ( 
.A(n_5654),
.Y(n_6052)
);

INVx1_ASAP7_75t_L g6053 ( 
.A(n_5663),
.Y(n_6053)
);

NAND2x1p5_ASAP7_75t_L g6054 ( 
.A(n_5691),
.B(n_504),
.Y(n_6054)
);

NAND3xp33_ASAP7_75t_L g6055 ( 
.A(n_5666),
.B(n_504),
.C(n_505),
.Y(n_6055)
);

INVx2_ASAP7_75t_L g6056 ( 
.A(n_5654),
.Y(n_6056)
);

INVxp67_ASAP7_75t_SL g6057 ( 
.A(n_5774),
.Y(n_6057)
);

INVx2_ASAP7_75t_L g6058 ( 
.A(n_5654),
.Y(n_6058)
);

OR2x2_ASAP7_75t_L g6059 ( 
.A(n_5685),
.B(n_505),
.Y(n_6059)
);

INVxp67_ASAP7_75t_L g6060 ( 
.A(n_5681),
.Y(n_6060)
);

INVx1_ASAP7_75t_L g6061 ( 
.A(n_5663),
.Y(n_6061)
);

NAND2xp5_ASAP7_75t_L g6062 ( 
.A(n_5742),
.B(n_506),
.Y(n_6062)
);

NAND2xp5_ASAP7_75t_L g6063 ( 
.A(n_5742),
.B(n_506),
.Y(n_6063)
);

INVx1_ASAP7_75t_L g6064 ( 
.A(n_5663),
.Y(n_6064)
);

INVx1_ASAP7_75t_L g6065 ( 
.A(n_5663),
.Y(n_6065)
);

AND2x2_ASAP7_75t_L g6066 ( 
.A(n_5681),
.B(n_507),
.Y(n_6066)
);

INVx2_ASAP7_75t_L g6067 ( 
.A(n_5654),
.Y(n_6067)
);

AND2x2_ASAP7_75t_L g6068 ( 
.A(n_5681),
.B(n_508),
.Y(n_6068)
);

AND2x2_ASAP7_75t_L g6069 ( 
.A(n_5681),
.B(n_508),
.Y(n_6069)
);

NAND2xp5_ASAP7_75t_L g6070 ( 
.A(n_5742),
.B(n_509),
.Y(n_6070)
);

AND2x2_ASAP7_75t_L g6071 ( 
.A(n_5681),
.B(n_510),
.Y(n_6071)
);

AND2x2_ASAP7_75t_L g6072 ( 
.A(n_5681),
.B(n_511),
.Y(n_6072)
);

AND2x2_ASAP7_75t_L g6073 ( 
.A(n_5681),
.B(n_512),
.Y(n_6073)
);

AND2x4_ASAP7_75t_L g6074 ( 
.A(n_5649),
.B(n_512),
.Y(n_6074)
);

BUFx2_ASAP7_75t_L g6075 ( 
.A(n_5646),
.Y(n_6075)
);

NAND2xp5_ASAP7_75t_L g6076 ( 
.A(n_5742),
.B(n_513),
.Y(n_6076)
);

AND2x2_ASAP7_75t_L g6077 ( 
.A(n_5681),
.B(n_513),
.Y(n_6077)
);

NAND2xp5_ASAP7_75t_L g6078 ( 
.A(n_5742),
.B(n_514),
.Y(n_6078)
);

HB1xp67_ASAP7_75t_L g6079 ( 
.A(n_5657),
.Y(n_6079)
);

AND2x2_ASAP7_75t_L g6080 ( 
.A(n_5681),
.B(n_514),
.Y(n_6080)
);

AND2x2_ASAP7_75t_L g6081 ( 
.A(n_5681),
.B(n_515),
.Y(n_6081)
);

INVx1_ASAP7_75t_L g6082 ( 
.A(n_5663),
.Y(n_6082)
);

NAND3xp33_ASAP7_75t_L g6083 ( 
.A(n_5666),
.B(n_516),
.C(n_517),
.Y(n_6083)
);

INVx2_ASAP7_75t_L g6084 ( 
.A(n_5654),
.Y(n_6084)
);

AND2x2_ASAP7_75t_L g6085 ( 
.A(n_5681),
.B(n_516),
.Y(n_6085)
);

AND2x2_ASAP7_75t_L g6086 ( 
.A(n_5681),
.B(n_518),
.Y(n_6086)
);

AND2x2_ASAP7_75t_L g6087 ( 
.A(n_5681),
.B(n_518),
.Y(n_6087)
);

AND2x2_ASAP7_75t_L g6088 ( 
.A(n_5681),
.B(n_519),
.Y(n_6088)
);

INVxp67_ASAP7_75t_L g6089 ( 
.A(n_5681),
.Y(n_6089)
);

INVxp67_ASAP7_75t_SL g6090 ( 
.A(n_5774),
.Y(n_6090)
);

NAND2xp5_ASAP7_75t_L g6091 ( 
.A(n_5742),
.B(n_519),
.Y(n_6091)
);

NAND2xp5_ASAP7_75t_L g6092 ( 
.A(n_5742),
.B(n_521),
.Y(n_6092)
);

INVx1_ASAP7_75t_L g6093 ( 
.A(n_5663),
.Y(n_6093)
);

OA21x2_ASAP7_75t_L g6094 ( 
.A1(n_5881),
.A2(n_521),
.B(n_522),
.Y(n_6094)
);

AOI22xp33_ASAP7_75t_L g6095 ( 
.A1(n_5928),
.A2(n_525),
.B1(n_522),
.B2(n_523),
.Y(n_6095)
);

INVx2_ASAP7_75t_L g6096 ( 
.A(n_6010),
.Y(n_6096)
);

OA21x2_ASAP7_75t_L g6097 ( 
.A1(n_5996),
.A2(n_525),
.B(n_527),
.Y(n_6097)
);

BUFx3_ASAP7_75t_L g6098 ( 
.A(n_5862),
.Y(n_6098)
);

INVx4_ASAP7_75t_L g6099 ( 
.A(n_6046),
.Y(n_6099)
);

INVx1_ASAP7_75t_L g6100 ( 
.A(n_5896),
.Y(n_6100)
);

AOI22xp33_ASAP7_75t_L g6101 ( 
.A1(n_6025),
.A2(n_6000),
.B1(n_5846),
.B2(n_5838),
.Y(n_6101)
);

NAND4xp25_ASAP7_75t_L g6102 ( 
.A(n_6060),
.B(n_529),
.C(n_527),
.D(n_528),
.Y(n_6102)
);

OAI21x1_ASAP7_75t_L g6103 ( 
.A1(n_5850),
.A2(n_528),
.B(n_529),
.Y(n_6103)
);

INVx1_ASAP7_75t_L g6104 ( 
.A(n_5946),
.Y(n_6104)
);

INVx2_ASAP7_75t_L g6105 ( 
.A(n_5869),
.Y(n_6105)
);

INVx1_ASAP7_75t_L g6106 ( 
.A(n_5886),
.Y(n_6106)
);

AND2x4_ASAP7_75t_L g6107 ( 
.A(n_5962),
.B(n_530),
.Y(n_6107)
);

AND2x4_ASAP7_75t_L g6108 ( 
.A(n_5957),
.B(n_530),
.Y(n_6108)
);

HB1xp67_ASAP7_75t_L g6109 ( 
.A(n_6020),
.Y(n_6109)
);

AND2x2_ASAP7_75t_L g6110 ( 
.A(n_5848),
.B(n_531),
.Y(n_6110)
);

OAI22xp33_ASAP7_75t_L g6111 ( 
.A1(n_6027),
.A2(n_6090),
.B1(n_6057),
.B2(n_6006),
.Y(n_6111)
);

AO21x2_ASAP7_75t_L g6112 ( 
.A1(n_5851),
.A2(n_532),
.B(n_533),
.Y(n_6112)
);

INVx1_ASAP7_75t_L g6113 ( 
.A(n_5902),
.Y(n_6113)
);

AO21x2_ASAP7_75t_L g6114 ( 
.A1(n_5843),
.A2(n_532),
.B(n_534),
.Y(n_6114)
);

OAI31xp33_ASAP7_75t_L g6115 ( 
.A1(n_6024),
.A2(n_536),
.A3(n_534),
.B(n_535),
.Y(n_6115)
);

INVx1_ASAP7_75t_L g6116 ( 
.A(n_5990),
.Y(n_6116)
);

INVx1_ASAP7_75t_L g6117 ( 
.A(n_5834),
.Y(n_6117)
);

AND2x2_ASAP7_75t_L g6118 ( 
.A(n_5981),
.B(n_535),
.Y(n_6118)
);

HB1xp67_ASAP7_75t_L g6119 ( 
.A(n_6089),
.Y(n_6119)
);

INVx3_ASAP7_75t_L g6120 ( 
.A(n_5866),
.Y(n_6120)
);

INVx1_ASAP7_75t_L g6121 ( 
.A(n_5835),
.Y(n_6121)
);

INVx2_ASAP7_75t_L g6122 ( 
.A(n_6022),
.Y(n_6122)
);

INVx2_ASAP7_75t_SL g6123 ( 
.A(n_5845),
.Y(n_6123)
);

AOI221xp5_ASAP7_75t_L g6124 ( 
.A1(n_6019),
.A2(n_538),
.B1(n_536),
.B2(n_537),
.C(n_539),
.Y(n_6124)
);

BUFx3_ASAP7_75t_L g6125 ( 
.A(n_5862),
.Y(n_6125)
);

INVx1_ASAP7_75t_L g6126 ( 
.A(n_5836),
.Y(n_6126)
);

OA21x2_ASAP7_75t_L g6127 ( 
.A1(n_5943),
.A2(n_5941),
.B(n_6023),
.Y(n_6127)
);

AO21x2_ASAP7_75t_L g6128 ( 
.A1(n_5839),
.A2(n_537),
.B(n_538),
.Y(n_6128)
);

AOI21x1_ASAP7_75t_L g6129 ( 
.A1(n_5864),
.A2(n_6075),
.B(n_5989),
.Y(n_6129)
);

INVx1_ASAP7_75t_L g6130 ( 
.A(n_5865),
.Y(n_6130)
);

OR2x2_ASAP7_75t_L g6131 ( 
.A(n_5997),
.B(n_539),
.Y(n_6131)
);

INVx2_ASAP7_75t_L g6132 ( 
.A(n_6016),
.Y(n_6132)
);

INVx1_ASAP7_75t_L g6133 ( 
.A(n_5868),
.Y(n_6133)
);

INVxp67_ASAP7_75t_SL g6134 ( 
.A(n_5905),
.Y(n_6134)
);

AND2x2_ASAP7_75t_L g6135 ( 
.A(n_5929),
.B(n_5912),
.Y(n_6135)
);

INVx1_ASAP7_75t_L g6136 ( 
.A(n_5872),
.Y(n_6136)
);

OR2x2_ASAP7_75t_L g6137 ( 
.A(n_5963),
.B(n_540),
.Y(n_6137)
);

INVx2_ASAP7_75t_L g6138 ( 
.A(n_6021),
.Y(n_6138)
);

AOI22xp33_ASAP7_75t_L g6139 ( 
.A1(n_6032),
.A2(n_542),
.B1(n_540),
.B2(n_541),
.Y(n_6139)
);

NAND2xp5_ASAP7_75t_SL g6140 ( 
.A(n_6034),
.B(n_541),
.Y(n_6140)
);

AOI22xp33_ASAP7_75t_L g6141 ( 
.A1(n_6043),
.A2(n_546),
.B1(n_543),
.B2(n_544),
.Y(n_6141)
);

INVx2_ASAP7_75t_L g6142 ( 
.A(n_5930),
.Y(n_6142)
);

AOI21xp5_ASAP7_75t_L g6143 ( 
.A1(n_5940),
.A2(n_543),
.B(n_544),
.Y(n_6143)
);

INVx1_ASAP7_75t_L g6144 ( 
.A(n_5874),
.Y(n_6144)
);

AOI22xp33_ASAP7_75t_L g6145 ( 
.A1(n_6048),
.A2(n_548),
.B1(n_546),
.B2(n_547),
.Y(n_6145)
);

INVx2_ASAP7_75t_L g6146 ( 
.A(n_5908),
.Y(n_6146)
);

INVx1_ASAP7_75t_L g6147 ( 
.A(n_5877),
.Y(n_6147)
);

NAND2xp5_ASAP7_75t_L g6148 ( 
.A(n_5958),
.B(n_547),
.Y(n_6148)
);

OAI31xp33_ASAP7_75t_L g6149 ( 
.A1(n_5966),
.A2(n_552),
.A3(n_548),
.B(n_549),
.Y(n_6149)
);

NAND2x1p5_ASAP7_75t_L g6150 ( 
.A(n_5982),
.B(n_549),
.Y(n_6150)
);

OR2x2_ASAP7_75t_L g6151 ( 
.A(n_5965),
.B(n_553),
.Y(n_6151)
);

INVx2_ASAP7_75t_L g6152 ( 
.A(n_6050),
.Y(n_6152)
);

NOR2x1_ASAP7_75t_L g6153 ( 
.A(n_6046),
.B(n_554),
.Y(n_6153)
);

AND2x2_ASAP7_75t_L g6154 ( 
.A(n_5922),
.B(n_556),
.Y(n_6154)
);

AND2x2_ASAP7_75t_L g6155 ( 
.A(n_5858),
.B(n_5891),
.Y(n_6155)
);

AND2x4_ASAP7_75t_L g6156 ( 
.A(n_5913),
.B(n_557),
.Y(n_6156)
);

AOI22xp33_ASAP7_75t_L g6157 ( 
.A1(n_6052),
.A2(n_559),
.B1(n_557),
.B2(n_558),
.Y(n_6157)
);

AND2x2_ASAP7_75t_L g6158 ( 
.A(n_5892),
.B(n_559),
.Y(n_6158)
);

OAI21xp33_ASAP7_75t_L g6159 ( 
.A1(n_5952),
.A2(n_560),
.B(n_561),
.Y(n_6159)
);

INVx1_ASAP7_75t_L g6160 ( 
.A(n_5879),
.Y(n_6160)
);

HB1xp67_ASAP7_75t_L g6161 ( 
.A(n_6079),
.Y(n_6161)
);

AOI21x1_ASAP7_75t_L g6162 ( 
.A1(n_5837),
.A2(n_6040),
.B(n_6036),
.Y(n_6162)
);

INVx1_ASAP7_75t_L g6163 ( 
.A(n_5880),
.Y(n_6163)
);

BUFx3_ASAP7_75t_L g6164 ( 
.A(n_5955),
.Y(n_6164)
);

NAND2xp5_ASAP7_75t_L g6165 ( 
.A(n_5916),
.B(n_560),
.Y(n_6165)
);

AOI221xp5_ASAP7_75t_L g6166 ( 
.A1(n_6056),
.A2(n_563),
.B1(n_561),
.B2(n_562),
.C(n_564),
.Y(n_6166)
);

INVx2_ASAP7_75t_L g6167 ( 
.A(n_6058),
.Y(n_6167)
);

NOR2xp33_ASAP7_75t_L g6168 ( 
.A(n_5857),
.B(n_565),
.Y(n_6168)
);

INVx1_ASAP7_75t_L g6169 ( 
.A(n_5882),
.Y(n_6169)
);

INVx2_ASAP7_75t_SL g6170 ( 
.A(n_6039),
.Y(n_6170)
);

AOI33xp33_ASAP7_75t_L g6171 ( 
.A1(n_6028),
.A2(n_568),
.A3(n_570),
.B1(n_566),
.B2(n_567),
.B3(n_569),
.Y(n_6171)
);

NAND3xp33_ASAP7_75t_L g6172 ( 
.A(n_6055),
.B(n_567),
.C(n_568),
.Y(n_6172)
);

AOI31xp33_ASAP7_75t_L g6173 ( 
.A1(n_6049),
.A2(n_578),
.A3(n_587),
.B(n_569),
.Y(n_6173)
);

INVxp67_ASAP7_75t_SL g6174 ( 
.A(n_6011),
.Y(n_6174)
);

NAND2xp5_ASAP7_75t_L g6175 ( 
.A(n_5841),
.B(n_570),
.Y(n_6175)
);

INVx1_ASAP7_75t_L g6176 ( 
.A(n_5883),
.Y(n_6176)
);

INVx2_ASAP7_75t_SL g6177 ( 
.A(n_5853),
.Y(n_6177)
);

AOI22xp33_ASAP7_75t_L g6178 ( 
.A1(n_6067),
.A2(n_573),
.B1(n_571),
.B2(n_572),
.Y(n_6178)
);

INVx2_ASAP7_75t_L g6179 ( 
.A(n_6084),
.Y(n_6179)
);

OAI221xp5_ASAP7_75t_SL g6180 ( 
.A1(n_6083),
.A2(n_575),
.B1(n_571),
.B2(n_573),
.C(n_576),
.Y(n_6180)
);

NAND2xp5_ASAP7_75t_L g6181 ( 
.A(n_5903),
.B(n_576),
.Y(n_6181)
);

INVx2_ASAP7_75t_L g6182 ( 
.A(n_5999),
.Y(n_6182)
);

INVx1_ASAP7_75t_L g6183 ( 
.A(n_5884),
.Y(n_6183)
);

OAI22xp33_ASAP7_75t_L g6184 ( 
.A1(n_6026),
.A2(n_586),
.B1(n_594),
.B2(n_577),
.Y(n_6184)
);

BUFx3_ASAP7_75t_L g6185 ( 
.A(n_5980),
.Y(n_6185)
);

INVx2_ASAP7_75t_L g6186 ( 
.A(n_5923),
.Y(n_6186)
);

BUFx2_ASAP7_75t_L g6187 ( 
.A(n_5910),
.Y(n_6187)
);

INVxp67_ASAP7_75t_L g6188 ( 
.A(n_5947),
.Y(n_6188)
);

AOI221xp5_ASAP7_75t_L g6189 ( 
.A1(n_6031),
.A2(n_579),
.B1(n_577),
.B2(n_578),
.C(n_580),
.Y(n_6189)
);

INVx1_ASAP7_75t_L g6190 ( 
.A(n_5895),
.Y(n_6190)
);

AND2x2_ASAP7_75t_L g6191 ( 
.A(n_5893),
.B(n_580),
.Y(n_6191)
);

NAND4xp25_ASAP7_75t_L g6192 ( 
.A(n_5840),
.B(n_584),
.C(n_581),
.D(n_583),
.Y(n_6192)
);

AND2x2_ASAP7_75t_L g6193 ( 
.A(n_5899),
.B(n_5901),
.Y(n_6193)
);

INVx2_ASAP7_75t_L g6194 ( 
.A(n_5854),
.Y(n_6194)
);

AOI22xp33_ASAP7_75t_L g6195 ( 
.A1(n_5863),
.A2(n_587),
.B1(n_585),
.B2(n_586),
.Y(n_6195)
);

AND2x4_ASAP7_75t_SL g6196 ( 
.A(n_5910),
.B(n_588),
.Y(n_6196)
);

AND2x4_ASAP7_75t_L g6197 ( 
.A(n_5939),
.B(n_588),
.Y(n_6197)
);

INVx1_ASAP7_75t_L g6198 ( 
.A(n_5904),
.Y(n_6198)
);

AND2x2_ASAP7_75t_L g6199 ( 
.A(n_5859),
.B(n_6042),
.Y(n_6199)
);

OAI21x1_ASAP7_75t_L g6200 ( 
.A1(n_5873),
.A2(n_589),
.B(n_590),
.Y(n_6200)
);

INVx2_ASAP7_75t_L g6201 ( 
.A(n_5876),
.Y(n_6201)
);

INVx2_ASAP7_75t_L g6202 ( 
.A(n_5878),
.Y(n_6202)
);

INVx3_ASAP7_75t_L g6203 ( 
.A(n_5927),
.Y(n_6203)
);

OAI322xp33_ASAP7_75t_L g6204 ( 
.A1(n_5856),
.A2(n_595),
.A3(n_594),
.B1(n_592),
.B2(n_589),
.C1(n_591),
.C2(n_593),
.Y(n_6204)
);

CKINVDCx20_ASAP7_75t_R g6205 ( 
.A(n_5994),
.Y(n_6205)
);

AND2x2_ASAP7_75t_L g6206 ( 
.A(n_6066),
.B(n_591),
.Y(n_6206)
);

NAND2xp5_ASAP7_75t_L g6207 ( 
.A(n_5987),
.B(n_593),
.Y(n_6207)
);

INVx2_ASAP7_75t_L g6208 ( 
.A(n_5889),
.Y(n_6208)
);

INVx3_ASAP7_75t_L g6209 ( 
.A(n_5927),
.Y(n_6209)
);

BUFx3_ASAP7_75t_L g6210 ( 
.A(n_5968),
.Y(n_6210)
);

NAND2xp5_ASAP7_75t_L g6211 ( 
.A(n_5911),
.B(n_595),
.Y(n_6211)
);

OAI31xp33_ASAP7_75t_L g6212 ( 
.A1(n_5909),
.A2(n_598),
.A3(n_596),
.B(n_597),
.Y(n_6212)
);

INVx2_ASAP7_75t_L g6213 ( 
.A(n_5897),
.Y(n_6213)
);

INVx2_ASAP7_75t_L g6214 ( 
.A(n_5898),
.Y(n_6214)
);

OA21x2_ASAP7_75t_L g6215 ( 
.A1(n_5900),
.A2(n_598),
.B(n_599),
.Y(n_6215)
);

INVx2_ASAP7_75t_L g6216 ( 
.A(n_5906),
.Y(n_6216)
);

INVx2_ASAP7_75t_L g6217 ( 
.A(n_5907),
.Y(n_6217)
);

AOI22xp33_ASAP7_75t_L g6218 ( 
.A1(n_6029),
.A2(n_602),
.B1(n_600),
.B2(n_601),
.Y(n_6218)
);

NAND3xp33_ASAP7_75t_L g6219 ( 
.A(n_6015),
.B(n_600),
.C(n_601),
.Y(n_6219)
);

AOI21xp33_ASAP7_75t_L g6220 ( 
.A1(n_5970),
.A2(n_602),
.B(n_603),
.Y(n_6220)
);

INVx1_ASAP7_75t_L g6221 ( 
.A(n_6038),
.Y(n_6221)
);

INVx2_ASAP7_75t_L g6222 ( 
.A(n_5950),
.Y(n_6222)
);

AND2x2_ASAP7_75t_L g6223 ( 
.A(n_6068),
.B(n_603),
.Y(n_6223)
);

INVx2_ASAP7_75t_L g6224 ( 
.A(n_6054),
.Y(n_6224)
);

OAI211xp5_ASAP7_75t_L g6225 ( 
.A1(n_5852),
.A2(n_606),
.B(n_604),
.C(n_605),
.Y(n_6225)
);

HB1xp67_ASAP7_75t_L g6226 ( 
.A(n_6041),
.Y(n_6226)
);

NOR2xp33_ASAP7_75t_L g6227 ( 
.A(n_5975),
.B(n_604),
.Y(n_6227)
);

INVx4_ASAP7_75t_L g6228 ( 
.A(n_5875),
.Y(n_6228)
);

INVx2_ASAP7_75t_SL g6229 ( 
.A(n_5860),
.Y(n_6229)
);

BUFx3_ASAP7_75t_L g6230 ( 
.A(n_5847),
.Y(n_6230)
);

BUFx2_ASAP7_75t_L g6231 ( 
.A(n_6069),
.Y(n_6231)
);

HB1xp67_ASAP7_75t_L g6232 ( 
.A(n_6044),
.Y(n_6232)
);

AND2x2_ASAP7_75t_L g6233 ( 
.A(n_6071),
.B(n_605),
.Y(n_6233)
);

INVx1_ASAP7_75t_L g6234 ( 
.A(n_6047),
.Y(n_6234)
);

BUFx3_ASAP7_75t_L g6235 ( 
.A(n_6074),
.Y(n_6235)
);

HB1xp67_ASAP7_75t_L g6236 ( 
.A(n_6051),
.Y(n_6236)
);

BUFx3_ASAP7_75t_L g6237 ( 
.A(n_5993),
.Y(n_6237)
);

OAI221xp5_ASAP7_75t_L g6238 ( 
.A1(n_5894),
.A2(n_609),
.B1(n_607),
.B2(n_608),
.C(n_610),
.Y(n_6238)
);

AND2x2_ASAP7_75t_L g6239 ( 
.A(n_6072),
.B(n_607),
.Y(n_6239)
);

BUFx2_ASAP7_75t_L g6240 ( 
.A(n_6073),
.Y(n_6240)
);

INVx1_ASAP7_75t_L g6241 ( 
.A(n_6053),
.Y(n_6241)
);

BUFx2_ASAP7_75t_L g6242 ( 
.A(n_6077),
.Y(n_6242)
);

INVx2_ASAP7_75t_L g6243 ( 
.A(n_5983),
.Y(n_6243)
);

INVx1_ASAP7_75t_L g6244 ( 
.A(n_6061),
.Y(n_6244)
);

OAI21x1_ASAP7_75t_L g6245 ( 
.A1(n_5921),
.A2(n_609),
.B(n_611),
.Y(n_6245)
);

BUFx3_ASAP7_75t_L g6246 ( 
.A(n_5995),
.Y(n_6246)
);

AOI221xp5_ASAP7_75t_L g6247 ( 
.A1(n_5971),
.A2(n_613),
.B1(n_611),
.B2(n_612),
.C(n_614),
.Y(n_6247)
);

INVx1_ASAP7_75t_SL g6248 ( 
.A(n_5967),
.Y(n_6248)
);

AOI221xp5_ASAP7_75t_L g6249 ( 
.A1(n_5890),
.A2(n_615),
.B1(n_612),
.B2(n_614),
.C(n_617),
.Y(n_6249)
);

INVx1_ASAP7_75t_L g6250 ( 
.A(n_6064),
.Y(n_6250)
);

AND2x4_ASAP7_75t_L g6251 ( 
.A(n_5870),
.B(n_615),
.Y(n_6251)
);

OAI21x1_ASAP7_75t_L g6252 ( 
.A1(n_5938),
.A2(n_617),
.B(n_618),
.Y(n_6252)
);

AO21x2_ASAP7_75t_L g6253 ( 
.A1(n_6037),
.A2(n_618),
.B(n_619),
.Y(n_6253)
);

BUFx6f_ASAP7_75t_L g6254 ( 
.A(n_5844),
.Y(n_6254)
);

AOI222xp33_ASAP7_75t_L g6255 ( 
.A1(n_5984),
.A2(n_647),
.B1(n_627),
.B2(n_655),
.C1(n_638),
.C2(n_619),
.Y(n_6255)
);

OAI221xp5_ASAP7_75t_L g6256 ( 
.A1(n_5925),
.A2(n_622),
.B1(n_620),
.B2(n_621),
.C(n_623),
.Y(n_6256)
);

OR2x2_ASAP7_75t_L g6257 ( 
.A(n_5991),
.B(n_622),
.Y(n_6257)
);

INVx2_ASAP7_75t_L g6258 ( 
.A(n_6001),
.Y(n_6258)
);

INVx2_ASAP7_75t_L g6259 ( 
.A(n_6005),
.Y(n_6259)
);

NAND4xp25_ASAP7_75t_L g6260 ( 
.A(n_6080),
.B(n_625),
.C(n_623),
.D(n_624),
.Y(n_6260)
);

INVx2_ASAP7_75t_L g6261 ( 
.A(n_6007),
.Y(n_6261)
);

AOI22xp5_ASAP7_75t_L g6262 ( 
.A1(n_6030),
.A2(n_627),
.B1(n_625),
.B2(n_626),
.Y(n_6262)
);

OAI221xp5_ASAP7_75t_L g6263 ( 
.A1(n_5973),
.A2(n_630),
.B1(n_628),
.B2(n_629),
.C(n_631),
.Y(n_6263)
);

AND2x2_ASAP7_75t_L g6264 ( 
.A(n_6081),
.B(n_630),
.Y(n_6264)
);

BUFx2_ASAP7_75t_L g6265 ( 
.A(n_6085),
.Y(n_6265)
);

OAI21x1_ASAP7_75t_L g6266 ( 
.A1(n_5926),
.A2(n_631),
.B(n_632),
.Y(n_6266)
);

OAI211xp5_ASAP7_75t_SL g6267 ( 
.A1(n_6002),
.A2(n_636),
.B(n_632),
.C(n_635),
.Y(n_6267)
);

INVx1_ASAP7_75t_L g6268 ( 
.A(n_6065),
.Y(n_6268)
);

INVx2_ASAP7_75t_L g6269 ( 
.A(n_6014),
.Y(n_6269)
);

INVx1_ASAP7_75t_L g6270 ( 
.A(n_6082),
.Y(n_6270)
);

OAI221xp5_ASAP7_75t_L g6271 ( 
.A1(n_5977),
.A2(n_640),
.B1(n_638),
.B2(n_639),
.C(n_641),
.Y(n_6271)
);

INVx2_ASAP7_75t_L g6272 ( 
.A(n_6017),
.Y(n_6272)
);

AOI21xp33_ASAP7_75t_SL g6273 ( 
.A1(n_6086),
.A2(n_651),
.B(n_641),
.Y(n_6273)
);

AND2x2_ASAP7_75t_L g6274 ( 
.A(n_6087),
.B(n_642),
.Y(n_6274)
);

AND2x2_ASAP7_75t_L g6275 ( 
.A(n_6088),
.B(n_642),
.Y(n_6275)
);

INVxp33_ASAP7_75t_SL g6276 ( 
.A(n_5849),
.Y(n_6276)
);

OAI321xp33_ASAP7_75t_L g6277 ( 
.A1(n_5998),
.A2(n_646),
.A3(n_649),
.B1(n_644),
.B2(n_645),
.C(n_648),
.Y(n_6277)
);

INVx2_ASAP7_75t_L g6278 ( 
.A(n_5949),
.Y(n_6278)
);

INVx1_ASAP7_75t_L g6279 ( 
.A(n_6093),
.Y(n_6279)
);

AOI22xp33_ASAP7_75t_L g6280 ( 
.A1(n_5992),
.A2(n_6008),
.B1(n_6018),
.B2(n_6004),
.Y(n_6280)
);

NAND2xp5_ASAP7_75t_L g6281 ( 
.A(n_6174),
.B(n_5954),
.Y(n_6281)
);

NAND2xp5_ASAP7_75t_L g6282 ( 
.A(n_6248),
.B(n_5861),
.Y(n_6282)
);

INVx1_ASAP7_75t_L g6283 ( 
.A(n_6161),
.Y(n_6283)
);

NAND2xp5_ASAP7_75t_L g6284 ( 
.A(n_6231),
.B(n_5867),
.Y(n_6284)
);

BUFx2_ASAP7_75t_L g6285 ( 
.A(n_6237),
.Y(n_6285)
);

AOI22xp33_ASAP7_75t_L g6286 ( 
.A1(n_6132),
.A2(n_5937),
.B1(n_5961),
.B2(n_5956),
.Y(n_6286)
);

AND2x2_ASAP7_75t_L g6287 ( 
.A(n_6099),
.B(n_5885),
.Y(n_6287)
);

INVx1_ASAP7_75t_L g6288 ( 
.A(n_6226),
.Y(n_6288)
);

INVx1_ASAP7_75t_L g6289 ( 
.A(n_6232),
.Y(n_6289)
);

NAND2xp5_ASAP7_75t_L g6290 ( 
.A(n_6240),
.B(n_5842),
.Y(n_6290)
);

INVx2_ASAP7_75t_L g6291 ( 
.A(n_6246),
.Y(n_6291)
);

NOR2xp33_ASAP7_75t_L g6292 ( 
.A(n_6123),
.B(n_6062),
.Y(n_6292)
);

INVx1_ASAP7_75t_L g6293 ( 
.A(n_6236),
.Y(n_6293)
);

INVx1_ASAP7_75t_L g6294 ( 
.A(n_6148),
.Y(n_6294)
);

AND2x2_ASAP7_75t_L g6295 ( 
.A(n_6242),
.B(n_5855),
.Y(n_6295)
);

AND2x2_ASAP7_75t_L g6296 ( 
.A(n_6265),
.B(n_5914),
.Y(n_6296)
);

INVx1_ASAP7_75t_L g6297 ( 
.A(n_6109),
.Y(n_6297)
);

INVx2_ASAP7_75t_L g6298 ( 
.A(n_6254),
.Y(n_6298)
);

INVx2_ASAP7_75t_L g6299 ( 
.A(n_6254),
.Y(n_6299)
);

OR2x2_ASAP7_75t_L g6300 ( 
.A(n_6119),
.B(n_5918),
.Y(n_6300)
);

NAND2xp5_ASAP7_75t_L g6301 ( 
.A(n_6188),
.B(n_5917),
.Y(n_6301)
);

INVx1_ASAP7_75t_L g6302 ( 
.A(n_6131),
.Y(n_6302)
);

AND2x2_ASAP7_75t_L g6303 ( 
.A(n_6199),
.B(n_5931),
.Y(n_6303)
);

AND2x2_ASAP7_75t_L g6304 ( 
.A(n_6120),
.B(n_5933),
.Y(n_6304)
);

INVx1_ASAP7_75t_L g6305 ( 
.A(n_6104),
.Y(n_6305)
);

INVx1_ASAP7_75t_L g6306 ( 
.A(n_6113),
.Y(n_6306)
);

AND2x2_ASAP7_75t_L g6307 ( 
.A(n_6135),
.B(n_5972),
.Y(n_6307)
);

AND2x2_ASAP7_75t_L g6308 ( 
.A(n_6155),
.B(n_5948),
.Y(n_6308)
);

NOR2xp33_ASAP7_75t_L g6309 ( 
.A(n_6276),
.B(n_6063),
.Y(n_6309)
);

NAND2xp5_ASAP7_75t_L g6310 ( 
.A(n_6112),
.B(n_6009),
.Y(n_6310)
);

INVx1_ASAP7_75t_L g6311 ( 
.A(n_6117),
.Y(n_6311)
);

NAND2xp5_ASAP7_75t_L g6312 ( 
.A(n_6128),
.B(n_5985),
.Y(n_6312)
);

INVx2_ASAP7_75t_L g6313 ( 
.A(n_6230),
.Y(n_6313)
);

INVx1_ASAP7_75t_L g6314 ( 
.A(n_6121),
.Y(n_6314)
);

OR2x2_ASAP7_75t_L g6315 ( 
.A(n_6182),
.B(n_6070),
.Y(n_6315)
);

INVx2_ASAP7_75t_SL g6316 ( 
.A(n_6098),
.Y(n_6316)
);

NAND2xp5_ASAP7_75t_L g6317 ( 
.A(n_6253),
.B(n_5986),
.Y(n_6317)
);

INVx1_ASAP7_75t_L g6318 ( 
.A(n_6126),
.Y(n_6318)
);

INVxp33_ASAP7_75t_L g6319 ( 
.A(n_6193),
.Y(n_6319)
);

AND2x2_ASAP7_75t_L g6320 ( 
.A(n_6142),
.B(n_5887),
.Y(n_6320)
);

INVx1_ASAP7_75t_L g6321 ( 
.A(n_6130),
.Y(n_6321)
);

INVx2_ASAP7_75t_L g6322 ( 
.A(n_6235),
.Y(n_6322)
);

AND2x4_ASAP7_75t_L g6323 ( 
.A(n_6185),
.B(n_5974),
.Y(n_6323)
);

HB1xp67_ASAP7_75t_L g6324 ( 
.A(n_6127),
.Y(n_6324)
);

AOI22xp33_ASAP7_75t_L g6325 ( 
.A1(n_6146),
.A2(n_5978),
.B1(n_5979),
.B2(n_5959),
.Y(n_6325)
);

INVx2_ASAP7_75t_L g6326 ( 
.A(n_6187),
.Y(n_6326)
);

INVx1_ASAP7_75t_L g6327 ( 
.A(n_6133),
.Y(n_6327)
);

HB1xp67_ASAP7_75t_L g6328 ( 
.A(n_6162),
.Y(n_6328)
);

INVx2_ASAP7_75t_L g6329 ( 
.A(n_6228),
.Y(n_6329)
);

OR2x2_ASAP7_75t_L g6330 ( 
.A(n_6116),
.B(n_6092),
.Y(n_6330)
);

OR2x2_ASAP7_75t_L g6331 ( 
.A(n_6106),
.B(n_6076),
.Y(n_6331)
);

NAND2xp5_ASAP7_75t_L g6332 ( 
.A(n_6114),
.B(n_5988),
.Y(n_6332)
);

INVx1_ASAP7_75t_L g6333 ( 
.A(n_6136),
.Y(n_6333)
);

AND2x4_ASAP7_75t_L g6334 ( 
.A(n_6210),
.B(n_5951),
.Y(n_6334)
);

INVxp33_ASAP7_75t_L g6335 ( 
.A(n_6227),
.Y(n_6335)
);

INVx1_ASAP7_75t_L g6336 ( 
.A(n_6144),
.Y(n_6336)
);

INVx1_ASAP7_75t_L g6337 ( 
.A(n_6147),
.Y(n_6337)
);

OR2x2_ASAP7_75t_L g6338 ( 
.A(n_6122),
.B(n_6078),
.Y(n_6338)
);

OR2x2_ASAP7_75t_L g6339 ( 
.A(n_6211),
.B(n_6091),
.Y(n_6339)
);

INVx1_ASAP7_75t_L g6340 ( 
.A(n_6160),
.Y(n_6340)
);

OR2x2_ASAP7_75t_L g6341 ( 
.A(n_6207),
.B(n_5915),
.Y(n_6341)
);

AND2x2_ASAP7_75t_L g6342 ( 
.A(n_6170),
.B(n_5871),
.Y(n_6342)
);

NAND2xp5_ASAP7_75t_L g6343 ( 
.A(n_6097),
.B(n_6033),
.Y(n_6343)
);

AND2x2_ASAP7_75t_L g6344 ( 
.A(n_6105),
.B(n_5976),
.Y(n_6344)
);

OR2x2_ASAP7_75t_L g6345 ( 
.A(n_6257),
.B(n_6035),
.Y(n_6345)
);

NAND2xp5_ASAP7_75t_L g6346 ( 
.A(n_6118),
.B(n_6045),
.Y(n_6346)
);

INVx2_ASAP7_75t_L g6347 ( 
.A(n_6129),
.Y(n_6347)
);

AND2x2_ASAP7_75t_L g6348 ( 
.A(n_6096),
.B(n_6059),
.Y(n_6348)
);

NOR2xp33_ASAP7_75t_L g6349 ( 
.A(n_6125),
.B(n_5964),
.Y(n_6349)
);

INVx3_ASAP7_75t_L g6350 ( 
.A(n_6164),
.Y(n_6350)
);

AND2x2_ASAP7_75t_L g6351 ( 
.A(n_6177),
.B(n_5924),
.Y(n_6351)
);

INVx2_ASAP7_75t_L g6352 ( 
.A(n_6215),
.Y(n_6352)
);

AND2x2_ASAP7_75t_L g6353 ( 
.A(n_6203),
.B(n_5934),
.Y(n_6353)
);

INVx2_ASAP7_75t_L g6354 ( 
.A(n_6209),
.Y(n_6354)
);

OR2x2_ASAP7_75t_L g6355 ( 
.A(n_6137),
.B(n_5953),
.Y(n_6355)
);

NAND2xp5_ASAP7_75t_L g6356 ( 
.A(n_6273),
.B(n_5935),
.Y(n_6356)
);

INVx3_ASAP7_75t_R g6357 ( 
.A(n_6156),
.Y(n_6357)
);

INVx1_ASAP7_75t_L g6358 ( 
.A(n_6163),
.Y(n_6358)
);

INVx2_ASAP7_75t_L g6359 ( 
.A(n_6224),
.Y(n_6359)
);

INVx2_ASAP7_75t_L g6360 ( 
.A(n_6151),
.Y(n_6360)
);

AND2x2_ASAP7_75t_L g6361 ( 
.A(n_6110),
.B(n_5936),
.Y(n_6361)
);

AND2x2_ASAP7_75t_L g6362 ( 
.A(n_6229),
.B(n_5942),
.Y(n_6362)
);

AOI21xp33_ASAP7_75t_L g6363 ( 
.A1(n_6111),
.A2(n_5932),
.B(n_5919),
.Y(n_6363)
);

NAND2xp5_ASAP7_75t_L g6364 ( 
.A(n_6094),
.B(n_5944),
.Y(n_6364)
);

AND2x2_ASAP7_75t_L g6365 ( 
.A(n_6108),
.B(n_5969),
.Y(n_6365)
);

INVx1_ASAP7_75t_L g6366 ( 
.A(n_6169),
.Y(n_6366)
);

OR2x2_ASAP7_75t_L g6367 ( 
.A(n_6181),
.B(n_5945),
.Y(n_6367)
);

HB1xp67_ASAP7_75t_L g6368 ( 
.A(n_6176),
.Y(n_6368)
);

INVx2_ASAP7_75t_L g6369 ( 
.A(n_6150),
.Y(n_6369)
);

INVx1_ASAP7_75t_SL g6370 ( 
.A(n_6205),
.Y(n_6370)
);

OR2x2_ASAP7_75t_L g6371 ( 
.A(n_6183),
.B(n_5960),
.Y(n_6371)
);

INVx1_ASAP7_75t_L g6372 ( 
.A(n_6190),
.Y(n_6372)
);

NAND2xp5_ASAP7_75t_L g6373 ( 
.A(n_6171),
.B(n_5888),
.Y(n_6373)
);

NOR2xp33_ASAP7_75t_L g6374 ( 
.A(n_6134),
.B(n_6173),
.Y(n_6374)
);

INVx3_ASAP7_75t_SL g6375 ( 
.A(n_6107),
.Y(n_6375)
);

INVx1_ASAP7_75t_L g6376 ( 
.A(n_6198),
.Y(n_6376)
);

INVx2_ASAP7_75t_L g6377 ( 
.A(n_6197),
.Y(n_6377)
);

INVx1_ASAP7_75t_L g6378 ( 
.A(n_6221),
.Y(n_6378)
);

AND2x2_ASAP7_75t_L g6379 ( 
.A(n_6154),
.B(n_6003),
.Y(n_6379)
);

INVx2_ASAP7_75t_L g6380 ( 
.A(n_6152),
.Y(n_6380)
);

NAND2xp5_ASAP7_75t_L g6381 ( 
.A(n_6206),
.B(n_6223),
.Y(n_6381)
);

AND2x2_ASAP7_75t_L g6382 ( 
.A(n_6233),
.B(n_6012),
.Y(n_6382)
);

INVx1_ASAP7_75t_L g6383 ( 
.A(n_6234),
.Y(n_6383)
);

AND2x2_ASAP7_75t_L g6384 ( 
.A(n_6239),
.B(n_5920),
.Y(n_6384)
);

OR2x2_ASAP7_75t_L g6385 ( 
.A(n_6241),
.B(n_6013),
.Y(n_6385)
);

NAND2xp5_ASAP7_75t_L g6386 ( 
.A(n_6264),
.B(n_645),
.Y(n_6386)
);

AND2x2_ASAP7_75t_L g6387 ( 
.A(n_6274),
.B(n_646),
.Y(n_6387)
);

INVx2_ASAP7_75t_L g6388 ( 
.A(n_6167),
.Y(n_6388)
);

HB1xp67_ASAP7_75t_L g6389 ( 
.A(n_6244),
.Y(n_6389)
);

AND2x4_ASAP7_75t_L g6390 ( 
.A(n_6153),
.B(n_648),
.Y(n_6390)
);

INVx1_ASAP7_75t_L g6391 ( 
.A(n_6250),
.Y(n_6391)
);

INVx1_ASAP7_75t_L g6392 ( 
.A(n_6268),
.Y(n_6392)
);

INVx1_ASAP7_75t_L g6393 ( 
.A(n_6270),
.Y(n_6393)
);

AOI22xp5_ASAP7_75t_L g6394 ( 
.A1(n_6267),
.A2(n_652),
.B1(n_649),
.B2(n_650),
.Y(n_6394)
);

AND2x2_ASAP7_75t_L g6395 ( 
.A(n_6275),
.B(n_650),
.Y(n_6395)
);

AND2x2_ASAP7_75t_L g6396 ( 
.A(n_6158),
.B(n_652),
.Y(n_6396)
);

OR2x2_ASAP7_75t_L g6397 ( 
.A(n_6279),
.B(n_653),
.Y(n_6397)
);

INVx2_ASAP7_75t_L g6398 ( 
.A(n_6179),
.Y(n_6398)
);

NAND2x1_ASAP7_75t_L g6399 ( 
.A(n_6100),
.B(n_6191),
.Y(n_6399)
);

NAND2xp5_ASAP7_75t_L g6400 ( 
.A(n_6138),
.B(n_653),
.Y(n_6400)
);

INVx2_ASAP7_75t_L g6401 ( 
.A(n_6196),
.Y(n_6401)
);

AND2x4_ASAP7_75t_L g6402 ( 
.A(n_6251),
.B(n_654),
.Y(n_6402)
);

NAND2xp5_ASAP7_75t_L g6403 ( 
.A(n_6115),
.B(n_655),
.Y(n_6403)
);

INVx2_ASAP7_75t_L g6404 ( 
.A(n_6200),
.Y(n_6404)
);

AND2x2_ASAP7_75t_L g6405 ( 
.A(n_6168),
.B(n_6140),
.Y(n_6405)
);

NAND2xp5_ASAP7_75t_L g6406 ( 
.A(n_6159),
.B(n_656),
.Y(n_6406)
);

INVx1_ASAP7_75t_L g6407 ( 
.A(n_6222),
.Y(n_6407)
);

INVx1_ASAP7_75t_L g6408 ( 
.A(n_6278),
.Y(n_6408)
);

INVx1_ASAP7_75t_L g6409 ( 
.A(n_6165),
.Y(n_6409)
);

NAND2xp67_ASAP7_75t_L g6410 ( 
.A(n_6143),
.B(n_656),
.Y(n_6410)
);

AND2x2_ASAP7_75t_L g6411 ( 
.A(n_6175),
.B(n_657),
.Y(n_6411)
);

NAND2xp5_ASAP7_75t_L g6412 ( 
.A(n_6255),
.B(n_657),
.Y(n_6412)
);

OR2x2_ASAP7_75t_L g6413 ( 
.A(n_6260),
.B(n_658),
.Y(n_6413)
);

INVx1_ASAP7_75t_L g6414 ( 
.A(n_6245),
.Y(n_6414)
);

OR2x2_ASAP7_75t_L g6415 ( 
.A(n_6102),
.B(n_658),
.Y(n_6415)
);

HB1xp67_ASAP7_75t_L g6416 ( 
.A(n_6103),
.Y(n_6416)
);

AOI22xp5_ASAP7_75t_L g6417 ( 
.A1(n_6412),
.A2(n_6192),
.B1(n_6262),
.B2(n_6225),
.Y(n_6417)
);

AND2x4_ASAP7_75t_SL g6418 ( 
.A(n_6323),
.B(n_6218),
.Y(n_6418)
);

NOR2xp33_ASAP7_75t_L g6419 ( 
.A(n_6370),
.B(n_6204),
.Y(n_6419)
);

INVx1_ASAP7_75t_L g6420 ( 
.A(n_6368),
.Y(n_6420)
);

INVx1_ASAP7_75t_L g6421 ( 
.A(n_6389),
.Y(n_6421)
);

INVx1_ASAP7_75t_L g6422 ( 
.A(n_6300),
.Y(n_6422)
);

NAND2xp5_ASAP7_75t_L g6423 ( 
.A(n_6382),
.B(n_6149),
.Y(n_6423)
);

O2A1O1Ixp33_ASAP7_75t_SL g6424 ( 
.A1(n_6328),
.A2(n_6220),
.B(n_6247),
.C(n_6249),
.Y(n_6424)
);

INVx1_ASAP7_75t_L g6425 ( 
.A(n_6297),
.Y(n_6425)
);

INVx1_ASAP7_75t_L g6426 ( 
.A(n_6283),
.Y(n_6426)
);

OR2x2_ASAP7_75t_L g6427 ( 
.A(n_6326),
.B(n_6385),
.Y(n_6427)
);

AND2x2_ASAP7_75t_L g6428 ( 
.A(n_6375),
.B(n_6280),
.Y(n_6428)
);

HB1xp67_ASAP7_75t_L g6429 ( 
.A(n_6324),
.Y(n_6429)
);

AND2x2_ASAP7_75t_L g6430 ( 
.A(n_6308),
.B(n_6101),
.Y(n_6430)
);

INVx1_ASAP7_75t_L g6431 ( 
.A(n_6301),
.Y(n_6431)
);

AND2x2_ASAP7_75t_L g6432 ( 
.A(n_6307),
.B(n_6285),
.Y(n_6432)
);

AND2x2_ASAP7_75t_L g6433 ( 
.A(n_6295),
.B(n_6095),
.Y(n_6433)
);

NAND2xp5_ASAP7_75t_L g6434 ( 
.A(n_6303),
.B(n_6189),
.Y(n_6434)
);

INVx2_ASAP7_75t_L g6435 ( 
.A(n_6334),
.Y(n_6435)
);

AND2x2_ASAP7_75t_L g6436 ( 
.A(n_6350),
.B(n_6362),
.Y(n_6436)
);

AND2x2_ASAP7_75t_L g6437 ( 
.A(n_6319),
.B(n_6194),
.Y(n_6437)
);

AOI22xp33_ASAP7_75t_L g6438 ( 
.A1(n_6352),
.A2(n_6201),
.B1(n_6208),
.B2(n_6202),
.Y(n_6438)
);

INVx1_ASAP7_75t_L g6439 ( 
.A(n_6302),
.Y(n_6439)
);

AOI22xp33_ASAP7_75t_L g6440 ( 
.A1(n_6335),
.A2(n_6213),
.B1(n_6216),
.B2(n_6214),
.Y(n_6440)
);

NOR2x1_ASAP7_75t_L g6441 ( 
.A(n_6397),
.B(n_6172),
.Y(n_6441)
);

AND2x4_ASAP7_75t_L g6442 ( 
.A(n_6316),
.B(n_6252),
.Y(n_6442)
);

OR2x2_ASAP7_75t_L g6443 ( 
.A(n_6284),
.B(n_6217),
.Y(n_6443)
);

INVx1_ASAP7_75t_L g6444 ( 
.A(n_6371),
.Y(n_6444)
);

INVxp67_ASAP7_75t_SL g6445 ( 
.A(n_6374),
.Y(n_6445)
);

AND2x2_ASAP7_75t_L g6446 ( 
.A(n_6342),
.B(n_6243),
.Y(n_6446)
);

AND2x2_ASAP7_75t_L g6447 ( 
.A(n_6287),
.B(n_6258),
.Y(n_6447)
);

AND2x2_ASAP7_75t_L g6448 ( 
.A(n_6353),
.B(n_6259),
.Y(n_6448)
);

NAND2xp5_ASAP7_75t_L g6449 ( 
.A(n_6344),
.B(n_6124),
.Y(n_6449)
);

INVx2_ASAP7_75t_L g6450 ( 
.A(n_6361),
.Y(n_6450)
);

OAI211xp5_ASAP7_75t_SL g6451 ( 
.A1(n_6363),
.A2(n_6212),
.B(n_6166),
.C(n_6263),
.Y(n_6451)
);

INVx1_ASAP7_75t_L g6452 ( 
.A(n_6400),
.Y(n_6452)
);

AND2x2_ASAP7_75t_L g6453 ( 
.A(n_6351),
.B(n_6261),
.Y(n_6453)
);

AND2x2_ASAP7_75t_L g6454 ( 
.A(n_6291),
.B(n_6269),
.Y(n_6454)
);

NAND2xp5_ASAP7_75t_L g6455 ( 
.A(n_6296),
.B(n_6184),
.Y(n_6455)
);

INVx1_ASAP7_75t_L g6456 ( 
.A(n_6305),
.Y(n_6456)
);

AOI22xp5_ASAP7_75t_L g6457 ( 
.A1(n_6394),
.A2(n_6390),
.B1(n_6405),
.B2(n_6364),
.Y(n_6457)
);

NAND2xp5_ASAP7_75t_L g6458 ( 
.A(n_6360),
.B(n_6139),
.Y(n_6458)
);

AND2x2_ASAP7_75t_L g6459 ( 
.A(n_6320),
.B(n_6272),
.Y(n_6459)
);

AND2x2_ASAP7_75t_L g6460 ( 
.A(n_6313),
.B(n_6186),
.Y(n_6460)
);

OAI21xp33_ASAP7_75t_SL g6461 ( 
.A1(n_6347),
.A2(n_6145),
.B(n_6141),
.Y(n_6461)
);

INVx2_ASAP7_75t_L g6462 ( 
.A(n_6365),
.Y(n_6462)
);

AND2x4_ASAP7_75t_L g6463 ( 
.A(n_6322),
.B(n_6266),
.Y(n_6463)
);

INVx1_ASAP7_75t_L g6464 ( 
.A(n_6306),
.Y(n_6464)
);

AND2x2_ASAP7_75t_L g6465 ( 
.A(n_6354),
.B(n_6157),
.Y(n_6465)
);

NAND2xp5_ASAP7_75t_L g6466 ( 
.A(n_6409),
.B(n_6178),
.Y(n_6466)
);

INVx3_ASAP7_75t_L g6467 ( 
.A(n_6402),
.Y(n_6467)
);

INVx2_ASAP7_75t_L g6468 ( 
.A(n_6384),
.Y(n_6468)
);

AND2x4_ASAP7_75t_L g6469 ( 
.A(n_6401),
.B(n_6219),
.Y(n_6469)
);

NAND2xp5_ASAP7_75t_L g6470 ( 
.A(n_6379),
.B(n_6195),
.Y(n_6470)
);

AOI22xp5_ASAP7_75t_L g6471 ( 
.A1(n_6312),
.A2(n_6238),
.B1(n_6271),
.B2(n_6256),
.Y(n_6471)
);

NOR2xp67_ASAP7_75t_L g6472 ( 
.A(n_6381),
.B(n_6277),
.Y(n_6472)
);

INVx1_ASAP7_75t_L g6473 ( 
.A(n_6311),
.Y(n_6473)
);

INVx1_ASAP7_75t_L g6474 ( 
.A(n_6314),
.Y(n_6474)
);

NAND2x1_ASAP7_75t_L g6475 ( 
.A(n_6349),
.B(n_6329),
.Y(n_6475)
);

BUFx2_ASAP7_75t_L g6476 ( 
.A(n_6282),
.Y(n_6476)
);

NAND2x1p5_ASAP7_75t_L g6477 ( 
.A(n_6387),
.B(n_6180),
.Y(n_6477)
);

INVx2_ASAP7_75t_SL g6478 ( 
.A(n_6399),
.Y(n_6478)
);

INVx1_ASAP7_75t_L g6479 ( 
.A(n_6318),
.Y(n_6479)
);

INVx2_ASAP7_75t_L g6480 ( 
.A(n_6355),
.Y(n_6480)
);

OR2x2_ASAP7_75t_L g6481 ( 
.A(n_6290),
.B(n_659),
.Y(n_6481)
);

NAND2xp5_ASAP7_75t_L g6482 ( 
.A(n_6416),
.B(n_6309),
.Y(n_6482)
);

INVx2_ASAP7_75t_L g6483 ( 
.A(n_6410),
.Y(n_6483)
);

INVx2_ASAP7_75t_L g6484 ( 
.A(n_6345),
.Y(n_6484)
);

OR2x2_ASAP7_75t_L g6485 ( 
.A(n_6331),
.B(n_659),
.Y(n_6485)
);

INVx2_ASAP7_75t_L g6486 ( 
.A(n_6377),
.Y(n_6486)
);

INVx1_ASAP7_75t_L g6487 ( 
.A(n_6321),
.Y(n_6487)
);

AOI211xp5_ASAP7_75t_L g6488 ( 
.A1(n_6343),
.A2(n_662),
.B(n_660),
.C(n_661),
.Y(n_6488)
);

INVx1_ASAP7_75t_L g6489 ( 
.A(n_6327),
.Y(n_6489)
);

INVx1_ASAP7_75t_L g6490 ( 
.A(n_6333),
.Y(n_6490)
);

AND2x2_ASAP7_75t_L g6491 ( 
.A(n_6298),
.B(n_660),
.Y(n_6491)
);

OAI22xp5_ASAP7_75t_L g6492 ( 
.A1(n_6281),
.A2(n_6346),
.B1(n_6332),
.B2(n_6310),
.Y(n_6492)
);

INVx1_ASAP7_75t_L g6493 ( 
.A(n_6336),
.Y(n_6493)
);

OAI31xp33_ASAP7_75t_L g6494 ( 
.A1(n_6317),
.A2(n_664),
.A3(n_662),
.B(n_663),
.Y(n_6494)
);

INVx1_ASAP7_75t_L g6495 ( 
.A(n_6337),
.Y(n_6495)
);

INVxp67_ASAP7_75t_L g6496 ( 
.A(n_6292),
.Y(n_6496)
);

AND2x2_ASAP7_75t_L g6497 ( 
.A(n_6299),
.B(n_665),
.Y(n_6497)
);

AND2x4_ASAP7_75t_L g6498 ( 
.A(n_6369),
.B(n_666),
.Y(n_6498)
);

INVx2_ASAP7_75t_L g6499 ( 
.A(n_6395),
.Y(n_6499)
);

INVx1_ASAP7_75t_L g6500 ( 
.A(n_6340),
.Y(n_6500)
);

INVx1_ASAP7_75t_SL g6501 ( 
.A(n_6396),
.Y(n_6501)
);

NAND2xp5_ASAP7_75t_L g6502 ( 
.A(n_6294),
.B(n_666),
.Y(n_6502)
);

INVx1_ASAP7_75t_L g6503 ( 
.A(n_6358),
.Y(n_6503)
);

INVx2_ASAP7_75t_L g6504 ( 
.A(n_6338),
.Y(n_6504)
);

OAI21xp5_ASAP7_75t_L g6505 ( 
.A1(n_6403),
.A2(n_667),
.B(n_668),
.Y(n_6505)
);

INVx1_ASAP7_75t_SL g6506 ( 
.A(n_6356),
.Y(n_6506)
);

NOR2xp33_ASAP7_75t_L g6507 ( 
.A(n_6357),
.B(n_668),
.Y(n_6507)
);

INVx2_ASAP7_75t_L g6508 ( 
.A(n_6404),
.Y(n_6508)
);

INVx1_ASAP7_75t_L g6509 ( 
.A(n_6366),
.Y(n_6509)
);

INVxp67_ASAP7_75t_SL g6510 ( 
.A(n_6367),
.Y(n_6510)
);

OAI21xp5_ASAP7_75t_L g6511 ( 
.A1(n_6413),
.A2(n_669),
.B(n_670),
.Y(n_6511)
);

INVx1_ASAP7_75t_L g6512 ( 
.A(n_6372),
.Y(n_6512)
);

INVx1_ASAP7_75t_L g6513 ( 
.A(n_6376),
.Y(n_6513)
);

AND2x2_ASAP7_75t_L g6514 ( 
.A(n_6304),
.B(n_669),
.Y(n_6514)
);

OAI211xp5_ASAP7_75t_SL g6515 ( 
.A1(n_6288),
.A2(n_674),
.B(n_672),
.C(n_673),
.Y(n_6515)
);

NAND2xp5_ASAP7_75t_L g6516 ( 
.A(n_6341),
.B(n_673),
.Y(n_6516)
);

INVx4_ASAP7_75t_L g6517 ( 
.A(n_6411),
.Y(n_6517)
);

INVx1_ASAP7_75t_L g6518 ( 
.A(n_6378),
.Y(n_6518)
);

AND2x4_ASAP7_75t_L g6519 ( 
.A(n_6348),
.B(n_674),
.Y(n_6519)
);

BUFx2_ASAP7_75t_L g6520 ( 
.A(n_6289),
.Y(n_6520)
);

NAND2xp5_ASAP7_75t_SL g6521 ( 
.A(n_6315),
.B(n_675),
.Y(n_6521)
);

AND2x2_ASAP7_75t_L g6522 ( 
.A(n_6293),
.B(n_677),
.Y(n_6522)
);

OAI21xp5_ASAP7_75t_SL g6523 ( 
.A1(n_6415),
.A2(n_677),
.B(n_678),
.Y(n_6523)
);

INVx1_ASAP7_75t_L g6524 ( 
.A(n_6383),
.Y(n_6524)
);

INVx1_ASAP7_75t_L g6525 ( 
.A(n_6391),
.Y(n_6525)
);

NAND2xp5_ASAP7_75t_L g6526 ( 
.A(n_6373),
.B(n_678),
.Y(n_6526)
);

INVx1_ASAP7_75t_L g6527 ( 
.A(n_6392),
.Y(n_6527)
);

AND2x4_ASAP7_75t_L g6528 ( 
.A(n_6359),
.B(n_679),
.Y(n_6528)
);

AND2x2_ASAP7_75t_L g6529 ( 
.A(n_6330),
.B(n_680),
.Y(n_6529)
);

INVx2_ASAP7_75t_L g6530 ( 
.A(n_6414),
.Y(n_6530)
);

NAND2xp5_ASAP7_75t_L g6531 ( 
.A(n_6339),
.B(n_681),
.Y(n_6531)
);

INVx1_ASAP7_75t_L g6532 ( 
.A(n_6393),
.Y(n_6532)
);

INVx1_ASAP7_75t_L g6533 ( 
.A(n_6407),
.Y(n_6533)
);

AOI33xp33_ASAP7_75t_L g6534 ( 
.A1(n_6325),
.A2(n_706),
.A3(n_689),
.B1(n_714),
.B2(n_698),
.B3(n_681),
.Y(n_6534)
);

OA21x2_ASAP7_75t_L g6535 ( 
.A1(n_6408),
.A2(n_682),
.B(n_683),
.Y(n_6535)
);

NOR2xp33_ASAP7_75t_L g6536 ( 
.A(n_6386),
.B(n_684),
.Y(n_6536)
);

AND2x2_ASAP7_75t_L g6537 ( 
.A(n_6406),
.B(n_684),
.Y(n_6537)
);

AND2x2_ASAP7_75t_L g6538 ( 
.A(n_6286),
.B(n_6380),
.Y(n_6538)
);

NAND2xp5_ASAP7_75t_L g6539 ( 
.A(n_6388),
.B(n_6398),
.Y(n_6539)
);

AND2x2_ASAP7_75t_L g6540 ( 
.A(n_6375),
.B(n_685),
.Y(n_6540)
);

NOR2x1_ASAP7_75t_SL g6541 ( 
.A(n_6381),
.B(n_685),
.Y(n_6541)
);

INVx2_ASAP7_75t_SL g6542 ( 
.A(n_6323),
.Y(n_6542)
);

HB1xp67_ASAP7_75t_L g6543 ( 
.A(n_6324),
.Y(n_6543)
);

INVx2_ASAP7_75t_L g6544 ( 
.A(n_6323),
.Y(n_6544)
);

AND2x2_ASAP7_75t_L g6545 ( 
.A(n_6375),
.B(n_686),
.Y(n_6545)
);

NAND2xp5_ASAP7_75t_L g6546 ( 
.A(n_6382),
.B(n_686),
.Y(n_6546)
);

AND2x2_ASAP7_75t_L g6547 ( 
.A(n_6375),
.B(n_687),
.Y(n_6547)
);

OR2x2_ASAP7_75t_L g6548 ( 
.A(n_6326),
.B(n_687),
.Y(n_6548)
);

INVx1_ASAP7_75t_L g6549 ( 
.A(n_6368),
.Y(n_6549)
);

INVx1_ASAP7_75t_L g6550 ( 
.A(n_6510),
.Y(n_6550)
);

NAND3xp33_ASAP7_75t_SL g6551 ( 
.A(n_6494),
.B(n_688),
.C(n_689),
.Y(n_6551)
);

AND2x2_ASAP7_75t_L g6552 ( 
.A(n_6432),
.B(n_688),
.Y(n_6552)
);

INVx2_ASAP7_75t_L g6553 ( 
.A(n_6517),
.Y(n_6553)
);

INVx1_ASAP7_75t_L g6554 ( 
.A(n_6516),
.Y(n_6554)
);

NAND2xp5_ASAP7_75t_L g6555 ( 
.A(n_6501),
.B(n_690),
.Y(n_6555)
);

O2A1O1Ixp33_ASAP7_75t_SL g6556 ( 
.A1(n_6475),
.A2(n_701),
.B(n_710),
.C(n_691),
.Y(n_6556)
);

NOR2xp33_ASAP7_75t_R g6557 ( 
.A(n_6542),
.B(n_691),
.Y(n_6557)
);

OR2x2_ASAP7_75t_L g6558 ( 
.A(n_6427),
.B(n_692),
.Y(n_6558)
);

INVx2_ASAP7_75t_L g6559 ( 
.A(n_6436),
.Y(n_6559)
);

INVx2_ASAP7_75t_L g6560 ( 
.A(n_6541),
.Y(n_6560)
);

NAND5xp2_ASAP7_75t_L g6561 ( 
.A(n_6445),
.B(n_694),
.C(n_692),
.D(n_693),
.E(n_695),
.Y(n_6561)
);

HB1xp67_ASAP7_75t_L g6562 ( 
.A(n_6540),
.Y(n_6562)
);

INVx2_ASAP7_75t_L g6563 ( 
.A(n_6519),
.Y(n_6563)
);

INVx2_ASAP7_75t_L g6564 ( 
.A(n_6545),
.Y(n_6564)
);

OR2x2_ASAP7_75t_L g6565 ( 
.A(n_6476),
.B(n_6482),
.Y(n_6565)
);

AND2x2_ASAP7_75t_L g6566 ( 
.A(n_6450),
.B(n_693),
.Y(n_6566)
);

OR2x2_ASAP7_75t_L g6567 ( 
.A(n_6444),
.B(n_694),
.Y(n_6567)
);

NAND2xp33_ASAP7_75t_L g6568 ( 
.A(n_6547),
.B(n_695),
.Y(n_6568)
);

AND2x2_ASAP7_75t_L g6569 ( 
.A(n_6435),
.B(n_697),
.Y(n_6569)
);

INVx1_ASAP7_75t_L g6570 ( 
.A(n_6531),
.Y(n_6570)
);

NAND2x1_ASAP7_75t_SL g6571 ( 
.A(n_6467),
.B(n_697),
.Y(n_6571)
);

NAND4xp25_ASAP7_75t_L g6572 ( 
.A(n_6496),
.B(n_701),
.C(n_699),
.D(n_700),
.Y(n_6572)
);

INVx1_ASAP7_75t_L g6573 ( 
.A(n_6529),
.Y(n_6573)
);

NAND4xp25_ASAP7_75t_L g6574 ( 
.A(n_6544),
.B(n_704),
.C(n_702),
.D(n_703),
.Y(n_6574)
);

AND2x2_ASAP7_75t_L g6575 ( 
.A(n_6468),
.B(n_702),
.Y(n_6575)
);

INVx2_ASAP7_75t_SL g6576 ( 
.A(n_6453),
.Y(n_6576)
);

NAND2x1_ASAP7_75t_SL g6577 ( 
.A(n_6447),
.B(n_705),
.Y(n_6577)
);

INVxp67_ASAP7_75t_L g6578 ( 
.A(n_6507),
.Y(n_6578)
);

INVx1_ASAP7_75t_L g6579 ( 
.A(n_6546),
.Y(n_6579)
);

AND2x2_ASAP7_75t_L g6580 ( 
.A(n_6462),
.B(n_707),
.Y(n_6580)
);

AND2x4_ASAP7_75t_L g6581 ( 
.A(n_6446),
.B(n_6499),
.Y(n_6581)
);

HB1xp67_ASAP7_75t_L g6582 ( 
.A(n_6429),
.Y(n_6582)
);

INVx1_ASAP7_75t_L g6583 ( 
.A(n_6485),
.Y(n_6583)
);

NAND2xp5_ASAP7_75t_L g6584 ( 
.A(n_6472),
.B(n_707),
.Y(n_6584)
);

AND2x2_ASAP7_75t_L g6585 ( 
.A(n_6522),
.B(n_6514),
.Y(n_6585)
);

AND2x2_ASAP7_75t_L g6586 ( 
.A(n_6478),
.B(n_708),
.Y(n_6586)
);

INVx1_ASAP7_75t_L g6587 ( 
.A(n_6520),
.Y(n_6587)
);

INVx3_ASAP7_75t_SL g6588 ( 
.A(n_6481),
.Y(n_6588)
);

NAND2x1_ASAP7_75t_L g6589 ( 
.A(n_6428),
.B(n_708),
.Y(n_6589)
);

INVx2_ASAP7_75t_L g6590 ( 
.A(n_6535),
.Y(n_6590)
);

INVx2_ASAP7_75t_L g6591 ( 
.A(n_6528),
.Y(n_6591)
);

NAND4xp25_ASAP7_75t_L g6592 ( 
.A(n_6492),
.B(n_712),
.C(n_709),
.D(n_711),
.Y(n_6592)
);

NOR3xp33_ASAP7_75t_SL g6593 ( 
.A(n_6431),
.B(n_709),
.C(n_713),
.Y(n_6593)
);

NAND3xp33_ASAP7_75t_L g6594 ( 
.A(n_6488),
.B(n_714),
.C(n_716),
.Y(n_6594)
);

NAND2xp5_ASAP7_75t_L g6595 ( 
.A(n_6477),
.B(n_717),
.Y(n_6595)
);

NAND3xp33_ASAP7_75t_L g6596 ( 
.A(n_6543),
.B(n_718),
.C(n_719),
.Y(n_6596)
);

NAND2xp5_ASAP7_75t_L g6597 ( 
.A(n_6419),
.B(n_718),
.Y(n_6597)
);

INVx1_ASAP7_75t_L g6598 ( 
.A(n_6480),
.Y(n_6598)
);

OR2x2_ASAP7_75t_L g6599 ( 
.A(n_6422),
.B(n_719),
.Y(n_6599)
);

OR2x2_ASAP7_75t_L g6600 ( 
.A(n_6484),
.B(n_6506),
.Y(n_6600)
);

INVx2_ASAP7_75t_SL g6601 ( 
.A(n_6448),
.Y(n_6601)
);

AND2x2_ASAP7_75t_L g6602 ( 
.A(n_6437),
.B(n_720),
.Y(n_6602)
);

NOR2x1_ASAP7_75t_L g6603 ( 
.A(n_6526),
.B(n_720),
.Y(n_6603)
);

INVxp33_ASAP7_75t_L g6604 ( 
.A(n_6441),
.Y(n_6604)
);

NAND2xp5_ASAP7_75t_L g6605 ( 
.A(n_6459),
.B(n_722),
.Y(n_6605)
);

INVx1_ASAP7_75t_L g6606 ( 
.A(n_6530),
.Y(n_6606)
);

NOR3xp33_ASAP7_75t_SL g6607 ( 
.A(n_6420),
.B(n_722),
.C(n_723),
.Y(n_6607)
);

INVx1_ASAP7_75t_L g6608 ( 
.A(n_6502),
.Y(n_6608)
);

NAND2xp33_ASAP7_75t_R g6609 ( 
.A(n_6548),
.B(n_723),
.Y(n_6609)
);

OAI211xp5_ASAP7_75t_SL g6610 ( 
.A1(n_6461),
.A2(n_726),
.B(n_724),
.C(n_725),
.Y(n_6610)
);

NAND2xp5_ASAP7_75t_SL g6611 ( 
.A(n_6457),
.B(n_724),
.Y(n_6611)
);

OR2x2_ASAP7_75t_L g6612 ( 
.A(n_6443),
.B(n_725),
.Y(n_6612)
);

INVx2_ASAP7_75t_L g6613 ( 
.A(n_6498),
.Y(n_6613)
);

NOR3xp33_ASAP7_75t_L g6614 ( 
.A(n_6523),
.B(n_726),
.C(n_727),
.Y(n_6614)
);

NOR2xp33_ASAP7_75t_R g6615 ( 
.A(n_6421),
.B(n_727),
.Y(n_6615)
);

NAND2xp5_ASAP7_75t_L g6616 ( 
.A(n_6417),
.B(n_728),
.Y(n_6616)
);

INVx1_ASAP7_75t_L g6617 ( 
.A(n_6504),
.Y(n_6617)
);

AOI211xp5_ASAP7_75t_L g6618 ( 
.A1(n_6424),
.A2(n_730),
.B(n_728),
.C(n_729),
.Y(n_6618)
);

AND2x2_ASAP7_75t_L g6619 ( 
.A(n_6433),
.B(n_730),
.Y(n_6619)
);

INVx1_ASAP7_75t_L g6620 ( 
.A(n_6486),
.Y(n_6620)
);

INVx3_ASAP7_75t_L g6621 ( 
.A(n_6469),
.Y(n_6621)
);

AND2x2_ASAP7_75t_L g6622 ( 
.A(n_6430),
.B(n_731),
.Y(n_6622)
);

INVx1_ASAP7_75t_L g6623 ( 
.A(n_6549),
.Y(n_6623)
);

AND2x4_ASAP7_75t_L g6624 ( 
.A(n_6454),
.B(n_731),
.Y(n_6624)
);

INVx1_ASAP7_75t_L g6625 ( 
.A(n_6539),
.Y(n_6625)
);

OAI21xp5_ASAP7_75t_SL g6626 ( 
.A1(n_6434),
.A2(n_732),
.B(n_733),
.Y(n_6626)
);

BUFx2_ASAP7_75t_L g6627 ( 
.A(n_6425),
.Y(n_6627)
);

INVx1_ASAP7_75t_L g6628 ( 
.A(n_6439),
.Y(n_6628)
);

INVx1_ASAP7_75t_L g6629 ( 
.A(n_6508),
.Y(n_6629)
);

OAI211xp5_ASAP7_75t_L g6630 ( 
.A1(n_6455),
.A2(n_735),
.B(n_733),
.C(n_734),
.Y(n_6630)
);

AND2x2_ASAP7_75t_L g6631 ( 
.A(n_6491),
.B(n_734),
.Y(n_6631)
);

OR2x2_ASAP7_75t_L g6632 ( 
.A(n_6426),
.B(n_735),
.Y(n_6632)
);

BUFx2_ASAP7_75t_L g6633 ( 
.A(n_6511),
.Y(n_6633)
);

NAND2xp5_ASAP7_75t_L g6634 ( 
.A(n_6460),
.B(n_736),
.Y(n_6634)
);

NOR2x1_ASAP7_75t_L g6635 ( 
.A(n_6515),
.B(n_737),
.Y(n_6635)
);

NOR2xp33_ASAP7_75t_R g6636 ( 
.A(n_6497),
.B(n_737),
.Y(n_6636)
);

NAND3xp33_ASAP7_75t_L g6637 ( 
.A(n_6451),
.B(n_738),
.C(n_739),
.Y(n_6637)
);

INVx2_ASAP7_75t_L g6638 ( 
.A(n_6463),
.Y(n_6638)
);

AND2x2_ASAP7_75t_L g6639 ( 
.A(n_6418),
.B(n_738),
.Y(n_6639)
);

INVx1_ASAP7_75t_L g6640 ( 
.A(n_6456),
.Y(n_6640)
);

INVx1_ASAP7_75t_L g6641 ( 
.A(n_6464),
.Y(n_6641)
);

INVx1_ASAP7_75t_L g6642 ( 
.A(n_6473),
.Y(n_6642)
);

INVx1_ASAP7_75t_L g6643 ( 
.A(n_6474),
.Y(n_6643)
);

NAND2xp33_ASAP7_75t_R g6644 ( 
.A(n_6423),
.B(n_740),
.Y(n_6644)
);

NAND2xp5_ASAP7_75t_L g6645 ( 
.A(n_6536),
.B(n_740),
.Y(n_6645)
);

INVx1_ASAP7_75t_L g6646 ( 
.A(n_6479),
.Y(n_6646)
);

INVx1_ASAP7_75t_L g6647 ( 
.A(n_6487),
.Y(n_6647)
);

INVx2_ASAP7_75t_L g6648 ( 
.A(n_6442),
.Y(n_6648)
);

AND2x2_ASAP7_75t_L g6649 ( 
.A(n_6465),
.B(n_741),
.Y(n_6649)
);

INVx2_ASAP7_75t_L g6650 ( 
.A(n_6537),
.Y(n_6650)
);

AND2x2_ASAP7_75t_L g6651 ( 
.A(n_6489),
.B(n_741),
.Y(n_6651)
);

NAND4xp25_ASAP7_75t_L g6652 ( 
.A(n_6490),
.B(n_6493),
.C(n_6500),
.D(n_6495),
.Y(n_6652)
);

OR2x2_ASAP7_75t_L g6653 ( 
.A(n_6449),
.B(n_742),
.Y(n_6653)
);

AND2x2_ASAP7_75t_L g6654 ( 
.A(n_6503),
.B(n_743),
.Y(n_6654)
);

INVx1_ASAP7_75t_SL g6655 ( 
.A(n_6470),
.Y(n_6655)
);

NAND2xp33_ASAP7_75t_R g6656 ( 
.A(n_6505),
.B(n_743),
.Y(n_6656)
);

INVx2_ASAP7_75t_L g6657 ( 
.A(n_6483),
.Y(n_6657)
);

OR2x2_ASAP7_75t_L g6658 ( 
.A(n_6452),
.B(n_745),
.Y(n_6658)
);

NAND2xp5_ASAP7_75t_L g6659 ( 
.A(n_6534),
.B(n_745),
.Y(n_6659)
);

OR2x2_ASAP7_75t_L g6660 ( 
.A(n_6509),
.B(n_746),
.Y(n_6660)
);

INVx2_ASAP7_75t_L g6661 ( 
.A(n_6538),
.Y(n_6661)
);

AND2x2_ASAP7_75t_L g6662 ( 
.A(n_6512),
.B(n_746),
.Y(n_6662)
);

INVx1_ASAP7_75t_L g6663 ( 
.A(n_6513),
.Y(n_6663)
);

AND2x2_ASAP7_75t_L g6664 ( 
.A(n_6518),
.B(n_747),
.Y(n_6664)
);

INVx2_ASAP7_75t_L g6665 ( 
.A(n_6521),
.Y(n_6665)
);

AND2x2_ASAP7_75t_L g6666 ( 
.A(n_6524),
.B(n_747),
.Y(n_6666)
);

AOI21xp33_ASAP7_75t_SL g6667 ( 
.A1(n_6471),
.A2(n_756),
.B(n_748),
.Y(n_6667)
);

NAND2xp5_ASAP7_75t_L g6668 ( 
.A(n_6533),
.B(n_748),
.Y(n_6668)
);

INVx1_ASAP7_75t_L g6669 ( 
.A(n_6525),
.Y(n_6669)
);

INVx2_ASAP7_75t_L g6670 ( 
.A(n_6527),
.Y(n_6670)
);

AOI22xp33_ASAP7_75t_L g6671 ( 
.A1(n_6458),
.A2(n_751),
.B1(n_749),
.B2(n_750),
.Y(n_6671)
);

AND2x2_ASAP7_75t_L g6672 ( 
.A(n_6532),
.B(n_749),
.Y(n_6672)
);

INVx1_ASAP7_75t_L g6673 ( 
.A(n_6466),
.Y(n_6673)
);

NOR2xp33_ASAP7_75t_R g6674 ( 
.A(n_6438),
.B(n_6440),
.Y(n_6674)
);

NAND2xp5_ASAP7_75t_L g6675 ( 
.A(n_6501),
.B(n_750),
.Y(n_6675)
);

INVx1_ASAP7_75t_L g6676 ( 
.A(n_6510),
.Y(n_6676)
);

INVx2_ASAP7_75t_SL g6677 ( 
.A(n_6436),
.Y(n_6677)
);

INVx1_ASAP7_75t_L g6678 ( 
.A(n_6510),
.Y(n_6678)
);

INVx1_ASAP7_75t_L g6679 ( 
.A(n_6510),
.Y(n_6679)
);

AND2x2_ASAP7_75t_L g6680 ( 
.A(n_6432),
.B(n_751),
.Y(n_6680)
);

AND2x2_ASAP7_75t_L g6681 ( 
.A(n_6432),
.B(n_752),
.Y(n_6681)
);

HB1xp67_ASAP7_75t_L g6682 ( 
.A(n_6562),
.Y(n_6682)
);

INVxp33_ASAP7_75t_L g6683 ( 
.A(n_6571),
.Y(n_6683)
);

AND2x2_ASAP7_75t_L g6684 ( 
.A(n_6552),
.B(n_752),
.Y(n_6684)
);

NAND2xp5_ASAP7_75t_L g6685 ( 
.A(n_6588),
.B(n_753),
.Y(n_6685)
);

INVx1_ASAP7_75t_L g6686 ( 
.A(n_6600),
.Y(n_6686)
);

NAND2xp5_ASAP7_75t_L g6687 ( 
.A(n_6624),
.B(n_753),
.Y(n_6687)
);

INVx1_ASAP7_75t_L g6688 ( 
.A(n_6653),
.Y(n_6688)
);

AND2x2_ASAP7_75t_L g6689 ( 
.A(n_6680),
.B(n_6681),
.Y(n_6689)
);

NAND4xp25_ASAP7_75t_L g6690 ( 
.A(n_6621),
.B(n_757),
.C(n_754),
.D(n_755),
.Y(n_6690)
);

INVx1_ASAP7_75t_L g6691 ( 
.A(n_6619),
.Y(n_6691)
);

BUFx2_ASAP7_75t_L g6692 ( 
.A(n_6581),
.Y(n_6692)
);

OR2x2_ASAP7_75t_L g6693 ( 
.A(n_6565),
.B(n_6550),
.Y(n_6693)
);

INVx1_ASAP7_75t_SL g6694 ( 
.A(n_6557),
.Y(n_6694)
);

INVx1_ASAP7_75t_L g6695 ( 
.A(n_6622),
.Y(n_6695)
);

INVx1_ASAP7_75t_L g6696 ( 
.A(n_6567),
.Y(n_6696)
);

OR2x2_ASAP7_75t_L g6697 ( 
.A(n_6676),
.B(n_754),
.Y(n_6697)
);

NAND2xp5_ASAP7_75t_SL g6698 ( 
.A(n_6560),
.B(n_755),
.Y(n_6698)
);

AND2x2_ASAP7_75t_L g6699 ( 
.A(n_6576),
.B(n_757),
.Y(n_6699)
);

INVx1_ASAP7_75t_L g6700 ( 
.A(n_6582),
.Y(n_6700)
);

INVx1_ASAP7_75t_L g6701 ( 
.A(n_6612),
.Y(n_6701)
);

INVxp67_ASAP7_75t_L g6702 ( 
.A(n_6644),
.Y(n_6702)
);

AOI22xp5_ASAP7_75t_L g6703 ( 
.A1(n_6610),
.A2(n_760),
.B1(n_758),
.B2(n_759),
.Y(n_6703)
);

NAND2xp5_ASAP7_75t_L g6704 ( 
.A(n_6624),
.B(n_758),
.Y(n_6704)
);

INVx1_ASAP7_75t_L g6705 ( 
.A(n_6558),
.Y(n_6705)
);

AND2x4_ASAP7_75t_L g6706 ( 
.A(n_6581),
.B(n_759),
.Y(n_6706)
);

INVx1_ASAP7_75t_L g6707 ( 
.A(n_6658),
.Y(n_6707)
);

INVx1_ASAP7_75t_L g6708 ( 
.A(n_6660),
.Y(n_6708)
);

INVx1_ASAP7_75t_L g6709 ( 
.A(n_6649),
.Y(n_6709)
);

NOR2xp33_ASAP7_75t_L g6710 ( 
.A(n_6604),
.B(n_760),
.Y(n_6710)
);

OR2x2_ASAP7_75t_L g6711 ( 
.A(n_6678),
.B(n_761),
.Y(n_6711)
);

OR2x2_ASAP7_75t_L g6712 ( 
.A(n_6679),
.B(n_761),
.Y(n_6712)
);

OR2x2_ASAP7_75t_L g6713 ( 
.A(n_6587),
.B(n_762),
.Y(n_6713)
);

INVx1_ASAP7_75t_L g6714 ( 
.A(n_6599),
.Y(n_6714)
);

INVx1_ASAP7_75t_L g6715 ( 
.A(n_6584),
.Y(n_6715)
);

INVx1_ASAP7_75t_L g6716 ( 
.A(n_6632),
.Y(n_6716)
);

INVx2_ASAP7_75t_SL g6717 ( 
.A(n_6677),
.Y(n_6717)
);

INVx2_ASAP7_75t_L g6718 ( 
.A(n_6577),
.Y(n_6718)
);

NOR2xp33_ASAP7_75t_L g6719 ( 
.A(n_6556),
.B(n_762),
.Y(n_6719)
);

AND2x2_ASAP7_75t_L g6720 ( 
.A(n_6601),
.B(n_763),
.Y(n_6720)
);

HB1xp67_ASAP7_75t_L g6721 ( 
.A(n_6585),
.Y(n_6721)
);

HB1xp67_ASAP7_75t_L g6722 ( 
.A(n_6615),
.Y(n_6722)
);

NAND2xp5_ASAP7_75t_L g6723 ( 
.A(n_6593),
.B(n_763),
.Y(n_6723)
);

AND2x2_ASAP7_75t_L g6724 ( 
.A(n_6559),
.B(n_764),
.Y(n_6724)
);

AND2x2_ASAP7_75t_L g6725 ( 
.A(n_6553),
.B(n_765),
.Y(n_6725)
);

AND2x2_ASAP7_75t_L g6726 ( 
.A(n_6586),
.B(n_766),
.Y(n_6726)
);

AND2x2_ASAP7_75t_L g6727 ( 
.A(n_6627),
.B(n_767),
.Y(n_6727)
);

AND2x2_ASAP7_75t_L g6728 ( 
.A(n_6564),
.B(n_767),
.Y(n_6728)
);

INVx1_ASAP7_75t_L g6729 ( 
.A(n_6590),
.Y(n_6729)
);

INVx1_ASAP7_75t_L g6730 ( 
.A(n_6651),
.Y(n_6730)
);

AND2x2_ASAP7_75t_L g6731 ( 
.A(n_6654),
.B(n_769),
.Y(n_6731)
);

INVx1_ASAP7_75t_SL g6732 ( 
.A(n_6631),
.Y(n_6732)
);

INVx1_ASAP7_75t_L g6733 ( 
.A(n_6662),
.Y(n_6733)
);

INVx1_ASAP7_75t_L g6734 ( 
.A(n_6664),
.Y(n_6734)
);

INVx1_ASAP7_75t_L g6735 ( 
.A(n_6666),
.Y(n_6735)
);

AND2x2_ASAP7_75t_L g6736 ( 
.A(n_6672),
.B(n_769),
.Y(n_6736)
);

INVx1_ASAP7_75t_L g6737 ( 
.A(n_6555),
.Y(n_6737)
);

AND2x2_ASAP7_75t_L g6738 ( 
.A(n_6566),
.B(n_770),
.Y(n_6738)
);

INVx2_ASAP7_75t_L g6739 ( 
.A(n_6589),
.Y(n_6739)
);

OAI31xp33_ASAP7_75t_SL g6740 ( 
.A1(n_6635),
.A2(n_774),
.A3(n_775),
.B(n_772),
.Y(n_6740)
);

INVx1_ASAP7_75t_L g6741 ( 
.A(n_6675),
.Y(n_6741)
);

NAND2xp5_ASAP7_75t_SL g6742 ( 
.A(n_6563),
.B(n_771),
.Y(n_6742)
);

AND2x2_ASAP7_75t_L g6743 ( 
.A(n_6602),
.B(n_777),
.Y(n_6743)
);

INVxp67_ASAP7_75t_SL g6744 ( 
.A(n_6618),
.Y(n_6744)
);

AND2x2_ASAP7_75t_L g6745 ( 
.A(n_6648),
.B(n_777),
.Y(n_6745)
);

NAND2xp5_ASAP7_75t_L g6746 ( 
.A(n_6639),
.B(n_778),
.Y(n_6746)
);

INVx1_ASAP7_75t_L g6747 ( 
.A(n_6583),
.Y(n_6747)
);

INVx1_ASAP7_75t_L g6748 ( 
.A(n_6634),
.Y(n_6748)
);

INVx1_ASAP7_75t_L g6749 ( 
.A(n_6616),
.Y(n_6749)
);

NAND2xp5_ASAP7_75t_L g6750 ( 
.A(n_6573),
.B(n_779),
.Y(n_6750)
);

INVx1_ASAP7_75t_L g6751 ( 
.A(n_6605),
.Y(n_6751)
);

HB1xp67_ASAP7_75t_L g6752 ( 
.A(n_6569),
.Y(n_6752)
);

AND2x4_ASAP7_75t_L g6753 ( 
.A(n_6580),
.B(n_780),
.Y(n_6753)
);

NAND2xp5_ASAP7_75t_L g6754 ( 
.A(n_6607),
.B(n_780),
.Y(n_6754)
);

OR2x2_ASAP7_75t_L g6755 ( 
.A(n_6592),
.B(n_781),
.Y(n_6755)
);

OR2x2_ASAP7_75t_L g6756 ( 
.A(n_6598),
.B(n_781),
.Y(n_6756)
);

OR2x2_ASAP7_75t_L g6757 ( 
.A(n_6668),
.B(n_782),
.Y(n_6757)
);

AND2x2_ASAP7_75t_L g6758 ( 
.A(n_6575),
.B(n_783),
.Y(n_6758)
);

INVx2_ASAP7_75t_L g6759 ( 
.A(n_6650),
.Y(n_6759)
);

AND2x2_ASAP7_75t_L g6760 ( 
.A(n_6670),
.B(n_784),
.Y(n_6760)
);

OR2x4_ASAP7_75t_L g6761 ( 
.A(n_6551),
.B(n_785),
.Y(n_6761)
);

OR2x2_ASAP7_75t_L g6762 ( 
.A(n_6652),
.B(n_6625),
.Y(n_6762)
);

OR2x2_ASAP7_75t_L g6763 ( 
.A(n_6596),
.B(n_785),
.Y(n_6763)
);

INVx1_ASAP7_75t_L g6764 ( 
.A(n_6645),
.Y(n_6764)
);

INVx1_ASAP7_75t_L g6765 ( 
.A(n_6597),
.Y(n_6765)
);

NAND2x1_ASAP7_75t_L g6766 ( 
.A(n_6628),
.B(n_786),
.Y(n_6766)
);

INVxp67_ASAP7_75t_L g6767 ( 
.A(n_6561),
.Y(n_6767)
);

INVx2_ASAP7_75t_L g6768 ( 
.A(n_6613),
.Y(n_6768)
);

AND2x2_ASAP7_75t_L g6769 ( 
.A(n_6623),
.B(n_786),
.Y(n_6769)
);

NAND2xp5_ASAP7_75t_L g6770 ( 
.A(n_6614),
.B(n_787),
.Y(n_6770)
);

NAND2xp5_ASAP7_75t_L g6771 ( 
.A(n_6626),
.B(n_787),
.Y(n_6771)
);

NAND2xp5_ASAP7_75t_L g6772 ( 
.A(n_6633),
.B(n_788),
.Y(n_6772)
);

AOI22xp33_ASAP7_75t_SL g6773 ( 
.A1(n_6674),
.A2(n_793),
.B1(n_789),
.B2(n_791),
.Y(n_6773)
);

INVx1_ASAP7_75t_L g6774 ( 
.A(n_6595),
.Y(n_6774)
);

INVx1_ASAP7_75t_L g6775 ( 
.A(n_6579),
.Y(n_6775)
);

NAND2xp5_ASAP7_75t_L g6776 ( 
.A(n_6603),
.B(n_6665),
.Y(n_6776)
);

AND2x2_ASAP7_75t_L g6777 ( 
.A(n_6640),
.B(n_6641),
.Y(n_6777)
);

INVxp67_ASAP7_75t_L g6778 ( 
.A(n_6609),
.Y(n_6778)
);

INVx1_ASAP7_75t_L g6779 ( 
.A(n_6617),
.Y(n_6779)
);

NAND2xp5_ASAP7_75t_L g6780 ( 
.A(n_6554),
.B(n_6667),
.Y(n_6780)
);

NAND2xp5_ASAP7_75t_L g6781 ( 
.A(n_6570),
.B(n_793),
.Y(n_6781)
);

INVxp67_ASAP7_75t_L g6782 ( 
.A(n_6656),
.Y(n_6782)
);

AND2x2_ASAP7_75t_L g6783 ( 
.A(n_6642),
.B(n_794),
.Y(n_6783)
);

OR2x2_ASAP7_75t_L g6784 ( 
.A(n_6608),
.B(n_795),
.Y(n_6784)
);

AND2x2_ASAP7_75t_L g6785 ( 
.A(n_6643),
.B(n_796),
.Y(n_6785)
);

INVx1_ASAP7_75t_L g6786 ( 
.A(n_6659),
.Y(n_6786)
);

CKINVDCx5p33_ASAP7_75t_R g6787 ( 
.A(n_6636),
.Y(n_6787)
);

NAND2xp5_ASAP7_75t_L g6788 ( 
.A(n_6673),
.B(n_796),
.Y(n_6788)
);

NAND2xp5_ASAP7_75t_L g6789 ( 
.A(n_6671),
.B(n_6638),
.Y(n_6789)
);

INVx1_ASAP7_75t_L g6790 ( 
.A(n_6620),
.Y(n_6790)
);

AND2x2_ASAP7_75t_L g6791 ( 
.A(n_6646),
.B(n_797),
.Y(n_6791)
);

AND2x2_ASAP7_75t_L g6792 ( 
.A(n_6647),
.B(n_6663),
.Y(n_6792)
);

OR2x6_ASAP7_75t_L g6793 ( 
.A(n_6578),
.B(n_798),
.Y(n_6793)
);

INVx2_ASAP7_75t_L g6794 ( 
.A(n_6591),
.Y(n_6794)
);

INVx1_ASAP7_75t_L g6795 ( 
.A(n_6629),
.Y(n_6795)
);

NAND2xp5_ASAP7_75t_L g6796 ( 
.A(n_6630),
.B(n_799),
.Y(n_6796)
);

HB1xp67_ASAP7_75t_L g6797 ( 
.A(n_6606),
.Y(n_6797)
);

INVx1_ASAP7_75t_L g6798 ( 
.A(n_6568),
.Y(n_6798)
);

AND2x2_ASAP7_75t_L g6799 ( 
.A(n_6669),
.B(n_800),
.Y(n_6799)
);

INVx1_ASAP7_75t_L g6800 ( 
.A(n_6661),
.Y(n_6800)
);

INVx1_ASAP7_75t_L g6801 ( 
.A(n_6574),
.Y(n_6801)
);

AND2x2_ASAP7_75t_L g6802 ( 
.A(n_6611),
.B(n_800),
.Y(n_6802)
);

NAND2xp5_ASAP7_75t_L g6803 ( 
.A(n_6655),
.B(n_6594),
.Y(n_6803)
);

BUFx2_ASAP7_75t_L g6804 ( 
.A(n_6572),
.Y(n_6804)
);

INVx2_ASAP7_75t_L g6805 ( 
.A(n_6657),
.Y(n_6805)
);

INVx1_ASAP7_75t_L g6806 ( 
.A(n_6637),
.Y(n_6806)
);

AND2x2_ASAP7_75t_L g6807 ( 
.A(n_6552),
.B(n_801),
.Y(n_6807)
);

NAND2xp5_ASAP7_75t_L g6808 ( 
.A(n_6588),
.B(n_802),
.Y(n_6808)
);

NAND2x1p5_ASAP7_75t_L g6809 ( 
.A(n_6624),
.B(n_802),
.Y(n_6809)
);

INVx1_ASAP7_75t_L g6810 ( 
.A(n_6600),
.Y(n_6810)
);

INVx2_ASAP7_75t_L g6811 ( 
.A(n_6577),
.Y(n_6811)
);

NAND2xp5_ASAP7_75t_L g6812 ( 
.A(n_6588),
.B(n_804),
.Y(n_6812)
);

INVx1_ASAP7_75t_L g6813 ( 
.A(n_6600),
.Y(n_6813)
);

INVx2_ASAP7_75t_SL g6814 ( 
.A(n_6581),
.Y(n_6814)
);

INVx2_ASAP7_75t_SL g6815 ( 
.A(n_6581),
.Y(n_6815)
);

NAND2xp5_ASAP7_75t_L g6816 ( 
.A(n_6588),
.B(n_804),
.Y(n_6816)
);

AND2x2_ASAP7_75t_L g6817 ( 
.A(n_6552),
.B(n_805),
.Y(n_6817)
);

NAND2xp5_ASAP7_75t_L g6818 ( 
.A(n_6588),
.B(n_806),
.Y(n_6818)
);

CKINVDCx16_ASAP7_75t_R g6819 ( 
.A(n_6557),
.Y(n_6819)
);

INVx1_ASAP7_75t_L g6820 ( 
.A(n_6600),
.Y(n_6820)
);

AND2x2_ASAP7_75t_L g6821 ( 
.A(n_6552),
.B(n_806),
.Y(n_6821)
);

INVx2_ASAP7_75t_SL g6822 ( 
.A(n_6581),
.Y(n_6822)
);

AOI222xp33_ASAP7_75t_L g6823 ( 
.A1(n_6604),
.A2(n_813),
.B1(n_815),
.B2(n_808),
.C1(n_810),
.C2(n_814),
.Y(n_6823)
);

INVx1_ASAP7_75t_SL g6824 ( 
.A(n_6571),
.Y(n_6824)
);

INVx2_ASAP7_75t_L g6825 ( 
.A(n_6577),
.Y(n_6825)
);

INVx2_ASAP7_75t_L g6826 ( 
.A(n_6577),
.Y(n_6826)
);

NAND2xp5_ASAP7_75t_L g6827 ( 
.A(n_6588),
.B(n_808),
.Y(n_6827)
);

INVx1_ASAP7_75t_L g6828 ( 
.A(n_6600),
.Y(n_6828)
);

INVx2_ASAP7_75t_L g6829 ( 
.A(n_6577),
.Y(n_6829)
);

AND2x2_ASAP7_75t_L g6830 ( 
.A(n_6552),
.B(n_810),
.Y(n_6830)
);

OR2x2_ASAP7_75t_L g6831 ( 
.A(n_6565),
.B(n_813),
.Y(n_6831)
);

AND2x2_ASAP7_75t_SL g6832 ( 
.A(n_6614),
.B(n_814),
.Y(n_6832)
);

INVx2_ASAP7_75t_L g6833 ( 
.A(n_6577),
.Y(n_6833)
);

AND2x2_ASAP7_75t_L g6834 ( 
.A(n_6552),
.B(n_815),
.Y(n_6834)
);

AND2x2_ASAP7_75t_L g6835 ( 
.A(n_6552),
.B(n_816),
.Y(n_6835)
);

INVx1_ASAP7_75t_L g6836 ( 
.A(n_6600),
.Y(n_6836)
);

INVx4_ASAP7_75t_L g6837 ( 
.A(n_6553),
.Y(n_6837)
);

NAND2xp33_ASAP7_75t_L g6838 ( 
.A(n_6565),
.B(n_816),
.Y(n_6838)
);

AND2x2_ASAP7_75t_L g6839 ( 
.A(n_6552),
.B(n_817),
.Y(n_6839)
);

AND2x2_ASAP7_75t_L g6840 ( 
.A(n_6552),
.B(n_817),
.Y(n_6840)
);

NOR2xp33_ASAP7_75t_L g6841 ( 
.A(n_6604),
.B(n_818),
.Y(n_6841)
);

AND2x4_ASAP7_75t_SL g6842 ( 
.A(n_6621),
.B(n_818),
.Y(n_6842)
);

INVx1_ASAP7_75t_L g6843 ( 
.A(n_6600),
.Y(n_6843)
);

OR2x2_ASAP7_75t_L g6844 ( 
.A(n_6565),
.B(n_819),
.Y(n_6844)
);

INVxp67_ASAP7_75t_L g6845 ( 
.A(n_6644),
.Y(n_6845)
);

INVx2_ASAP7_75t_L g6846 ( 
.A(n_6577),
.Y(n_6846)
);

INVx2_ASAP7_75t_L g6847 ( 
.A(n_6577),
.Y(n_6847)
);

OR2x2_ASAP7_75t_L g6848 ( 
.A(n_6565),
.B(n_819),
.Y(n_6848)
);

NAND2xp33_ASAP7_75t_L g6849 ( 
.A(n_6565),
.B(n_820),
.Y(n_6849)
);

NOR2x1_ASAP7_75t_L g6850 ( 
.A(n_6592),
.B(n_821),
.Y(n_6850)
);

INVx1_ASAP7_75t_L g6851 ( 
.A(n_6600),
.Y(n_6851)
);

INVx1_ASAP7_75t_SL g6852 ( 
.A(n_6571),
.Y(n_6852)
);

AOI22xp5_ASAP7_75t_L g6853 ( 
.A1(n_6644),
.A2(n_823),
.B1(n_821),
.B2(n_822),
.Y(n_6853)
);

INVx2_ASAP7_75t_L g6854 ( 
.A(n_6577),
.Y(n_6854)
);

BUFx3_ASAP7_75t_L g6855 ( 
.A(n_6621),
.Y(n_6855)
);

NAND2x1p5_ASAP7_75t_L g6856 ( 
.A(n_6624),
.B(n_822),
.Y(n_6856)
);

INVxp67_ASAP7_75t_SL g6857 ( 
.A(n_6604),
.Y(n_6857)
);

NAND2xp5_ASAP7_75t_L g6858 ( 
.A(n_6588),
.B(n_823),
.Y(n_6858)
);

OR2x2_ASAP7_75t_L g6859 ( 
.A(n_6565),
.B(n_824),
.Y(n_6859)
);

INVx3_ASAP7_75t_L g6860 ( 
.A(n_6581),
.Y(n_6860)
);

NOR2xp33_ASAP7_75t_L g6861 ( 
.A(n_6604),
.B(n_824),
.Y(n_6861)
);

AND2x2_ASAP7_75t_L g6862 ( 
.A(n_6552),
.B(n_825),
.Y(n_6862)
);

AND2x2_ASAP7_75t_L g6863 ( 
.A(n_6552),
.B(n_825),
.Y(n_6863)
);

INVx2_ASAP7_75t_L g6864 ( 
.A(n_6577),
.Y(n_6864)
);

INVx1_ASAP7_75t_L g6865 ( 
.A(n_6600),
.Y(n_6865)
);

NOR2x1_ASAP7_75t_L g6866 ( 
.A(n_6592),
.B(n_826),
.Y(n_6866)
);

INVx1_ASAP7_75t_SL g6867 ( 
.A(n_6571),
.Y(n_6867)
);

INVx1_ASAP7_75t_L g6868 ( 
.A(n_6600),
.Y(n_6868)
);

INVx1_ASAP7_75t_L g6869 ( 
.A(n_6600),
.Y(n_6869)
);

INVx1_ASAP7_75t_SL g6870 ( 
.A(n_6571),
.Y(n_6870)
);

AND2x4_ASAP7_75t_L g6871 ( 
.A(n_6581),
.B(n_826),
.Y(n_6871)
);

NAND4xp25_ASAP7_75t_L g6872 ( 
.A(n_6621),
.B(n_829),
.C(n_827),
.D(n_828),
.Y(n_6872)
);

AND2x2_ASAP7_75t_L g6873 ( 
.A(n_6552),
.B(n_828),
.Y(n_6873)
);

NOR2xp33_ASAP7_75t_R g6874 ( 
.A(n_6855),
.B(n_830),
.Y(n_6874)
);

OAI21xp33_ASAP7_75t_L g6875 ( 
.A1(n_6857),
.A2(n_830),
.B(n_831),
.Y(n_6875)
);

INVx1_ASAP7_75t_L g6876 ( 
.A(n_6692),
.Y(n_6876)
);

INVxp67_ASAP7_75t_L g6877 ( 
.A(n_6721),
.Y(n_6877)
);

OAI21xp5_ASAP7_75t_L g6878 ( 
.A1(n_6850),
.A2(n_831),
.B(n_832),
.Y(n_6878)
);

INVx2_ASAP7_75t_L g6879 ( 
.A(n_6809),
.Y(n_6879)
);

INVx1_ASAP7_75t_L g6880 ( 
.A(n_6682),
.Y(n_6880)
);

INVx1_ASAP7_75t_L g6881 ( 
.A(n_6752),
.Y(n_6881)
);

AOI221xp5_ASAP7_75t_L g6882 ( 
.A1(n_6729),
.A2(n_835),
.B1(n_833),
.B2(n_834),
.C(n_837),
.Y(n_6882)
);

INVx1_ASAP7_75t_L g6883 ( 
.A(n_6860),
.Y(n_6883)
);

HB1xp67_ASAP7_75t_L g6884 ( 
.A(n_6689),
.Y(n_6884)
);

NOR2xp33_ASAP7_75t_L g6885 ( 
.A(n_6819),
.B(n_834),
.Y(n_6885)
);

AOI22xp33_ASAP7_75t_L g6886 ( 
.A1(n_6786),
.A2(n_840),
.B1(n_837),
.B2(n_838),
.Y(n_6886)
);

INVx1_ASAP7_75t_L g6887 ( 
.A(n_6814),
.Y(n_6887)
);

NAND2xp5_ASAP7_75t_L g6888 ( 
.A(n_6702),
.B(n_838),
.Y(n_6888)
);

AND2x2_ASAP7_75t_L g6889 ( 
.A(n_6815),
.B(n_840),
.Y(n_6889)
);

INVx1_ASAP7_75t_L g6890 ( 
.A(n_6822),
.Y(n_6890)
);

INVx1_ASAP7_75t_L g6891 ( 
.A(n_6727),
.Y(n_6891)
);

INVx1_ASAP7_75t_L g6892 ( 
.A(n_6831),
.Y(n_6892)
);

AOI21xp33_ASAP7_75t_L g6893 ( 
.A1(n_6683),
.A2(n_841),
.B(n_842),
.Y(n_6893)
);

OAI22xp5_ASAP7_75t_L g6894 ( 
.A1(n_6686),
.A2(n_843),
.B1(n_841),
.B2(n_842),
.Y(n_6894)
);

OR2x2_ASAP7_75t_L g6895 ( 
.A(n_6693),
.B(n_843),
.Y(n_6895)
);

INVx2_ASAP7_75t_L g6896 ( 
.A(n_6856),
.Y(n_6896)
);

INVx1_ASAP7_75t_SL g6897 ( 
.A(n_6824),
.Y(n_6897)
);

OAI322xp33_ASAP7_75t_L g6898 ( 
.A1(n_6762),
.A2(n_849),
.A3(n_848),
.B1(n_846),
.B2(n_844),
.C1(n_845),
.C2(n_847),
.Y(n_6898)
);

AOI22xp5_ASAP7_75t_L g6899 ( 
.A1(n_6852),
.A2(n_6870),
.B1(n_6867),
.B2(n_6694),
.Y(n_6899)
);

OAI22xp33_ASAP7_75t_SL g6900 ( 
.A1(n_6845),
.A2(n_849),
.B1(n_847),
.B2(n_848),
.Y(n_6900)
);

INVx1_ASAP7_75t_SL g6901 ( 
.A(n_6732),
.Y(n_6901)
);

NAND2xp5_ASAP7_75t_L g6902 ( 
.A(n_6767),
.B(n_850),
.Y(n_6902)
);

INVx1_ASAP7_75t_L g6903 ( 
.A(n_6844),
.Y(n_6903)
);

INVx2_ASAP7_75t_L g6904 ( 
.A(n_6718),
.Y(n_6904)
);

OAI21xp33_ASAP7_75t_L g6905 ( 
.A1(n_6810),
.A2(n_850),
.B(n_851),
.Y(n_6905)
);

INVxp33_ASAP7_75t_L g6906 ( 
.A(n_6722),
.Y(n_6906)
);

NAND2xp5_ASAP7_75t_L g6907 ( 
.A(n_6684),
.B(n_851),
.Y(n_6907)
);

A2O1A1Ixp33_ASAP7_75t_L g6908 ( 
.A1(n_6740),
.A2(n_854),
.B(n_852),
.C(n_853),
.Y(n_6908)
);

AOI21xp5_ASAP7_75t_L g6909 ( 
.A1(n_6838),
.A2(n_852),
.B(n_853),
.Y(n_6909)
);

NAND2xp5_ASAP7_75t_L g6910 ( 
.A(n_6807),
.B(n_855),
.Y(n_6910)
);

OAI22xp5_ASAP7_75t_L g6911 ( 
.A1(n_6813),
.A2(n_858),
.B1(n_856),
.B2(n_857),
.Y(n_6911)
);

OAI211xp5_ASAP7_75t_L g6912 ( 
.A1(n_6820),
.A2(n_860),
.B(n_856),
.C(n_858),
.Y(n_6912)
);

NAND2x1p5_ASAP7_75t_L g6913 ( 
.A(n_6837),
.B(n_862),
.Y(n_6913)
);

INVx2_ASAP7_75t_L g6914 ( 
.A(n_6811),
.Y(n_6914)
);

INVx1_ASAP7_75t_L g6915 ( 
.A(n_6848),
.Y(n_6915)
);

AOI311xp33_ASAP7_75t_L g6916 ( 
.A1(n_6700),
.A2(n_6828),
.A3(n_6851),
.B(n_6843),
.C(n_6836),
.Y(n_6916)
);

AOI33xp33_ASAP7_75t_L g6917 ( 
.A1(n_6865),
.A2(n_863),
.A3(n_865),
.B1(n_861),
.B2(n_862),
.B3(n_864),
.Y(n_6917)
);

AND2x2_ASAP7_75t_L g6918 ( 
.A(n_6868),
.B(n_863),
.Y(n_6918)
);

OAI33xp33_ASAP7_75t_L g6919 ( 
.A1(n_6800),
.A2(n_866),
.A3(n_869),
.B1(n_864),
.B2(n_865),
.B3(n_868),
.Y(n_6919)
);

NAND2xp5_ASAP7_75t_L g6920 ( 
.A(n_6817),
.B(n_866),
.Y(n_6920)
);

INVx2_ASAP7_75t_L g6921 ( 
.A(n_6825),
.Y(n_6921)
);

NAND2xp5_ASAP7_75t_L g6922 ( 
.A(n_6821),
.B(n_868),
.Y(n_6922)
);

INVx2_ASAP7_75t_L g6923 ( 
.A(n_6826),
.Y(n_6923)
);

OAI21xp5_ASAP7_75t_SL g6924 ( 
.A1(n_6869),
.A2(n_6717),
.B(n_6804),
.Y(n_6924)
);

OR2x2_ASAP7_75t_L g6925 ( 
.A(n_6859),
.B(n_869),
.Y(n_6925)
);

NAND2xp5_ASAP7_75t_L g6926 ( 
.A(n_6830),
.B(n_870),
.Y(n_6926)
);

AND2x2_ASAP7_75t_L g6927 ( 
.A(n_6699),
.B(n_871),
.Y(n_6927)
);

INVx1_ASAP7_75t_L g6928 ( 
.A(n_6834),
.Y(n_6928)
);

INVx3_ASAP7_75t_L g6929 ( 
.A(n_6706),
.Y(n_6929)
);

INVxp67_ASAP7_75t_SL g6930 ( 
.A(n_6766),
.Y(n_6930)
);

NAND3xp33_ASAP7_75t_L g6931 ( 
.A(n_6849),
.B(n_872),
.C(n_873),
.Y(n_6931)
);

INVx1_ASAP7_75t_SL g6932 ( 
.A(n_6842),
.Y(n_6932)
);

INVx1_ASAP7_75t_L g6933 ( 
.A(n_6835),
.Y(n_6933)
);

INVx1_ASAP7_75t_L g6934 ( 
.A(n_6839),
.Y(n_6934)
);

XOR2x2_ASAP7_75t_L g6935 ( 
.A(n_6866),
.B(n_872),
.Y(n_6935)
);

NAND2xp5_ASAP7_75t_L g6936 ( 
.A(n_6840),
.B(n_874),
.Y(n_6936)
);

INVx1_ASAP7_75t_L g6937 ( 
.A(n_6862),
.Y(n_6937)
);

AOI22xp5_ASAP7_75t_L g6938 ( 
.A1(n_6778),
.A2(n_876),
.B1(n_874),
.B2(n_875),
.Y(n_6938)
);

OAI22xp33_ASAP7_75t_L g6939 ( 
.A1(n_6761),
.A2(n_879),
.B1(n_877),
.B2(n_878),
.Y(n_6939)
);

AND2x2_ASAP7_75t_L g6940 ( 
.A(n_6720),
.B(n_880),
.Y(n_6940)
);

INVx1_ASAP7_75t_L g6941 ( 
.A(n_6863),
.Y(n_6941)
);

AOI221xp5_ASAP7_75t_L g6942 ( 
.A1(n_6806),
.A2(n_883),
.B1(n_881),
.B2(n_882),
.C(n_884),
.Y(n_6942)
);

INVxp33_ASAP7_75t_L g6943 ( 
.A(n_6829),
.Y(n_6943)
);

OAI22xp33_ASAP7_75t_L g6944 ( 
.A1(n_6853),
.A2(n_884),
.B1(n_881),
.B2(n_882),
.Y(n_6944)
);

OAI21xp33_ASAP7_75t_L g6945 ( 
.A1(n_6801),
.A2(n_886),
.B(n_887),
.Y(n_6945)
);

AOI222xp33_ASAP7_75t_L g6946 ( 
.A1(n_6744),
.A2(n_888),
.B1(n_891),
.B2(n_886),
.C1(n_887),
.C2(n_889),
.Y(n_6946)
);

INVx1_ASAP7_75t_L g6947 ( 
.A(n_6873),
.Y(n_6947)
);

OAI32xp33_ASAP7_75t_L g6948 ( 
.A1(n_6776),
.A2(n_893),
.A3(n_888),
.B1(n_892),
.B2(n_894),
.Y(n_6948)
);

O2A1O1Ixp5_ASAP7_75t_L g6949 ( 
.A1(n_6739),
.A2(n_897),
.B(n_895),
.C(n_896),
.Y(n_6949)
);

OAI21xp33_ASAP7_75t_L g6950 ( 
.A1(n_6730),
.A2(n_895),
.B(n_896),
.Y(n_6950)
);

INVx1_ASAP7_75t_L g6951 ( 
.A(n_6743),
.Y(n_6951)
);

NOR2xp33_ASAP7_75t_L g6952 ( 
.A(n_6690),
.B(n_6872),
.Y(n_6952)
);

AOI21xp33_ASAP7_75t_L g6953 ( 
.A1(n_6833),
.A2(n_897),
.B(n_898),
.Y(n_6953)
);

INVx1_ASAP7_75t_L g6954 ( 
.A(n_6731),
.Y(n_6954)
);

INVx1_ASAP7_75t_L g6955 ( 
.A(n_6736),
.Y(n_6955)
);

AOI221xp5_ASAP7_75t_L g6956 ( 
.A1(n_6782),
.A2(n_6749),
.B1(n_6803),
.B2(n_6797),
.C(n_6774),
.Y(n_6956)
);

INVx1_ASAP7_75t_L g6957 ( 
.A(n_6691),
.Y(n_6957)
);

OAI21xp5_ASAP7_75t_L g6958 ( 
.A1(n_6710),
.A2(n_898),
.B(n_899),
.Y(n_6958)
);

INVx1_ASAP7_75t_L g6959 ( 
.A(n_6695),
.Y(n_6959)
);

OAI21xp33_ASAP7_75t_L g6960 ( 
.A1(n_6733),
.A2(n_900),
.B(n_901),
.Y(n_6960)
);

A2O1A1Ixp33_ASAP7_75t_L g6961 ( 
.A1(n_6719),
.A2(n_903),
.B(n_901),
.C(n_902),
.Y(n_6961)
);

OAI222xp33_ASAP7_75t_L g6962 ( 
.A1(n_6846),
.A2(n_6854),
.B1(n_6864),
.B2(n_6847),
.C1(n_6773),
.C2(n_6798),
.Y(n_6962)
);

AO22x1_ASAP7_75t_L g6963 ( 
.A1(n_6841),
.A2(n_906),
.B1(n_902),
.B2(n_905),
.Y(n_6963)
);

AO22x1_ASAP7_75t_L g6964 ( 
.A1(n_6861),
.A2(n_909),
.B1(n_907),
.B2(n_908),
.Y(n_6964)
);

INVx1_ASAP7_75t_L g6965 ( 
.A(n_6709),
.Y(n_6965)
);

AOI22xp5_ASAP7_75t_L g6966 ( 
.A1(n_6737),
.A2(n_910),
.B1(n_907),
.B2(n_909),
.Y(n_6966)
);

INVx1_ASAP7_75t_L g6967 ( 
.A(n_6685),
.Y(n_6967)
);

OR2x2_ASAP7_75t_L g6968 ( 
.A(n_6713),
.B(n_911),
.Y(n_6968)
);

NAND2xp5_ASAP7_75t_SL g6969 ( 
.A(n_6832),
.B(n_911),
.Y(n_6969)
);

OAI22xp5_ASAP7_75t_L g6970 ( 
.A1(n_6759),
.A2(n_914),
.B1(n_912),
.B2(n_913),
.Y(n_6970)
);

NAND2xp5_ASAP7_75t_SL g6971 ( 
.A(n_6871),
.B(n_912),
.Y(n_6971)
);

OR2x2_ASAP7_75t_L g6972 ( 
.A(n_6808),
.B(n_915),
.Y(n_6972)
);

AOI22xp5_ASAP7_75t_L g6973 ( 
.A1(n_6741),
.A2(n_917),
.B1(n_915),
.B2(n_916),
.Y(n_6973)
);

INVx2_ASAP7_75t_SL g6974 ( 
.A(n_6725),
.Y(n_6974)
);

O2A1O1Ixp33_ASAP7_75t_L g6975 ( 
.A1(n_6772),
.A2(n_918),
.B(n_916),
.C(n_917),
.Y(n_6975)
);

INVxp67_ASAP7_75t_L g6976 ( 
.A(n_6726),
.Y(n_6976)
);

OAI21xp33_ASAP7_75t_L g6977 ( 
.A1(n_6734),
.A2(n_918),
.B(n_920),
.Y(n_6977)
);

INVx2_ASAP7_75t_L g6978 ( 
.A(n_6753),
.Y(n_6978)
);

NAND2xp5_ASAP7_75t_L g6979 ( 
.A(n_6738),
.B(n_920),
.Y(n_6979)
);

INVx1_ASAP7_75t_L g6980 ( 
.A(n_6812),
.Y(n_6980)
);

NOR2xp33_ASAP7_75t_L g6981 ( 
.A(n_6698),
.B(n_921),
.Y(n_6981)
);

AOI21xp33_ASAP7_75t_SL g6982 ( 
.A1(n_6816),
.A2(n_924),
.B(n_923),
.Y(n_6982)
);

INVx1_ASAP7_75t_L g6983 ( 
.A(n_6818),
.Y(n_6983)
);

NAND2xp5_ASAP7_75t_L g6984 ( 
.A(n_6758),
.B(n_921),
.Y(n_6984)
);

OAI222xp33_ASAP7_75t_L g6985 ( 
.A1(n_6780),
.A2(n_6703),
.B1(n_6789),
.B2(n_6688),
.C1(n_6705),
.C2(n_6701),
.Y(n_6985)
);

O2A1O1Ixp33_ASAP7_75t_L g6986 ( 
.A1(n_6770),
.A2(n_925),
.B(n_923),
.C(n_924),
.Y(n_6986)
);

OR2x2_ASAP7_75t_L g6987 ( 
.A(n_6827),
.B(n_925),
.Y(n_6987)
);

INVx1_ASAP7_75t_L g6988 ( 
.A(n_6858),
.Y(n_6988)
);

NAND2xp5_ASAP7_75t_L g6989 ( 
.A(n_6724),
.B(n_926),
.Y(n_6989)
);

INVx1_ASAP7_75t_SL g6990 ( 
.A(n_6728),
.Y(n_6990)
);

INVx1_ASAP7_75t_L g6991 ( 
.A(n_6783),
.Y(n_6991)
);

AOI22xp5_ASAP7_75t_L g6992 ( 
.A1(n_6715),
.A2(n_931),
.B1(n_927),
.B2(n_930),
.Y(n_6992)
);

OR2x2_ASAP7_75t_L g6993 ( 
.A(n_6779),
.B(n_927),
.Y(n_6993)
);

NAND2x1_ASAP7_75t_L g6994 ( 
.A(n_6777),
.B(n_930),
.Y(n_6994)
);

AOI22xp5_ASAP7_75t_L g6995 ( 
.A1(n_6787),
.A2(n_6696),
.B1(n_6714),
.B2(n_6707),
.Y(n_6995)
);

NOR2xp33_ASAP7_75t_L g6996 ( 
.A(n_6742),
.B(n_931),
.Y(n_6996)
);

CKINVDCx14_ASAP7_75t_R g6997 ( 
.A(n_6745),
.Y(n_6997)
);

NAND2xp5_ASAP7_75t_SL g6998 ( 
.A(n_6735),
.B(n_932),
.Y(n_6998)
);

AND2x2_ASAP7_75t_L g6999 ( 
.A(n_6792),
.B(n_6747),
.Y(n_6999)
);

INVx1_ASAP7_75t_L g7000 ( 
.A(n_6785),
.Y(n_7000)
);

NAND2x1p5_ASAP7_75t_L g7001 ( 
.A(n_6760),
.B(n_6802),
.Y(n_7001)
);

INVx1_ASAP7_75t_L g7002 ( 
.A(n_6791),
.Y(n_7002)
);

OAI221xp5_ASAP7_75t_L g7003 ( 
.A1(n_6708),
.A2(n_934),
.B1(n_932),
.B2(n_933),
.C(n_935),
.Y(n_7003)
);

BUFx2_ASAP7_75t_L g7004 ( 
.A(n_6769),
.Y(n_7004)
);

INVx1_ASAP7_75t_L g7005 ( 
.A(n_6799),
.Y(n_7005)
);

INVx1_ASAP7_75t_L g7006 ( 
.A(n_6756),
.Y(n_7006)
);

AOI22xp5_ASAP7_75t_L g7007 ( 
.A1(n_6765),
.A2(n_935),
.B1(n_933),
.B2(n_934),
.Y(n_7007)
);

XOR2x2_ASAP7_75t_L g7008 ( 
.A(n_6723),
.B(n_936),
.Y(n_7008)
);

AOI21xp33_ASAP7_75t_L g7009 ( 
.A1(n_6716),
.A2(n_936),
.B(n_937),
.Y(n_7009)
);

AOI22xp33_ASAP7_75t_L g7010 ( 
.A1(n_6805),
.A2(n_939),
.B1(n_937),
.B2(n_938),
.Y(n_7010)
);

NOR2xp33_ASAP7_75t_L g7011 ( 
.A(n_6771),
.B(n_938),
.Y(n_7011)
);

OAI221xp5_ASAP7_75t_L g7012 ( 
.A1(n_6751),
.A2(n_941),
.B1(n_939),
.B2(n_940),
.C(n_942),
.Y(n_7012)
);

INVx1_ASAP7_75t_L g7013 ( 
.A(n_6784),
.Y(n_7013)
);

INVx1_ASAP7_75t_L g7014 ( 
.A(n_6697),
.Y(n_7014)
);

AOI22xp5_ASAP7_75t_L g7015 ( 
.A1(n_6748),
.A2(n_945),
.B1(n_941),
.B2(n_944),
.Y(n_7015)
);

A2O1A1Ixp33_ASAP7_75t_L g7016 ( 
.A1(n_6796),
.A2(n_948),
.B(n_944),
.C(n_946),
.Y(n_7016)
);

OAI22xp5_ASAP7_75t_L g7017 ( 
.A1(n_6755),
.A2(n_950),
.B1(n_946),
.B2(n_948),
.Y(n_7017)
);

NAND2xp5_ASAP7_75t_L g7018 ( 
.A(n_6823),
.B(n_952),
.Y(n_7018)
);

INVx1_ASAP7_75t_L g7019 ( 
.A(n_6711),
.Y(n_7019)
);

INVx1_ASAP7_75t_L g7020 ( 
.A(n_6884),
.Y(n_7020)
);

NAND2xp5_ASAP7_75t_L g7021 ( 
.A(n_7004),
.B(n_6764),
.Y(n_7021)
);

NAND2xp5_ASAP7_75t_L g7022 ( 
.A(n_6963),
.B(n_6793),
.Y(n_7022)
);

INVx1_ASAP7_75t_L g7023 ( 
.A(n_6925),
.Y(n_7023)
);

INVx1_ASAP7_75t_L g7024 ( 
.A(n_6999),
.Y(n_7024)
);

AND2x2_ASAP7_75t_L g7025 ( 
.A(n_6901),
.B(n_6775),
.Y(n_7025)
);

NAND2xp5_ASAP7_75t_L g7026 ( 
.A(n_6964),
.B(n_6793),
.Y(n_7026)
);

AND2x2_ASAP7_75t_L g7027 ( 
.A(n_6897),
.B(n_6790),
.Y(n_7027)
);

INVx1_ASAP7_75t_L g7028 ( 
.A(n_6895),
.Y(n_7028)
);

INVxp67_ASAP7_75t_L g7029 ( 
.A(n_6885),
.Y(n_7029)
);

INVx1_ASAP7_75t_L g7030 ( 
.A(n_6979),
.Y(n_7030)
);

INVx1_ASAP7_75t_L g7031 ( 
.A(n_6984),
.Y(n_7031)
);

INVx1_ASAP7_75t_L g7032 ( 
.A(n_6968),
.Y(n_7032)
);

OR2x2_ASAP7_75t_L g7033 ( 
.A(n_6876),
.B(n_6712),
.Y(n_7033)
);

INVx1_ASAP7_75t_L g7034 ( 
.A(n_6907),
.Y(n_7034)
);

INVx1_ASAP7_75t_L g7035 ( 
.A(n_6910),
.Y(n_7035)
);

INVx1_ASAP7_75t_L g7036 ( 
.A(n_6920),
.Y(n_7036)
);

NAND2xp5_ASAP7_75t_L g7037 ( 
.A(n_6929),
.B(n_6746),
.Y(n_7037)
);

NAND2xp5_ASAP7_75t_L g7038 ( 
.A(n_6929),
.B(n_6795),
.Y(n_7038)
);

INVx1_ASAP7_75t_SL g7039 ( 
.A(n_6874),
.Y(n_7039)
);

NAND3xp33_ASAP7_75t_L g7040 ( 
.A(n_6899),
.B(n_6794),
.C(n_6768),
.Y(n_7040)
);

INVx1_ASAP7_75t_L g7041 ( 
.A(n_6922),
.Y(n_7041)
);

NOR2xp33_ASAP7_75t_L g7042 ( 
.A(n_6962),
.B(n_6757),
.Y(n_7042)
);

HB1xp67_ASAP7_75t_L g7043 ( 
.A(n_6994),
.Y(n_7043)
);

NAND2xp5_ASAP7_75t_L g7044 ( 
.A(n_6974),
.B(n_6754),
.Y(n_7044)
);

NOR2xp33_ASAP7_75t_R g7045 ( 
.A(n_6887),
.B(n_6750),
.Y(n_7045)
);

AND2x2_ASAP7_75t_L g7046 ( 
.A(n_6916),
.B(n_6788),
.Y(n_7046)
);

NAND2xp5_ASAP7_75t_L g7047 ( 
.A(n_6927),
.B(n_6687),
.Y(n_7047)
);

INVx1_ASAP7_75t_L g7048 ( 
.A(n_6926),
.Y(n_7048)
);

INVx1_ASAP7_75t_L g7049 ( 
.A(n_6936),
.Y(n_7049)
);

NAND2xp5_ASAP7_75t_SL g7050 ( 
.A(n_6900),
.B(n_6932),
.Y(n_7050)
);

OR2x2_ASAP7_75t_L g7051 ( 
.A(n_6877),
.B(n_6781),
.Y(n_7051)
);

AOI22xp33_ASAP7_75t_L g7052 ( 
.A1(n_6997),
.A2(n_6763),
.B1(n_6704),
.B2(n_954),
.Y(n_7052)
);

INVx2_ASAP7_75t_L g7053 ( 
.A(n_6913),
.Y(n_7053)
);

INVx1_ASAP7_75t_L g7054 ( 
.A(n_6917),
.Y(n_7054)
);

NAND2xp5_ASAP7_75t_L g7055 ( 
.A(n_6940),
.B(n_952),
.Y(n_7055)
);

NAND2xp5_ASAP7_75t_L g7056 ( 
.A(n_6954),
.B(n_953),
.Y(n_7056)
);

INVx1_ASAP7_75t_L g7057 ( 
.A(n_6918),
.Y(n_7057)
);

NOR2xp33_ASAP7_75t_L g7058 ( 
.A(n_6919),
.B(n_956),
.Y(n_7058)
);

NOR2xp33_ASAP7_75t_L g7059 ( 
.A(n_6906),
.B(n_957),
.Y(n_7059)
);

INVx1_ASAP7_75t_L g7060 ( 
.A(n_6955),
.Y(n_7060)
);

INVx1_ASAP7_75t_L g7061 ( 
.A(n_6928),
.Y(n_7061)
);

NAND2xp33_ASAP7_75t_L g7062 ( 
.A(n_6880),
.B(n_957),
.Y(n_7062)
);

INVx1_ASAP7_75t_L g7063 ( 
.A(n_6933),
.Y(n_7063)
);

INVx2_ASAP7_75t_SL g7064 ( 
.A(n_6889),
.Y(n_7064)
);

OR2x2_ASAP7_75t_L g7065 ( 
.A(n_6881),
.B(n_958),
.Y(n_7065)
);

INVx1_ASAP7_75t_L g7066 ( 
.A(n_6934),
.Y(n_7066)
);

INVx1_ASAP7_75t_L g7067 ( 
.A(n_6937),
.Y(n_7067)
);

INVx2_ASAP7_75t_L g7068 ( 
.A(n_7001),
.Y(n_7068)
);

INVx1_ASAP7_75t_L g7069 ( 
.A(n_6941),
.Y(n_7069)
);

INVx1_ASAP7_75t_L g7070 ( 
.A(n_6947),
.Y(n_7070)
);

HB1xp67_ASAP7_75t_L g7071 ( 
.A(n_6935),
.Y(n_7071)
);

OAI21xp33_ASAP7_75t_SL g7072 ( 
.A1(n_6930),
.A2(n_6890),
.B(n_6883),
.Y(n_7072)
);

INVx2_ASAP7_75t_L g7073 ( 
.A(n_7008),
.Y(n_7073)
);

NAND2xp5_ASAP7_75t_L g7074 ( 
.A(n_6951),
.B(n_959),
.Y(n_7074)
);

AND2x2_ASAP7_75t_L g7075 ( 
.A(n_6943),
.B(n_959),
.Y(n_7075)
);

NOR2xp33_ASAP7_75t_L g7076 ( 
.A(n_6976),
.B(n_6898),
.Y(n_7076)
);

NAND2xp5_ASAP7_75t_SL g7077 ( 
.A(n_6939),
.B(n_960),
.Y(n_7077)
);

NAND2xp5_ASAP7_75t_L g7078 ( 
.A(n_6990),
.B(n_961),
.Y(n_7078)
);

NAND2xp5_ASAP7_75t_L g7079 ( 
.A(n_6946),
.B(n_962),
.Y(n_7079)
);

AOI22xp5_ASAP7_75t_L g7080 ( 
.A1(n_6967),
.A2(n_970),
.B1(n_978),
.B2(n_962),
.Y(n_7080)
);

NAND2xp5_ASAP7_75t_L g7081 ( 
.A(n_6892),
.B(n_6903),
.Y(n_7081)
);

INVx1_ASAP7_75t_SL g7082 ( 
.A(n_6972),
.Y(n_7082)
);

NAND2xp5_ASAP7_75t_L g7083 ( 
.A(n_6915),
.B(n_963),
.Y(n_7083)
);

NAND2xp5_ASAP7_75t_L g7084 ( 
.A(n_6909),
.B(n_964),
.Y(n_7084)
);

INVx1_ASAP7_75t_L g7085 ( 
.A(n_6989),
.Y(n_7085)
);

NOR3xp33_ASAP7_75t_L g7086 ( 
.A(n_6956),
.B(n_965),
.C(n_966),
.Y(n_7086)
);

INVx3_ASAP7_75t_L g7087 ( 
.A(n_6904),
.Y(n_7087)
);

INVx1_ASAP7_75t_L g7088 ( 
.A(n_6993),
.Y(n_7088)
);

INVx1_ASAP7_75t_L g7089 ( 
.A(n_6987),
.Y(n_7089)
);

NAND2xp5_ASAP7_75t_SL g7090 ( 
.A(n_6879),
.B(n_965),
.Y(n_7090)
);

HB1xp67_ASAP7_75t_L g7091 ( 
.A(n_6896),
.Y(n_7091)
);

NAND2xp5_ASAP7_75t_L g7092 ( 
.A(n_6891),
.B(n_966),
.Y(n_7092)
);

AND2x2_ASAP7_75t_L g7093 ( 
.A(n_6957),
.B(n_967),
.Y(n_7093)
);

INVx1_ASAP7_75t_L g7094 ( 
.A(n_6991),
.Y(n_7094)
);

NAND2x1_ASAP7_75t_L g7095 ( 
.A(n_6914),
.B(n_968),
.Y(n_7095)
);

OR2x2_ASAP7_75t_L g7096 ( 
.A(n_6959),
.B(n_969),
.Y(n_7096)
);

INVx2_ASAP7_75t_L g7097 ( 
.A(n_6978),
.Y(n_7097)
);

NAND2xp5_ASAP7_75t_SL g7098 ( 
.A(n_6921),
.B(n_969),
.Y(n_7098)
);

NAND2xp5_ASAP7_75t_L g7099 ( 
.A(n_7000),
.B(n_970),
.Y(n_7099)
);

INVx2_ASAP7_75t_L g7100 ( 
.A(n_6949),
.Y(n_7100)
);

INVx1_ASAP7_75t_L g7101 ( 
.A(n_7002),
.Y(n_7101)
);

INVx1_ASAP7_75t_L g7102 ( 
.A(n_7005),
.Y(n_7102)
);

NAND2xp5_ASAP7_75t_L g7103 ( 
.A(n_6908),
.B(n_7014),
.Y(n_7103)
);

INVxp67_ASAP7_75t_L g7104 ( 
.A(n_6969),
.Y(n_7104)
);

INVx1_ASAP7_75t_L g7105 ( 
.A(n_7019),
.Y(n_7105)
);

INVx1_ASAP7_75t_L g7106 ( 
.A(n_7006),
.Y(n_7106)
);

NOR2xp33_ASAP7_75t_L g7107 ( 
.A(n_6912),
.B(n_971),
.Y(n_7107)
);

OR2x6_ASAP7_75t_L g7108 ( 
.A(n_6923),
.B(n_6888),
.Y(n_7108)
);

AND2x2_ASAP7_75t_L g7109 ( 
.A(n_6965),
.B(n_972),
.Y(n_7109)
);

NOR4xp25_ASAP7_75t_L g7110 ( 
.A(n_6985),
.B(n_6924),
.C(n_6983),
.D(n_6980),
.Y(n_7110)
);

AND2x2_ASAP7_75t_L g7111 ( 
.A(n_6995),
.B(n_972),
.Y(n_7111)
);

CKINVDCx16_ASAP7_75t_R g7112 ( 
.A(n_6878),
.Y(n_7112)
);

AND2x2_ASAP7_75t_L g7113 ( 
.A(n_6952),
.B(n_973),
.Y(n_7113)
);

AND2x2_ASAP7_75t_L g7114 ( 
.A(n_6988),
.B(n_974),
.Y(n_7114)
);

NAND2xp5_ASAP7_75t_L g7115 ( 
.A(n_7013),
.B(n_974),
.Y(n_7115)
);

INVx1_ASAP7_75t_SL g7116 ( 
.A(n_6971),
.Y(n_7116)
);

NAND2xp5_ASAP7_75t_L g7117 ( 
.A(n_6961),
.B(n_975),
.Y(n_7117)
);

NAND2xp5_ASAP7_75t_L g7118 ( 
.A(n_6982),
.B(n_976),
.Y(n_7118)
);

NAND2xp5_ASAP7_75t_L g7119 ( 
.A(n_6981),
.B(n_976),
.Y(n_7119)
);

NOR2xp33_ASAP7_75t_L g7120 ( 
.A(n_6948),
.B(n_977),
.Y(n_7120)
);

INVx1_ASAP7_75t_L g7121 ( 
.A(n_6902),
.Y(n_7121)
);

NAND2xp5_ASAP7_75t_L g7122 ( 
.A(n_6996),
.B(n_7011),
.Y(n_7122)
);

INVx2_ASAP7_75t_SL g7123 ( 
.A(n_6998),
.Y(n_7123)
);

OR2x2_ASAP7_75t_L g7124 ( 
.A(n_7018),
.B(n_978),
.Y(n_7124)
);

AND2x2_ASAP7_75t_L g7125 ( 
.A(n_6958),
.B(n_979),
.Y(n_7125)
);

NAND2x1_ASAP7_75t_L g7126 ( 
.A(n_6938),
.B(n_979),
.Y(n_7126)
);

AND2x2_ASAP7_75t_L g7127 ( 
.A(n_6875),
.B(n_980),
.Y(n_7127)
);

OR2x2_ASAP7_75t_L g7128 ( 
.A(n_6905),
.B(n_980),
.Y(n_7128)
);

INVx1_ASAP7_75t_L g7129 ( 
.A(n_6975),
.Y(n_7129)
);

NAND2xp5_ASAP7_75t_L g7130 ( 
.A(n_7016),
.B(n_981),
.Y(n_7130)
);

INVx1_ASAP7_75t_SL g7131 ( 
.A(n_6893),
.Y(n_7131)
);

NAND2xp5_ASAP7_75t_L g7132 ( 
.A(n_6944),
.B(n_981),
.Y(n_7132)
);

NAND2xp5_ASAP7_75t_L g7133 ( 
.A(n_6950),
.B(n_982),
.Y(n_7133)
);

INVx1_ASAP7_75t_L g7134 ( 
.A(n_6986),
.Y(n_7134)
);

INVx1_ASAP7_75t_L g7135 ( 
.A(n_6894),
.Y(n_7135)
);

NAND3x1_ASAP7_75t_L g7136 ( 
.A(n_7015),
.B(n_984),
.C(n_983),
.Y(n_7136)
);

INVx1_ASAP7_75t_L g7137 ( 
.A(n_6911),
.Y(n_7137)
);

INVx2_ASAP7_75t_L g7138 ( 
.A(n_6931),
.Y(n_7138)
);

NOR2xp67_ASAP7_75t_L g7139 ( 
.A(n_7007),
.B(n_982),
.Y(n_7139)
);

INVx2_ASAP7_75t_L g7140 ( 
.A(n_7003),
.Y(n_7140)
);

INVxp67_ASAP7_75t_L g7141 ( 
.A(n_7012),
.Y(n_7141)
);

NOR2x1_ASAP7_75t_L g7142 ( 
.A(n_6970),
.B(n_983),
.Y(n_7142)
);

INVx1_ASAP7_75t_L g7143 ( 
.A(n_7017),
.Y(n_7143)
);

INVxp67_ASAP7_75t_L g7144 ( 
.A(n_6992),
.Y(n_7144)
);

NAND2xp5_ASAP7_75t_SL g7145 ( 
.A(n_6882),
.B(n_984),
.Y(n_7145)
);

INVx1_ASAP7_75t_L g7146 ( 
.A(n_6966),
.Y(n_7146)
);

NAND2xp5_ASAP7_75t_L g7147 ( 
.A(n_6960),
.B(n_985),
.Y(n_7147)
);

INVx4_ASAP7_75t_L g7148 ( 
.A(n_6945),
.Y(n_7148)
);

AND2x2_ASAP7_75t_L g7149 ( 
.A(n_6977),
.B(n_985),
.Y(n_7149)
);

NOR2xp33_ASAP7_75t_L g7150 ( 
.A(n_6953),
.B(n_987),
.Y(n_7150)
);

INVx3_ASAP7_75t_L g7151 ( 
.A(n_6942),
.Y(n_7151)
);

INVx1_ASAP7_75t_L g7152 ( 
.A(n_6973),
.Y(n_7152)
);

INVxp67_ASAP7_75t_L g7153 ( 
.A(n_7009),
.Y(n_7153)
);

NOR3xp33_ASAP7_75t_SL g7154 ( 
.A(n_6886),
.B(n_987),
.C(n_988),
.Y(n_7154)
);

OR2x2_ASAP7_75t_L g7155 ( 
.A(n_7010),
.B(n_989),
.Y(n_7155)
);

AND2x2_ASAP7_75t_L g7156 ( 
.A(n_6884),
.B(n_989),
.Y(n_7156)
);

INVx1_ASAP7_75t_L g7157 ( 
.A(n_6884),
.Y(n_7157)
);

INVx1_ASAP7_75t_L g7158 ( 
.A(n_6884),
.Y(n_7158)
);

AND2x2_ASAP7_75t_L g7159 ( 
.A(n_6884),
.B(n_990),
.Y(n_7159)
);

NAND2xp5_ASAP7_75t_L g7160 ( 
.A(n_7004),
.B(n_990),
.Y(n_7160)
);

NAND2xp5_ASAP7_75t_L g7161 ( 
.A(n_7004),
.B(n_992),
.Y(n_7161)
);

NOR2xp33_ASAP7_75t_L g7162 ( 
.A(n_6962),
.B(n_993),
.Y(n_7162)
);

NAND2xp5_ASAP7_75t_L g7163 ( 
.A(n_7004),
.B(n_993),
.Y(n_7163)
);

INVx2_ASAP7_75t_L g7164 ( 
.A(n_6913),
.Y(n_7164)
);

OR2x2_ASAP7_75t_L g7165 ( 
.A(n_6884),
.B(n_994),
.Y(n_7165)
);

OR2x2_ASAP7_75t_L g7166 ( 
.A(n_6884),
.B(n_994),
.Y(n_7166)
);

INVx1_ASAP7_75t_L g7167 ( 
.A(n_6884),
.Y(n_7167)
);

NAND2xp5_ASAP7_75t_L g7168 ( 
.A(n_7004),
.B(n_995),
.Y(n_7168)
);

HB1xp67_ASAP7_75t_L g7169 ( 
.A(n_6884),
.Y(n_7169)
);

INVx1_ASAP7_75t_L g7170 ( 
.A(n_6884),
.Y(n_7170)
);

NAND2xp5_ASAP7_75t_L g7171 ( 
.A(n_7004),
.B(n_996),
.Y(n_7171)
);

AND2x2_ASAP7_75t_L g7172 ( 
.A(n_6884),
.B(n_996),
.Y(n_7172)
);

NAND2xp5_ASAP7_75t_L g7173 ( 
.A(n_7004),
.B(n_997),
.Y(n_7173)
);

NAND2xp5_ASAP7_75t_L g7174 ( 
.A(n_7004),
.B(n_997),
.Y(n_7174)
);

AND2x2_ASAP7_75t_L g7175 ( 
.A(n_6884),
.B(n_998),
.Y(n_7175)
);

INVx2_ASAP7_75t_L g7176 ( 
.A(n_6913),
.Y(n_7176)
);

INVx1_ASAP7_75t_L g7177 ( 
.A(n_6884),
.Y(n_7177)
);

INVx1_ASAP7_75t_L g7178 ( 
.A(n_6884),
.Y(n_7178)
);

HB1xp67_ASAP7_75t_L g7179 ( 
.A(n_6884),
.Y(n_7179)
);

OAI31xp33_ASAP7_75t_L g7180 ( 
.A1(n_6897),
.A2(n_1001),
.A3(n_998),
.B(n_1000),
.Y(n_7180)
);

AND2x2_ASAP7_75t_L g7181 ( 
.A(n_6884),
.B(n_1000),
.Y(n_7181)
);

OR2x2_ASAP7_75t_L g7182 ( 
.A(n_6884),
.B(n_1001),
.Y(n_7182)
);

INVx1_ASAP7_75t_L g7183 ( 
.A(n_6884),
.Y(n_7183)
);

NAND2xp5_ASAP7_75t_L g7184 ( 
.A(n_7043),
.B(n_1002),
.Y(n_7184)
);

XOR2xp5_ASAP7_75t_L g7185 ( 
.A(n_7071),
.B(n_1003),
.Y(n_7185)
);

XOR2x2_ASAP7_75t_L g7186 ( 
.A(n_7040),
.B(n_1002),
.Y(n_7186)
);

NOR2xp33_ASAP7_75t_L g7187 ( 
.A(n_7039),
.B(n_1003),
.Y(n_7187)
);

XOR2x2_ASAP7_75t_L g7188 ( 
.A(n_7042),
.B(n_1004),
.Y(n_7188)
);

AND2x2_ASAP7_75t_L g7189 ( 
.A(n_7027),
.B(n_1005),
.Y(n_7189)
);

NOR2xp33_ASAP7_75t_L g7190 ( 
.A(n_7087),
.B(n_1005),
.Y(n_7190)
);

INVx1_ASAP7_75t_L g7191 ( 
.A(n_7169),
.Y(n_7191)
);

INVx2_ASAP7_75t_SL g7192 ( 
.A(n_7179),
.Y(n_7192)
);

AND3x2_ASAP7_75t_L g7193 ( 
.A(n_7110),
.B(n_1006),
.C(n_1007),
.Y(n_7193)
);

INVx2_ASAP7_75t_L g7194 ( 
.A(n_7165),
.Y(n_7194)
);

AND2x2_ASAP7_75t_L g7195 ( 
.A(n_7025),
.B(n_1006),
.Y(n_7195)
);

INVxp67_ASAP7_75t_L g7196 ( 
.A(n_7162),
.Y(n_7196)
);

NOR2x1_ASAP7_75t_L g7197 ( 
.A(n_7166),
.B(n_1007),
.Y(n_7197)
);

NAND2xp5_ASAP7_75t_SL g7198 ( 
.A(n_7100),
.B(n_1008),
.Y(n_7198)
);

INVx1_ASAP7_75t_L g7199 ( 
.A(n_7156),
.Y(n_7199)
);

OAI22xp5_ASAP7_75t_L g7200 ( 
.A1(n_7020),
.A2(n_1010),
.B1(n_1008),
.B2(n_1009),
.Y(n_7200)
);

OR2x2_ASAP7_75t_L g7201 ( 
.A(n_7182),
.B(n_1010),
.Y(n_7201)
);

NOR3xp33_ASAP7_75t_L g7202 ( 
.A(n_7072),
.B(n_1012),
.C(n_1013),
.Y(n_7202)
);

NAND2xp5_ASAP7_75t_L g7203 ( 
.A(n_7159),
.B(n_1013),
.Y(n_7203)
);

AOI211x1_ASAP7_75t_SL g7204 ( 
.A1(n_7050),
.A2(n_1018),
.B(n_1015),
.C(n_1016),
.Y(n_7204)
);

NOR2x1_ASAP7_75t_L g7205 ( 
.A(n_7157),
.B(n_1015),
.Y(n_7205)
);

NAND2xp5_ASAP7_75t_L g7206 ( 
.A(n_7172),
.B(n_1016),
.Y(n_7206)
);

AND2x2_ASAP7_75t_L g7207 ( 
.A(n_7024),
.B(n_1018),
.Y(n_7207)
);

AND2x2_ASAP7_75t_L g7208 ( 
.A(n_7158),
.B(n_1019),
.Y(n_7208)
);

INVx1_ASAP7_75t_L g7209 ( 
.A(n_7175),
.Y(n_7209)
);

INVx1_ASAP7_75t_L g7210 ( 
.A(n_7181),
.Y(n_7210)
);

NOR4xp25_ASAP7_75t_SL g7211 ( 
.A(n_7167),
.B(n_1023),
.C(n_1020),
.D(n_1021),
.Y(n_7211)
);

INVx2_ASAP7_75t_L g7212 ( 
.A(n_7095),
.Y(n_7212)
);

XOR2x2_ASAP7_75t_L g7213 ( 
.A(n_7136),
.B(n_1020),
.Y(n_7213)
);

NAND2xp5_ASAP7_75t_L g7214 ( 
.A(n_7112),
.B(n_1023),
.Y(n_7214)
);

INVx1_ASAP7_75t_L g7215 ( 
.A(n_7055),
.Y(n_7215)
);

AND2x2_ASAP7_75t_L g7216 ( 
.A(n_7170),
.B(n_1024),
.Y(n_7216)
);

NAND2xp5_ASAP7_75t_SL g7217 ( 
.A(n_7177),
.B(n_1024),
.Y(n_7217)
);

XNOR2xp5_ASAP7_75t_L g7218 ( 
.A(n_7091),
.B(n_1026),
.Y(n_7218)
);

NOR2xp33_ASAP7_75t_L g7219 ( 
.A(n_7116),
.B(n_1026),
.Y(n_7219)
);

INVx1_ASAP7_75t_L g7220 ( 
.A(n_7047),
.Y(n_7220)
);

AOI22xp5_ASAP7_75t_L g7221 ( 
.A1(n_7058),
.A2(n_1029),
.B1(n_1027),
.B2(n_1028),
.Y(n_7221)
);

BUFx2_ASAP7_75t_L g7222 ( 
.A(n_7045),
.Y(n_7222)
);

OR2x2_ASAP7_75t_L g7223 ( 
.A(n_7178),
.B(n_1028),
.Y(n_7223)
);

INVx1_ASAP7_75t_L g7224 ( 
.A(n_7183),
.Y(n_7224)
);

NOR2xp33_ASAP7_75t_L g7225 ( 
.A(n_7064),
.B(n_1029),
.Y(n_7225)
);

NAND2xp5_ASAP7_75t_L g7226 ( 
.A(n_7082),
.B(n_1031),
.Y(n_7226)
);

AND3x2_ASAP7_75t_L g7227 ( 
.A(n_7029),
.B(n_1032),
.C(n_1033),
.Y(n_7227)
);

NOR2xp33_ASAP7_75t_R g7228 ( 
.A(n_7060),
.B(n_1034),
.Y(n_7228)
);

NOR3x1_ASAP7_75t_L g7229 ( 
.A(n_7123),
.B(n_1032),
.C(n_1034),
.Y(n_7229)
);

INVxp67_ASAP7_75t_L g7230 ( 
.A(n_7022),
.Y(n_7230)
);

INVx1_ASAP7_75t_L g7231 ( 
.A(n_7114),
.Y(n_7231)
);

OAI21x1_ASAP7_75t_L g7232 ( 
.A1(n_7026),
.A2(n_1035),
.B(n_1036),
.Y(n_7232)
);

OR2x2_ASAP7_75t_L g7233 ( 
.A(n_7033),
.B(n_1036),
.Y(n_7233)
);

NAND4xp25_ASAP7_75t_L g7234 ( 
.A(n_7076),
.B(n_1039),
.C(n_1037),
.D(n_1038),
.Y(n_7234)
);

INVx1_ASAP7_75t_L g7235 ( 
.A(n_7093),
.Y(n_7235)
);

INVx1_ASAP7_75t_SL g7236 ( 
.A(n_7109),
.Y(n_7236)
);

INVx1_ASAP7_75t_L g7237 ( 
.A(n_7160),
.Y(n_7237)
);

NAND2xp5_ASAP7_75t_SL g7238 ( 
.A(n_7068),
.B(n_1037),
.Y(n_7238)
);

INVx2_ASAP7_75t_L g7239 ( 
.A(n_7096),
.Y(n_7239)
);

INVx1_ASAP7_75t_L g7240 ( 
.A(n_7161),
.Y(n_7240)
);

INVx1_ASAP7_75t_L g7241 ( 
.A(n_7163),
.Y(n_7241)
);

INVxp33_ASAP7_75t_SL g7242 ( 
.A(n_7021),
.Y(n_7242)
);

OAI21xp5_ASAP7_75t_SL g7243 ( 
.A1(n_7046),
.A2(n_1038),
.B(n_1039),
.Y(n_7243)
);

OAI21xp33_ASAP7_75t_L g7244 ( 
.A1(n_7044),
.A2(n_1040),
.B(n_1042),
.Y(n_7244)
);

NAND2xp5_ASAP7_75t_L g7245 ( 
.A(n_7028),
.B(n_1043),
.Y(n_7245)
);

AOI21xp33_ASAP7_75t_L g7246 ( 
.A1(n_7131),
.A2(n_1044),
.B(n_1045),
.Y(n_7246)
);

NOR2xp33_ASAP7_75t_L g7247 ( 
.A(n_7057),
.B(n_1049),
.Y(n_7247)
);

NAND2xp5_ASAP7_75t_L g7248 ( 
.A(n_7073),
.B(n_1050),
.Y(n_7248)
);

INVx2_ASAP7_75t_L g7249 ( 
.A(n_7108),
.Y(n_7249)
);

INVx1_ASAP7_75t_L g7250 ( 
.A(n_7168),
.Y(n_7250)
);

NAND3xp33_ASAP7_75t_L g7251 ( 
.A(n_7062),
.B(n_1058),
.C(n_1050),
.Y(n_7251)
);

INVx1_ASAP7_75t_L g7252 ( 
.A(n_7171),
.Y(n_7252)
);

NOR4xp25_ASAP7_75t_SL g7253 ( 
.A(n_7105),
.B(n_1053),
.C(n_1051),
.D(n_1052),
.Y(n_7253)
);

NAND2xp5_ASAP7_75t_L g7254 ( 
.A(n_7089),
.B(n_1051),
.Y(n_7254)
);

INVx2_ASAP7_75t_L g7255 ( 
.A(n_7108),
.Y(n_7255)
);

NAND2xp5_ASAP7_75t_L g7256 ( 
.A(n_7053),
.B(n_1052),
.Y(n_7256)
);

AND2x2_ASAP7_75t_L g7257 ( 
.A(n_7111),
.B(n_1053),
.Y(n_7257)
);

NOR2x1_ASAP7_75t_L g7258 ( 
.A(n_7038),
.B(n_1054),
.Y(n_7258)
);

NAND2xp33_ASAP7_75t_SL g7259 ( 
.A(n_7051),
.B(n_1054),
.Y(n_7259)
);

NAND2x1_ASAP7_75t_L g7260 ( 
.A(n_7164),
.B(n_1055),
.Y(n_7260)
);

INVx1_ASAP7_75t_L g7261 ( 
.A(n_7173),
.Y(n_7261)
);

INVx1_ASAP7_75t_L g7262 ( 
.A(n_7174),
.Y(n_7262)
);

INVx1_ASAP7_75t_L g7263 ( 
.A(n_7037),
.Y(n_7263)
);

INVx3_ASAP7_75t_L g7264 ( 
.A(n_7176),
.Y(n_7264)
);

AOI21xp5_ASAP7_75t_L g7265 ( 
.A1(n_7098),
.A2(n_1056),
.B(n_1057),
.Y(n_7265)
);

AND2x2_ASAP7_75t_L g7266 ( 
.A(n_7061),
.B(n_1056),
.Y(n_7266)
);

INVx1_ASAP7_75t_L g7267 ( 
.A(n_7118),
.Y(n_7267)
);

AOI322xp5_ASAP7_75t_L g7268 ( 
.A1(n_7052),
.A2(n_1065),
.A3(n_1064),
.B1(n_1060),
.B2(n_1058),
.C1(n_1059),
.C2(n_1062),
.Y(n_7268)
);

AND2x2_ASAP7_75t_L g7269 ( 
.A(n_7063),
.B(n_1059),
.Y(n_7269)
);

INVx1_ASAP7_75t_L g7270 ( 
.A(n_7032),
.Y(n_7270)
);

INVx1_ASAP7_75t_L g7271 ( 
.A(n_7075),
.Y(n_7271)
);

INVx1_ASAP7_75t_SL g7272 ( 
.A(n_7065),
.Y(n_7272)
);

INVx1_ASAP7_75t_L g7273 ( 
.A(n_7023),
.Y(n_7273)
);

INVx1_ASAP7_75t_L g7274 ( 
.A(n_7097),
.Y(n_7274)
);

NAND2xp5_ASAP7_75t_SL g7275 ( 
.A(n_7180),
.B(n_1060),
.Y(n_7275)
);

OA22x2_ASAP7_75t_L g7276 ( 
.A1(n_7054),
.A2(n_1065),
.B1(n_1062),
.B2(n_1064),
.Y(n_7276)
);

NAND2xp5_ASAP7_75t_L g7277 ( 
.A(n_7088),
.B(n_1066),
.Y(n_7277)
);

INVx2_ASAP7_75t_L g7278 ( 
.A(n_7125),
.Y(n_7278)
);

OR2x2_ASAP7_75t_L g7279 ( 
.A(n_7081),
.B(n_1066),
.Y(n_7279)
);

NAND3xp33_ASAP7_75t_SL g7280 ( 
.A(n_7204),
.B(n_7086),
.C(n_7103),
.Y(n_7280)
);

O2A1O1Ixp33_ASAP7_75t_L g7281 ( 
.A1(n_7243),
.A2(n_7079),
.B(n_7106),
.C(n_7066),
.Y(n_7281)
);

NOR2xp33_ASAP7_75t_L g7282 ( 
.A(n_7242),
.B(n_7148),
.Y(n_7282)
);

AOI221xp5_ASAP7_75t_L g7283 ( 
.A1(n_7230),
.A2(n_7134),
.B1(n_7034),
.B2(n_7035),
.C(n_7031),
.Y(n_7283)
);

O2A1O1Ixp33_ASAP7_75t_SL g7284 ( 
.A1(n_7192),
.A2(n_7069),
.B(n_7070),
.C(n_7067),
.Y(n_7284)
);

NOR2xp33_ASAP7_75t_L g7285 ( 
.A(n_7236),
.B(n_7148),
.Y(n_7285)
);

NOR2x1_ASAP7_75t_L g7286 ( 
.A(n_7222),
.B(n_7094),
.Y(n_7286)
);

NOR4xp25_ASAP7_75t_L g7287 ( 
.A(n_7198),
.B(n_7102),
.C(n_7101),
.D(n_7036),
.Y(n_7287)
);

NOR3xp33_ASAP7_75t_L g7288 ( 
.A(n_7264),
.B(n_7078),
.C(n_7083),
.Y(n_7288)
);

OAI21xp5_ASAP7_75t_L g7289 ( 
.A1(n_7274),
.A2(n_7104),
.B(n_7059),
.Y(n_7289)
);

AOI221xp5_ASAP7_75t_L g7290 ( 
.A1(n_7199),
.A2(n_7048),
.B1(n_7049),
.B2(n_7041),
.C(n_7030),
.Y(n_7290)
);

AND2x2_ASAP7_75t_L g7291 ( 
.A(n_7189),
.B(n_7195),
.Y(n_7291)
);

AOI211xp5_ASAP7_75t_SL g7292 ( 
.A1(n_7191),
.A2(n_7074),
.B(n_7056),
.C(n_7141),
.Y(n_7292)
);

AOI222xp33_ASAP7_75t_L g7293 ( 
.A1(n_7259),
.A2(n_7153),
.B1(n_7129),
.B2(n_7144),
.C1(n_7121),
.C2(n_7085),
.Y(n_7293)
);

NAND2xp5_ASAP7_75t_L g7294 ( 
.A(n_7193),
.B(n_7107),
.Y(n_7294)
);

INVx1_ASAP7_75t_L g7295 ( 
.A(n_7218),
.Y(n_7295)
);

AOI21xp5_ASAP7_75t_L g7296 ( 
.A1(n_7238),
.A2(n_7090),
.B(n_7092),
.Y(n_7296)
);

NAND2xp5_ASAP7_75t_L g7297 ( 
.A(n_7227),
.B(n_7139),
.Y(n_7297)
);

INVx1_ASAP7_75t_SL g7298 ( 
.A(n_7228),
.Y(n_7298)
);

NOR3x1_ASAP7_75t_L g7299 ( 
.A(n_7234),
.B(n_7217),
.C(n_7184),
.Y(n_7299)
);

INVx1_ASAP7_75t_L g7300 ( 
.A(n_7185),
.Y(n_7300)
);

INVx1_ASAP7_75t_L g7301 ( 
.A(n_7197),
.Y(n_7301)
);

AOI22xp5_ASAP7_75t_L g7302 ( 
.A1(n_7221),
.A2(n_7210),
.B1(n_7209),
.B2(n_7267),
.Y(n_7302)
);

NOR3xp33_ASAP7_75t_L g7303 ( 
.A(n_7264),
.B(n_7115),
.C(n_7099),
.Y(n_7303)
);

NAND5xp2_ASAP7_75t_L g7304 ( 
.A(n_7220),
.B(n_7143),
.C(n_7137),
.D(n_7135),
.E(n_7146),
.Y(n_7304)
);

NOR3xp33_ASAP7_75t_L g7305 ( 
.A(n_7214),
.B(n_7124),
.C(n_7113),
.Y(n_7305)
);

NAND2xp5_ASAP7_75t_SL g7306 ( 
.A(n_7202),
.B(n_7138),
.Y(n_7306)
);

INVx1_ASAP7_75t_L g7307 ( 
.A(n_7205),
.Y(n_7307)
);

AND2x2_ASAP7_75t_L g7308 ( 
.A(n_7270),
.B(n_7127),
.Y(n_7308)
);

NAND2xp33_ASAP7_75t_R g7309 ( 
.A(n_7211),
.B(n_7120),
.Y(n_7309)
);

INVx1_ASAP7_75t_L g7310 ( 
.A(n_7188),
.Y(n_7310)
);

INVx1_ASAP7_75t_SL g7311 ( 
.A(n_7233),
.Y(n_7311)
);

NAND2xp5_ASAP7_75t_SL g7312 ( 
.A(n_7194),
.B(n_7084),
.Y(n_7312)
);

NOR2xp67_ASAP7_75t_L g7313 ( 
.A(n_7273),
.B(n_7128),
.Y(n_7313)
);

NOR2x1_ASAP7_75t_L g7314 ( 
.A(n_7279),
.B(n_7119),
.Y(n_7314)
);

NOR4xp25_ASAP7_75t_L g7315 ( 
.A(n_7272),
.B(n_7122),
.C(n_7140),
.D(n_7152),
.Y(n_7315)
);

INVx1_ASAP7_75t_L g7316 ( 
.A(n_7276),
.Y(n_7316)
);

NAND2xp5_ASAP7_75t_L g7317 ( 
.A(n_7258),
.B(n_7142),
.Y(n_7317)
);

NAND3xp33_ASAP7_75t_SL g7318 ( 
.A(n_7253),
.B(n_7260),
.C(n_7255),
.Y(n_7318)
);

NAND3xp33_ASAP7_75t_L g7319 ( 
.A(n_7219),
.B(n_7150),
.C(n_7130),
.Y(n_7319)
);

NAND4xp25_ASAP7_75t_SL g7320 ( 
.A(n_7224),
.B(n_7080),
.C(n_7147),
.D(n_7133),
.Y(n_7320)
);

INVx1_ASAP7_75t_L g7321 ( 
.A(n_7201),
.Y(n_7321)
);

HB1xp67_ASAP7_75t_L g7322 ( 
.A(n_7229),
.Y(n_7322)
);

NOR2xp33_ASAP7_75t_L g7323 ( 
.A(n_7231),
.B(n_7126),
.Y(n_7323)
);

AND2x2_ASAP7_75t_L g7324 ( 
.A(n_7208),
.B(n_7149),
.Y(n_7324)
);

INVx1_ASAP7_75t_L g7325 ( 
.A(n_7213),
.Y(n_7325)
);

AOI211xp5_ASAP7_75t_L g7326 ( 
.A1(n_7225),
.A2(n_7145),
.B(n_7077),
.C(n_7155),
.Y(n_7326)
);

NAND2xp5_ASAP7_75t_L g7327 ( 
.A(n_7207),
.B(n_7154),
.Y(n_7327)
);

NAND3xp33_ASAP7_75t_L g7328 ( 
.A(n_7187),
.B(n_7117),
.C(n_7132),
.Y(n_7328)
);

INVx1_ASAP7_75t_L g7329 ( 
.A(n_7203),
.Y(n_7329)
);

NAND4xp25_ASAP7_75t_L g7330 ( 
.A(n_7263),
.B(n_7275),
.C(n_7196),
.D(n_7151),
.Y(n_7330)
);

NAND2xp5_ASAP7_75t_L g7331 ( 
.A(n_7257),
.B(n_1068),
.Y(n_7331)
);

INVx1_ASAP7_75t_L g7332 ( 
.A(n_7206),
.Y(n_7332)
);

INVx2_ASAP7_75t_L g7333 ( 
.A(n_7212),
.Y(n_7333)
);

NAND2xp5_ASAP7_75t_L g7334 ( 
.A(n_7266),
.B(n_1068),
.Y(n_7334)
);

NAND2xp33_ASAP7_75t_L g7335 ( 
.A(n_7216),
.B(n_1070),
.Y(n_7335)
);

BUFx4f_ASAP7_75t_SL g7336 ( 
.A(n_7223),
.Y(n_7336)
);

INVx1_ASAP7_75t_L g7337 ( 
.A(n_7269),
.Y(n_7337)
);

AOI221x1_ASAP7_75t_L g7338 ( 
.A1(n_7226),
.A2(n_1073),
.B1(n_1071),
.B2(n_1072),
.C(n_1074),
.Y(n_7338)
);

NOR3xp33_ASAP7_75t_L g7339 ( 
.A(n_7249),
.B(n_1071),
.C(n_1072),
.Y(n_7339)
);

OAI31xp33_ASAP7_75t_SL g7340 ( 
.A1(n_7235),
.A2(n_1077),
.A3(n_1075),
.B(n_1076),
.Y(n_7340)
);

AOI211xp5_ASAP7_75t_L g7341 ( 
.A1(n_7190),
.A2(n_7247),
.B(n_7244),
.C(n_7265),
.Y(n_7341)
);

NAND2xp5_ASAP7_75t_SL g7342 ( 
.A(n_7268),
.B(n_1075),
.Y(n_7342)
);

NOR3xp33_ASAP7_75t_L g7343 ( 
.A(n_7318),
.B(n_7248),
.C(n_7254),
.Y(n_7343)
);

NAND3xp33_ASAP7_75t_L g7344 ( 
.A(n_7293),
.B(n_7215),
.C(n_7237),
.Y(n_7344)
);

NOR3xp33_ASAP7_75t_L g7345 ( 
.A(n_7330),
.B(n_7256),
.C(n_7245),
.Y(n_7345)
);

NOR3xp33_ASAP7_75t_L g7346 ( 
.A(n_7325),
.B(n_7286),
.C(n_7283),
.Y(n_7346)
);

NOR3xp33_ASAP7_75t_L g7347 ( 
.A(n_7298),
.B(n_7277),
.C(n_7241),
.Y(n_7347)
);

NOR2x1_ASAP7_75t_L g7348 ( 
.A(n_7282),
.B(n_7285),
.Y(n_7348)
);

AOI221xp5_ASAP7_75t_L g7349 ( 
.A1(n_7281),
.A2(n_7252),
.B1(n_7261),
.B2(n_7250),
.C(n_7240),
.Y(n_7349)
);

NOR3xp33_ASAP7_75t_L g7350 ( 
.A(n_7300),
.B(n_7262),
.C(n_7232),
.Y(n_7350)
);

AOI221xp5_ASAP7_75t_L g7351 ( 
.A1(n_7307),
.A2(n_7271),
.B1(n_7239),
.B2(n_7278),
.C(n_7251),
.Y(n_7351)
);

NAND3xp33_ASAP7_75t_L g7352 ( 
.A(n_7292),
.B(n_7246),
.C(n_7200),
.Y(n_7352)
);

OAI21xp33_ASAP7_75t_SL g7353 ( 
.A1(n_7287),
.A2(n_7186),
.B(n_1078),
.Y(n_7353)
);

NAND4xp25_ASAP7_75t_L g7354 ( 
.A(n_7304),
.B(n_1080),
.C(n_1078),
.D(n_1079),
.Y(n_7354)
);

NAND4xp25_ASAP7_75t_L g7355 ( 
.A(n_7290),
.B(n_1082),
.C(n_1080),
.D(n_1081),
.Y(n_7355)
);

NAND4xp25_ASAP7_75t_L g7356 ( 
.A(n_7299),
.B(n_1084),
.C(n_1081),
.D(n_1083),
.Y(n_7356)
);

NOR4xp75_ASAP7_75t_L g7357 ( 
.A(n_7289),
.B(n_1086),
.C(n_1083),
.D(n_1085),
.Y(n_7357)
);

NAND2xp5_ASAP7_75t_L g7358 ( 
.A(n_7340),
.B(n_1085),
.Y(n_7358)
);

NAND4xp25_ASAP7_75t_L g7359 ( 
.A(n_7341),
.B(n_1088),
.C(n_1086),
.D(n_1087),
.Y(n_7359)
);

NOR3xp33_ASAP7_75t_L g7360 ( 
.A(n_7310),
.B(n_1089),
.C(n_1090),
.Y(n_7360)
);

NAND4xp25_ASAP7_75t_L g7361 ( 
.A(n_7313),
.B(n_1091),
.C(n_1089),
.D(n_1090),
.Y(n_7361)
);

NOR3xp33_ASAP7_75t_L g7362 ( 
.A(n_7295),
.B(n_1093),
.C(n_1094),
.Y(n_7362)
);

AOI32xp33_ASAP7_75t_L g7363 ( 
.A1(n_7308),
.A2(n_1098),
.A3(n_1094),
.B1(n_1096),
.B2(n_1099),
.Y(n_7363)
);

NAND4xp25_ASAP7_75t_SL g7364 ( 
.A(n_7296),
.B(n_1100),
.C(n_1096),
.D(n_1099),
.Y(n_7364)
);

NOR2xp33_ASAP7_75t_L g7365 ( 
.A(n_7322),
.B(n_1100),
.Y(n_7365)
);

NOR2xp33_ASAP7_75t_L g7366 ( 
.A(n_7336),
.B(n_1101),
.Y(n_7366)
);

NAND2xp5_ASAP7_75t_L g7367 ( 
.A(n_7291),
.B(n_1102),
.Y(n_7367)
);

NAND5xp2_ASAP7_75t_L g7368 ( 
.A(n_7326),
.B(n_1104),
.C(n_1106),
.D(n_1103),
.E(n_1105),
.Y(n_7368)
);

BUFx4f_ASAP7_75t_SL g7369 ( 
.A(n_7333),
.Y(n_7369)
);

AOI21xp33_ASAP7_75t_L g7370 ( 
.A1(n_7309),
.A2(n_1102),
.B(n_1103),
.Y(n_7370)
);

INVx1_ASAP7_75t_L g7371 ( 
.A(n_7301),
.Y(n_7371)
);

NAND4xp25_ASAP7_75t_L g7372 ( 
.A(n_7302),
.B(n_7303),
.C(n_7280),
.D(n_7323),
.Y(n_7372)
);

NAND2xp5_ASAP7_75t_L g7373 ( 
.A(n_7311),
.B(n_1104),
.Y(n_7373)
);

NOR3x1_ASAP7_75t_SL g7374 ( 
.A(n_7320),
.B(n_1105),
.C(n_1106),
.Y(n_7374)
);

A2O1A1Ixp33_ASAP7_75t_L g7375 ( 
.A1(n_7288),
.A2(n_7316),
.B(n_7294),
.C(n_7328),
.Y(n_7375)
);

AOI211xp5_ASAP7_75t_SL g7376 ( 
.A1(n_7284),
.A2(n_7337),
.B(n_7317),
.C(n_7335),
.Y(n_7376)
);

OAI211xp5_ASAP7_75t_SL g7377 ( 
.A1(n_7306),
.A2(n_1109),
.B(n_1107),
.C(n_1108),
.Y(n_7377)
);

NAND4xp75_ASAP7_75t_SL g7378 ( 
.A(n_7324),
.B(n_1110),
.C(n_1107),
.D(n_1108),
.Y(n_7378)
);

AOI211xp5_ASAP7_75t_L g7379 ( 
.A1(n_7315),
.A2(n_1113),
.B(n_1111),
.C(n_1112),
.Y(n_7379)
);

NOR3x1_ASAP7_75t_L g7380 ( 
.A(n_7319),
.B(n_1111),
.C(n_1113),
.Y(n_7380)
);

AND3x2_ASAP7_75t_L g7381 ( 
.A(n_7339),
.B(n_1124),
.C(n_1114),
.Y(n_7381)
);

NAND4xp25_ASAP7_75t_SL g7382 ( 
.A(n_7305),
.B(n_1117),
.C(n_1115),
.D(n_1116),
.Y(n_7382)
);

CKINVDCx20_ASAP7_75t_R g7383 ( 
.A(n_7369),
.Y(n_7383)
);

NOR2x1_ASAP7_75t_L g7384 ( 
.A(n_7348),
.B(n_7334),
.Y(n_7384)
);

NOR2x1_ASAP7_75t_L g7385 ( 
.A(n_7372),
.B(n_7331),
.Y(n_7385)
);

INVx1_ASAP7_75t_L g7386 ( 
.A(n_7374),
.Y(n_7386)
);

AOI221xp5_ASAP7_75t_L g7387 ( 
.A1(n_7370),
.A2(n_7343),
.B1(n_7353),
.B2(n_7345),
.C(n_7346),
.Y(n_7387)
);

INVx1_ASAP7_75t_L g7388 ( 
.A(n_7358),
.Y(n_7388)
);

NAND2xp5_ASAP7_75t_L g7389 ( 
.A(n_7379),
.B(n_7338),
.Y(n_7389)
);

NOR2xp33_ASAP7_75t_L g7390 ( 
.A(n_7368),
.B(n_7312),
.Y(n_7390)
);

INVx1_ASAP7_75t_L g7391 ( 
.A(n_7357),
.Y(n_7391)
);

OAI22xp5_ASAP7_75t_L g7392 ( 
.A1(n_7371),
.A2(n_7327),
.B1(n_7314),
.B2(n_7342),
.Y(n_7392)
);

AOI221xp5_ASAP7_75t_L g7393 ( 
.A1(n_7347),
.A2(n_7329),
.B1(n_7332),
.B2(n_7321),
.C(n_7297),
.Y(n_7393)
);

OR2x2_ASAP7_75t_L g7394 ( 
.A(n_7354),
.B(n_1115),
.Y(n_7394)
);

NOR2x1p5_ASAP7_75t_L g7395 ( 
.A(n_7355),
.B(n_7361),
.Y(n_7395)
);

OAI211xp5_ASAP7_75t_L g7396 ( 
.A1(n_7376),
.A2(n_1120),
.B(n_1117),
.C(n_1118),
.Y(n_7396)
);

NAND3xp33_ASAP7_75t_SL g7397 ( 
.A(n_7350),
.B(n_7351),
.C(n_7375),
.Y(n_7397)
);

OR2x2_ASAP7_75t_L g7398 ( 
.A(n_7356),
.B(n_7359),
.Y(n_7398)
);

OAI21xp5_ASAP7_75t_SL g7399 ( 
.A1(n_7344),
.A2(n_1121),
.B(n_1122),
.Y(n_7399)
);

INVx1_ASAP7_75t_L g7400 ( 
.A(n_7367),
.Y(n_7400)
);

NAND3xp33_ASAP7_75t_L g7401 ( 
.A(n_7349),
.B(n_1121),
.C(n_1122),
.Y(n_7401)
);

AND2x2_ASAP7_75t_L g7402 ( 
.A(n_7365),
.B(n_1124),
.Y(n_7402)
);

CKINVDCx16_ASAP7_75t_R g7403 ( 
.A(n_7366),
.Y(n_7403)
);

AOI22xp5_ASAP7_75t_L g7404 ( 
.A1(n_7373),
.A2(n_1129),
.B1(n_1126),
.B2(n_1127),
.Y(n_7404)
);

AOI221xp5_ASAP7_75t_L g7405 ( 
.A1(n_7352),
.A2(n_1131),
.B1(n_1126),
.B2(n_1127),
.C(n_1132),
.Y(n_7405)
);

NOR3xp33_ASAP7_75t_L g7406 ( 
.A(n_7382),
.B(n_7364),
.C(n_7360),
.Y(n_7406)
);

NOR2x1_ASAP7_75t_L g7407 ( 
.A(n_7383),
.B(n_7378),
.Y(n_7407)
);

NAND2xp5_ASAP7_75t_L g7408 ( 
.A(n_7386),
.B(n_7381),
.Y(n_7408)
);

AND2x2_ASAP7_75t_L g7409 ( 
.A(n_7384),
.B(n_7380),
.Y(n_7409)
);

NOR2x1_ASAP7_75t_L g7410 ( 
.A(n_7397),
.B(n_7377),
.Y(n_7410)
);

NAND3xp33_ASAP7_75t_SL g7411 ( 
.A(n_7387),
.B(n_7362),
.C(n_7363),
.Y(n_7411)
);

NAND2xp5_ASAP7_75t_L g7412 ( 
.A(n_7391),
.B(n_1131),
.Y(n_7412)
);

NAND2xp5_ASAP7_75t_L g7413 ( 
.A(n_7390),
.B(n_1133),
.Y(n_7413)
);

HB1xp67_ASAP7_75t_L g7414 ( 
.A(n_7385),
.Y(n_7414)
);

INVx2_ASAP7_75t_L g7415 ( 
.A(n_7402),
.Y(n_7415)
);

AND2x2_ASAP7_75t_L g7416 ( 
.A(n_7395),
.B(n_1133),
.Y(n_7416)
);

AND3x4_ASAP7_75t_L g7417 ( 
.A(n_7406),
.B(n_1134),
.C(n_1135),
.Y(n_7417)
);

NAND3xp33_ASAP7_75t_L g7418 ( 
.A(n_7393),
.B(n_1134),
.C(n_1136),
.Y(n_7418)
);

OAI22xp5_ASAP7_75t_L g7419 ( 
.A1(n_7398),
.A2(n_1139),
.B1(n_1137),
.B2(n_1138),
.Y(n_7419)
);

NAND3xp33_ASAP7_75t_SL g7420 ( 
.A(n_7396),
.B(n_1138),
.C(n_1139),
.Y(n_7420)
);

NOR2x1_ASAP7_75t_L g7421 ( 
.A(n_7401),
.B(n_1140),
.Y(n_7421)
);

NAND2xp33_ASAP7_75t_SL g7422 ( 
.A(n_7394),
.B(n_1141),
.Y(n_7422)
);

NOR3xp33_ASAP7_75t_L g7423 ( 
.A(n_7403),
.B(n_7392),
.C(n_7388),
.Y(n_7423)
);

NOR3x1_ASAP7_75t_L g7424 ( 
.A(n_7399),
.B(n_1140),
.C(n_1142),
.Y(n_7424)
);

INVxp67_ASAP7_75t_L g7425 ( 
.A(n_7389),
.Y(n_7425)
);

AND2x4_ASAP7_75t_L g7426 ( 
.A(n_7407),
.B(n_7400),
.Y(n_7426)
);

NOR2x1_ASAP7_75t_L g7427 ( 
.A(n_7418),
.B(n_7405),
.Y(n_7427)
);

NOR4xp75_ASAP7_75t_L g7428 ( 
.A(n_7408),
.B(n_7404),
.C(n_1145),
.D(n_1143),
.Y(n_7428)
);

AND3x2_ASAP7_75t_L g7429 ( 
.A(n_7414),
.B(n_1143),
.C(n_1144),
.Y(n_7429)
);

AND2x2_ASAP7_75t_SL g7430 ( 
.A(n_7409),
.B(n_1146),
.Y(n_7430)
);

NOR3xp33_ASAP7_75t_L g7431 ( 
.A(n_7425),
.B(n_7423),
.C(n_7413),
.Y(n_7431)
);

NOR2xp33_ASAP7_75t_R g7432 ( 
.A(n_7411),
.B(n_1146),
.Y(n_7432)
);

NAND3xp33_ASAP7_75t_SL g7433 ( 
.A(n_7417),
.B(n_1155),
.C(n_1147),
.Y(n_7433)
);

OR2x2_ASAP7_75t_L g7434 ( 
.A(n_7420),
.B(n_7422),
.Y(n_7434)
);

HB1xp67_ASAP7_75t_L g7435 ( 
.A(n_7410),
.Y(n_7435)
);

INVx1_ASAP7_75t_L g7436 ( 
.A(n_7415),
.Y(n_7436)
);

OAI21xp5_ASAP7_75t_L g7437 ( 
.A1(n_7421),
.A2(n_1148),
.B(n_1149),
.Y(n_7437)
);

NAND4xp75_ASAP7_75t_L g7438 ( 
.A(n_7424),
.B(n_1151),
.C(n_1149),
.D(n_1150),
.Y(n_7438)
);

NAND3x1_ASAP7_75t_SL g7439 ( 
.A(n_7416),
.B(n_1150),
.C(n_1151),
.Y(n_7439)
);

NAND2xp5_ASAP7_75t_L g7440 ( 
.A(n_7430),
.B(n_7419),
.Y(n_7440)
);

INVx1_ASAP7_75t_L g7441 ( 
.A(n_7435),
.Y(n_7441)
);

OR2x2_ASAP7_75t_L g7442 ( 
.A(n_7433),
.B(n_7412),
.Y(n_7442)
);

INVxp67_ASAP7_75t_SL g7443 ( 
.A(n_7436),
.Y(n_7443)
);

NAND2xp5_ASAP7_75t_L g7444 ( 
.A(n_7429),
.B(n_1152),
.Y(n_7444)
);

AOI22xp33_ASAP7_75t_L g7445 ( 
.A1(n_7441),
.A2(n_7431),
.B1(n_7426),
.B2(n_7434),
.Y(n_7445)
);

OA22x2_ASAP7_75t_L g7446 ( 
.A1(n_7443),
.A2(n_7437),
.B1(n_7439),
.B2(n_7428),
.Y(n_7446)
);

AOI22xp5_ASAP7_75t_L g7447 ( 
.A1(n_7440),
.A2(n_7427),
.B1(n_7444),
.B2(n_7438),
.Y(n_7447)
);

INVxp67_ASAP7_75t_L g7448 ( 
.A(n_7442),
.Y(n_7448)
);

INVx1_ASAP7_75t_L g7449 ( 
.A(n_7446),
.Y(n_7449)
);

NOR3xp33_ASAP7_75t_L g7450 ( 
.A(n_7448),
.B(n_7432),
.C(n_1152),
.Y(n_7450)
);

NAND4xp25_ASAP7_75t_L g7451 ( 
.A(n_7450),
.B(n_7445),
.C(n_7447),
.D(n_1155),
.Y(n_7451)
);

HB1xp67_ASAP7_75t_L g7452 ( 
.A(n_7449),
.Y(n_7452)
);

HB1xp67_ASAP7_75t_L g7453 ( 
.A(n_7452),
.Y(n_7453)
);

OAI22xp5_ASAP7_75t_L g7454 ( 
.A1(n_7451),
.A2(n_1156),
.B1(n_1153),
.B2(n_1154),
.Y(n_7454)
);

INVx1_ASAP7_75t_SL g7455 ( 
.A(n_7453),
.Y(n_7455)
);

INVx1_ASAP7_75t_L g7456 ( 
.A(n_7454),
.Y(n_7456)
);

INVx1_ASAP7_75t_L g7457 ( 
.A(n_7455),
.Y(n_7457)
);

NAND2x1p5_ASAP7_75t_L g7458 ( 
.A(n_7457),
.B(n_7456),
.Y(n_7458)
);

INVxp67_ASAP7_75t_SL g7459 ( 
.A(n_7457),
.Y(n_7459)
);

NAND2xp5_ASAP7_75t_L g7460 ( 
.A(n_7459),
.B(n_1153),
.Y(n_7460)
);

OAI21xp5_ASAP7_75t_SL g7461 ( 
.A1(n_7458),
.A2(n_1154),
.B(n_1157),
.Y(n_7461)
);

BUFx6f_ASAP7_75t_L g7462 ( 
.A(n_7460),
.Y(n_7462)
);

OAI222xp33_ASAP7_75t_L g7463 ( 
.A1(n_7461),
.A2(n_1161),
.B1(n_1164),
.B2(n_1158),
.C1(n_1159),
.C2(n_1162),
.Y(n_7463)
);

OR2x6_ASAP7_75t_L g7464 ( 
.A(n_7462),
.B(n_1158),
.Y(n_7464)
);

AOI21xp5_ASAP7_75t_L g7465 ( 
.A1(n_7463),
.A2(n_1159),
.B(n_1164),
.Y(n_7465)
);

AOI221xp5_ASAP7_75t_L g7466 ( 
.A1(n_7465),
.A2(n_1167),
.B1(n_1165),
.B2(n_1166),
.C(n_1169),
.Y(n_7466)
);

AOI211xp5_ASAP7_75t_L g7467 ( 
.A1(n_7466),
.A2(n_7464),
.B(n_1167),
.C(n_1165),
.Y(n_7467)
);


endmodule