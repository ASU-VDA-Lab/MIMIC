module fake_jpeg_18119_n_31 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_31);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_31;

wire n_13;
wire n_21;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_11;
wire n_17;
wire n_25;
wire n_29;
wire n_12;
wire n_15;

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_9),
.B(n_0),
.Y(n_10)
);

HAxp5_ASAP7_75t_SL g11 ( 
.A(n_1),
.B(n_2),
.CON(n_11),
.SN(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

AND2x2_ASAP7_75t_L g13 ( 
.A(n_6),
.B(n_5),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_1),
.B(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_4),
.B(n_3),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_14),
.A2(n_7),
.B1(n_16),
.B2(n_12),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_24),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_17),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_23),
.Y(n_26)
);

NAND3xp33_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_10),
.C(n_19),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_25),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_19),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_13),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_16),
.A2(n_11),
.B1(n_13),
.B2(n_18),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_20),
.C(n_21),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_29),
.A2(n_26),
.B1(n_28),
.B2(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);


endmodule