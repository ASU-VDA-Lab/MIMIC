module fake_jpeg_16839_n_356 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_356);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_356;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_43),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_22),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_48),
.Y(n_58)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_26),
.B(n_0),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_34),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_67),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_34),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_69),
.B(n_36),
.Y(n_106)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_75),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_55),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_78),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_44),
.B(n_32),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_71),
.A2(n_52),
.B1(n_49),
.B2(n_56),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_88),
.A2(n_74),
.B1(n_64),
.B2(n_65),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_44),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_94),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_71),
.A2(n_29),
.B1(n_20),
.B2(n_28),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_91),
.A2(n_92),
.B1(n_115),
.B2(n_116),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_29),
.B1(n_20),
.B2(n_28),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_43),
.Y(n_94)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_62),
.B(n_37),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_101),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_30),
.Y(n_99)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_86),
.A2(n_37),
.B(n_35),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_100),
.A2(n_25),
.B(n_51),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_20),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_57),
.A2(n_29),
.B1(n_53),
.B2(n_26),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_104),
.A2(n_105),
.B1(n_113),
.B2(n_25),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_57),
.A2(n_53),
.B1(n_32),
.B2(n_30),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_106),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_86),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_111),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_33),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_70),
.A2(n_31),
.B1(n_24),
.B2(n_23),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_45),
.B1(n_38),
.B2(n_36),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_85),
.A2(n_45),
.B1(n_31),
.B2(n_23),
.Y(n_116)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_93),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_118),
.B(n_134),
.Y(n_164)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_123),
.Y(n_152)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_126),
.A2(n_145),
.B1(n_63),
.B2(n_107),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_90),
.A2(n_24),
.B(n_25),
.C(n_21),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_127),
.A2(n_141),
.B(n_147),
.Y(n_171)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_95),
.Y(n_129)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_130),
.A2(n_140),
.B1(n_114),
.B2(n_108),
.Y(n_159)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

FAx1_ASAP7_75t_SL g134 ( 
.A(n_94),
.B(n_50),
.CI(n_51),
.CON(n_134),
.SN(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_93),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_139),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_50),
.C(n_81),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_100),
.C(n_82),
.Y(n_157)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_96),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_89),
.B(n_21),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_142),
.Y(n_165)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_108),
.A2(n_63),
.B1(n_25),
.B2(n_38),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_101),
.B(n_64),
.Y(n_146)
);

AND2x2_ASAP7_75t_SL g158 ( 
.A(n_146),
.B(n_110),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_111),
.A2(n_82),
.B(n_61),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_115),
.A2(n_68),
.B1(n_65),
.B2(n_38),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_114),
.B1(n_95),
.B2(n_88),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_149),
.A2(n_159),
.B1(n_129),
.B2(n_117),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_150),
.B(n_151),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_121),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_173),
.C(n_148),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_134),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_123),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_167),
.A2(n_120),
.B1(n_126),
.B2(n_129),
.Y(n_180)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_172),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_97),
.C(n_80),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_154),
.Y(n_174)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_174),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_171),
.A2(n_131),
.B1(n_147),
.B2(n_124),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_134),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_197),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_119),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_180),
.A2(n_191),
.B(n_167),
.Y(n_216)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_171),
.A2(n_131),
.B1(n_124),
.B2(n_146),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_182),
.B(n_187),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_188),
.Y(n_209)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_185),
.Y(n_198)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_122),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_122),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_195),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_157),
.A2(n_149),
.B1(n_164),
.B2(n_130),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_190),
.B(n_192),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_165),
.A2(n_141),
.B(n_137),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_119),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_153),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_194),
.B(n_150),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_127),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_97),
.Y(n_197)
);

OR2x4_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_89),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_199),
.A2(n_216),
.B(n_215),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_221),
.C(n_178),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_161),
.Y(n_205)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_195),
.B(n_125),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_207),
.B(n_214),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_151),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_217),
.Y(n_232)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_197),
.B(n_99),
.Y(n_214)
);

XNOR2x2_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_106),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_215),
.B(n_178),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_179),
.B(n_163),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_176),
.B(n_170),
.Y(n_218)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_170),
.Y(n_219)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_156),
.Y(n_220)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_155),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_166),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_203),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_163),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_174),
.Y(n_235)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_224),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_219),
.B(n_185),
.Y(n_225)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

NAND3xp33_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_191),
.C(n_106),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_SL g261 ( 
.A(n_227),
.B(n_238),
.C(n_107),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_198),
.B(n_194),
.Y(n_228)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_228),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_206),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_240),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_235),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_236),
.B(n_144),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_212),
.Y(n_237)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_152),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_201),
.B(n_183),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_183),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_242),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_174),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_154),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_246),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_154),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_208),
.B(n_181),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_248),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_204),
.B(n_166),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_248),
.A2(n_204),
.B1(n_224),
.B2(n_233),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_249),
.A2(n_250),
.B1(n_251),
.B2(n_255),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_233),
.A2(n_205),
.B1(n_218),
.B2(n_202),
.Y(n_250)
);

XOR2x2_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_226),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_259),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_234),
.A2(n_216),
.B1(n_221),
.B2(n_205),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_243),
.B(n_162),
.Y(n_256)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_256),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_234),
.A2(n_218),
.B1(n_208),
.B2(n_211),
.Y(n_257)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_257),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_243),
.B(n_211),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_245),
.A2(n_153),
.B1(n_162),
.B2(n_172),
.Y(n_260)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_260),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_266),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_232),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_262),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_236),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_239),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_278),
.C(n_284),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_251),
.A2(n_226),
.B1(n_230),
.B2(n_229),
.Y(n_276)
);

XNOR2x1_ASAP7_75t_L g304 ( 
.A(n_276),
.B(n_287),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_268),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_277),
.B(n_1),
.Y(n_300)
);

AOI21xp33_ASAP7_75t_L g281 ( 
.A1(n_263),
.A2(n_229),
.B(n_231),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_281),
.A2(n_270),
.B(n_2),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_254),
.A2(n_245),
.B1(n_225),
.B2(n_230),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_282),
.A2(n_38),
.B1(n_59),
.B2(n_60),
.Y(n_305)
);

NOR3xp33_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_232),
.C(n_237),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_264),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_250),
.B(n_228),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_252),
.B(n_247),
.Y(n_285)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_285),
.Y(n_292)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_267),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_289),
.Y(n_291)
);

OAI21xp33_ASAP7_75t_L g287 ( 
.A1(n_253),
.A2(n_152),
.B(n_103),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_260),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_265),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_262),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_273),
.B(n_266),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_293),
.B(n_306),
.Y(n_316)
);

OA21x2_ASAP7_75t_L g294 ( 
.A1(n_276),
.A2(n_249),
.B(n_288),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_294),
.B(n_60),
.Y(n_317)
);

AOI221xp5_ASAP7_75t_L g295 ( 
.A1(n_279),
.A2(n_255),
.B1(n_257),
.B2(n_287),
.C(n_271),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_295),
.A2(n_272),
.B1(n_5),
.B2(n_6),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_300),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_297),
.A2(n_299),
.B1(n_302),
.B2(n_303),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_132),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_7),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_280),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_284),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_305),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_272),
.B(n_4),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_304),
.A2(n_291),
.B1(n_292),
.B2(n_294),
.Y(n_307)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_307),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_274),
.C(n_278),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_309),
.C(n_314),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_274),
.C(n_282),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_9),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_311),
.B(n_315),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_304),
.A2(n_5),
.B(n_7),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_312),
.A2(n_10),
.B(n_11),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_59),
.C(n_61),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_318),
.Y(n_323)
);

INVx11_ASAP7_75t_L g318 ( 
.A(n_294),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_303),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_320),
.B(n_306),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_329),
.Y(n_334)
);

AO21x1_ASAP7_75t_L g324 ( 
.A1(n_313),
.A2(n_8),
.B(n_9),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_324),
.B(n_325),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_326),
.A2(n_10),
.B(n_11),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_309),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_308),
.B(n_39),
.C(n_61),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_330),
.B(n_314),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_307),
.B(n_10),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_331),
.B(n_12),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_332),
.B(n_339),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_321),
.B(n_316),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_333),
.B(n_323),
.C(n_39),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_329),
.A2(n_318),
.B(n_319),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_336),
.A2(n_323),
.B(n_15),
.Y(n_344)
);

OAI21x1_ASAP7_75t_L g337 ( 
.A1(n_327),
.A2(n_317),
.B(n_316),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_337),
.B(n_338),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_328),
.B(n_13),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_340),
.B(n_14),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_341),
.B(n_345),
.Y(n_349)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_343),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_344),
.Y(n_348)
);

AOI21xp33_ASAP7_75t_L g345 ( 
.A1(n_334),
.A2(n_39),
.B(n_15),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_349),
.B(n_334),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_350),
.B(n_351),
.C(n_335),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_348),
.A2(n_342),
.B(n_346),
.Y(n_351)
);

AOI322xp5_ASAP7_75t_L g353 ( 
.A1(n_352),
.A2(n_347),
.A3(n_21),
.B1(n_17),
.B2(n_16),
.C1(n_14),
.C2(n_83),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_353),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_354),
.B(n_14),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_355),
.B(n_83),
.Y(n_356)
);


endmodule