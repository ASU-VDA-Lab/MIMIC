module fake_jpeg_1776_n_91 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_91);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_91;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NAND2xp33_ASAP7_75t_SL g38 ( 
.A(n_35),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_28),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_50),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_34),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_27),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_36),
.C(n_31),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_36),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_55),
.B(n_56),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_1),
.Y(n_56)
);

AND2x6_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_14),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_57),
.B(n_58),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_2),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_43),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_61),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_67),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_57),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_55),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_63),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_33),
.B1(n_32),
.B2(n_30),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_69),
.A2(n_30),
.B1(n_33),
.B2(n_32),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_71),
.B(n_72),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g74 ( 
.A1(n_64),
.A2(n_12),
.B(n_25),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_74),
.A2(n_77),
.B(n_78),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_76),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_66),
.B(n_2),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_3),
.B(n_4),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_4),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_17),
.C(n_26),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_79),
.A2(n_74),
.B(n_19),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_84),
.C(n_82),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_80),
.A2(n_70),
.B1(n_61),
.B2(n_78),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_85),
.A2(n_81),
.B1(n_11),
.B2(n_7),
.Y(n_86)
);

OAI31xp33_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_13),
.A3(n_23),
.B(n_9),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_10),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_21),
.C(n_24),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_5),
.Y(n_90)
);

BUFx24_ASAP7_75t_SL g91 ( 
.A(n_90),
.Y(n_91)
);


endmodule