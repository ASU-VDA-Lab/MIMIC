module fake_jpeg_1940_n_44 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_44);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;
wire n_15;

BUFx10_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_0),
.B(n_8),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_9),
.A2(n_0),
.B1(n_8),
.B2(n_2),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_5),
.B(n_1),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_L g18 ( 
.A1(n_13),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_22),
.A2(n_13),
.B1(n_14),
.B2(n_17),
.Y(n_25)
);

OAI22x1_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_13),
.B1(n_15),
.B2(n_5),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_17),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_12),
.Y(n_29)
);

AOI32xp33_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_16),
.A3(n_21),
.B1(n_13),
.B2(n_15),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_28),
.B(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_13),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_28),
.B(n_26),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_35),
.A2(n_36),
.B(n_11),
.Y(n_39)
);

OR2x6_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_30),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_38),
.Y(n_41)
);

FAx1_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_15),
.CI(n_26),
.CON(n_38),
.SN(n_38)
);

AOI322xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_33),
.A3(n_7),
.B1(n_9),
.B2(n_10),
.C1(n_6),
.C2(n_36),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_6),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_42),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_41),
.Y(n_44)
);


endmodule