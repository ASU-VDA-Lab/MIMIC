module fake_netlist_6_4776_n_807 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_807);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_807;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_698;
wire n_617;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_683;
wire n_620;
wire n_420;
wire n_608;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_25),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_105),
.Y(n_167)
);

INVxp33_ASAP7_75t_SL g168 ( 
.A(n_51),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_102),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_87),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_82),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_118),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_130),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_50),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_122),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_81),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_20),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_72),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_127),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_31),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_28),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_108),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_126),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_159),
.Y(n_189)
);

BUFx2_ASAP7_75t_SL g190 ( 
.A(n_69),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_61),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_80),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_84),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_35),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_53),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_146),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_76),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_147),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_111),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_67),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_19),
.Y(n_201)
);

BUFx10_ASAP7_75t_L g202 ( 
.A(n_26),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_10),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_66),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_17),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_63),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_38),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_137),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_160),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_65),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_52),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_20),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_40),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_27),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_59),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_134),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_148),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_34),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_154),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_151),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_123),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_62),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_142),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_144),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_1),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_145),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_129),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_121),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_136),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_98),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_104),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_128),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_132),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_97),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_54),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_150),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_114),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_201),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

AND2x6_ASAP7_75t_L g240 ( 
.A(n_178),
.B(n_22),
.Y(n_240)
);

BUFx12f_ASAP7_75t_L g241 ( 
.A(n_202),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_169),
.B(n_192),
.Y(n_242)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_178),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_212),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_184),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_0),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_178),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_205),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_180),
.Y(n_250)
);

OAI22x1_ASAP7_75t_R g251 ( 
.A1(n_180),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_184),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_211),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_253)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_202),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_178),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_232),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_232),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_219),
.B(n_3),
.Y(n_258)
);

NAND2xp33_ASAP7_75t_L g259 ( 
.A(n_222),
.B(n_4),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_222),
.Y(n_260)
);

AND2x6_ASAP7_75t_L g261 ( 
.A(n_222),
.B(n_23),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_171),
.B(n_176),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_222),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_202),
.B(n_5),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_213),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_211),
.B(n_6),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_213),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_171),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_176),
.Y(n_269)
);

AND2x4_ASAP7_75t_L g270 ( 
.A(n_182),
.B(n_199),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_218),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_182),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_199),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_207),
.Y(n_274)
);

BUFx8_ASAP7_75t_SL g275 ( 
.A(n_218),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_166),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_207),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_208),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_208),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_167),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_166),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_170),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_172),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_173),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_174),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_175),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_183),
.B(n_223),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_268),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_275),
.Y(n_289)
);

OR2x6_ASAP7_75t_L g290 ( 
.A(n_241),
.B(n_190),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_264),
.B(n_168),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_266),
.B(n_168),
.Y(n_292)
);

NAND2xp33_ASAP7_75t_L g293 ( 
.A(n_258),
.B(n_172),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_254),
.B(n_177),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_263),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_252),
.B(n_7),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_268),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_254),
.B(n_221),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_250),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_250),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_268),
.Y(n_301)
);

INVxp33_ASAP7_75t_L g302 ( 
.A(n_276),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_L g303 ( 
.A1(n_242),
.A2(n_253),
.B1(n_249),
.B2(n_281),
.Y(n_303)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_248),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_263),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_283),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_268),
.Y(n_307)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_248),
.Y(n_308)
);

BUFx6f_ASAP7_75t_SL g309 ( 
.A(n_252),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_275),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_179),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_273),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_273),
.Y(n_313)
);

NOR2x1p5_ASAP7_75t_L g314 ( 
.A(n_241),
.B(n_221),
.Y(n_314)
);

AND2x2_ASAP7_75t_SL g315 ( 
.A(n_259),
.B(n_181),
.Y(n_315)
);

OR2x6_ASAP7_75t_L g316 ( 
.A(n_265),
.B(n_186),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_273),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_247),
.B(n_224),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_239),
.Y(n_319)
);

OR2x6_ASAP7_75t_L g320 ( 
.A(n_267),
.B(n_237),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_273),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_277),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_287),
.B(n_187),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_277),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_277),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_246),
.Y(n_326)
);

NAND3xp33_ASAP7_75t_L g327 ( 
.A(n_247),
.B(n_231),
.C(n_224),
.Y(n_327)
);

AND2x6_ASAP7_75t_L g328 ( 
.A(n_270),
.B(n_248),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_270),
.B(n_227),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_277),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_279),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_248),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_262),
.B(n_189),
.Y(n_333)
);

AO21x2_ASAP7_75t_L g334 ( 
.A1(n_259),
.A2(n_210),
.B(n_235),
.Y(n_334)
);

NOR3xp33_ASAP7_75t_L g335 ( 
.A(n_271),
.B(n_236),
.C(n_234),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_256),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_333),
.B(n_270),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_312),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_279),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_292),
.B(n_281),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_326),
.Y(n_341)
);

INVxp33_ASAP7_75t_L g342 ( 
.A(n_302),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_326),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_312),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_336),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_313),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_292),
.B(n_227),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_306),
.B(n_231),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_291),
.A2(n_185),
.B1(n_188),
.B2(n_193),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_336),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_291),
.A2(n_198),
.B1(n_196),
.B2(n_195),
.Y(n_351)
);

O2A1O1Ixp33_ASAP7_75t_L g352 ( 
.A1(n_311),
.A2(n_245),
.B(n_238),
.C(n_244),
.Y(n_352)
);

NAND3xp33_ASAP7_75t_L g353 ( 
.A(n_323),
.B(n_257),
.C(n_280),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_295),
.B(n_279),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_289),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_288),
.Y(n_356)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_328),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_295),
.B(n_269),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_335),
.A2(n_191),
.B1(n_228),
.B2(n_229),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_289),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_319),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_297),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_298),
.B(n_280),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_299),
.B(n_194),
.Y(n_364)
);

OR2x2_ASAP7_75t_L g365 ( 
.A(n_329),
.B(n_284),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_305),
.B(n_301),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_302),
.B(n_284),
.Y(n_367)
);

INVx8_ASAP7_75t_L g368 ( 
.A(n_290),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_318),
.A2(n_197),
.B1(n_200),
.B2(n_204),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_305),
.B(n_269),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_328),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_300),
.B(n_206),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_298),
.B(n_285),
.Y(n_373)
);

NAND3xp33_ASAP7_75t_L g374 ( 
.A(n_318),
.B(n_285),
.C(n_286),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_332),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_307),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_313),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_320),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_327),
.B(n_209),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g380 ( 
.A(n_329),
.B(n_238),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_321),
.Y(n_381)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_328),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_303),
.B(n_215),
.Y(n_383)
);

OAI22xp33_ASAP7_75t_L g384 ( 
.A1(n_316),
.A2(n_216),
.B1(n_217),
.B2(n_220),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_315),
.B(n_243),
.Y(n_385)
);

INVxp67_ASAP7_75t_SL g386 ( 
.A(n_304),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_293),
.A2(n_226),
.B1(n_230),
.B2(n_233),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_303),
.B(n_282),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_294),
.B(n_282),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_317),
.B(n_272),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_293),
.A2(n_261),
.B1(n_240),
.B2(n_244),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_320),
.A2(n_261),
.B1(n_240),
.B2(n_286),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_320),
.B(n_282),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_322),
.B(n_272),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_315),
.B(n_296),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_L g396 ( 
.A1(n_334),
.A2(n_286),
.B1(n_282),
.B2(n_261),
.Y(n_396)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_290),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_330),
.Y(n_398)
);

NOR2xp67_ASAP7_75t_L g399 ( 
.A(n_349),
.B(n_310),
.Y(n_399)
);

BUFx12f_ASAP7_75t_L g400 ( 
.A(n_355),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_339),
.B(n_334),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_339),
.B(n_324),
.Y(n_402)
);

NOR2x1_ASAP7_75t_L g403 ( 
.A(n_385),
.B(n_290),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_338),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_337),
.B(n_325),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_337),
.B(n_325),
.Y(n_406)
);

AO32x1_ASAP7_75t_L g407 ( 
.A1(n_344),
.A2(n_274),
.A3(n_278),
.B1(n_331),
.B2(n_240),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_367),
.B(n_274),
.Y(n_408)
);

AO21x1_ASAP7_75t_L g409 ( 
.A1(n_395),
.A2(n_278),
.B(n_251),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_363),
.B(n_304),
.Y(n_410)
);

OR2x6_ASAP7_75t_L g411 ( 
.A(n_368),
.B(n_316),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_346),
.Y(n_412)
);

A2O1A1Ixp33_ASAP7_75t_L g413 ( 
.A1(n_373),
.A2(n_314),
.B(n_308),
.C(n_255),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_361),
.B(n_332),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_390),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_342),
.B(n_380),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_377),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_365),
.B(n_332),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_389),
.B(n_308),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_386),
.B(n_332),
.Y(n_420)
);

O2A1O1Ixp33_ASAP7_75t_L g421 ( 
.A1(n_388),
.A2(n_316),
.B(n_261),
.C(n_240),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_356),
.B(n_240),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_362),
.B(n_261),
.Y(n_423)
);

NAND3xp33_ASAP7_75t_SL g424 ( 
.A(n_359),
.B(n_309),
.C(n_9),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_376),
.B(n_255),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_374),
.A2(n_309),
.B(n_260),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_390),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_394),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_383),
.A2(n_260),
.B1(n_9),
.B2(n_10),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_357),
.A2(n_86),
.B(n_165),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_371),
.A2(n_85),
.B(n_163),
.Y(n_431)
);

O2A1O1Ixp5_ASAP7_75t_L g432 ( 
.A1(n_379),
.A2(n_371),
.B(n_347),
.C(n_382),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_382),
.A2(n_83),
.B(n_162),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_398),
.B(n_396),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_366),
.A2(n_79),
.B(n_161),
.Y(n_435)
);

O2A1O1Ixp5_ASAP7_75t_L g436 ( 
.A1(n_364),
.A2(n_78),
.B(n_157),
.C(n_156),
.Y(n_436)
);

BUFx8_ASAP7_75t_L g437 ( 
.A(n_378),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_381),
.Y(n_438)
);

NOR2xp67_ASAP7_75t_L g439 ( 
.A(n_351),
.B(n_24),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_348),
.B(n_8),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_341),
.B(n_8),
.Y(n_441)
);

A2O1A1Ixp33_ASAP7_75t_L g442 ( 
.A1(n_369),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_366),
.A2(n_88),
.B(n_153),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_343),
.B(n_345),
.Y(n_444)
);

A2O1A1Ixp33_ASAP7_75t_L g445 ( 
.A1(n_393),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_350),
.B(n_14),
.Y(n_446)
);

O2A1O1Ixp33_ASAP7_75t_L g447 ( 
.A1(n_352),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_340),
.B(n_15),
.Y(n_448)
);

NAND2x1p5_ASAP7_75t_L g449 ( 
.A(n_392),
.B(n_29),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_394),
.B(n_30),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_353),
.B(n_375),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_391),
.A2(n_91),
.B(n_152),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_372),
.Y(n_453)
);

AOI22xp33_ASAP7_75t_L g454 ( 
.A1(n_387),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_384),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_455)
);

O2A1O1Ixp33_ASAP7_75t_L g456 ( 
.A1(n_358),
.A2(n_21),
.B(n_32),
.C(n_33),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_397),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_375),
.B(n_41),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_368),
.B(n_42),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_375),
.B(n_43),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_368),
.B(n_44),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_358),
.B(n_45),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_354),
.B(n_46),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_370),
.A2(n_47),
.B(n_48),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_360),
.B(n_49),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_415),
.B(n_55),
.Y(n_466)
);

INVxp67_ASAP7_75t_SL g467 ( 
.A(n_434),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_404),
.Y(n_468)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_417),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_401),
.A2(n_56),
.B(n_57),
.Y(n_470)
);

AO21x1_ASAP7_75t_L g471 ( 
.A1(n_452),
.A2(n_58),
.B(n_60),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_417),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_412),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_416),
.B(n_64),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_453),
.B(n_68),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_403),
.B(n_70),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_448),
.B(n_71),
.Y(n_477)
);

AOI211x1_ASAP7_75t_L g478 ( 
.A1(n_409),
.A2(n_143),
.B(n_74),
.C(n_75),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_400),
.Y(n_479)
);

OAI21x1_ASAP7_75t_L g480 ( 
.A1(n_422),
.A2(n_423),
.B(n_432),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_440),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_438),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_405),
.A2(n_406),
.B(n_428),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_427),
.A2(n_73),
.B(n_77),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_458),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_402),
.B(n_89),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_408),
.B(n_90),
.Y(n_487)
);

INVxp67_ASAP7_75t_SL g488 ( 
.A(n_420),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_410),
.B(n_92),
.Y(n_489)
);

NAND3xp33_ASAP7_75t_L g490 ( 
.A(n_421),
.B(n_93),
.C(n_94),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_419),
.A2(n_95),
.B(n_96),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_444),
.Y(n_492)
);

O2A1O1Ixp33_ASAP7_75t_L g493 ( 
.A1(n_445),
.A2(n_99),
.B(n_100),
.C(n_101),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_418),
.A2(n_103),
.B(n_106),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_451),
.A2(n_107),
.B(n_109),
.Y(n_495)
);

AO21x1_ASAP7_75t_L g496 ( 
.A1(n_452),
.A2(n_112),
.B(n_113),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_463),
.A2(n_115),
.B(n_116),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_425),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_399),
.B(n_117),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_441),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_462),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_414),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_450),
.A2(n_119),
.B(n_120),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_460),
.A2(n_124),
.B(n_125),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_413),
.B(n_131),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_465),
.B(n_133),
.Y(n_506)
);

NOR2xp67_ASAP7_75t_L g507 ( 
.A(n_459),
.B(n_135),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_449),
.A2(n_138),
.B(n_139),
.Y(n_508)
);

AOI221xp5_ASAP7_75t_SL g509 ( 
.A1(n_429),
.A2(n_140),
.B1(n_141),
.B2(n_454),
.C(n_442),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_R g510 ( 
.A(n_424),
.B(n_437),
.Y(n_510)
);

OAI21x1_ASAP7_75t_L g511 ( 
.A1(n_433),
.A2(n_431),
.B(n_430),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_446),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_426),
.B(n_449),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_426),
.B(n_439),
.Y(n_514)
);

OAI21x1_ASAP7_75t_L g515 ( 
.A1(n_436),
.A2(n_435),
.B(n_443),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_461),
.B(n_429),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_455),
.A2(n_411),
.B1(n_457),
.B2(n_447),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_492),
.B(n_455),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_472),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_477),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_469),
.Y(n_521)
);

NOR2x1_ASAP7_75t_SL g522 ( 
.A(n_501),
.B(n_411),
.Y(n_522)
);

NAND2x1p5_ASAP7_75t_L g523 ( 
.A(n_469),
.B(n_464),
.Y(n_523)
);

AOI21x1_ASAP7_75t_L g524 ( 
.A1(n_489),
.A2(n_407),
.B(n_411),
.Y(n_524)
);

AO31x2_ASAP7_75t_L g525 ( 
.A1(n_471),
.A2(n_407),
.A3(n_456),
.B(n_437),
.Y(n_525)
);

OA21x2_ASAP7_75t_L g526 ( 
.A1(n_483),
.A2(n_407),
.B(n_509),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_472),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_467),
.B(n_500),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_481),
.B(n_483),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_468),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_488),
.A2(n_486),
.B(n_466),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_466),
.A2(n_513),
.B(n_514),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_510),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_473),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_482),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_474),
.B(n_512),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_502),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_516),
.B(n_475),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_516),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_507),
.A2(n_505),
.B(n_498),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_477),
.B(n_487),
.Y(n_541)
);

OAI21x1_ASAP7_75t_L g542 ( 
.A1(n_508),
.A2(n_470),
.B(n_491),
.Y(n_542)
);

AO21x1_ASAP7_75t_L g543 ( 
.A1(n_484),
.A2(n_517),
.B(n_493),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_479),
.Y(n_544)
);

AO31x2_ASAP7_75t_L g545 ( 
.A1(n_496),
.A2(n_517),
.A3(n_495),
.B(n_503),
.Y(n_545)
);

OAI21x1_ASAP7_75t_L g546 ( 
.A1(n_504),
.A2(n_494),
.B(n_497),
.Y(n_546)
);

AO21x2_ASAP7_75t_L g547 ( 
.A1(n_484),
.A2(n_490),
.B(n_476),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_506),
.B(n_499),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_485),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_SL g550 ( 
.A1(n_485),
.A2(n_479),
.B(n_478),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_485),
.Y(n_551)
);

CKINVDCx6p67_ASAP7_75t_R g552 ( 
.A(n_479),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_468),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_480),
.A2(n_511),
.B(n_515),
.Y(n_554)
);

AOI21xp33_ASAP7_75t_L g555 ( 
.A1(n_516),
.A2(n_340),
.B(n_481),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_492),
.B(n_467),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_474),
.A2(n_477),
.B1(n_481),
.B2(n_475),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_468),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_539),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_521),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_539),
.B(n_538),
.Y(n_561)
);

AND2x2_ASAP7_75t_SL g562 ( 
.A(n_548),
.B(n_557),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_520),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_541),
.B(n_549),
.Y(n_564)
);

OR2x2_ASAP7_75t_L g565 ( 
.A(n_529),
.B(n_556),
.Y(n_565)
);

INVx1_ASAP7_75t_SL g566 ( 
.A(n_544),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_519),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_519),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_528),
.B(n_518),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_527),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_527),
.Y(n_571)
);

OR2x2_ASAP7_75t_L g572 ( 
.A(n_536),
.B(n_555),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_537),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_530),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_521),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_534),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_526),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_544),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_548),
.B(n_535),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_553),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_533),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_558),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_551),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_526),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_526),
.Y(n_585)
);

NOR2x1_ASAP7_75t_SL g586 ( 
.A(n_547),
.B(n_524),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_543),
.Y(n_587)
);

OR2x6_ASAP7_75t_L g588 ( 
.A(n_550),
.B(n_532),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_545),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_547),
.B(n_545),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_522),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_545),
.B(n_532),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_545),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_523),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_561),
.B(n_525),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_559),
.Y(n_596)
);

INVx5_ASAP7_75t_L g597 ( 
.A(n_588),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_563),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_563),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_578),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_583),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_561),
.B(n_531),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_578),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_569),
.B(n_531),
.Y(n_604)
);

OR2x2_ASAP7_75t_L g605 ( 
.A(n_572),
.B(n_525),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_565),
.B(n_540),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_583),
.Y(n_607)
);

INVx1_ASAP7_75t_SL g608 ( 
.A(n_566),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_559),
.Y(n_609)
);

BUFx5_ASAP7_75t_L g610 ( 
.A(n_584),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_584),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_578),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_562),
.B(n_525),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_567),
.Y(n_614)
);

INVx5_ASAP7_75t_L g615 ( 
.A(n_588),
.Y(n_615)
);

NOR2x1_ASAP7_75t_L g616 ( 
.A(n_572),
.B(n_540),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_567),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_580),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_585),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_585),
.Y(n_620)
);

NOR2x2_ASAP7_75t_L g621 ( 
.A(n_580),
.B(n_533),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_562),
.B(n_525),
.Y(n_622)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_587),
.B(n_554),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_577),
.Y(n_624)
);

HB1xp67_ASAP7_75t_L g625 ( 
.A(n_564),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_560),
.Y(n_626)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_564),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_587),
.B(n_523),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_568),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_565),
.B(n_579),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_564),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_577),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_562),
.B(n_542),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_564),
.B(n_546),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_568),
.B(n_552),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_560),
.B(n_575),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_560),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_570),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_570),
.B(n_571),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_601),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_595),
.B(n_590),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_607),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_626),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_595),
.B(n_590),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_605),
.B(n_611),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_613),
.B(n_592),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_596),
.Y(n_647)
);

OR2x6_ASAP7_75t_L g648 ( 
.A(n_633),
.B(n_588),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_613),
.B(n_592),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_622),
.B(n_593),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_625),
.B(n_582),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_596),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_609),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_611),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_622),
.B(n_593),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_619),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_598),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_605),
.B(n_589),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_609),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_610),
.Y(n_660)
);

BUFx6f_ASAP7_75t_SL g661 ( 
.A(n_600),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_610),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_610),
.Y(n_663)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_619),
.B(n_589),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_610),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_626),
.Y(n_666)
);

NAND2x1_ASAP7_75t_L g667 ( 
.A(n_616),
.B(n_588),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_620),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_620),
.Y(n_669)
);

NOR2x1_ASAP7_75t_L g670 ( 
.A(n_630),
.B(n_612),
.Y(n_670)
);

NAND2x1_ASAP7_75t_L g671 ( 
.A(n_616),
.B(n_594),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_610),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_633),
.B(n_627),
.Y(n_673)
);

BUFx2_ASAP7_75t_L g674 ( 
.A(n_610),
.Y(n_674)
);

AND2x4_ASAP7_75t_SL g675 ( 
.A(n_599),
.B(n_591),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_610),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_624),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_610),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_624),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_654),
.Y(n_680)
);

NAND2x1p5_ASAP7_75t_L g681 ( 
.A(n_670),
.B(n_597),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_651),
.B(n_597),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_654),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_657),
.B(n_602),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_640),
.B(n_642),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_651),
.B(n_606),
.Y(n_686)
);

NAND2x1p5_ASAP7_75t_L g687 ( 
.A(n_667),
.B(n_615),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_656),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_651),
.B(n_631),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_656),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_647),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_641),
.B(n_604),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_641),
.B(n_628),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_652),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_653),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_644),
.B(n_673),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_644),
.B(n_618),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_673),
.B(n_634),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_646),
.B(n_634),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_659),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_668),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_648),
.B(n_615),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_669),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_646),
.B(n_618),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_677),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_649),
.B(n_650),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_649),
.B(n_632),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_658),
.B(n_650),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_677),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_664),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_645),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_679),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_658),
.B(n_639),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_706),
.B(n_648),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_684),
.B(n_655),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_690),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_690),
.Y(n_717)
);

OR2x2_ASAP7_75t_L g718 ( 
.A(n_696),
.B(n_645),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_692),
.B(n_675),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_680),
.Y(n_720)
);

OR2x2_ASAP7_75t_L g721 ( 
.A(n_708),
.B(n_648),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_712),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_686),
.B(n_655),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_683),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_693),
.B(n_648),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_706),
.B(n_674),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_711),
.B(n_662),
.Y(n_727)
);

OR2x2_ASAP7_75t_L g728 ( 
.A(n_685),
.B(n_662),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_688),
.Y(n_729)
);

INVx1_ASAP7_75t_SL g730 ( 
.A(n_697),
.Y(n_730)
);

NAND2x1p5_ASAP7_75t_L g731 ( 
.A(n_702),
.B(n_597),
.Y(n_731)
);

INVxp67_ASAP7_75t_SL g732 ( 
.A(n_710),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_691),
.Y(n_733)
);

OAI221xp5_ASAP7_75t_L g734 ( 
.A1(n_731),
.A2(n_681),
.B1(n_687),
.B2(n_608),
.C(n_682),
.Y(n_734)
);

OR2x2_ASAP7_75t_L g735 ( 
.A(n_718),
.B(n_710),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_720),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_731),
.A2(n_667),
.B(n_615),
.Y(n_737)
);

NAND3xp33_ASAP7_75t_SL g738 ( 
.A(n_730),
.B(n_681),
.C(n_687),
.Y(n_738)
);

OAI21xp5_ASAP7_75t_L g739 ( 
.A1(n_719),
.A2(n_682),
.B(n_671),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_724),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_729),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_719),
.B(n_704),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_723),
.B(n_699),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_SL g744 ( 
.A(n_732),
.B(n_597),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_722),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_714),
.B(n_699),
.Y(n_746)
);

AOI211xp5_ASAP7_75t_L g747 ( 
.A1(n_734),
.A2(n_728),
.B(n_721),
.C(n_733),
.Y(n_747)
);

AOI222xp33_ASAP7_75t_L g748 ( 
.A1(n_738),
.A2(n_715),
.B1(n_732),
.B2(n_689),
.C1(n_702),
.C2(n_726),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_SL g749 ( 
.A1(n_739),
.A2(n_581),
.B1(n_621),
.B2(n_702),
.Y(n_749)
);

OAI221xp5_ASAP7_75t_SL g750 ( 
.A1(n_737),
.A2(n_725),
.B1(n_727),
.B2(n_726),
.C(n_703),
.Y(n_750)
);

AOI221x1_ASAP7_75t_L g751 ( 
.A1(n_739),
.A2(n_722),
.B1(n_717),
.B2(n_716),
.C(n_694),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_742),
.A2(n_661),
.B1(n_698),
.B2(n_707),
.Y(n_752)
);

NAND4xp25_ASAP7_75t_L g753 ( 
.A(n_744),
.B(n_635),
.C(n_695),
.D(n_701),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_736),
.Y(n_754)
);

AOI221xp5_ASAP7_75t_L g755 ( 
.A1(n_747),
.A2(n_740),
.B1(n_741),
.B2(n_735),
.C(n_745),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_754),
.Y(n_756)
);

OAI22xp5_ASAP7_75t_L g757 ( 
.A1(n_749),
.A2(n_743),
.B1(n_661),
.B2(n_713),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_748),
.B(n_746),
.Y(n_758)
);

AOI221xp5_ASAP7_75t_L g759 ( 
.A1(n_750),
.A2(n_753),
.B1(n_752),
.B2(n_744),
.C(n_700),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_751),
.B(n_635),
.Y(n_760)
);

NOR3xp33_ASAP7_75t_L g761 ( 
.A(n_757),
.B(n_671),
.C(n_573),
.Y(n_761)
);

NAND3xp33_ASAP7_75t_L g762 ( 
.A(n_755),
.B(n_705),
.C(n_709),
.Y(n_762)
);

NAND4xp25_ASAP7_75t_L g763 ( 
.A(n_759),
.B(n_573),
.C(n_600),
.D(n_612),
.Y(n_763)
);

NOR4xp25_ASAP7_75t_L g764 ( 
.A(n_758),
.B(n_574),
.C(n_576),
.D(n_717),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_760),
.B(n_716),
.Y(n_765)
);

NAND4xp25_ASAP7_75t_L g766 ( 
.A(n_756),
.B(n_603),
.C(n_574),
.D(n_576),
.Y(n_766)
);

NOR3x1_ASAP7_75t_L g767 ( 
.A(n_763),
.B(n_674),
.C(n_628),
.Y(n_767)
);

NAND4xp75_ASAP7_75t_L g768 ( 
.A(n_765),
.B(n_707),
.C(n_594),
.D(n_639),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_764),
.B(n_675),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_762),
.B(n_712),
.Y(n_770)
);

NAND4xp25_ASAP7_75t_L g771 ( 
.A(n_761),
.B(n_603),
.C(n_582),
.D(n_660),
.Y(n_771)
);

NOR2x1_ASAP7_75t_L g772 ( 
.A(n_769),
.B(n_766),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_768),
.B(n_663),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_770),
.Y(n_774)
);

NOR4xp25_ASAP7_75t_L g775 ( 
.A(n_771),
.B(n_571),
.C(n_678),
.D(n_672),
.Y(n_775)
);

O2A1O1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_767),
.A2(n_663),
.B(n_678),
.C(n_676),
.Y(n_776)
);

NOR2x1_ASAP7_75t_L g777 ( 
.A(n_772),
.B(n_560),
.Y(n_777)
);

XOR2x1_ASAP7_75t_L g778 ( 
.A(n_774),
.B(n_661),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_773),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_775),
.B(n_665),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_776),
.B(n_665),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_774),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_772),
.B(n_636),
.Y(n_783)
);

OA22x2_ASAP7_75t_L g784 ( 
.A1(n_779),
.A2(n_660),
.B1(n_676),
.B2(n_672),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_782),
.B(n_636),
.Y(n_785)
);

OAI21xp33_ASAP7_75t_L g786 ( 
.A1(n_783),
.A2(n_664),
.B(n_679),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_777),
.Y(n_787)
);

AO21x2_ASAP7_75t_L g788 ( 
.A1(n_780),
.A2(n_617),
.B(n_638),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_L g789 ( 
.A1(n_781),
.A2(n_615),
.B1(n_597),
.B2(n_666),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_778),
.Y(n_790)
);

AO22x2_ASAP7_75t_L g791 ( 
.A1(n_779),
.A2(n_617),
.B1(n_638),
.B2(n_629),
.Y(n_791)
);

AOI221xp5_ASAP7_75t_L g792 ( 
.A1(n_790),
.A2(n_636),
.B1(n_666),
.B2(n_643),
.C(n_615),
.Y(n_792)
);

INVxp67_ASAP7_75t_L g793 ( 
.A(n_787),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_789),
.A2(n_785),
.B1(n_786),
.B2(n_788),
.Y(n_794)
);

INVxp67_ASAP7_75t_SL g795 ( 
.A(n_791),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_784),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_793),
.A2(n_615),
.B1(n_597),
.B2(n_666),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_796),
.A2(n_643),
.B1(n_623),
.B2(n_636),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_795),
.A2(n_643),
.B1(n_637),
.B2(n_626),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_L g800 ( 
.A1(n_794),
.A2(n_623),
.B1(n_637),
.B2(n_632),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_800),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_798),
.A2(n_792),
.B1(n_637),
.B2(n_629),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_799),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_801),
.A2(n_797),
.B(n_586),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_803),
.B(n_614),
.Y(n_805)
);

AO21x2_ASAP7_75t_L g806 ( 
.A1(n_805),
.A2(n_802),
.B(n_614),
.Y(n_806)
);

AOI21xp33_ASAP7_75t_L g807 ( 
.A1(n_806),
.A2(n_804),
.B(n_575),
.Y(n_807)
);


endmodule