module real_jpeg_7398_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g74 ( 
.A(n_0),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_1),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_1),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_1),
.B(n_187),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_1),
.B(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_1),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_1),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_1),
.B(n_384),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_2),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_2),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_2),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_2),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_2),
.B(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_2),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_2),
.B(n_459),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_3),
.B(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_3),
.B(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_3),
.B(n_106),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_3),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_3),
.B(n_145),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_3),
.B(n_176),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_4),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_5),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_5),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_5),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_5),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_5),
.B(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_5),
.B(n_347),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_5),
.B(n_388),
.Y(n_387)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_7),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_7),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_7),
.B(n_14),
.Y(n_294)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_8),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_8),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g229 ( 
.A(n_8),
.Y(n_229)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_8),
.Y(n_460)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_10),
.B(n_154),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_10),
.A2(n_229),
.B(n_230),
.Y(n_228)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_10),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_10),
.B(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_10),
.B(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_10),
.B(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_10),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_10),
.B(n_390),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_11),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_11),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_11),
.Y(n_154)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_11),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_12),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_12),
.B(n_82),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_12),
.B(n_114),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_12),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_12),
.B(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_12),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_12),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_12),
.B(n_405),
.Y(n_404)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_13),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_13),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_14),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_14),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_14),
.B(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_14),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_14),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_14),
.B(n_462),
.Y(n_461)
);

AND2x2_ASAP7_75t_SL g25 ( 
.A(n_15),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_15),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_15),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_15),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_15),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_15),
.B(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_15),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_441),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_195),
.B(n_439),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_162),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_20),
.B(n_162),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_96),
.C(n_126),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_21),
.B(n_96),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_62),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_44),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_23),
.B(n_44),
.C(n_62),
.Y(n_163)
);

MAJx2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_35),
.C(n_41),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_24),
.B(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.C(n_31),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_25),
.B(n_54),
.C(n_58),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_25),
.A2(n_58),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_25),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_25),
.A2(n_31),
.B1(n_92),
.B2(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_25),
.A2(n_92),
.B1(n_360),
.B2(n_365),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_25),
.B(n_365),
.Y(n_407)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_27),
.Y(n_358)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_27),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_28),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_28),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_28),
.A2(n_129),
.B1(n_191),
.B2(n_194),
.Y(n_190)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_30),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_30),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_31),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_31),
.B(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_31),
.A2(n_132),
.B1(n_254),
.B2(n_255),
.Y(n_326)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_33),
.Y(n_364)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g355 ( 
.A(n_34),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_35),
.A2(n_41),
.B1(n_52),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_35),
.Y(n_161)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_39),
.Y(n_251)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_40),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_46),
.B1(n_47),
.B2(n_52),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_53),
.B1(n_60),
.B2(n_61),
.Y(n_44)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_47),
.B(n_52),
.C(n_61),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_50),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_50),
.Y(n_316)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g193 ( 
.A(n_51),
.Y(n_193)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_54),
.A2(n_91),
.B1(n_94),
.B2(n_95),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_54),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_54),
.B(n_220),
.C(n_223),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_54),
.A2(n_94),
.B1(n_220),
.B2(n_284),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_56),
.Y(n_370)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_56),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_58),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_80),
.C(n_90),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_63),
.B(n_80),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_68),
.B2(n_69),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_71),
.C(n_75),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_64),
.A2(n_65),
.B1(n_120),
.B2(n_122),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_64),
.B(n_120),
.C(n_125),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_64),
.A2(n_65),
.B1(n_143),
.B2(n_144),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_65),
.B(n_144),
.Y(n_292)
);

INVx3_ASAP7_75t_SL g138 ( 
.A(n_66),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_67),
.Y(n_382)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_75),
.B2(n_79),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_74),
.Y(n_156)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_74),
.Y(n_344)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_74),
.Y(n_375)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_75),
.A2(n_79),
.B1(n_453),
.B2(n_454),
.Y(n_452)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.C(n_87),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_81),
.B(n_140),
.Y(n_139)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_84),
.B(n_87),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_86),
.Y(n_236)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_90),
.B(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_117),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_98),
.B(n_99),
.C(n_117),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_112),
.B2(n_113),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_105),
.B1(n_110),
.B2(n_111),
.Y(n_101)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_105),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_105),
.B(n_110),
.C(n_113),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_105),
.B(n_135),
.Y(n_204)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_109),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_109),
.Y(n_249)
);

INVx6_ASAP7_75t_L g321 ( 
.A(n_109),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_134),
.C(n_136),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_123),
.B2(n_125),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_120),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_123),
.A2(n_125),
.B1(n_175),
.B2(n_178),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_123),
.B(n_248),
.C(n_250),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_123),
.A2(n_125),
.B1(n_250),
.B2(n_310),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_125),
.B(n_170),
.C(n_175),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_126),
.B(n_275),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_141),
.C(n_159),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_127),
.B(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_133),
.C(n_139),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_128),
.B(n_242),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_129),
.B(n_186),
.C(n_191),
.Y(n_451)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_133),
.B(n_139),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_136),
.B(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_141),
.B(n_159),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_155),
.C(n_157),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_142),
.B(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_147),
.C(n_153),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_143),
.A2(n_144),
.B1(n_153),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_147),
.A2(n_259),
.B1(n_260),
.B2(n_261),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_147),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_147),
.A2(n_169),
.B1(n_170),
.B2(n_259),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_152),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_153),
.Y(n_262)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_154),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_155),
.A2(n_157),
.B1(n_158),
.B2(n_240),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_155),
.Y(n_240)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx24_ASAP7_75t_SL g467 ( 
.A(n_162),
.Y(n_467)
);

FAx1_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_164),
.CI(n_179),
.CON(n_162),
.SN(n_162)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_163),
.B(n_164),
.C(n_179),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_166),
.B(n_167),
.C(n_168),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_173),
.B2(n_174),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_206),
.C(n_211),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_169),
.A2(n_170),
.B1(n_206),
.B2(n_207),
.Y(n_246)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx11_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_175),
.Y(n_178)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_177),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_180),
.B(n_182),
.C(n_185),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_190),
.Y(n_185)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_189),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_189),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_191),
.Y(n_194)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

AOI221xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_332),
.B1(n_432),
.B2(n_437),
.C(n_438),
.Y(n_196)
);

NOR3xp33_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_272),
.C(n_276),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_198),
.A2(n_433),
.B(n_436),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_265),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g436 ( 
.A(n_199),
.B(n_265),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_241),
.C(n_243),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_200),
.B(n_241),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_226),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_201),
.B(n_227),
.C(n_238),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.C(n_218),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_203),
.B(n_219),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_205),
.B(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_210),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_211),
.B(n_246),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_220),
.Y(n_284)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_223),
.B(n_283),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_238),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_234),
.C(n_237),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_264),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_228),
.A2(n_230),
.B(n_286),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_237),
.Y(n_264)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_243),
.B(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_258),
.C(n_263),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_244),
.B(n_280),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.C(n_252),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_245),
.B(n_328),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_247),
.A2(n_252),
.B1(n_253),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_247),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_248),
.B(n_309),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_250),
.Y(n_310)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_263),
.Y(n_280)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_271),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_269),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_269),
.C(n_271),
.Y(n_273)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_272),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_273),
.B(n_274),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_303),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_277),
.A2(n_434),
.B(n_435),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_301),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_278),
.B(n_301),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_281),
.C(n_299),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_279),
.B(n_331),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_281),
.B(n_299),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_285),
.C(n_290),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_285),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_287),
.B(n_369),
.Y(n_368)
);

INVx8_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_293),
.C(n_295),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_291),
.A2(n_292),
.B1(n_420),
.B2(n_421),
.Y(n_419)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_293),
.A2(n_294),
.B1(n_295),
.B2(n_296),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx5_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_330),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_304),
.B(n_330),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_307),
.C(n_327),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_305),
.B(n_430),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_307),
.B(n_327),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_311),
.C(n_325),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_308),
.B(n_423),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_311),
.A2(n_325),
.B1(n_326),
.B2(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_311),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_317),
.C(n_322),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_312),
.A2(n_313),
.B1(n_322),
.B2(n_323),
.Y(n_411)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_317),
.B(n_411),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_318),
.B(n_354),
.Y(n_353)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx5_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_333),
.A2(n_427),
.B(n_431),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_413),
.B(n_426),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_400),
.B(n_412),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_376),
.B(n_399),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_337),
.B(n_366),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_337),
.B(n_366),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_351),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_338),
.B(n_352),
.C(n_359),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_345),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_339),
.B(n_346),
.C(n_348),
.Y(n_409)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_348),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_359),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_356),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_353),
.B(n_356),
.Y(n_367)
);

CKINVDCx14_ASAP7_75t_R g388 ( 
.A(n_354),
.Y(n_388)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_360),
.Y(n_365)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_368),
.C(n_371),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_367),
.B(n_396),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_368),
.A2(n_371),
.B1(n_372),
.B2(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_368),
.Y(n_397)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx5_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_377),
.A2(n_393),
.B(n_398),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_378),
.A2(n_386),
.B(n_392),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_379),
.B(n_385),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_379),
.B(n_385),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_383),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_380),
.B(n_383),
.Y(n_394)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_384),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_389),
.Y(n_386)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_395),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_394),
.B(n_395),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_402),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_401),
.B(n_402),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_408),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_403),
.B(n_409),
.C(n_410),
.Y(n_425)
);

BUFx24_ASAP7_75t_SL g466 ( 
.A(n_403),
.Y(n_466)
);

FAx1_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_406),
.CI(n_407),
.CON(n_403),
.SN(n_403)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_404),
.B(n_406),
.C(n_407),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_414),
.B(n_425),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_414),
.B(n_425),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_422),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_416),
.A2(n_417),
.B1(n_418),
.B2(n_419),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_416),
.B(n_419),
.C(n_422),
.Y(n_428)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_420),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_429),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_428),
.B(n_429),
.Y(n_431)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_465),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_445),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_444),
.B(n_445),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_447),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_449),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_455),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_452),
.Y(n_450)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_457),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_458),
.A2(n_461),
.B1(n_463),
.B2(n_464),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_458),
.Y(n_463)
);

INVx6_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_461),
.Y(n_464)
);


endmodule