module fake_jpeg_25539_n_308 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_308);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_308;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

CKINVDCx6p67_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_8),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_18),
.B(n_7),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_12),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_35),
.A2(n_32),
.B1(n_24),
.B2(n_26),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_55),
.B1(n_19),
.B2(n_32),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_49),
.Y(n_66)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_51),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_16),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_32),
.B1(n_24),
.B2(n_26),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_52),
.A2(n_41),
.B1(n_25),
.B2(n_28),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_53),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_32),
.B1(n_24),
.B2(n_19),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_59),
.Y(n_78)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_58),
.Y(n_69)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_62),
.Y(n_84)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_45),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_65),
.B(n_79),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_42),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_68),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_42),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_82),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_56),
.A2(n_39),
.B(n_25),
.C(n_28),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_71),
.A2(n_86),
.B(n_21),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_44),
.A2(n_41),
.B1(n_40),
.B2(n_19),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_73),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_47),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_56),
.B(n_39),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_76),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_17),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_64),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_54),
.B1(n_20),
.B2(n_28),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_17),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_63),
.A2(n_30),
.B1(n_31),
.B2(n_25),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_85),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_50),
.B(n_31),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_60),
.A2(n_62),
.B(n_52),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_57),
.A2(n_27),
.B1(n_17),
.B2(n_23),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_58),
.B1(n_54),
.B2(n_20),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_16),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_95),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_94),
.B1(n_109),
.B2(n_110),
.Y(n_118)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_30),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_107),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_97),
.A2(n_111),
.B1(n_22),
.B2(n_69),
.Y(n_139)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_102),
.Y(n_128)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_73),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_106),
.Y(n_141)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_31),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_112),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_70),
.A2(n_54),
.B1(n_20),
.B2(n_21),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_70),
.A2(n_86),
.B1(n_68),
.B2(n_77),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_87),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_113),
.Y(n_134)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_115),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_65),
.B(n_27),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_88),
.A2(n_21),
.B1(n_22),
.B2(n_30),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_116),
.A2(n_81),
.B1(n_66),
.B2(n_77),
.Y(n_120)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_87),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_120),
.A2(n_124),
.B1(n_137),
.B2(n_102),
.Y(n_147)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_121),
.B(n_130),
.Y(n_156)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_66),
.C(n_78),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_129),
.C(n_138),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_78),
.B1(n_80),
.B2(n_72),
.Y(n_124)
);

BUFx12_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_117),
.Y(n_155)
);

MAJx2_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_71),
.C(n_89),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_132),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_83),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_83),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_140),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_106),
.A2(n_80),
.B1(n_79),
.B2(n_72),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_121),
.B1(n_130),
.B2(n_140),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_93),
.A2(n_101),
.B1(n_104),
.B2(n_112),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_136),
.A2(n_139),
.B(n_22),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_93),
.A2(n_72),
.B1(n_69),
.B2(n_71),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_47),
.C(n_53),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_89),
.Y(n_142)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_53),
.C(n_23),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_23),
.C(n_33),
.Y(n_169)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_146),
.B(n_153),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_163),
.B1(n_167),
.B2(n_138),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_149),
.A2(n_33),
.B1(n_29),
.B2(n_9),
.Y(n_192)
);

OA22x2_ASAP7_75t_L g152 ( 
.A1(n_118),
.A2(n_111),
.B1(n_101),
.B2(n_109),
.Y(n_152)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_158),
.Y(n_186)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_134),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_161),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_141),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_165),
.Y(n_197)
);

AO22x2_ASAP7_75t_L g163 ( 
.A1(n_118),
.A2(n_120),
.B1(n_93),
.B2(n_133),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_123),
.B(n_107),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_168),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_99),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_137),
.A2(n_104),
.B(n_1),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_166),
.A2(n_172),
.B(n_132),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_124),
.A2(n_69),
.B1(n_96),
.B2(n_90),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_90),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_125),
.C(n_33),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_126),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_170),
.Y(n_200)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_126),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_174),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_119),
.A2(n_69),
.B1(n_27),
.B2(n_29),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_173),
.A2(n_27),
.B1(n_33),
.B2(n_29),
.Y(n_189)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_127),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_175),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_150),
.B(n_142),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_180),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_178),
.A2(n_166),
.B(n_172),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_179),
.A2(n_194),
.B1(n_163),
.B2(n_159),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_129),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_156),
.A2(n_136),
.B1(n_145),
.B2(n_131),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_181),
.A2(n_196),
.B1(n_13),
.B2(n_12),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_185),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_150),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_193),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_190),
.C(n_199),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_189),
.B(n_192),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_33),
.C(n_29),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_148),
.B(n_0),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_147),
.A2(n_33),
.B1(n_29),
.B2(n_9),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_195),
.B(n_0),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_163),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_157),
.B(n_29),
.C(n_7),
.Y(n_199)
);

AO21x1_ASAP7_75t_L g235 ( 
.A1(n_203),
.A2(n_202),
.B(n_200),
.Y(n_235)
);

AO22x1_ASAP7_75t_L g204 ( 
.A1(n_183),
.A2(n_163),
.B1(n_152),
.B2(n_148),
.Y(n_204)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_204),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_205),
.A2(n_206),
.B1(n_208),
.B2(n_212),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_187),
.A2(n_152),
.B1(n_159),
.B2(n_171),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_184),
.A2(n_152),
.B1(n_174),
.B2(n_154),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_198),
.Y(n_210)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_210),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_168),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_216),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_184),
.A2(n_151),
.B1(n_167),
.B2(n_169),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_178),
.A2(n_151),
.B(n_1),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_214),
.A2(n_176),
.B(n_201),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_179),
.A2(n_196),
.B1(n_185),
.B2(n_195),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_215),
.A2(n_221),
.B1(n_225),
.B2(n_214),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_164),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_219),
.Y(n_246)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_177),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_181),
.B(n_14),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_188),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_198),
.B(n_13),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_222),
.B(n_226),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_223),
.A2(n_197),
.B(n_202),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_180),
.A2(n_186),
.B1(n_194),
.B2(n_193),
.Y(n_225)
);

NAND3xp33_ASAP7_75t_L g226 ( 
.A(n_182),
.B(n_13),
.C(n_12),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_210),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_234),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_190),
.C(n_199),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_239),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_231),
.A2(n_232),
.B1(n_207),
.B2(n_225),
.Y(n_253)
);

XOR2x2_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_200),
.Y(n_232)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_233),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_203),
.Y(n_248)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_201),
.Y(n_236)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_238),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_189),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_11),
.C(n_10),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_210),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_242),
.B(n_244),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_215),
.Y(n_244)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_245),
.Y(n_256)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_248),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_234),
.A2(n_204),
.B1(n_218),
.B2(n_205),
.Y(n_249)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_253),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_235),
.B(n_228),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_254),
.B(n_246),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_232),
.A2(n_212),
.B1(n_206),
.B2(n_213),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_255),
.A2(n_260),
.B1(n_243),
.B2(n_251),
.Y(n_263)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_236),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_258),
.B(n_231),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_220),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_237),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_243),
.A2(n_224),
.B1(n_2),
.B2(n_3),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_257),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_265),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_261),
.B(n_239),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_230),
.C(n_229),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_271),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_270),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_229),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_247),
.B(n_244),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_227),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_272),
.B(n_273),
.Y(n_285)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_257),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_280),
.Y(n_286)
);

INVx6_ASAP7_75t_L g279 ( 
.A(n_267),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_279),
.B(n_1),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_262),
.A2(n_256),
.B(n_240),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_274),
.A2(n_260),
.B1(n_249),
.B2(n_248),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_282),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_259),
.Y(n_282)
);

OAI21x1_ASAP7_75t_SL g283 ( 
.A1(n_266),
.A2(n_255),
.B(n_241),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_283),
.A2(n_10),
.B(n_11),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_266),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_290),
.Y(n_298)
);

MAJx2_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_268),
.C(n_270),
.Y(n_289)
);

OAI21x1_ASAP7_75t_SL g300 ( 
.A1(n_289),
.A2(n_291),
.B(n_275),
.Y(n_300)
);

OAI21x1_ASAP7_75t_L g291 ( 
.A1(n_281),
.A2(n_11),
.B(n_2),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_293),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_4),
.C(n_5),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_278),
.B(n_4),
.Y(n_294)
);

A2O1A1Ixp33_ASAP7_75t_L g299 ( 
.A1(n_294),
.A2(n_5),
.B(n_6),
.C(n_282),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_286),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_297),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_288),
.A2(n_279),
.B1(n_285),
.B2(n_280),
.Y(n_297)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_299),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_300),
.A2(n_286),
.B(n_275),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_302),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_304),
.B(n_301),
.Y(n_305)
);

OAI321xp33_ASAP7_75t_L g306 ( 
.A1(n_305),
.A2(n_298),
.A3(n_296),
.B1(n_295),
.B2(n_303),
.C(n_6),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_306),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_6),
.B(n_304),
.Y(n_308)
);


endmodule