module fake_jpeg_1913_n_339 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_17),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_22),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_50),
.B(n_51),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_1),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_53),
.Y(n_132)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx11_ASAP7_75t_L g143 ( 
.A(n_54),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_23),
.B(n_1),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_56),
.B(n_72),
.Y(n_109)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_59),
.Y(n_142)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_26),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_61),
.B(n_63),
.Y(n_128)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_42),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_64),
.Y(n_152)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_68),
.Y(n_144)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_48),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_71),
.B(n_73),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_24),
.B(n_14),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

BUFx16f_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVxp67_ASAP7_75t_SL g115 ( 
.A(n_76),
.Y(n_115)
);

INVx3_ASAP7_75t_SL g77 ( 
.A(n_39),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

INVx2_ASAP7_75t_R g80 ( 
.A(n_20),
.Y(n_80)
);

NAND2xp33_ASAP7_75t_SL g145 ( 
.A(n_80),
.B(n_93),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_18),
.B(n_2),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_81),
.B(n_85),
.Y(n_130)
);

BUFx24_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_49),
.Y(n_83)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_18),
.A2(n_4),
.B(n_6),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_L g118 ( 
.A1(n_84),
.A2(n_95),
.B(n_9),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_4),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_7),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_86),
.B(n_96),
.Y(n_135)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_88),
.Y(n_151)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_21),
.Y(n_89)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_92),
.B(n_94),
.Y(n_140)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_24),
.Y(n_94)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_30),
.B(n_8),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_27),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_97),
.A2(n_45),
.B1(n_43),
.B2(n_41),
.Y(n_102)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_99),
.Y(n_137)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_83),
.A2(n_45),
.B1(n_43),
.B2(n_41),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_100),
.A2(n_105),
.B1(n_114),
.B2(n_111),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_102),
.A2(n_104),
.B1(n_119),
.B2(n_122),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_74),
.A2(n_27),
.B1(n_37),
.B2(n_29),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_76),
.A2(n_44),
.B1(n_37),
.B2(n_33),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_54),
.A2(n_69),
.B1(n_87),
.B2(n_60),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_118),
.B(n_141),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_75),
.A2(n_44),
.B1(n_33),
.B2(n_36),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_77),
.A2(n_68),
.B1(n_59),
.B2(n_55),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_L g125 ( 
.A1(n_88),
.A2(n_36),
.B1(n_38),
.B2(n_40),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_125),
.A2(n_131),
.B1(n_149),
.B2(n_40),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_90),
.A2(n_79),
.B1(n_70),
.B2(n_36),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_78),
.B(n_10),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_138),
.B(n_139),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_70),
.B(n_12),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_80),
.A2(n_53),
.B1(n_64),
.B2(n_38),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_82),
.B(n_36),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_147),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_95),
.A2(n_38),
.B1(n_40),
.B2(n_12),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_82),
.A2(n_38),
.B1(n_40),
.B2(n_51),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_142),
.Y(n_187)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_154),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_SL g199 ( 
.A1(n_155),
.A2(n_158),
.B(n_163),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_148),
.C(n_123),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_156),
.B(n_159),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_147),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_157),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_109),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_128),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_162),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_111),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_177),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_134),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_150),
.A2(n_125),
.B1(n_119),
.B2(n_146),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_164),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_101),
.A2(n_103),
.B1(n_117),
.B2(n_116),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_165),
.A2(n_187),
.B1(n_173),
.B2(n_157),
.Y(n_212)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_124),
.B(n_120),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_167),
.A2(n_171),
.B(n_175),
.Y(n_220)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_108),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_169),
.B(n_184),
.Y(n_208)
);

CKINVDCx12_ASAP7_75t_R g170 ( 
.A(n_115),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_170),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_136),
.A2(n_127),
.B1(n_110),
.B2(n_126),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_132),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_174),
.B(n_185),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_126),
.B(n_115),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_129),
.A2(n_152),
.B1(n_151),
.B2(n_143),
.Y(n_176)
);

INVx11_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_152),
.B(n_113),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_100),
.A2(n_105),
.B(n_114),
.Y(n_179)
);

NOR2x1_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_173),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_113),
.B(n_106),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_186),
.Y(n_202)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_107),
.Y(n_181)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_107),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_106),
.Y(n_183)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_183),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_112),
.B(n_121),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_112),
.B(n_121),
.Y(n_185)
);

BUFx16f_ASAP7_75t_L g186 ( 
.A(n_143),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_142),
.B(n_144),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_188),
.B(n_187),
.Y(n_201)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_137),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_192),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_147),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_137),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_194),
.Y(n_213)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_137),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_194),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_200),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_156),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_204),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_188),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_161),
.B(n_157),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_215),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_212),
.A2(n_199),
.B1(n_213),
.B2(n_200),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_178),
.B(n_190),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_214),
.B(n_167),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_190),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_216),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_218),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_228),
.Y(n_261)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_222),
.Y(n_225)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

AO32x1_ASAP7_75t_L g227 ( 
.A1(n_198),
.A2(n_179),
.A3(n_186),
.B1(n_175),
.B2(n_166),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_227),
.A2(n_248),
.B(n_220),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_218),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_208),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_212),
.A2(n_181),
.B1(n_182),
.B2(n_189),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_231),
.A2(n_240),
.B1(n_242),
.B2(n_244),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_218),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_238),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_233),
.B(n_236),
.Y(n_249)
);

O2A1O1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_216),
.A2(n_186),
.B(n_164),
.C(n_175),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_234),
.A2(n_227),
.B(n_230),
.Y(n_267)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_222),
.Y(n_235)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_235),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_208),
.B(n_167),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_202),
.Y(n_237)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_195),
.B(n_213),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_216),
.A2(n_183),
.B1(n_168),
.B2(n_154),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_201),
.B(n_204),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_246),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_196),
.B(n_206),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_243),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_215),
.A2(n_214),
.B1(n_198),
.B2(n_211),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_209),
.Y(n_245)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_245),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_217),
.B(n_205),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_209),
.Y(n_247)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_247),
.Y(n_268)
);

A2O1A1Ixp33_ASAP7_75t_SL g248 ( 
.A1(n_207),
.A2(n_202),
.B(n_220),
.C(n_210),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_205),
.C(n_203),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_264),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_257),
.A2(n_263),
.B(n_267),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_237),
.Y(n_259)
);

NOR3xp33_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_260),
.C(n_227),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_234),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_230),
.A2(n_203),
.B(n_207),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_226),
.B(n_219),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_224),
.B(n_219),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_224),
.Y(n_274)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_251),
.Y(n_270)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_271),
.Y(n_293)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_258),
.A2(n_242),
.B1(n_240),
.B2(n_231),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_273),
.A2(n_280),
.B1(n_282),
.B2(n_283),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_281),
.Y(n_292)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_253),
.Y(n_276)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_276),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_267),
.A2(n_248),
.B(n_239),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_278),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_239),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_259),
.A2(n_248),
.B1(n_244),
.B2(n_241),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_253),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_250),
.B(n_235),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_256),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_285),
.Y(n_287)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_256),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_257),
.A2(n_248),
.B(n_232),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_250),
.C(n_248),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_273),
.A2(n_258),
.B1(n_254),
.B2(n_260),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_289),
.A2(n_281),
.B1(n_274),
.B2(n_265),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_275),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_280),
.A2(n_265),
.B1(n_252),
.B2(n_262),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_297),
.A2(n_277),
.B1(n_283),
.B2(n_278),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_264),
.C(n_255),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_300),
.C(n_249),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_264),
.C(n_255),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_301),
.A2(n_309),
.B(n_297),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_302),
.A2(n_305),
.B1(n_308),
.B2(n_310),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_292),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_303),
.Y(n_317)
);

INVxp33_ASAP7_75t_L g319 ( 
.A(n_304),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_289),
.A2(n_292),
.B1(n_298),
.B2(n_288),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_311),
.C(n_287),
.Y(n_314)
);

INVx6_ASAP7_75t_L g307 ( 
.A(n_293),
.Y(n_307)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_307),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_294),
.A2(n_286),
.B1(n_275),
.B2(n_249),
.Y(n_308)
);

NAND3xp33_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_262),
.C(n_268),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_287),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_268),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_314),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_296),
.C(n_271),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_306),
.C(n_310),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_308),
.A2(n_261),
.B(n_291),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_302),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_323),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_305),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_321),
.B(n_322),
.Y(n_328)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_313),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_293),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_307),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_315),
.C(n_316),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_330),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_329),
.B(n_322),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_318),
.C(n_319),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_328),
.Y(n_331)
);

NOR2xp67_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_332),
.Y(n_334)
);

AOI322xp5_ASAP7_75t_L g335 ( 
.A1(n_333),
.A2(n_317),
.A3(n_328),
.B1(n_327),
.B2(n_295),
.C1(n_290),
.C2(n_261),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_335),
.A2(n_247),
.B1(n_245),
.B2(n_225),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_334),
.B(n_223),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_228),
.B1(n_197),
.B2(n_221),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_221),
.Y(n_339)
);


endmodule