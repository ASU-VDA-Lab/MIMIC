module real_aes_3345_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_908;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_941;
wire n_453;
wire n_374;
wire n_379;
wire n_932;
wire n_235;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_298;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_925;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_936;
wire n_610;
wire n_581;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_649;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_397;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_914;
wire n_203;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_662;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_922;
wire n_633;
wire n_926;
wire n_679;
wire n_149;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
NAND2xp5_ASAP7_75t_L g216 ( .A(n_0), .B(n_196), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_1), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_SL g268 ( .A1(n_2), .A2(n_139), .B(n_269), .C(n_270), .Y(n_268) );
OAI22xp33_ASAP7_75t_L g221 ( .A1(n_3), .A2(n_79), .B1(n_137), .B2(n_168), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_4), .A2(n_29), .B1(n_545), .B2(n_546), .Y(n_544) );
INVxp67_ASAP7_75t_L g113 ( .A(n_5), .Y(n_113) );
INVx1_ASAP7_75t_L g920 ( .A(n_5), .Y(n_920) );
INVx1_ASAP7_75t_L g924 ( .A(n_5), .Y(n_924) );
NAND3xp33_ASAP7_75t_SL g940 ( .A(n_5), .B(n_941), .C(n_942), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_6), .A2(n_87), .B1(n_598), .B2(n_599), .Y(n_597) );
CKINVDCx5p33_ASAP7_75t_R g247 ( .A(n_7), .Y(n_247) );
OAI22xp5_ASAP7_75t_L g165 ( .A1(n_8), .A2(n_65), .B1(n_166), .B2(n_168), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_9), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_10), .A2(n_30), .B1(n_567), .B2(n_568), .Y(n_566) );
INVx2_ASAP7_75t_L g692 ( .A(n_11), .Y(n_692) );
CKINVDCx5p33_ASAP7_75t_R g930 ( .A(n_12), .Y(n_930) );
AOI22xp5_ASAP7_75t_L g163 ( .A1(n_13), .A2(n_57), .B1(n_137), .B2(n_164), .Y(n_163) );
OA21x2_ASAP7_75t_L g153 ( .A1(n_14), .A2(n_64), .B(n_154), .Y(n_153) );
OA21x2_ASAP7_75t_L g158 ( .A1(n_14), .A2(n_64), .B(n_154), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_15), .B(n_634), .Y(n_633) );
INVx1_ASAP7_75t_SL g690 ( .A(n_16), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_17), .B(n_172), .Y(n_637) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_18), .Y(n_242) );
BUFx8_ASAP7_75t_SL g107 ( .A(n_19), .Y(n_107) );
BUFx3_ASAP7_75t_L g935 ( .A(n_19), .Y(n_935) );
O2A1O1Ixp33_ASAP7_75t_L g274 ( .A1(n_20), .A2(n_222), .B(n_275), .C(n_276), .Y(n_274) );
OAI22xp33_ASAP7_75t_SL g219 ( .A1(n_21), .A2(n_45), .B1(n_137), .B2(n_186), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g206 ( .A1(n_22), .A2(n_28), .B1(n_186), .B2(n_191), .Y(n_206) );
O2A1O1Ixp5_ASAP7_75t_L g641 ( .A1(n_23), .A2(n_548), .B(n_642), .C(n_645), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_24), .B(n_552), .Y(n_631) );
O2A1O1Ixp5_ASAP7_75t_L g132 ( .A1(n_25), .A2(n_133), .B(n_136), .C(n_139), .Y(n_132) );
INVx1_ASAP7_75t_L g118 ( .A(n_26), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_26), .B(n_76), .Y(n_939) );
INVx1_ASAP7_75t_SL g650 ( .A(n_27), .Y(n_650) );
AND2x2_ASAP7_75t_L g942 ( .A(n_31), .B(n_943), .Y(n_942) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_32), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_33), .B(n_212), .Y(n_211) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_34), .A2(n_38), .B1(n_551), .B2(n_553), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_35), .A2(n_63), .B1(n_553), .B2(n_586), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g630 ( .A(n_36), .B(n_547), .Y(n_630) );
INVx2_ASAP7_75t_L g579 ( .A(n_37), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_39), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_40), .B(n_259), .Y(n_604) );
OAI22xp33_ASAP7_75t_SL g121 ( .A1(n_41), .A2(n_92), .B1(n_122), .B2(n_123), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_41), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g684 ( .A(n_42), .Y(n_684) );
O2A1O1Ixp33_ASAP7_75t_L g687 ( .A1(n_43), .A2(n_222), .B(n_688), .C(n_689), .Y(n_687) );
INVx1_ASAP7_75t_L g671 ( .A(n_44), .Y(n_671) );
INVx2_ASAP7_75t_L g651 ( .A(n_46), .Y(n_651) );
INVx1_ASAP7_75t_L g154 ( .A(n_47), .Y(n_154) );
AND2x4_ASAP7_75t_L g149 ( .A(n_48), .B(n_150), .Y(n_149) );
AND2x4_ASAP7_75t_L g171 ( .A(n_48), .B(n_150), .Y(n_171) );
INVx2_ASAP7_75t_L g587 ( .A(n_49), .Y(n_587) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_50), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_51), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_52), .Y(n_146) );
INVx2_ASAP7_75t_L g192 ( .A(n_53), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g244 ( .A1(n_54), .A2(n_139), .B(n_245), .C(n_246), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_55), .Y(n_229) );
INVx1_ASAP7_75t_SL g646 ( .A(n_56), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g207 ( .A1(n_58), .A2(n_73), .B1(n_208), .B2(n_209), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_59), .B(n_172), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g590 ( .A(n_60), .Y(n_590) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_61), .Y(n_233) );
NAND2xp33_ASAP7_75t_R g173 ( .A(n_62), .B(n_158), .Y(n_173) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_62), .A2(n_102), .B1(n_212), .B2(n_395), .Y(n_394) );
O2A1O1Ixp33_ASAP7_75t_L g588 ( .A1(n_66), .A2(n_222), .B(n_545), .C(n_589), .Y(n_588) );
OR2x6_ASAP7_75t_L g115 ( .A(n_67), .B(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g941 ( .A(n_67), .Y(n_941) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_68), .Y(n_190) );
CKINVDCx16_ASAP7_75t_R g657 ( .A(n_69), .Y(n_657) );
INVx1_ASAP7_75t_L g667 ( .A(n_70), .Y(n_667) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_71), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_72), .B(n_567), .Y(n_635) );
NOR2xp67_ASAP7_75t_L g685 ( .A(n_74), .B(n_133), .Y(n_685) );
O2A1O1Ixp33_ASAP7_75t_L g582 ( .A1(n_75), .A2(n_139), .B(n_583), .C(n_585), .Y(n_582) );
O2A1O1Ixp33_ASAP7_75t_L g616 ( .A1(n_75), .A2(n_139), .B(n_583), .C(n_585), .Y(n_616) );
INVx1_ASAP7_75t_L g117 ( .A(n_76), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_77), .B(n_524), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_78), .A2(n_91), .B1(n_532), .B2(n_533), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_78), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_80), .A2(n_94), .B1(n_571), .B2(n_573), .Y(n_570) );
INVx1_ASAP7_75t_L g943 ( .A(n_81), .Y(n_943) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_82), .Y(n_135) );
BUFx5_ASAP7_75t_L g137 ( .A(n_82), .Y(n_137) );
INVx1_ASAP7_75t_L g167 ( .A(n_82), .Y(n_167) );
INVx2_ASAP7_75t_L g280 ( .A(n_83), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_84), .B(n_662), .Y(n_661) );
INVx2_ASAP7_75t_L g249 ( .A(n_85), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_86), .A2(n_104), .B1(n_936), .B2(n_944), .Y(n_103) );
AOI22xp5_ASAP7_75t_SL g528 ( .A1(n_88), .A2(n_529), .B1(n_530), .B2(n_531), .Y(n_528) );
CKINVDCx5p33_ASAP7_75t_R g529 ( .A(n_88), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_89), .Y(n_277) );
INVx2_ASAP7_75t_SL g150 ( .A(n_90), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_91), .Y(n_533) );
INVx1_ASAP7_75t_L g123 ( .A(n_92), .Y(n_123) );
INVx1_ASAP7_75t_L g144 ( .A(n_93), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_95), .B(n_158), .Y(n_668) );
INVx1_ASAP7_75t_SL g560 ( .A(n_96), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_97), .B(n_591), .Y(n_653) );
INVx2_ASAP7_75t_L g156 ( .A(n_98), .Y(n_156) );
AND2x2_ASAP7_75t_L g575 ( .A(n_99), .B(n_183), .Y(n_575) );
OAI21xp33_ASAP7_75t_SL g240 ( .A1(n_100), .A2(n_137), .B(n_241), .Y(n_240) );
OAI311xp33_ASAP7_75t_L g108 ( .A1(n_101), .A2(n_109), .A3(n_119), .B1(n_520), .C1(n_523), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g522 ( .A(n_101), .Y(n_522) );
INVxp67_ASAP7_75t_SL g194 ( .A(n_102), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_102), .B(n_212), .Y(n_303) );
OA21x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_108), .B(n_526), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_109), .B(n_522), .Y(n_521) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
BUFx12f_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx8_ASAP7_75t_L g525 ( .A(n_111), .Y(n_525) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
OR2x6_ASAP7_75t_L g919 ( .A(n_114), .B(n_920), .Y(n_919) );
INVx8_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g923 ( .A(n_115), .B(n_924), .Y(n_923) );
OR2x6_ASAP7_75t_L g931 ( .A(n_115), .B(n_924), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_119), .B(n_521), .Y(n_520) );
OA22x2_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_121), .B1(n_124), .B2(n_519), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g519 ( .A(n_124), .Y(n_519) );
NAND4xp75_ASAP7_75t_L g124 ( .A(n_125), .B(n_377), .C(n_448), .D(n_486), .Y(n_124) );
AND4x2_ASAP7_75t_L g921 ( .A(n_125), .B(n_377), .C(n_448), .D(n_486), .Y(n_921) );
NOR2x1_ASAP7_75t_L g125 ( .A(n_126), .B(n_315), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g126 ( .A(n_127), .B(n_295), .Y(n_126) );
O2A1O1Ixp33_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_174), .B(n_198), .C(n_250), .Y(n_127) );
AND2x2_ASAP7_75t_L g309 ( .A(n_128), .B(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_128), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g363 ( .A(n_128), .Y(n_363) );
AND2x2_ASAP7_75t_L g447 ( .A(n_128), .B(n_427), .Y(n_447) );
AND2x2_ASAP7_75t_L g454 ( .A(n_128), .B(n_252), .Y(n_454) );
AND2x4_ASAP7_75t_L g128 ( .A(n_129), .B(n_159), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_129), .B(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g511 ( .A(n_129), .B(n_411), .Y(n_511) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g282 ( .A(n_130), .B(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g289 ( .A(n_130), .Y(n_289) );
BUFx2_ASAP7_75t_R g349 ( .A(n_130), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_130), .B(n_266), .Y(n_419) );
AND2x2_ASAP7_75t_L g423 ( .A(n_130), .B(n_265), .Y(n_423) );
AO21x2_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_151), .B(n_155), .Y(n_130) );
NOR3xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_141), .C(n_148), .Y(n_131) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g142 ( .A(n_134), .Y(n_142) );
INVx1_ASAP7_75t_L g245 ( .A(n_134), .Y(n_245) );
INVx2_ASAP7_75t_L g547 ( .A(n_134), .Y(n_547) );
INVx2_ASAP7_75t_L g599 ( .A(n_134), .Y(n_599) );
INVx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g164 ( .A(n_135), .Y(n_164) );
INVx2_ASAP7_75t_L g168 ( .A(n_135), .Y(n_168) );
INVx6_ASAP7_75t_L g186 ( .A(n_135), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_137), .B(n_146), .Y(n_145) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_137), .A2(n_186), .B1(n_187), .B2(n_188), .Y(n_185) );
AOI22xp33_ASAP7_75t_SL g228 ( .A1(n_137), .A2(n_186), .B1(n_229), .B2(n_230), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g231 ( .A1(n_137), .A2(n_164), .B1(n_232), .B2(n_233), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_137), .B(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g552 ( .A(n_137), .Y(n_552) );
INVx2_ASAP7_75t_L g567 ( .A(n_137), .Y(n_567) );
INVx2_ASAP7_75t_L g573 ( .A(n_137), .Y(n_573) );
INVx1_ASAP7_75t_L g584 ( .A(n_137), .Y(n_584) );
INVx2_ASAP7_75t_L g598 ( .A(n_137), .Y(n_598) );
NAND2xp33_ASAP7_75t_L g683 ( .A(n_137), .B(n_684), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g162 ( .A1(n_139), .A2(n_147), .B1(n_163), .B2(n_165), .Y(n_162) );
OAI22xp33_ASAP7_75t_L g184 ( .A1(n_139), .A2(n_147), .B1(n_185), .B2(n_189), .Y(n_184) );
OAI221xp5_ASAP7_75t_L g227 ( .A1(n_139), .A2(n_171), .B1(n_222), .B2(n_228), .C(n_231), .Y(n_227) );
INVx1_ASAP7_75t_L g308 ( .A(n_139), .Y(n_308) );
INVx2_ASAP7_75t_SL g603 ( .A(n_139), .Y(n_603) );
INVx1_ASAP7_75t_L g636 ( .A(n_139), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_139), .B(n_667), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_139), .B(n_671), .Y(n_670) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_140), .B(n_144), .Y(n_143) );
INVx4_ASAP7_75t_L g147 ( .A(n_140), .Y(n_147) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_140), .Y(n_205) );
INVx1_ASAP7_75t_L g210 ( .A(n_140), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_140), .B(n_219), .Y(n_218) );
INVx3_ASAP7_75t_L g222 ( .A(n_140), .Y(n_222) );
INVxp67_ASAP7_75t_L g601 ( .A(n_140), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B1(n_145), .B2(n_147), .Y(n_141) );
INVx2_ASAP7_75t_L g243 ( .A(n_147), .Y(n_243) );
O2A1O1Ixp5_ASAP7_75t_SL g656 ( .A1(n_147), .A2(n_657), .B(n_658), .C(n_661), .Y(n_656) );
NOR2xp33_ASAP7_75t_SL g278 ( .A(n_148), .B(n_196), .Y(n_278) );
AOI221xp5_ASAP7_75t_L g305 ( .A1(n_148), .A2(n_243), .B1(n_306), .B2(n_307), .C(n_308), .Y(n_305) );
NOR4xp25_ASAP7_75t_L g581 ( .A(n_148), .B(n_582), .C(n_588), .D(n_591), .Y(n_581) );
NOR2x1_ASAP7_75t_SL g680 ( .A(n_148), .B(n_226), .Y(n_680) );
INVx4_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_149), .B(n_182), .Y(n_203) );
AND2x2_ASAP7_75t_L g237 ( .A(n_149), .B(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g304 ( .A(n_151), .B(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g627 ( .A(n_151), .Y(n_627) );
BUFx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx3_ASAP7_75t_L g172 ( .A(n_152), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_152), .B(n_249), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_152), .B(n_692), .Y(n_691) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx4_ASAP7_75t_L g197 ( .A(n_153), .Y(n_197) );
BUFx3_ASAP7_75t_L g259 ( .A(n_153), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx3_ASAP7_75t_L g183 ( .A(n_158), .Y(n_183) );
INVx1_ASAP7_75t_L g238 ( .A(n_158), .Y(n_238) );
INVx2_ASAP7_75t_L g396 ( .A(n_158), .Y(n_396) );
INVx1_ASAP7_75t_L g580 ( .A(n_158), .Y(n_580) );
INVx1_ASAP7_75t_SL g176 ( .A(n_159), .Y(n_176) );
INVx1_ASAP7_75t_L g290 ( .A(n_159), .Y(n_290) );
AND2x2_ASAP7_75t_L g372 ( .A(n_159), .B(n_265), .Y(n_372) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g283 ( .A(n_160), .Y(n_283) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_160), .Y(n_299) );
AND2x2_ASAP7_75t_L g420 ( .A(n_160), .B(n_179), .Y(n_420) );
AND2x2_ASAP7_75t_L g458 ( .A(n_160), .B(n_289), .Y(n_458) );
AND2x2_ASAP7_75t_L g160 ( .A(n_161), .B(n_173), .Y(n_160) );
AND2x2_ASAP7_75t_L g393 ( .A(n_161), .B(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_162), .B(n_169), .Y(n_161) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_164), .A2(n_190), .B1(n_191), .B2(n_192), .Y(n_189) );
INVx1_ASAP7_75t_L g275 ( .A(n_164), .Y(n_275) );
INVx2_ASAP7_75t_L g568 ( .A(n_164), .Y(n_568) );
INVxp67_ASAP7_75t_SL g688 ( .A(n_164), .Y(n_688) );
INVx2_ASAP7_75t_L g208 ( .A(n_166), .Y(n_208) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g191 ( .A(n_167), .Y(n_191) );
INVx2_ASAP7_75t_L g586 ( .A(n_168), .Y(n_586) );
INVx1_ASAP7_75t_L g662 ( .A(n_168), .Y(n_662) );
NOR2xp67_ASAP7_75t_L g169 ( .A(n_170), .B(n_172), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_170), .B(n_259), .Y(n_652) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_171), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_171), .B(n_197), .Y(n_223) );
INVx3_ASAP7_75t_L g558 ( .A(n_171), .Y(n_558) );
AND2x2_ASAP7_75t_L g574 ( .A(n_171), .B(n_258), .Y(n_574) );
INVxp67_ASAP7_75t_SL g174 ( .A(n_175), .Y(n_174) );
OR2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_177), .B(n_281), .Y(n_508) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x4_ASAP7_75t_L g374 ( .A(n_179), .B(n_266), .Y(n_374) );
OAI21x1_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_184), .B(n_193), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_181), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_181), .B(n_258), .Y(n_613) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g306 ( .A(n_185), .Y(n_306) );
INVx2_ASAP7_75t_SL g209 ( .A(n_186), .Y(n_209) );
INVx2_ASAP7_75t_L g271 ( .A(n_186), .Y(n_271) );
INVx1_ASAP7_75t_L g634 ( .A(n_186), .Y(n_634) );
INVx2_ASAP7_75t_L g644 ( .A(n_186), .Y(n_644) );
INVx1_ASAP7_75t_L g660 ( .A(n_186), .Y(n_660) );
INVx1_ASAP7_75t_L g307 ( .A(n_189), .Y(n_307) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_191), .B(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_191), .B(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g553 ( .A(n_191), .Y(n_553) );
INVx2_ASAP7_75t_L g572 ( .A(n_191), .Y(n_572) );
OR2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
INVx2_ASAP7_75t_L g226 ( .A(n_195), .Y(n_226) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx2_ASAP7_75t_L g212 ( .A(n_197), .Y(n_212) );
NOR2xp33_ASAP7_75t_SL g279 ( .A(n_197), .B(n_280), .Y(n_279) );
INVxp67_ASAP7_75t_SL g198 ( .A(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_200), .B(n_213), .Y(n_199) );
AND2x4_ASAP7_75t_L g292 ( .A(n_200), .B(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g376 ( .A(n_201), .B(n_345), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_201), .B(n_370), .Y(n_460) );
OR2x2_ASAP7_75t_L g493 ( .A(n_201), .B(n_410), .Y(n_493) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g329 ( .A(n_202), .Y(n_329) );
OAI21x1_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_211), .Y(n_202) );
INVx1_ASAP7_75t_L g257 ( .A(n_204), .Y(n_257) );
OA22x2_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B1(n_207), .B2(n_210), .Y(n_204) );
INVx4_ASAP7_75t_L g548 ( .A(n_205), .Y(n_548) );
INVx1_ASAP7_75t_L g269 ( .A(n_208), .Y(n_269) );
INVx3_ASAP7_75t_L g545 ( .A(n_208), .Y(n_545) );
INVx1_ASAP7_75t_L g260 ( .A(n_211), .Y(n_260) );
INVx2_ASAP7_75t_L g556 ( .A(n_212), .Y(n_556) );
BUFx2_ASAP7_75t_SL g357 ( .A(n_213), .Y(n_357) );
NOR2xp67_ASAP7_75t_L g213 ( .A(n_214), .B(n_224), .Y(n_213) );
INVx1_ASAP7_75t_L g312 ( .A(n_214), .Y(n_312) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g294 ( .A(n_215), .Y(n_294) );
INVx3_ASAP7_75t_L g331 ( .A(n_215), .Y(n_331) );
AND2x2_ASAP7_75t_L g366 ( .A(n_215), .B(n_332), .Y(n_366) );
AND2x2_ASAP7_75t_L g466 ( .A(n_215), .B(n_235), .Y(n_466) );
AND2x4_ASAP7_75t_L g215 ( .A(n_216), .B(n_217), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_218), .B(n_220), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_223), .Y(n_220) );
INVx3_ASAP7_75t_L g554 ( .A(n_222), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_235), .Y(n_224) );
INVx2_ASAP7_75t_L g261 ( .A(n_225), .Y(n_261) );
INVx2_ASAP7_75t_L g314 ( .A(n_225), .Y(n_314) );
OA21x2_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_234), .Y(n_225) );
OA21x2_ASAP7_75t_L g332 ( .A1(n_226), .A2(n_227), .B(n_234), .Y(n_332) );
INVx1_ASAP7_75t_L g253 ( .A(n_235), .Y(n_253) );
AND2x2_ASAP7_75t_L g313 ( .A(n_235), .B(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g339 ( .A(n_235), .B(n_294), .Y(n_339) );
INVx2_ASAP7_75t_L g345 ( .A(n_235), .Y(n_345) );
AND2x2_ASAP7_75t_L g370 ( .A(n_235), .B(n_331), .Y(n_370) );
BUFx2_ASAP7_75t_L g400 ( .A(n_235), .Y(n_400) );
INVx2_ASAP7_75t_L g411 ( .A(n_235), .Y(n_411) );
INVx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AOI21x1_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_239), .B(n_248), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_243), .B(n_244), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g629 ( .A1(n_243), .A2(n_630), .B(n_631), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_262), .B1(n_284), .B2(n_291), .Y(n_250) );
OR2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g351 ( .A(n_255), .B(n_344), .Y(n_351) );
INVx2_ASAP7_75t_SL g406 ( .A(n_255), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_255), .B(n_466), .Y(n_465) );
AND2x4_ASAP7_75t_L g255 ( .A(n_256), .B(n_261), .Y(n_255) );
OR2x2_ASAP7_75t_L g337 ( .A(n_256), .B(n_332), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_258), .B(n_260), .Y(n_256) );
INVx3_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x4_ASAP7_75t_L g293 ( .A(n_261), .B(n_294), .Y(n_293) );
NAND3xp33_ASAP7_75t_L g317 ( .A(n_262), .B(n_318), .C(n_322), .Y(n_317) );
OR2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_281), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g300 ( .A(n_264), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g310 ( .A(n_266), .B(n_302), .Y(n_310) );
INVx1_ASAP7_75t_L g321 ( .A(n_266), .Y(n_321) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_266), .Y(n_325) );
OR2x2_ASAP7_75t_L g354 ( .A(n_266), .B(n_302), .Y(n_354) );
INVx1_ASAP7_75t_L g428 ( .A(n_266), .Y(n_428) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_266), .Y(n_513) );
AO31x2_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_273), .A3(n_278), .B(n_279), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_271), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_275), .A2(n_649), .B1(n_650), .B2(n_651), .Y(n_648) );
OR2x2_ASAP7_75t_L g340 ( .A(n_281), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g352 ( .A(n_282), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g361 ( .A(n_282), .B(n_310), .Y(n_361) );
AND2x4_ASAP7_75t_L g467 ( .A(n_282), .B(n_374), .Y(n_467) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
BUFx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g403 ( .A(n_287), .B(n_325), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_288), .B(n_302), .Y(n_444) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g429 ( .A(n_289), .B(n_392), .Y(n_429) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_289), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_291), .B(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g436 ( .A(n_292), .B(n_387), .Y(n_436) );
NAND2x1p5_ASAP7_75t_L g399 ( .A(n_293), .B(n_400), .Y(n_399) );
NAND2x1p5_ASAP7_75t_L g446 ( .A(n_293), .B(n_441), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_293), .B(n_376), .Y(n_497) );
AND2x2_ASAP7_75t_L g359 ( .A(n_294), .B(n_329), .Y(n_359) );
OAI21xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_309), .B(n_311), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_300), .Y(n_297) );
AND2x2_ASAP7_75t_L g319 ( .A(n_298), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_298), .B(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_298), .B(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g470 ( .A(n_298), .B(n_471), .Y(n_470) );
INVx2_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g407 ( .A(n_300), .Y(n_407) );
INVx1_ASAP7_75t_L g517 ( .A(n_301), .Y(n_517) );
AND2x2_ASAP7_75t_L g320 ( .A(n_302), .B(n_321), .Y(n_320) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_302), .Y(n_476) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
AND2x2_ASAP7_75t_L g392 ( .A(n_304), .B(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_310), .B(n_349), .Y(n_348) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_310), .Y(n_414) );
AOI22xp5_ASAP7_75t_SL g462 ( .A1(n_311), .A2(n_463), .B1(n_464), .B2(n_467), .Y(n_462) );
AND2x4_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_350), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_326), .B(n_333), .Y(n_316) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g364 ( .A(n_320), .Y(n_364) );
OR2x2_ASAP7_75t_L g390 ( .A(n_321), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g502 ( .A(n_321), .B(n_420), .Y(n_502) );
INVxp67_ASAP7_75t_SL g463 ( .A(n_322), .Y(n_463) );
BUFx3_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVxp67_ASAP7_75t_L g341 ( .A(n_324), .Y(n_341) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_330), .Y(n_326) );
OR2x2_ASAP7_75t_L g433 ( .A(n_327), .B(n_339), .Y(n_433) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_327), .A2(n_466), .B(n_469), .C(n_472), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_327), .B(n_330), .Y(n_505) );
AND2x2_ASAP7_75t_L g518 ( .A(n_327), .B(n_366), .Y(n_518) );
INVx3_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x4_ASAP7_75t_L g386 ( .A(n_328), .B(n_330), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_328), .B(n_366), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_328), .B(n_370), .Y(n_489) );
AND2x2_ASAP7_75t_L g494 ( .A(n_328), .B(n_466), .Y(n_494) );
INVx3_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g453 ( .A(n_329), .Y(n_453) );
AND2x2_ASAP7_75t_L g500 ( .A(n_329), .B(n_332), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_330), .B(n_400), .Y(n_432) );
AND2x2_ASAP7_75t_L g477 ( .A(n_330), .B(n_376), .Y(n_477) );
AND2x4_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_331), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g452 ( .A(n_332), .B(n_453), .Y(n_452) );
OAI22xp5_ASAP7_75t_SL g333 ( .A1(n_334), .A2(n_340), .B1(n_342), .B2(n_346), .Y(n_333) );
INVx2_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
AND2x2_ASAP7_75t_L g343 ( .A(n_336), .B(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_336), .B(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g368 ( .A(n_337), .Y(n_368) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g387 ( .A(n_344), .Y(n_387) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g397 ( .A(n_345), .B(n_366), .Y(n_397) );
INVx1_ASAP7_75t_L g442 ( .A(n_345), .Y(n_442) );
AND2x2_ASAP7_75t_L g480 ( .A(n_345), .B(n_359), .Y(n_480) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_347), .A2(n_447), .B1(n_492), .B2(n_494), .Y(n_491) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g382 ( .A(n_349), .Y(n_382) );
AOI211xp5_ASAP7_75t_SL g350 ( .A1(n_351), .A2(n_352), .B(n_355), .C(n_362), .Y(n_350) );
NOR2x1_ASAP7_75t_L g490 ( .A(n_352), .B(n_417), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_353), .B(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AOI21xp33_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_358), .B(n_360), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OAI332xp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .A3(n_365), .B1(n_367), .B2(n_369), .B3(n_371), .C1(n_373), .C2(n_375), .Y(n_362) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_366), .A2(n_417), .B1(n_421), .B2(n_422), .Y(n_416) );
INVxp67_ASAP7_75t_SL g421 ( .A(n_367), .Y(n_421) );
INVx2_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
INVx2_ASAP7_75t_SL g515 ( .A(n_369), .Y(n_515) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g443 ( .A(n_372), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g516 ( .A(n_372), .B(n_517), .Y(n_516) );
INVx2_ASAP7_75t_SL g471 ( .A(n_374), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_374), .B(n_458), .Y(n_472) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NOR2x1_ASAP7_75t_L g377 ( .A(n_378), .B(n_415), .Y(n_377) );
OAI211xp5_ASAP7_75t_SL g378 ( .A1(n_379), .A2(n_383), .B(n_388), .C(n_404), .Y(n_378) );
INVxp67_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
OR2x2_ASAP7_75t_L g498 ( .A(n_387), .B(n_499), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_397), .B1(n_398), .B2(n_401), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_390), .B(n_505), .Y(n_504) );
OR2x2_ASAP7_75t_L g512 ( .A(n_391), .B(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g435 ( .A(n_392), .Y(n_435) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_396), .B(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g591 ( .A(n_396), .Y(n_591) );
INVx1_ASAP7_75t_L g481 ( .A(n_397), .Y(n_481) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AOI32xp33_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_407), .A3(n_408), .B1(n_409), .B2(n_412), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OAI321xp33_ASAP7_75t_L g506 ( .A1(n_408), .A2(n_421), .A3(n_451), .B1(n_507), .B2(n_509), .C(n_514), .Y(n_506) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND3xp33_ASAP7_75t_SL g415 ( .A(n_416), .B(n_424), .C(n_437), .Y(n_415) );
AND2x4_ASAP7_75t_L g417 ( .A(n_418), .B(n_420), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g422 ( .A(n_420), .B(n_423), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_420), .A2(n_515), .B1(n_516), .B2(n_518), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_430), .B1(n_434), .B2(n_436), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NAND2x1p5_ASAP7_75t_SL g426 ( .A(n_427), .B(n_429), .Y(n_426) );
INVx2_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g461 ( .A(n_428), .Y(n_461) );
NAND3xp33_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .C(n_433), .Y(n_430) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_433), .A2(n_488), .B(n_490), .C(n_491), .Y(n_487) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_443), .B1(n_445), .B2(n_447), .Y(n_437) );
BUFx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AND4x1_ASAP7_75t_L g448 ( .A(n_449), .B(n_462), .C(n_468), .D(n_473), .Y(n_448) );
A2O1A1Ixp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_454), .B(n_455), .C(n_461), .Y(n_449) );
INVxp67_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
INVx3_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVxp67_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_459), .Y(n_456) );
BUFx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_471), .A2(n_479), .B(n_481), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_477), .B(n_478), .C(n_482), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVxp67_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVxp67_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
NOR3xp33_ASAP7_75t_L g486 ( .A(n_487), .B(n_495), .C(n_506), .Y(n_486) );
BUFx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_498), .B(n_501), .C(n_503), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVxp67_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NOR2x1_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
NAND3xp33_ASAP7_75t_L g526 ( .A(n_523), .B(n_527), .C(n_932), .Y(n_526) );
INVxp67_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OA21x2_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_534), .B(n_925), .Y(n_527) );
AOI21x1_ASAP7_75t_L g925 ( .A1(n_528), .A2(n_926), .B(n_929), .Y(n_925) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AOI22x1_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_914), .B1(n_921), .B2(n_922), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g927 ( .A(n_536), .Y(n_927) );
OR2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_804), .Y(n_536) );
NAND4xp25_ASAP7_75t_L g537 ( .A(n_538), .B(n_730), .C(n_764), .D(n_773), .Y(n_537) );
O2A1O1Ixp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_605), .B(n_621), .C(n_673), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_561), .Y(n_539) );
INVxp67_ASAP7_75t_L g738 ( .A(n_540), .Y(n_738) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g607 ( .A(n_541), .B(n_608), .Y(n_607) );
NAND2x1_ASAP7_75t_L g753 ( .A(n_541), .B(n_620), .Y(n_753) );
NOR2x1_ASAP7_75t_L g762 ( .A(n_541), .B(n_612), .Y(n_762) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g701 ( .A(n_542), .Y(n_701) );
AOI21x1_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_549), .B(n_559), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_548), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_545), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_548), .B(n_570), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_554), .B(n_555), .Y(n_549) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_554), .B(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
AOI21x1_ASAP7_75t_L g608 ( .A1(n_556), .A2(n_609), .B(n_610), .Y(n_608) );
OAI21x1_ASAP7_75t_L g628 ( .A1(n_557), .A2(n_629), .B(n_632), .Y(n_628) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
OAI21x1_ASAP7_75t_L g672 ( .A1(n_558), .A2(n_627), .B(n_668), .Y(n_672) );
AOI21xp33_ASAP7_75t_L g807 ( .A1(n_561), .A2(n_749), .B(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g811 ( .A(n_561), .Y(n_811) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_576), .Y(n_561) );
INVx1_ASAP7_75t_L g721 ( .A(n_562), .Y(n_721) );
AND2x6_ASAP7_75t_SL g736 ( .A(n_562), .B(n_607), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_562), .B(n_741), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_562), .B(n_762), .Y(n_761) );
BUFx3_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_563), .B(n_593), .Y(n_696) );
AND2x2_ASAP7_75t_L g841 ( .A(n_563), .B(n_577), .Y(n_841) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx2_ASAP7_75t_SL g620 ( .A(n_564), .Y(n_620) );
AO31x2_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_569), .A3(n_574), .B(n_575), .Y(n_564) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g665 ( .A(n_573), .Y(n_665) );
INVx1_ASAP7_75t_L g856 ( .A(n_576), .Y(n_856) );
NOR2x1_ASAP7_75t_L g576 ( .A(n_577), .B(n_592), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_577), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g741 ( .A(n_577), .Y(n_741) );
AND2x4_ASAP7_75t_L g767 ( .A(n_577), .B(n_619), .Y(n_767) );
INVx1_ASAP7_75t_L g777 ( .A(n_577), .Y(n_777) );
OR2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_581), .Y(n_577) );
INVxp67_ASAP7_75t_SL g618 ( .A(n_578), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
INVx1_ASAP7_75t_L g594 ( .A(n_580), .Y(n_594) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_586), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g649 ( .A(n_586), .Y(n_649) );
INVxp67_ASAP7_75t_SL g617 ( .A(n_588), .Y(n_617) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g720 ( .A(n_593), .B(n_707), .Y(n_720) );
BUFx6f_ASAP7_75t_L g729 ( .A(n_593), .Y(n_729) );
INVx1_ASAP7_75t_L g896 ( .A(n_593), .Y(n_896) );
OA21x2_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_595), .B(n_604), .Y(n_593) );
OAI21x1_ASAP7_75t_L g718 ( .A1(n_594), .A2(n_628), .B(n_637), .Y(n_718) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_596), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_600), .B1(n_602), .B2(n_603), .Y(n_596) );
OAI21xp5_ASAP7_75t_SL g647 ( .A1(n_600), .A2(n_648), .B(n_652), .Y(n_647) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g610 ( .A(n_604), .Y(n_610) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_611), .Y(n_606) );
AND2x2_ASAP7_75t_L g827 ( .A(n_607), .B(n_746), .Y(n_827) );
HB1xp67_ASAP7_75t_L g835 ( .A(n_607), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_607), .B(n_890), .Y(n_889) );
OR2x2_ASAP7_75t_L g706 ( .A(n_608), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g798 ( .A(n_608), .Y(n_798) );
AND2x2_ASAP7_75t_L g727 ( .A(n_611), .B(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g750 ( .A(n_611), .B(n_738), .Y(n_750) );
AND2x4_ASAP7_75t_L g913 ( .A(n_611), .B(n_766), .Y(n_913) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_619), .Y(n_611) );
AND2x4_ASAP7_75t_L g747 ( .A(n_612), .B(n_707), .Y(n_747) );
INVxp67_ASAP7_75t_SL g893 ( .A(n_612), .Y(n_893) );
OA21x2_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_614), .B(n_618), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_617), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g705 ( .A(n_619), .Y(n_705) );
BUFx2_ASAP7_75t_SL g746 ( .A(n_619), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_619), .B(n_798), .Y(n_878) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g764 ( .A1(n_621), .A2(n_747), .B1(n_765), .B2(n_768), .C(n_771), .Y(n_764) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND2x1p5_ASAP7_75t_L g622 ( .A(n_623), .B(n_638), .Y(n_622) );
INVx2_ASAP7_75t_L g770 ( .A(n_623), .Y(n_770) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g783 ( .A(n_624), .B(n_716), .Y(n_783) );
HB1xp67_ASAP7_75t_L g800 ( .A(n_624), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_624), .B(n_654), .Y(n_825) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g744 ( .A(n_625), .B(n_655), .Y(n_744) );
AND2x2_ASAP7_75t_L g787 ( .A(n_625), .B(n_639), .Y(n_787) );
AND2x2_ASAP7_75t_L g862 ( .A(n_625), .B(n_726), .Y(n_862) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OAI21x1_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_628), .B(n_637), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_635), .B(n_636), .Y(n_632) );
OAI21xp5_ASAP7_75t_L g681 ( .A1(n_636), .A2(n_682), .B(n_685), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_638), .B(n_800), .Y(n_799) );
AND2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_654), .Y(n_638) );
INVx2_ASAP7_75t_SL g711 ( .A(n_639), .Y(n_711) );
BUFx2_ASAP7_75t_L g890 ( .A(n_639), .Y(n_890) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g677 ( .A(n_640), .Y(n_677) );
INVx3_ASAP7_75t_L g719 ( .A(n_640), .Y(n_719) );
OA21x2_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_647), .B(n_653), .Y(n_640) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x4_ASAP7_75t_L g678 ( .A(n_654), .B(n_679), .Y(n_678) );
OR2x2_ASAP7_75t_L g848 ( .A(n_654), .B(n_679), .Y(n_848) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g734 ( .A(n_655), .B(n_718), .Y(n_734) );
OAI21x1_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_663), .B(n_672), .Y(n_655) );
OAI21xp5_ASAP7_75t_L g713 ( .A1(n_656), .A2(n_663), .B(n_672), .Y(n_713) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_659), .B(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND3x1_ASAP7_75t_L g663 ( .A(n_664), .B(n_668), .C(n_669), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
OAI211xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_693), .B(n_702), .C(n_714), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .Y(n_675) );
AND2x2_ASAP7_75t_L g823 ( .A(n_676), .B(n_824), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_676), .B(n_843), .Y(n_842) );
OR2x2_ASAP7_75t_L g847 ( .A(n_676), .B(n_848), .Y(n_847) );
INVx2_ASAP7_75t_R g676 ( .A(n_677), .Y(n_676) );
BUFx2_ASAP7_75t_L g792 ( .A(n_677), .Y(n_792) );
INVx2_ASAP7_75t_L g763 ( .A(n_678), .Y(n_763) );
AND2x2_ASAP7_75t_L g769 ( .A(n_678), .B(n_770), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_678), .B(n_792), .Y(n_791) );
OAI322xp33_ASAP7_75t_L g819 ( .A1(n_678), .A2(n_749), .A3(n_820), .B1(n_822), .B2(n_826), .C1(n_828), .C2(n_834), .Y(n_819) );
AND2x2_ASAP7_75t_L g907 ( .A(n_678), .B(n_862), .Y(n_907) );
OR2x2_ASAP7_75t_L g712 ( .A(n_679), .B(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g716 ( .A(n_679), .Y(n_716) );
INVx1_ASAP7_75t_L g724 ( .A(n_679), .Y(n_724) );
AND2x2_ASAP7_75t_L g898 ( .A(n_679), .B(n_713), .Y(n_898) );
HB1xp67_ASAP7_75t_L g910 ( .A(n_679), .Y(n_910) );
AO31x2_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_681), .A3(n_686), .B(n_691), .Y(n_679) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_697), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g797 ( .A(n_700), .B(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g803 ( .A(n_700), .Y(n_803) );
HB1xp67_ASAP7_75t_L g902 ( .A(n_700), .Y(n_902) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g707 ( .A(n_701), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_703), .B(n_708), .Y(n_702) );
NOR3xp33_ASAP7_75t_L g735 ( .A(n_703), .B(n_736), .C(n_737), .Y(n_735) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
OR2x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
AND2x2_ASAP7_75t_L g796 ( .A(n_705), .B(n_797), .Y(n_796) );
INVx2_ASAP7_75t_L g866 ( .A(n_705), .Y(n_866) );
INVx2_ASAP7_75t_L g766 ( .A(n_706), .Y(n_766) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OR2x2_ASAP7_75t_L g709 ( .A(n_710), .B(n_712), .Y(n_709) );
AND2x2_ASAP7_75t_L g912 ( .A(n_710), .B(n_744), .Y(n_912) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g743 ( .A(n_711), .B(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_L g768 ( .A(n_711), .B(n_769), .Y(n_768) );
OR2x2_ASAP7_75t_L g818 ( .A(n_711), .B(n_712), .Y(n_818) );
NOR3xp33_ASAP7_75t_L g892 ( .A(n_711), .B(n_866), .C(n_893), .Y(n_892) );
OAI21xp5_ASAP7_75t_L g806 ( .A1(n_712), .A2(n_807), .B(n_809), .Y(n_806) );
OAI31xp33_ASAP7_75t_L g810 ( .A1(n_712), .A2(n_811), .A3(n_812), .B(n_813), .Y(n_810) );
AOI32xp33_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_720), .A3(n_721), .B1(n_722), .B2(n_727), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
AND2x2_ASAP7_75t_L g780 ( .A(n_716), .B(n_726), .Y(n_780) );
INVx1_ASAP7_75t_L g832 ( .A(n_716), .Y(n_832) );
INVx1_ASAP7_75t_L g844 ( .A(n_716), .Y(n_844) );
AND2x2_ASAP7_75t_L g857 ( .A(n_716), .B(n_744), .Y(n_857) );
INVx1_ASAP7_75t_L g861 ( .A(n_716), .Y(n_861) );
OR2x2_ASAP7_75t_L g864 ( .A(n_716), .B(n_830), .Y(n_864) );
INVx1_ASAP7_75t_L g754 ( .A(n_717), .Y(n_754) );
INVx1_ASAP7_75t_L g885 ( .A(n_717), .Y(n_885) );
AND2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
AND2x2_ASAP7_75t_L g725 ( .A(n_718), .B(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_719), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_719), .B(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g789 ( .A(n_720), .Y(n_789) );
AND2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_725), .Y(n_722) );
INVx2_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
AND2x4_ASAP7_75t_L g733 ( .A(n_724), .B(n_734), .Y(n_733) );
OR2x2_ASAP7_75t_L g884 ( .A(n_724), .B(n_885), .Y(n_884) );
INVx1_ASAP7_75t_L g749 ( .A(n_725), .Y(n_749) );
HB1xp67_ASAP7_75t_L g812 ( .A(n_725), .Y(n_812) );
AND2x2_ASAP7_75t_L g782 ( .A(n_726), .B(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g793 ( .A(n_727), .Y(n_793) );
INVx1_ASAP7_75t_L g840 ( .A(n_728), .Y(n_840) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g759 ( .A(n_729), .Y(n_759) );
NOR2x1p5_ASAP7_75t_L g816 ( .A(n_729), .B(n_753), .Y(n_816) );
NAND2x1p5_ASAP7_75t_L g868 ( .A(n_729), .B(n_747), .Y(n_868) );
NOR2xp33_ASAP7_75t_SL g730 ( .A(n_731), .B(n_751), .Y(n_730) );
OAI21xp33_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_735), .B(n_742), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_733), .B(n_745), .Y(n_772) );
AND2x2_ASAP7_75t_L g779 ( .A(n_734), .B(n_780), .Y(n_779) );
AND2x4_ASAP7_75t_L g843 ( .A(n_734), .B(n_844), .Y(n_843) );
NAND2xp5_ASAP7_75t_SL g863 ( .A(n_734), .B(n_792), .Y(n_863) );
INVx1_ASAP7_75t_L g813 ( .A(n_736), .Y(n_813) );
AND2x2_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
NOR2xp33_ASAP7_75t_SL g894 ( .A(n_738), .B(n_895), .Y(n_894) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g833 ( .A(n_740), .B(n_830), .Y(n_833) );
INVx1_ASAP7_75t_L g815 ( .A(n_741), .Y(n_815) );
AND2x2_ASAP7_75t_L g821 ( .A(n_741), .B(n_803), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_745), .B1(n_748), .B2(n_750), .Y(n_742) );
OAI21xp5_ASAP7_75t_SL g781 ( .A1(n_743), .A2(n_782), .B(n_784), .Y(n_781) );
INVx2_ASAP7_75t_L g830 ( .A(n_744), .Y(n_830) );
AND2x4_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
O2A1O1Ixp33_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_754), .B(n_755), .C(n_763), .Y(n_751) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
OR2x2_ASAP7_75t_L g855 ( .A(n_753), .B(n_856), .Y(n_855) );
INVx2_ASAP7_75t_L g853 ( .A(n_754), .Y(n_853) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
AND2x4_ASAP7_75t_L g756 ( .A(n_757), .B(n_760), .Y(n_756) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_757), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_757), .B(n_821), .Y(n_820) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g851 ( .A(n_761), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_762), .A2(n_853), .B1(n_854), .B2(n_857), .Y(n_852) );
AND2x2_ASAP7_75t_L g876 ( .A(n_762), .B(n_877), .Y(n_876) );
AND2x4_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_767), .Y(n_784) );
INVx2_ASAP7_75t_SL g790 ( .A(n_767), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_767), .B(n_803), .Y(n_802) );
AND2x2_ASAP7_75t_L g901 ( .A(n_767), .B(n_902), .Y(n_901) );
INVx2_ASAP7_75t_L g809 ( .A(n_769), .Y(n_809) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
AOI211xp5_ASAP7_75t_SL g773 ( .A1(n_774), .A2(n_775), .B(n_785), .C(n_794), .Y(n_773) );
OAI21xp5_ASAP7_75t_SL g775 ( .A1(n_776), .A2(n_778), .B(n_781), .Y(n_775) );
INVxp67_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx2_ASAP7_75t_L g801 ( .A(n_780), .Y(n_801) );
OAI21xp5_ASAP7_75t_L g911 ( .A1(n_783), .A2(n_912), .B(n_913), .Y(n_911) );
OAI22xp33_ASAP7_75t_SL g785 ( .A1(n_786), .A2(n_788), .B1(n_791), .B2(n_793), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
BUFx2_ASAP7_75t_L g808 ( .A(n_787), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_787), .B(n_904), .Y(n_903) );
NAND2x1_ASAP7_75t_SL g909 ( .A(n_787), .B(n_910), .Y(n_909) );
OR2x2_ASAP7_75t_L g788 ( .A(n_789), .B(n_790), .Y(n_788) );
OAI22xp33_ASAP7_75t_L g794 ( .A1(n_795), .A2(n_799), .B1(n_801), .B2(n_802), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g871 ( .A(n_797), .Y(n_871) );
NOR2x1_ASAP7_75t_L g849 ( .A(n_801), .B(n_850), .Y(n_849) );
NAND3xp33_ASAP7_75t_L g804 ( .A(n_805), .B(n_836), .C(n_879), .Y(n_804) );
AOI221xp5_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_810), .B1(n_814), .B2(n_817), .C(n_819), .Y(n_805) );
OAI221xp5_ASAP7_75t_L g869 ( .A1(n_809), .A2(n_870), .B1(n_872), .B2(n_873), .C(n_874), .Y(n_869) );
INVx1_ASAP7_75t_L g881 ( .A(n_814), .Y(n_881) );
AND2x2_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .Y(n_814) );
HB1xp67_ASAP7_75t_L g906 ( .A(n_816), .Y(n_906) );
INVxp67_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g873 ( .A(n_821), .Y(n_873) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g850 ( .A(n_824), .Y(n_850) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
AOI22xp5_ASAP7_75t_L g905 ( .A1(n_827), .A2(n_906), .B1(n_907), .B2(n_908), .Y(n_905) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_829), .B(n_833), .Y(n_828) );
INVx2_ASAP7_75t_SL g872 ( .A(n_829), .Y(n_872) );
NOR2x1_ASAP7_75t_L g829 ( .A(n_830), .B(n_831), .Y(n_829) );
INVx1_ASAP7_75t_L g875 ( .A(n_830), .Y(n_875) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
NOR3xp33_ASAP7_75t_L g836 ( .A(n_837), .B(n_858), .C(n_869), .Y(n_836) );
OAI211xp5_ASAP7_75t_SL g837 ( .A1(n_838), .A2(n_842), .B(n_845), .C(n_852), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
AND2x2_ASAP7_75t_L g839 ( .A(n_840), .B(n_841), .Y(n_839) );
INVx1_ASAP7_75t_L g904 ( .A(n_844), .Y(n_904) );
OAI21xp5_ASAP7_75t_L g845 ( .A1(n_846), .A2(n_849), .B(n_851), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx2_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
AOI31xp33_ASAP7_75t_L g858 ( .A1(n_859), .A2(n_863), .A3(n_864), .B(n_865), .Y(n_858) );
NAND2xp5_ASAP7_75t_SL g883 ( .A(n_859), .B(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
AND2x2_ASAP7_75t_L g860 ( .A(n_861), .B(n_862), .Y(n_860) );
NAND2x1p5_ASAP7_75t_L g865 ( .A(n_866), .B(n_867), .Y(n_865) );
HB1xp67_ASAP7_75t_L g888 ( .A(n_866), .Y(n_888) );
INVx2_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
HB1xp67_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_875), .B(n_876), .Y(n_874) );
INVx1_ASAP7_75t_L g882 ( .A(n_876), .Y(n_882) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
AOI211xp5_ASAP7_75t_SL g879 ( .A1(n_880), .A2(n_883), .B(n_886), .C(n_899), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_881), .B(n_882), .Y(n_880) );
O2A1O1Ixp33_ASAP7_75t_SL g886 ( .A1(n_887), .A2(n_889), .B(n_891), .C(n_897), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_892), .B(n_894), .Y(n_891) );
INVx1_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
INVx2_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
OAI211xp5_ASAP7_75t_L g899 ( .A1(n_900), .A2(n_903), .B(n_905), .C(n_911), .Y(n_899) );
INVx2_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
INVx1_ASAP7_75t_SL g908 ( .A(n_909), .Y(n_908) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
BUFx3_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
OAI22x1_ASAP7_75t_L g926 ( .A1(n_916), .A2(n_921), .B1(n_927), .B2(n_928), .Y(n_926) );
BUFx12f_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
CKINVDCx11_ASAP7_75t_R g917 ( .A(n_918), .Y(n_917) );
INVx2_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
CKINVDCx20_ASAP7_75t_R g928 ( .A(n_922), .Y(n_928) );
BUFx8_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
NOR2xp33_ASAP7_75t_L g929 ( .A(n_930), .B(n_931), .Y(n_929) );
BUFx4_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
CKINVDCx6p67_ASAP7_75t_R g934 ( .A(n_935), .Y(n_934) );
BUFx4_ASAP7_75t_SL g936 ( .A(n_937), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
BUFx4_ASAP7_75t_SL g944 ( .A(n_938), .Y(n_944) );
OR2x2_ASAP7_75t_L g938 ( .A(n_939), .B(n_940), .Y(n_938) );
endmodule