module fake_netlist_5_547_n_16249 (n_924, n_1263, n_3304, n_977, n_1378, n_2253, n_2417, n_611, n_2756, n_3912, n_1126, n_1423, n_1729, n_2739, n_1166, n_2380, n_1751, n_469, n_1508, n_82, n_2771, n_785, n_3241, n_549, n_2617, n_2200, n_3261, n_3006, n_532, n_1161, n_3795, n_3863, n_3027, n_1859, n_2746, n_1677, n_1150, n_2327, n_3179, n_3127, n_226, n_1780, n_3256, n_3732, n_1488, n_667, n_2899, n_2955, n_790, n_3619, n_1055, n_3541, n_3622, n_2386, n_3596, n_1501, n_111, n_2395, n_3906, n_880, n_3086, n_3297, n_544, n_1007, n_2369, n_155, n_2927, n_552, n_1528, n_2683, n_1370, n_1292, n_2347, n_2520, n_2821, n_1198, n_1360, n_2388, n_1099, n_2568, n_3641, n_956, n_564, n_423, n_1738, n_2021, n_3728, n_21, n_2134, n_3064, n_2391, n_105, n_3088, n_1021, n_1960, n_2843, n_2185, n_4, n_3270, n_551, n_2143, n_3713, n_2853, n_3615, n_2059, n_1323, n_3663, n_1466, n_688, n_1695, n_2487, n_3766, n_1353, n_800, n_3595, n_3246, n_3202, n_1347, n_2495, n_2880, n_1535, n_3813, n_1789, n_1666, n_3350, n_2389, n_671, n_819, n_1451, n_1022, n_4038, n_2302, n_915, n_1545, n_2374, n_864, n_173, n_859, n_951, n_3341, n_1947, n_1264, n_3587, n_2114, n_3445, n_447, n_247, n_2001, n_1494, n_3407, n_3571, n_3599, n_292, n_3785, n_625, n_854, n_1462, n_1799, n_2069, n_2396, n_3621, n_1580, n_674, n_417, n_1939, n_2486, n_3434, n_1806, n_516, n_933, n_2244, n_3815, n_2257, n_1152, n_3501, n_3448, n_497, n_1869, n_1607, n_1563, n_606, n_3019, n_275, n_3039, n_2011, n_2096, n_4013, n_26, n_4033, n_877, n_2105, n_2538, n_3776, n_2024, n_2, n_2530, n_1696, n_2483, n_3163, n_755, n_1118, n_6, n_1686, n_947, n_1285, n_373, n_3710, n_307, n_3851, n_1860, n_2543, n_1359, n_530, n_87, n_150, n_1107, n_1728, n_556, n_2031, n_2076, n_2482, n_3036, n_3891, n_2677, n_1230, n_668, n_375, n_301, n_1896, n_2165, n_2147, n_929, n_3010, n_3180, n_3379, n_3832, n_3532, n_2770, n_1124, n_3987, n_4061, n_1818, n_2127, n_902, n_1576, n_191, n_1104, n_1294, n_659, n_51, n_1705, n_2584, n_1257, n_2639, n_171, n_1182, n_3188, n_3325, n_3107, n_3531, n_3403, n_4021, n_579, n_1698, n_3880, n_1261, n_2329, n_938, n_1098, n_2963, n_3624, n_3834, n_2142, n_3186, n_3461, n_3082, n_320, n_1154, n_2189, n_3796, n_3332, n_1242, n_3283, n_1135, n_3048, n_3258, n_3937, n_3696, n_24, n_406, n_519, n_2323, n_2203, n_2597, n_1016, n_1243, n_546, n_2959, n_101, n_3340, n_2047, n_1280, n_3277, n_3782, n_1845, n_281, n_240, n_2052, n_2193, n_2978, n_2058, n_2458, n_2478, n_3650, n_291, n_3786, n_231, n_257, n_2761, n_731, n_371, n_1483, n_2888, n_3638, n_1314, n_1512, n_3157, n_709, n_1490, n_317, n_1236, n_1633, n_2537, n_2983, n_3763, n_569, n_2669, n_2144, n_1778, n_3214, n_227, n_2306, n_920, n_2515, n_3022, n_3810, n_1289, n_1517, n_2091, n_2466, n_2635, n_2652, n_94, n_335, n_3631, n_2715, n_3806, n_3087, n_2085, n_3489, n_1669, n_2566, n_370, n_976, n_1949, n_343, n_1449, n_308, n_1946, n_2936, n_1566, n_2032, n_297, n_2587, n_156, n_2149, n_1078, n_2782, n_1670, n_2672, n_775, n_219, n_3060, n_157, n_2651, n_3947, n_3490, n_3656, n_600, n_1484, n_2071, n_2561, n_1374, n_1328, n_2643, n_223, n_2141, n_1948, n_3013, n_3183, n_1984, n_3437, n_3868, n_2099, n_2408, n_3446, n_3353, n_264, n_1877, n_3687, n_1831, n_1598, n_3049, n_1723, n_955, n_1850, n_163, n_3028, n_339, n_1146, n_882, n_183, n_243, n_2384, n_1036, n_1097, n_1749, n_347, n_3156, n_59, n_550, n_696, n_3101, n_3669, n_897, n_215, n_350, n_196, n_798, n_3376, n_646, n_1428, n_2663, n_436, n_1394, n_2659, n_3653, n_1414, n_1216, n_290, n_580, n_2693, n_3798, n_3702, n_1040, n_4065, n_3836, n_2202, n_2648, n_3963, n_1872, n_3389, n_1852, n_2159, n_578, n_2976, n_3876, n_926, n_2180, n_2249, n_344, n_2353, n_1218, n_1931, n_2439, n_2632, n_2276, n_3089, n_422, n_475, n_777, n_1070, n_1547, n_2089, n_3420, n_1030, n_72, n_2470, n_1755, n_3222, n_415, n_1071, n_485, n_1165, n_1267, n_1561, n_496, n_1801, n_3985, n_1391, n_958, n_1034, n_670, n_1513, n_2908, n_2970, n_3361, n_1600, n_48, n_521, n_3744, n_663, n_845, n_2235, n_1862, n_673, n_837, n_3980, n_1239, n_2915, n_528, n_2300, n_2791, n_1796, n_2551, n_3291, n_680, n_1473, n_1587, n_2682, n_395, n_164, n_553, n_901, n_3755, n_2432, n_3668, n_813, n_1521, n_1284, n_1590, n_3440, n_3405, n_214, n_2174, n_2714, n_1748, n_3563, n_2934, n_1672, n_2506, n_675, n_2699, n_4064, n_888, n_1880, n_2769, n_3542, n_2337, n_3436, n_1167, n_1626, n_3550, n_637, n_2615, n_3940, n_1384, n_1556, n_184, n_446, n_3907, n_1863, n_1064, n_144, n_858, n_2079, n_3841, n_2238, n_114, n_96, n_923, n_2118, n_691, n_1151, n_2985, n_2944, n_881, n_1405, n_2407, n_1706, n_468, n_3418, n_213, n_129, n_342, n_2932, n_2753, n_464, n_2980, n_363, n_1582, n_197, n_3637, n_1069, n_3306, n_1784, n_2859, n_2842, n_1075, n_3262, n_3136, n_1836, n_2868, n_3395, n_1450, n_4080, n_4006, n_3141, n_1322, n_2101, n_1471, n_1986, n_2863, n_2072, n_3164, n_2738, n_1750, n_3570, n_3690, n_1459, n_460, n_889, n_2358, n_973, n_3986, n_3716, n_4025, n_2968, n_1700, n_2833, n_477, n_3191, n_571, n_1585, n_461, n_2684, n_2712, n_3593, n_3193, n_3837, n_3885, n_1971, n_1599, n_3936, n_3252, n_2275, n_2855, n_3507, n_3273, n_3821, n_2713, n_3544, n_2644, n_2700, n_1211, n_1197, n_3367, n_4020, n_2951, n_1523, n_2730, n_1950, n_3008, n_3709, n_907, n_1447, n_2251, n_3096, n_1377, n_3915, n_2370, n_190, n_3496, n_3954, n_989, n_2544, n_1039, n_2214, n_3339, n_34, n_2055, n_3427, n_228, n_283, n_3025, n_3349, n_1403, n_3735, n_4067, n_2248, n_4042, n_2356, n_488, n_736, n_892, n_3320, n_3007, n_2688, n_1000, n_1202, n_2750, n_3899, n_2620, n_1278, n_2622, n_2062, n_2668, n_3714, n_1002, n_1463, n_1581, n_2100, n_49, n_3071, n_3739, n_4089, n_3651, n_310, n_3310, n_54, n_593, n_3487, n_2258, n_4069, n_12, n_748, n_586, n_1058, n_1667, n_3359, n_838, n_2784, n_3718, n_3983, n_2919, n_332, n_3092, n_1053, n_3470, n_1224, n_2865, n_349, n_2557, n_1926, n_2706, n_1248, n_230, n_1331, n_953, n_279, n_1014, n_1241, n_3676, n_70, n_2150, n_3146, n_2241, n_2757, n_3789, n_2152, n_3598, n_289, n_963, n_1052, n_954, n_627, n_3781, n_1385, n_440, n_793, n_478, n_2590, n_2776, n_2140, n_2385, n_3580, n_1819, n_2330, n_2139, n_2942, n_476, n_2987, n_1527, n_2042, n_534, n_3106, n_1882, n_884, n_3328, n_345, n_944, n_1754, n_3889, n_3611, n_1623, n_2862, n_2175, n_2921, n_2720, n_2324, n_1854, n_91, n_2606, n_2674, n_3187, n_1565, n_4088, n_3508, n_2828, n_3682, n_3371, n_1809, n_1856, n_182, n_143, n_647, n_3433, n_237, n_4024, n_407, n_1072, n_2218, n_2267, n_832, n_857, n_2305, n_3392, n_3430, n_3975, n_2636, n_2450, n_3208, n_207, n_561, n_1319, n_2379, n_3331, n_3447, n_2616, n_2911, n_3992, n_3305, n_2154, n_1825, n_1951, n_1883, n_1906, n_2759, n_1712, n_1387, n_3528, n_3649, n_2262, n_2462, n_2514, n_1532, n_2322, n_2271, n_2625, n_18, n_3257, n_3625, n_1027, n_971, n_1156, n_117, n_326, n_794, n_404, n_2798, n_2331, n_2945, n_2293, n_686, n_3989, n_2837, n_847, n_3804, n_4051, n_1393, n_2319, n_596, n_1775, n_2979, n_3296, n_2028, n_1368, n_3481, n_2762, n_558, n_3655, n_2808, n_702, n_1276, n_3009, n_2548, n_822, n_1412, n_2676, n_1709, n_2679, n_3981, n_2108, n_3640, n_728, n_266, n_1162, n_272, n_1538, n_2930, n_1838, n_1199, n_1847, n_1779, n_2767, n_2777, n_2603, n_3514, n_3116, n_352, n_1884, n_2434, n_2660, n_53, n_3602, n_1038, n_2967, n_520, n_1369, n_3909, n_409, n_2611, n_1841, n_1660, n_887, n_1905, n_2553, n_154, n_3706, n_3207, n_2581, n_71, n_3944, n_2195, n_2529, n_3224, n_300, n_2698, n_3752, n_4090, n_809, n_3923, n_870, n_931, n_599, n_1711, n_1662, n_1891, n_1481, n_2626, n_3441, n_3042, n_1942, n_434, n_1978, n_1544, n_4001, n_2510, n_3047, n_3526, n_868, n_2454, n_639, n_2804, n_914, n_3659, n_2120, n_411, n_414, n_2546, n_1629, n_1293, n_2801, n_3120, n_965, n_1876, n_1743, n_4007, n_3790, n_4011, n_3491, n_935, n_121, n_1175, n_817, n_2763, n_360, n_36, n_1479, n_1810, n_2350, n_2813, n_64, n_2825, n_1888, n_2009, n_759, n_3643, n_3895, n_2222, n_1892, n_3510, n_28, n_3745, n_806, n_2990, n_1997, n_2667, n_1766, n_3218, n_3748, n_1477, n_3142, n_324, n_1635, n_1963, n_2226, n_1571, n_2891, n_3119, n_187, n_1189, n_2690, n_4028, n_103, n_4082, n_97, n_3370, n_11, n_2215, n_3479, n_4085, n_7, n_1259, n_4073, n_1690, n_3819, n_706, n_746, n_1649, n_3150, n_747, n_2064, n_52, n_784, n_3978, n_110, n_2449, n_3867, n_1733, n_1244, n_3500, n_2413, n_431, n_1194, n_1925, n_3660, n_2297, n_1815, n_3279, n_2621, n_615, n_851, n_1759, n_843, n_1788, n_2177, n_2491, n_3747, n_523, n_913, n_1537, n_705, n_3833, n_865, n_61, n_2227, n_3775, n_678, n_2671, n_697, n_127, n_1222, n_75, n_1679, n_2190, n_3346, n_776, n_1798, n_2022, n_3814, n_1790, n_2518, n_2876, n_1415, n_367, n_2629, n_2592, n_3416, n_452, n_525, n_3484, n_3620, n_1260, n_1746, n_1647, n_2181, n_2479, n_2838, n_1829, n_1464, n_3133, n_3513, n_649, n_547, n_2563, n_43, n_1444, n_4030, n_1191, n_2387, n_2992, n_1674, n_3725, n_1833, n_116, n_3138, n_1830, n_2517, n_2073, n_1710, n_284, n_1128, n_2928, n_3128, n_139, n_1734, n_3038, n_744, n_590, n_629, n_3770, n_4014, n_2631, n_1308, n_2871, n_2178, n_3068, n_1767, n_3144, n_2943, n_2913, n_2336, n_3143, n_3168, n_254, n_1680, n_1233, n_3469, n_2607, n_3994, n_23, n_1615, n_1529, n_2005, n_526, n_1916, n_3317, n_293, n_372, n_677, n_244, n_47, n_1333, n_2469, n_1121, n_2723, n_3355, n_314, n_368, n_433, n_604, n_2007, n_8, n_3220, n_949, n_2539, n_3917, n_3942, n_3263, n_100, n_2582, n_1443, n_1008, n_3855, n_946, n_1539, n_2736, n_1001, n_1503, n_2054, n_3765, n_498, n_1468, n_1559, n_3823, n_1765, n_3455, n_1866, n_689, n_3158, n_738, n_1624, n_3000, n_640, n_3452, n_1510, n_252, n_624, n_1380, n_1744, n_2623, n_1617, n_295, n_133, n_1010, n_1994, n_1231, n_739, n_1279, n_1406, n_3108, n_3113, n_3111, n_2718, n_1195, n_1837, n_1839, n_610, n_2577, n_3760, n_4078, n_1760, n_2875, n_936, n_568, n_1500, n_2960, n_39, n_1090, n_2796, n_757, n_3844, n_3280, n_2342, n_633, n_2856, n_4054, n_439, n_3471, n_106, n_1832, n_259, n_448, n_1851, n_758, n_999, n_3205, n_2046, n_2848, n_2741, n_2937, n_3666, n_3003, n_3610, n_1933, n_3828, n_2290, n_93, n_1656, n_3564, n_3288, n_1158, n_3095, n_2045, n_3369, n_3783, n_3988, n_1509, n_1874, n_2040, n_563, n_2060, n_3199, n_2613, n_1987, n_2805, n_3667, n_1145, n_878, n_524, n_3843, n_3457, n_204, n_394, n_1678, n_1049, n_1153, n_3856, n_2145, n_741, n_1639, n_1306, n_3703, n_1068, n_3030, n_3558, n_1871, n_2580, n_3630, n_2545, n_2787, n_3685, n_2914, n_1964, n_2869, n_122, n_4002, n_331, n_10, n_906, n_1163, n_3271, n_2039, n_1207, n_919, n_908, n_4086, n_2412, n_2406, n_3623, n_90, n_2846, n_724, n_3753, n_1781, n_2084, n_2925, n_3648, n_2035, n_658, n_2061, n_3773, n_3555, n_3579, n_3918, n_3075, n_3173, n_2378, n_2509, n_1740, n_3236, n_2398, n_1362, n_3969, n_2857, n_3932, n_1586, n_456, n_959, n_2459, n_3031, n_535, n_152, n_3396, n_3701, n_940, n_1445, n_9, n_3516, n_4023, n_1492, n_2155, n_2516, n_3797, n_1923, n_1773, n_592, n_3243, n_1169, n_45, n_1596, n_1692, n_2666, n_2982, n_3385, n_1017, n_2481, n_2947, n_3545, n_2171, n_123, n_978, n_2768, n_2116, n_2314, n_1434, n_1054, n_2507, n_1474, n_1665, n_1269, n_4019, n_2420, n_2900, n_1095, n_3343, n_3515, n_1828, n_1614, n_2886, n_267, n_514, n_457, n_1079, n_1045, n_1208, n_2093, n_2038, n_2320, n_2339, n_2473, n_3287, n_2137, n_3378, n_603, n_1431, n_2583, n_484, n_1593, n_1033, n_3767, n_442, n_3426, n_3454, n_2299, n_131, n_2540, n_2873, n_3820, n_636, n_3741, n_660, n_3410, n_2087, n_1640, n_2162, n_1732, n_1009, n_2847, n_1148, n_2051, n_109, n_742, n_750, n_2029, n_995, n_454, n_3221, n_2168, n_2790, n_1609, n_374, n_3629, n_3021, n_1989, n_3818, n_185, n_2359, n_2941, n_3674, n_396, n_1887, n_3502, n_2523, n_1383, n_3098, n_1073, n_255, n_2346, n_2457, n_662, n_459, n_2312, n_3990, n_218, n_962, n_3475, n_1215, n_3015, n_1171, n_1578, n_723, n_1920, n_1065, n_1592, n_2536, n_1336, n_2882, n_3719, n_1721, n_1959, n_1758, n_2338, n_3681, n_2952, n_2737, n_1574, n_3672, n_2399, n_3058, n_2812, n_473, n_2048, n_3197, n_3109, n_3607, n_2355, n_2133, n_1921, n_2721, n_1309, n_1878, n_1426, n_3830, n_1043, n_2585, n_355, n_3505, n_486, n_3002, n_1800, n_1548, n_2725, n_614, n_337, n_1421, n_88, n_2571, n_1286, n_3730, n_3883, n_1177, n_3276, n_1355, n_168, n_974, n_2565, n_727, n_3897, n_1159, n_3845, n_957, n_3787, n_773, n_208, n_142, n_2124, n_743, n_3001, n_2081, n_299, n_303, n_3945, n_3149, n_296, n_613, n_1119, n_2156, n_1240, n_2261, n_1820, n_2729, n_3268, n_3597, n_2418, n_3827, n_65, n_829, n_2519, n_3354, n_2724, n_1612, n_2179, n_1416, n_2077, n_2897, n_3614, n_2909, n_1724, n_2111, n_2521, n_3301, n_361, n_3466, n_3458, n_700, n_1237, n_573, n_69, n_1420, n_3185, n_1132, n_3330, n_388, n_1366, n_1300, n_3960, n_2595, n_1127, n_3248, n_2277, n_761, n_2477, n_3523, n_1785, n_1568, n_2829, n_3905, n_1006, n_3411, n_3887, n_4087, n_2110, n_329, n_3811, n_274, n_4093, n_1270, n_1664, n_3200, n_1486, n_582, n_3586, n_1332, n_3519, n_2231, n_1390, n_2017, n_73, n_2474, n_2879, n_2604, n_19, n_2090, n_3374, n_3153, n_3045, n_1870, n_309, n_30, n_512, n_2367, n_1591, n_2033, n_4071, n_84, n_3453, n_130, n_322, n_1682, n_1980, n_2390, n_2628, n_1249, n_3399, n_2896, n_652, n_1111, n_3213, n_1365, n_4074, n_1927, n_25, n_3065, n_2132, n_1349, n_1093, n_288, n_2400, n_1031, n_3645, n_263, n_609, n_1041, n_1265, n_3223, n_1909, n_3838, n_44, n_224, n_3077, n_3929, n_2681, n_1562, n_383, n_3103, n_834, n_3474, n_112, n_765, n_3675, n_2255, n_2424, n_2272, n_893, n_3984, n_1015, n_1140, n_891, n_1651, n_1965, n_239, n_3387, n_630, n_1902, n_2151, n_1941, n_55, n_2106, n_2775, n_2716, n_3938, n_1913, n_2878, n_504, n_1823, n_511, n_3679, n_3779, n_874, n_2464, n_358, n_3422, n_3888, n_1101, n_2831, n_77, n_102, n_1106, n_1456, n_3557, n_2230, n_3498, n_2015, n_2365, n_1875, n_1982, n_1304, n_2803, n_1324, n_2851, n_3707, n_987, n_3189, n_1846, n_3037, n_261, n_174, n_2066, n_1885, n_1455, n_3429, n_767, n_993, n_1903, n_2490, n_1407, n_3849, n_3946, n_2452, n_1551, n_3154, n_545, n_441, n_860, n_3229, n_450, n_2849, n_1805, n_3925, n_2176, n_2204, n_2905, n_1816, n_3692, n_429, n_948, n_3965, n_3566, n_1217, n_2220, n_4059, n_2455, n_628, n_365, n_1849, n_3788, n_4084, n_2410, n_729, n_1131, n_1084, n_1961, n_970, n_4037, n_1935, n_911, n_2922, n_1430, n_83, n_3275, n_3499, n_2645, n_2467, n_513, n_3366, n_2727, n_1094, n_1354, n_560, n_1534, n_340, n_2288, n_3421, n_1351, n_2240, n_2696, n_4063, n_1044, n_1205, n_2436, n_346, n_1209, n_3029, n_1552, n_2508, n_3242, n_3592, n_3618, n_4031, n_495, n_602, n_3525, n_574, n_2593, n_3486, n_1435, n_879, n_3394, n_3793, n_16, n_3683, n_2416, n_58, n_2405, n_3642, n_623, n_3995, n_3286, n_2088, n_405, n_2953, n_3808, n_824, n_4036, n_359, n_1645, n_3881, n_4041, n_2461, n_490, n_1327, n_2858, n_2243, n_4060, n_996, n_921, n_1684, n_233, n_2658, n_3590, n_1717, n_572, n_366, n_2895, n_815, n_1795, n_2128, n_2578, n_3097, n_3483, n_128, n_1821, n_3894, n_120, n_2929, n_3424, n_327, n_3478, n_135, n_1381, n_2555, n_3751, n_2662, n_2740, n_3824, n_3890, n_1611, n_1037, n_2368, n_3388, n_2656, n_1080, n_2301, n_1274, n_3583, n_2890, n_3560, n_3059, n_3524, n_4076, n_2554, n_3465, n_1316, n_1708, n_2419, n_3215, n_426, n_1438, n_3698, n_3927, n_1082, n_1840, n_589, n_3961, n_716, n_1630, n_2122, n_2512, n_3589, n_562, n_1436, n_62, n_3549, n_1691, n_952, n_2786, n_2534, n_2092, n_3171, n_1229, n_391, n_701, n_1437, n_1023, n_2075, n_645, n_539, n_3658, n_3449, n_803, n_1092, n_2694, n_238, n_1776, n_3559, n_2198, n_2610, n_2661, n_2572, n_2989, n_2281, n_2131, n_2789, n_3026, n_3993, n_2216, n_531, n_3020, n_3677, n_1757, n_890, n_1897, n_764, n_1919, n_1056, n_1424, n_162, n_960, n_3462, n_3588, n_2933, n_2308, n_3468, n_1893, n_2910, n_222, n_3419, n_3886, n_1290, n_1123, n_1467, n_1047, n_2053, n_2163, n_634, n_2328, n_199, n_1958, n_32, n_2254, n_1252, n_348, n_3860, n_1382, n_1029, n_925, n_3546, n_1206, n_424, n_2647, n_3784, n_3160, n_1311, n_2191, n_2864, n_2969, n_3941, n_3195, n_1519, n_256, n_950, n_3190, n_2428, n_1553, n_3678, n_3847, n_2664, n_1811, n_2443, n_2624, n_3012, n_3456, n_380, n_419, n_1346, n_3053, n_444, n_1299, n_3244, n_2158, n_1808, n_3893, n_3290, n_1060, n_1141, n_316, n_2266, n_389, n_3130, n_2465, n_2824, n_3033, n_2650, n_3298, n_418, n_248, n_136, n_86, n_146, n_912, n_315, n_968, n_3548, n_451, n_619, n_408, n_2440, n_1386, n_1699, n_376, n_3334, n_967, n_1442, n_2923, n_3665, n_3494, n_2541, n_74, n_1139, n_2731, n_3264, n_515, n_2333, n_57, n_351, n_3953, n_885, n_2916, n_3166, n_397, n_1432, n_3875, n_3976, n_1357, n_483, n_2125, n_3771, n_3979, n_683, n_1632, n_3110, n_2998, n_1057, n_1051, n_1085, n_1066, n_4003, n_3800, n_721, n_2402, n_1157, n_3073, n_2403, n_841, n_1050, n_22, n_802, n_1954, n_4048, n_4026, n_2265, n_46, n_3162, n_1608, n_983, n_1844, n_2760, n_2792, n_3554, n_38, n_3377, n_2870, n_3777, n_280, n_1305, n_3749, n_3178, n_873, n_1826, n_3962, n_3991, n_378, n_1112, n_3134, n_2304, n_2999, n_762, n_1283, n_1644, n_17, n_2334, n_2637, n_3695, n_690, n_33, n_4046, n_1974, n_2463, n_583, n_2086, n_3537, n_2289, n_3080, n_3051, n_302, n_4096, n_1343, n_2701, n_2783, n_2263, n_3362, n_2881, n_1203, n_1631, n_3750, n_3282, n_2472, n_821, n_3816, n_1763, n_2341, n_3105, n_3231, n_1966, n_3632, n_1768, n_321, n_2294, n_1179, n_621, n_753, n_2475, n_2733, n_455, n_1048, n_1719, n_2993, n_3864, n_1288, n_212, n_385, n_2785, n_2556, n_507, n_2269, n_2732, n_3569, n_2309, n_2415, n_2948, n_3274, n_3041, n_3299, n_2646, n_1560, n_3715, n_1605, n_2236, n_330, n_1228, n_2816, n_2123, n_3209, n_972, n_3504, n_692, n_2037, n_2685, n_3920, n_3040, n_1953, n_1938, n_820, n_1200, n_2499, n_1911, n_3616, n_2460, n_4058, n_3568, n_3664, n_2589, n_3203, n_1301, n_1363, n_1668, n_3737, n_3913, n_1185, n_991, n_2903, n_3417, n_3482, n_3866, n_828, n_1967, n_779, n_576, n_1143, n_1579, n_2233, n_3717, n_4034, n_1329, n_2743, n_2675, n_3255, n_1312, n_1439, n_804, n_537, n_2827, n_1688, n_3052, n_945, n_2997, n_492, n_3743, n_3327, n_153, n_1504, n_943, n_3326, n_3956, n_341, n_3572, n_250, n_992, n_3067, n_1932, n_3375, n_2755, n_4047, n_543, n_260, n_842, n_3734, n_650, n_984, n_694, n_3237, n_2082, n_286, n_1992, n_2429, n_1643, n_883, n_1983, n_3167, n_4029, n_3400, n_470, n_325, n_449, n_1594, n_132, n_1214, n_1342, n_1400, n_3423, n_900, n_2362, n_856, n_2609, n_3870, n_1793, n_3382, n_1976, n_2223, n_3044, n_3574, n_918, n_3529, n_3854, n_942, n_2169, n_1804, n_189, n_1147, n_1557, n_1977, n_2153, n_2468, n_1610, n_13, n_1077, n_1422, n_3196, n_4095, n_3078, n_2364, n_2533, n_540, n_3492, n_618, n_3094, n_896, n_2310, n_2780, n_323, n_3952, n_2287, n_2860, n_3316, n_195, n_356, n_2291, n_3099, n_4043, n_3704, n_2596, n_894, n_1636, n_2056, n_3253, n_1730, n_3601, n_3603, n_4027, n_831, n_2280, n_2192, n_964, n_3633, n_3363, n_1373, n_1350, n_1511, n_1865, n_2973, n_1470, n_1096, n_2094, n_2670, n_234, n_1575, n_1697, n_1735, n_833, n_2318, n_2393, n_3689, n_2020, n_3831, n_5, n_1646, n_2502, n_3801, n_225, n_2504, n_1307, n_1881, n_2974, n_988, n_2749, n_2043, n_2901, n_1940, n_814, n_2707, n_2751, n_2793, n_3372, n_3451, n_192, n_2971, n_3442, n_1549, n_1934, n_2311, n_1201, n_1114, n_3950, n_4000, n_655, n_3240, n_2025, n_1616, n_3998, n_1446, n_2285, n_3147, n_2758, n_669, n_472, n_1458, n_1176, n_1472, n_2298, n_2471, n_1807, n_387, n_3869, n_1149, n_2618, n_398, n_1671, n_635, n_2559, n_763, n_3230, n_1020, n_1062, n_3342, n_211, n_2303, n_1824, n_1917, n_2295, n_1219, n_3386, n_3931, n_3, n_3708, n_1204, n_4010, n_2840, n_3729, n_2810, n_2325, n_178, n_2747, n_2446, n_3488, n_1814, n_1035, n_2822, n_3861, n_287, n_3780, n_555, n_783, n_1848, n_1928, n_2126, n_2893, n_3636, n_1188, n_2588, n_2962, n_4004, n_1722, n_3957, n_661, n_2441, n_3848, n_41, n_1802, n_3083, n_2600, n_3919, n_4079, n_3898, n_849, n_2795, n_15, n_4091, n_336, n_584, n_681, n_1638, n_1786, n_2981, n_50, n_430, n_2002, n_2282, n_3608, n_510, n_2800, n_216, n_3712, n_2371, n_2935, n_311, n_3233, n_3829, n_3380, n_3177, n_4053, n_830, n_2098, n_1296, n_2627, n_3409, n_3460, n_2352, n_3538, n_1413, n_801, n_4040, n_2207, n_2080, n_2377, n_2619, n_2340, n_3085, n_2444, n_2068, n_241, n_3552, n_875, n_357, n_1110, n_1655, n_445, n_2641, n_3198, n_749, n_1895, n_3123, n_3684, n_3137, n_2574, n_1134, n_1358, n_717, n_165, n_939, n_3697, n_482, n_2361, n_1088, n_588, n_1173, n_789, n_3393, n_1232, n_1603, n_734, n_638, n_2638, n_866, n_107, n_969, n_1401, n_4018, n_4044, n_3900, n_4062, n_3520, n_3971, n_2492, n_1019, n_1105, n_249, n_1998, n_304, n_3759, n_1338, n_577, n_4005, n_2016, n_1522, n_3872, n_2949, n_1687, n_1637, n_2034, n_1419, n_2711, n_3933, n_338, n_149, n_1653, n_693, n_2270, n_1506, n_3206, n_2653, n_3578, n_3966, n_14, n_836, n_990, n_2867, n_3812, n_2496, n_1886, n_1389, n_1894, n_975, n_1908, n_1256, n_1702, n_2259, n_2794, n_567, n_1465, n_3145, n_3124, n_778, n_1122, n_4068, n_151, n_3192, n_2608, n_3877, n_306, n_3764, n_2657, n_458, n_770, n_2995, n_1375, n_2494, n_3547, n_2649, n_3977, n_1102, n_3727, n_2852, n_3774, n_4052, n_2392, n_3459, n_3093, n_1843, n_711, n_1499, n_3061, n_3155, n_85, n_1187, n_3517, n_2633, n_1441, n_3100, n_2522, n_2435, n_1392, n_1597, n_1929, n_2807, n_1164, n_1659, n_1834, n_2097, n_2313, n_2542, n_489, n_1174, n_2431, n_3324, n_3356, n_3758, n_2835, n_3914, n_3911, n_2558, n_1371, n_617, n_1303, n_2206, n_2063, n_3803, n_3182, n_1572, n_1968, n_3742, n_3269, n_2564, n_2252, n_876, n_1516, n_3736, n_1190, n_3506, n_3896, n_1736, n_3605, n_1685, n_3958, n_118, n_2409, n_601, n_917, n_3450, n_1714, n_966, n_253, n_1116, n_2000, n_1661, n_3402, n_1212, n_2074, n_1541, n_2576, n_3565, n_172, n_206, n_217, n_726, n_3174, n_982, n_2575, n_2988, n_3390, n_1573, n_1453, n_1731, n_2217, n_3746, n_818, n_2373, n_1970, n_861, n_1713, n_1183, n_3398, n_2307, n_2766, n_3817, n_1658, n_899, n_1253, n_210, n_1737, n_2201, n_2722, n_2117, n_2745, n_3408, n_1904, n_2640, n_1993, n_774, n_3835, n_1628, n_2493, n_2205, n_3432, n_1335, n_1514, n_1777, n_1957, n_1059, n_1345, n_3967, n_176, n_1133, n_1771, n_1912, n_3401, n_1899, n_3226, n_557, n_1410, n_1005, n_607, n_1003, n_679, n_710, n_3090, n_2067, n_527, n_1168, n_707, n_2219, n_2437, n_2885, n_3762, n_3902, n_3533, n_2877, n_3318, n_4070, n_2148, n_937, n_2445, n_1427, n_2779, n_3485, n_393, n_108, n_487, n_1584, n_665, n_1726, n_1835, n_3035, n_3654, n_66, n_1440, n_177, n_3839, n_2164, n_421, n_1988, n_3333, n_2115, n_1853, n_1356, n_2845, n_1787, n_2634, n_910, n_2232, n_3034, n_2212, n_2602, n_1657, n_768, n_1475, n_1302, n_1774, n_1725, n_205, n_1136, n_1313, n_1491, n_754, n_3972, n_2811, n_1496, n_3348, n_179, n_1125, n_125, n_410, n_2547, n_3014, n_3639, n_708, n_529, n_1812, n_735, n_2501, n_3079, n_232, n_1915, n_1109, n_126, n_895, n_2532, n_1310, n_2605, n_3358, n_2121, n_1803, n_202, n_3791, n_3308, n_2665, n_427, n_1399, n_1543, n_1991, n_1979, n_791, n_732, n_1533, n_2224, n_193, n_3368, n_2924, n_3467, n_808, n_2484, n_797, n_3530, n_1025, n_1930, n_1955, n_3731, n_2765, n_3329, n_500, n_2994, n_1067, n_3805, n_3825, n_2946, n_1720, n_148, n_2830, n_2401, n_3135, n_435, n_3657, n_2003, n_159, n_766, n_1457, n_3928, n_541, n_2692, n_3573, n_3148, n_538, n_2354, n_2246, n_2008, n_1117, n_799, n_2264, n_2754, n_687, n_3534, n_715, n_3901, n_1742, n_1480, n_1482, n_1213, n_2489, n_1266, n_3970, n_3757, n_536, n_3438, n_872, n_2012, n_594, n_3792, n_200, n_1291, n_3974, n_3381, n_3871, n_4094, n_3503, n_1297, n_1753, n_2283, n_2866, n_3278, n_1782, n_2245, n_3561, n_1155, n_1418, n_89, n_1972, n_1524, n_1689, n_1485, n_2806, n_115, n_1011, n_1184, n_2184, n_985, n_1855, n_2425, n_2917, n_869, n_810, n_2965, n_3536, n_3661, n_416, n_3635, n_827, n_3217, n_3404, n_3425, n_401, n_1703, n_3312, n_4055, n_1352, n_2926, n_626, n_2197, n_2199, n_3540, n_1650, n_3670, n_1144, n_3973, n_1137, n_1570, n_2814, n_3046, n_3882, n_3934, n_1170, n_305, n_2023, n_2213, n_3826, n_3249, n_3211, n_3285, n_2351, n_2211, n_2095, n_3121, n_3922, n_137, n_3846, n_676, n_294, n_318, n_2103, n_653, n_3968, n_2160, n_642, n_3337, n_2228, n_2527, n_1602, n_2498, n_194, n_855, n_1178, n_1461, n_2697, n_850, n_684, n_3074, n_124, n_3204, n_268, n_2421, n_2286, n_2902, n_664, n_1999, n_503, n_2372, n_2065, n_2136, n_3673, n_2480, n_4017, n_235, n_3768, n_1372, n_2861, n_605, n_2630, n_1273, n_3943, n_1822, n_3397, n_353, n_3740, n_620, n_643, n_2363, n_2430, n_4072, n_916, n_1081, n_2549, n_493, n_2705, n_3005, n_2332, n_1235, n_703, n_698, n_980, n_1115, n_2433, n_3293, n_3129, n_1282, n_1318, n_1783, n_780, n_2977, n_3606, n_2601, n_3043, n_4022, n_998, n_3802, n_2375, n_2550, n_1454, n_3723, n_467, n_1227, n_1531, n_840, n_1334, n_1907, n_3600, n_501, n_823, n_245, n_2686, n_2528, n_725, n_2344, n_3892, n_1388, n_1417, n_1295, n_2836, n_4035, n_2316, n_672, n_1985, n_3055, n_1898, n_2107, n_3294, n_3219, n_3711, n_3315, n_581, n_2906, n_382, n_554, n_1625, n_2130, n_3415, n_2187, n_2284, n_898, n_2817, n_3172, n_3139, n_2773, n_3239, n_3292, n_2598, n_3878, n_1762, n_1013, n_3365, n_3476, n_3686, n_1452, n_718, n_2687, n_265, n_3023, n_3553, n_1120, n_719, n_443, n_1791, n_198, n_1890, n_1747, n_714, n_2850, n_1683, n_1817, n_909, n_1944, n_1497, n_1530, n_4075, n_3982, n_2654, n_997, n_3431, n_3104, n_932, n_3169, n_3151, n_612, n_3822, n_3131, n_2078, n_1409, n_3850, n_788, n_1326, n_3070, n_3284, n_4066, n_3647, n_119, n_3176, n_2884, n_1268, n_2996, n_559, n_825, n_2819, n_3126, n_1981, n_508, n_2186, n_506, n_1320, n_1663, n_737, n_1718, n_4050, n_3700, n_3609, n_986, n_2315, n_509, n_3228, n_1317, n_147, n_1518, n_1715, n_2102, n_3581, n_2562, n_1281, n_67, n_1952, n_4077, n_1192, n_2221, n_1024, n_3576, n_1063, n_3720, n_1889, n_209, n_1792, n_1564, n_1868, n_1613, n_733, n_1489, n_1922, n_2966, n_4049, n_1376, n_941, n_2326, n_981, n_2560, n_3862, n_1569, n_2188, n_68, n_3495, n_3879, n_867, n_186, n_2348, n_2422, n_3959, n_134, n_2239, n_587, n_2950, n_63, n_792, n_756, n_1429, n_399, n_1238, n_2448, n_3140, n_3852, n_548, n_3170, n_3724, n_812, n_298, n_2104, n_2748, n_3311, n_518, n_505, n_2057, n_3272, n_4008, n_3011, n_1772, n_282, n_752, n_905, n_1476, n_1108, n_2898, n_782, n_2717, n_2818, n_1100, n_3646, n_1861, n_2129, n_1395, n_3345, n_862, n_3584, n_1425, n_760, n_3858, n_1901, n_3069, n_3756, n_1900, n_1620, n_3032, n_381, n_3628, n_2889, n_3691, n_220, n_390, n_1330, n_1867, n_31, n_1945, n_2772, n_481, n_3018, n_1675, n_3072, n_1924, n_2573, n_3084, n_3081, n_3313, n_1727, n_2710, n_1554, n_2939, n_1745, n_3924, n_2735, n_769, n_2497, n_2006, n_3412, n_3999, n_42, n_2844, n_1995, n_2411, n_3807, n_2138, n_1046, n_271, n_934, n_1618, n_2260, n_826, n_2343, n_1813, n_2447, n_3761, n_886, n_3439, n_2014, n_3056, n_1221, n_2345, n_2986, n_654, n_1172, n_167, n_2535, n_379, n_428, n_1341, n_2726, n_570, n_2774, n_3295, n_1641, n_1361, n_3184, n_2382, n_1707, n_853, n_3062, n_3161, n_377, n_2317, n_751, n_3289, n_2799, n_2172, n_1973, n_786, n_1083, n_1142, n_2376, n_2488, n_1129, n_392, n_2579, n_3477, n_3017, n_158, n_3626, n_2476, n_704, n_787, n_1770, n_138, n_2781, n_2456, n_3904, n_961, n_2250, n_2678, n_1756, n_771, n_2778, n_276, n_95, n_1716, n_2788, n_2872, n_1225, n_2984, n_1520, n_2451, n_169, n_2887, n_522, n_3364, n_1287, n_1262, n_2691, n_400, n_930, n_181, n_4092, n_3908, n_1873, n_1411, n_3926, n_3201, n_3054, n_221, n_622, n_1962, n_3996, n_1577, n_2423, n_3671, n_1087, n_3472, n_2526, n_2854, n_386, n_994, n_1701, n_3344, n_2194, n_848, n_1550, n_2874, n_2764, n_2703, n_1498, n_2167, n_3302, n_3235, n_1223, n_1272, n_2680, n_3391, n_104, n_682, n_1567, n_56, n_141, n_2567, n_3949, n_3543, n_1247, n_2709, n_3102, n_922, n_3122, n_816, n_1648, n_4015, n_591, n_3842, n_145, n_1536, n_3050, n_3265, n_1857, n_4056, n_1344, n_2041, n_313, n_631, n_3627, n_479, n_1246, n_3840, n_1339, n_1478, n_1797, n_432, n_1769, n_2957, n_839, n_3551, n_3903, n_1210, n_3518, n_2964, n_3769, n_1364, n_2956, n_2357, n_3733, n_2183, n_2673, n_2742, n_3314, n_2360, n_3254, n_328, n_140, n_2292, n_1250, n_2173, n_3859, n_369, n_3722, n_3865, n_1842, n_871, n_2442, n_3309, n_3738, n_4045, n_598, n_685, n_928, n_608, n_1367, n_78, n_1943, n_3634, n_1460, n_772, n_2018, n_3464, n_3260, n_1555, n_3117, n_2834, n_3245, n_3357, n_499, n_2531, n_1589, n_517, n_3428, n_98, n_2961, n_402, n_413, n_1086, n_2570, n_2702, n_796, n_1858, n_3351, n_1619, n_3527, n_2815, n_236, n_2119, n_1502, n_2157, n_2552, n_3754, n_1469, n_1012, n_1, n_1396, n_2744, n_1348, n_2030, n_903, n_2453, n_1525, n_1752, n_2397, n_740, n_2883, n_3115, n_203, n_3509, n_3352, n_384, n_2208, n_3076, n_1404, n_80, n_3063, n_3617, n_2912, n_1794, n_3535, n_2182, n_35, n_1315, n_2234, n_277, n_1061, n_3251, n_92, n_1910, n_333, n_1298, n_3955, n_2931, n_1652, n_2209, n_3794, n_462, n_2050, n_2809, n_1193, n_2797, n_1676, n_1255, n_258, n_1113, n_3118, n_29, n_79, n_4039, n_3227, n_3300, n_2321, n_3511, n_1226, n_722, n_1277, n_3680, n_2591, n_3443, n_188, n_2146, n_844, n_201, n_3384, n_471, n_852, n_3497, n_1487, n_40, n_1864, n_3644, n_1028, n_1601, n_4016, n_3336, n_3935, n_781, n_474, n_2940, n_542, n_3435, n_3521, n_463, n_3575, n_1546, n_595, n_502, n_3562, n_3948, n_466, n_2612, n_420, n_1337, n_1495, n_632, n_699, n_979, n_1515, n_2841, n_3165, n_1627, n_2918, n_3232, n_3322, n_3652, n_1245, n_846, n_2427, n_2438, n_2505, n_1673, n_465, n_2832, n_76, n_362, n_1321, n_170, n_1975, n_27, n_2296, n_2070, n_161, n_273, n_1937, n_585, n_2112, n_3250, n_4083, n_1739, n_3181, n_270, n_2958, n_616, n_2278, n_81, n_2594, n_3114, n_3125, n_2394, n_3234, n_1914, n_3612, n_2954, n_2135, n_2335, n_2904, n_3493, n_745, n_2381, n_3303, n_1654, n_3004, n_3323, n_3916, n_2569, n_3112, n_2349, n_1103, n_3921, n_4081, n_3132, n_3556, n_648, n_1379, n_2734, n_3874, n_312, n_2196, n_3591, n_3951, n_3024, n_2170, n_1076, n_2823, n_1091, n_1408, n_3512, n_494, n_1761, n_641, n_3238, n_3210, n_3930, n_730, n_3175, n_3522, n_2036, n_1325, n_3267, n_1595, n_2161, n_354, n_575, n_480, n_425, n_795, n_2404, n_2083, n_695, n_180, n_3281, n_656, n_3307, n_1606, n_2503, n_1220, n_37, n_1694, n_1540, n_3964, n_3266, n_2485, n_3772, n_229, n_1936, n_1956, n_437, n_1642, n_2279, n_3373, n_2655, n_2027, n_3884, n_60, n_403, n_453, n_2642, n_1130, n_720, n_0, n_2500, n_2366, n_1918, n_1526, n_863, n_3726, n_2210, n_805, n_3247, n_3997, n_1604, n_1275, n_2513, n_2525, n_3091, n_2695, n_1764, n_3480, n_2892, n_4032, n_3057, n_3194, n_3582, n_3066, n_113, n_712, n_2414, n_2907, n_246, n_1583, n_2426, n_2826, n_3577, n_3539, n_1042, n_1402, n_2820, n_269, n_3662, n_2049, n_2273, n_285, n_412, n_2719, n_1493, n_657, n_644, n_1741, n_2229, n_1160, n_1397, n_4057, n_491, n_1258, n_1074, n_3347, n_2004, n_3216, n_1621, n_2708, n_3809, n_2113, n_251, n_160, n_566, n_565, n_2586, n_3694, n_1448, n_2225, n_3567, n_3613, n_1507, n_1398, n_2383, n_1879, n_597, n_1996, n_3406, n_3604, n_3444, n_3853, n_1181, n_1505, n_1634, n_3939, n_1196, n_4012, n_2019, n_651, n_1340, n_2274, n_2972, n_334, n_811, n_1558, n_3225, n_807, n_3321, n_2166, n_3910, n_2938, n_3212, n_835, n_175, n_666, n_3319, n_262, n_1433, n_3594, n_1704, n_2256, n_3152, n_3721, n_3335, n_99, n_1254, n_3799, n_1026, n_3413, n_2026, n_1969, n_1234, n_2109, n_319, n_364, n_1138, n_927, n_20, n_1089, n_2013, n_1990, n_2044, n_2689, n_2920, n_3259, n_1004, n_1186, n_1032, n_242, n_2614, n_2511, n_1681, n_2010, n_2991, n_3688, n_3383, n_1018, n_2242, n_2247, n_2752, n_2894, n_3016, n_1693, n_3585, n_2975, n_3473, n_438, n_2599, n_713, n_2704, n_904, n_2839, n_3338, n_1588, n_1622, n_2237, n_3414, n_3463, n_3699, n_166, n_1180, n_1827, n_3360, n_2524, n_3873, n_1271, n_3705, n_2802, n_533, n_1542, n_1251, n_3693, n_4009, n_3159, n_278, n_2728, n_3857, n_2268, n_3778, n_16249);

input n_924;
input n_1263;
input n_3304;
input n_977;
input n_1378;
input n_2253;
input n_2417;
input n_611;
input n_2756;
input n_3912;
input n_1126;
input n_1423;
input n_1729;
input n_2739;
input n_1166;
input n_2380;
input n_1751;
input n_469;
input n_1508;
input n_82;
input n_2771;
input n_785;
input n_3241;
input n_549;
input n_2617;
input n_2200;
input n_3261;
input n_3006;
input n_532;
input n_1161;
input n_3795;
input n_3863;
input n_3027;
input n_1859;
input n_2746;
input n_1677;
input n_1150;
input n_2327;
input n_3179;
input n_3127;
input n_226;
input n_1780;
input n_3256;
input n_3732;
input n_1488;
input n_667;
input n_2899;
input n_2955;
input n_790;
input n_3619;
input n_1055;
input n_3541;
input n_3622;
input n_2386;
input n_3596;
input n_1501;
input n_111;
input n_2395;
input n_3906;
input n_880;
input n_3086;
input n_3297;
input n_544;
input n_1007;
input n_2369;
input n_155;
input n_2927;
input n_552;
input n_1528;
input n_2683;
input n_1370;
input n_1292;
input n_2347;
input n_2520;
input n_2821;
input n_1198;
input n_1360;
input n_2388;
input n_1099;
input n_2568;
input n_3641;
input n_956;
input n_564;
input n_423;
input n_1738;
input n_2021;
input n_3728;
input n_21;
input n_2134;
input n_3064;
input n_2391;
input n_105;
input n_3088;
input n_1021;
input n_1960;
input n_2843;
input n_2185;
input n_4;
input n_3270;
input n_551;
input n_2143;
input n_3713;
input n_2853;
input n_3615;
input n_2059;
input n_1323;
input n_3663;
input n_1466;
input n_688;
input n_1695;
input n_2487;
input n_3766;
input n_1353;
input n_800;
input n_3595;
input n_3246;
input n_3202;
input n_1347;
input n_2495;
input n_2880;
input n_1535;
input n_3813;
input n_1789;
input n_1666;
input n_3350;
input n_2389;
input n_671;
input n_819;
input n_1451;
input n_1022;
input n_4038;
input n_2302;
input n_915;
input n_1545;
input n_2374;
input n_864;
input n_173;
input n_859;
input n_951;
input n_3341;
input n_1947;
input n_1264;
input n_3587;
input n_2114;
input n_3445;
input n_447;
input n_247;
input n_2001;
input n_1494;
input n_3407;
input n_3571;
input n_3599;
input n_292;
input n_3785;
input n_625;
input n_854;
input n_1462;
input n_1799;
input n_2069;
input n_2396;
input n_3621;
input n_1580;
input n_674;
input n_417;
input n_1939;
input n_2486;
input n_3434;
input n_1806;
input n_516;
input n_933;
input n_2244;
input n_3815;
input n_2257;
input n_1152;
input n_3501;
input n_3448;
input n_497;
input n_1869;
input n_1607;
input n_1563;
input n_606;
input n_3019;
input n_275;
input n_3039;
input n_2011;
input n_2096;
input n_4013;
input n_26;
input n_4033;
input n_877;
input n_2105;
input n_2538;
input n_3776;
input n_2024;
input n_2;
input n_2530;
input n_1696;
input n_2483;
input n_3163;
input n_755;
input n_1118;
input n_6;
input n_1686;
input n_947;
input n_1285;
input n_373;
input n_3710;
input n_307;
input n_3851;
input n_1860;
input n_2543;
input n_1359;
input n_530;
input n_87;
input n_150;
input n_1107;
input n_1728;
input n_556;
input n_2031;
input n_2076;
input n_2482;
input n_3036;
input n_3891;
input n_2677;
input n_1230;
input n_668;
input n_375;
input n_301;
input n_1896;
input n_2165;
input n_2147;
input n_929;
input n_3010;
input n_3180;
input n_3379;
input n_3832;
input n_3532;
input n_2770;
input n_1124;
input n_3987;
input n_4061;
input n_1818;
input n_2127;
input n_902;
input n_1576;
input n_191;
input n_1104;
input n_1294;
input n_659;
input n_51;
input n_1705;
input n_2584;
input n_1257;
input n_2639;
input n_171;
input n_1182;
input n_3188;
input n_3325;
input n_3107;
input n_3531;
input n_3403;
input n_4021;
input n_579;
input n_1698;
input n_3880;
input n_1261;
input n_2329;
input n_938;
input n_1098;
input n_2963;
input n_3624;
input n_3834;
input n_2142;
input n_3186;
input n_3461;
input n_3082;
input n_320;
input n_1154;
input n_2189;
input n_3796;
input n_3332;
input n_1242;
input n_3283;
input n_1135;
input n_3048;
input n_3258;
input n_3937;
input n_3696;
input n_24;
input n_406;
input n_519;
input n_2323;
input n_2203;
input n_2597;
input n_1016;
input n_1243;
input n_546;
input n_2959;
input n_101;
input n_3340;
input n_2047;
input n_1280;
input n_3277;
input n_3782;
input n_1845;
input n_281;
input n_240;
input n_2052;
input n_2193;
input n_2978;
input n_2058;
input n_2458;
input n_2478;
input n_3650;
input n_291;
input n_3786;
input n_231;
input n_257;
input n_2761;
input n_731;
input n_371;
input n_1483;
input n_2888;
input n_3638;
input n_1314;
input n_1512;
input n_3157;
input n_709;
input n_1490;
input n_317;
input n_1236;
input n_1633;
input n_2537;
input n_2983;
input n_3763;
input n_569;
input n_2669;
input n_2144;
input n_1778;
input n_3214;
input n_227;
input n_2306;
input n_920;
input n_2515;
input n_3022;
input n_3810;
input n_1289;
input n_1517;
input n_2091;
input n_2466;
input n_2635;
input n_2652;
input n_94;
input n_335;
input n_3631;
input n_2715;
input n_3806;
input n_3087;
input n_2085;
input n_3489;
input n_1669;
input n_2566;
input n_370;
input n_976;
input n_1949;
input n_343;
input n_1449;
input n_308;
input n_1946;
input n_2936;
input n_1566;
input n_2032;
input n_297;
input n_2587;
input n_156;
input n_2149;
input n_1078;
input n_2782;
input n_1670;
input n_2672;
input n_775;
input n_219;
input n_3060;
input n_157;
input n_2651;
input n_3947;
input n_3490;
input n_3656;
input n_600;
input n_1484;
input n_2071;
input n_2561;
input n_1374;
input n_1328;
input n_2643;
input n_223;
input n_2141;
input n_1948;
input n_3013;
input n_3183;
input n_1984;
input n_3437;
input n_3868;
input n_2099;
input n_2408;
input n_3446;
input n_3353;
input n_264;
input n_1877;
input n_3687;
input n_1831;
input n_1598;
input n_3049;
input n_1723;
input n_955;
input n_1850;
input n_163;
input n_3028;
input n_339;
input n_1146;
input n_882;
input n_183;
input n_243;
input n_2384;
input n_1036;
input n_1097;
input n_1749;
input n_347;
input n_3156;
input n_59;
input n_550;
input n_696;
input n_3101;
input n_3669;
input n_897;
input n_215;
input n_350;
input n_196;
input n_798;
input n_3376;
input n_646;
input n_1428;
input n_2663;
input n_436;
input n_1394;
input n_2659;
input n_3653;
input n_1414;
input n_1216;
input n_290;
input n_580;
input n_2693;
input n_3798;
input n_3702;
input n_1040;
input n_4065;
input n_3836;
input n_2202;
input n_2648;
input n_3963;
input n_1872;
input n_3389;
input n_1852;
input n_2159;
input n_578;
input n_2976;
input n_3876;
input n_926;
input n_2180;
input n_2249;
input n_344;
input n_2353;
input n_1218;
input n_1931;
input n_2439;
input n_2632;
input n_2276;
input n_3089;
input n_422;
input n_475;
input n_777;
input n_1070;
input n_1547;
input n_2089;
input n_3420;
input n_1030;
input n_72;
input n_2470;
input n_1755;
input n_3222;
input n_415;
input n_1071;
input n_485;
input n_1165;
input n_1267;
input n_1561;
input n_496;
input n_1801;
input n_3985;
input n_1391;
input n_958;
input n_1034;
input n_670;
input n_1513;
input n_2908;
input n_2970;
input n_3361;
input n_1600;
input n_48;
input n_521;
input n_3744;
input n_663;
input n_845;
input n_2235;
input n_1862;
input n_673;
input n_837;
input n_3980;
input n_1239;
input n_2915;
input n_528;
input n_2300;
input n_2791;
input n_1796;
input n_2551;
input n_3291;
input n_680;
input n_1473;
input n_1587;
input n_2682;
input n_395;
input n_164;
input n_553;
input n_901;
input n_3755;
input n_2432;
input n_3668;
input n_813;
input n_1521;
input n_1284;
input n_1590;
input n_3440;
input n_3405;
input n_214;
input n_2174;
input n_2714;
input n_1748;
input n_3563;
input n_2934;
input n_1672;
input n_2506;
input n_675;
input n_2699;
input n_4064;
input n_888;
input n_1880;
input n_2769;
input n_3542;
input n_2337;
input n_3436;
input n_1167;
input n_1626;
input n_3550;
input n_637;
input n_2615;
input n_3940;
input n_1384;
input n_1556;
input n_184;
input n_446;
input n_3907;
input n_1863;
input n_1064;
input n_144;
input n_858;
input n_2079;
input n_3841;
input n_2238;
input n_114;
input n_96;
input n_923;
input n_2118;
input n_691;
input n_1151;
input n_2985;
input n_2944;
input n_881;
input n_1405;
input n_2407;
input n_1706;
input n_468;
input n_3418;
input n_213;
input n_129;
input n_342;
input n_2932;
input n_2753;
input n_464;
input n_2980;
input n_363;
input n_1582;
input n_197;
input n_3637;
input n_1069;
input n_3306;
input n_1784;
input n_2859;
input n_2842;
input n_1075;
input n_3262;
input n_3136;
input n_1836;
input n_2868;
input n_3395;
input n_1450;
input n_4080;
input n_4006;
input n_3141;
input n_1322;
input n_2101;
input n_1471;
input n_1986;
input n_2863;
input n_2072;
input n_3164;
input n_2738;
input n_1750;
input n_3570;
input n_3690;
input n_1459;
input n_460;
input n_889;
input n_2358;
input n_973;
input n_3986;
input n_3716;
input n_4025;
input n_2968;
input n_1700;
input n_2833;
input n_477;
input n_3191;
input n_571;
input n_1585;
input n_461;
input n_2684;
input n_2712;
input n_3593;
input n_3193;
input n_3837;
input n_3885;
input n_1971;
input n_1599;
input n_3936;
input n_3252;
input n_2275;
input n_2855;
input n_3507;
input n_3273;
input n_3821;
input n_2713;
input n_3544;
input n_2644;
input n_2700;
input n_1211;
input n_1197;
input n_3367;
input n_4020;
input n_2951;
input n_1523;
input n_2730;
input n_1950;
input n_3008;
input n_3709;
input n_907;
input n_1447;
input n_2251;
input n_3096;
input n_1377;
input n_3915;
input n_2370;
input n_190;
input n_3496;
input n_3954;
input n_989;
input n_2544;
input n_1039;
input n_2214;
input n_3339;
input n_34;
input n_2055;
input n_3427;
input n_228;
input n_283;
input n_3025;
input n_3349;
input n_1403;
input n_3735;
input n_4067;
input n_2248;
input n_4042;
input n_2356;
input n_488;
input n_736;
input n_892;
input n_3320;
input n_3007;
input n_2688;
input n_1000;
input n_1202;
input n_2750;
input n_3899;
input n_2620;
input n_1278;
input n_2622;
input n_2062;
input n_2668;
input n_3714;
input n_1002;
input n_1463;
input n_1581;
input n_2100;
input n_49;
input n_3071;
input n_3739;
input n_4089;
input n_3651;
input n_310;
input n_3310;
input n_54;
input n_593;
input n_3487;
input n_2258;
input n_4069;
input n_12;
input n_748;
input n_586;
input n_1058;
input n_1667;
input n_3359;
input n_838;
input n_2784;
input n_3718;
input n_3983;
input n_2919;
input n_332;
input n_3092;
input n_1053;
input n_3470;
input n_1224;
input n_2865;
input n_349;
input n_2557;
input n_1926;
input n_2706;
input n_1248;
input n_230;
input n_1331;
input n_953;
input n_279;
input n_1014;
input n_1241;
input n_3676;
input n_70;
input n_2150;
input n_3146;
input n_2241;
input n_2757;
input n_3789;
input n_2152;
input n_3598;
input n_289;
input n_963;
input n_1052;
input n_954;
input n_627;
input n_3781;
input n_1385;
input n_440;
input n_793;
input n_478;
input n_2590;
input n_2776;
input n_2140;
input n_2385;
input n_3580;
input n_1819;
input n_2330;
input n_2139;
input n_2942;
input n_476;
input n_2987;
input n_1527;
input n_2042;
input n_534;
input n_3106;
input n_1882;
input n_884;
input n_3328;
input n_345;
input n_944;
input n_1754;
input n_3889;
input n_3611;
input n_1623;
input n_2862;
input n_2175;
input n_2921;
input n_2720;
input n_2324;
input n_1854;
input n_91;
input n_2606;
input n_2674;
input n_3187;
input n_1565;
input n_4088;
input n_3508;
input n_2828;
input n_3682;
input n_3371;
input n_1809;
input n_1856;
input n_182;
input n_143;
input n_647;
input n_3433;
input n_237;
input n_4024;
input n_407;
input n_1072;
input n_2218;
input n_2267;
input n_832;
input n_857;
input n_2305;
input n_3392;
input n_3430;
input n_3975;
input n_2636;
input n_2450;
input n_3208;
input n_207;
input n_561;
input n_1319;
input n_2379;
input n_3331;
input n_3447;
input n_2616;
input n_2911;
input n_3992;
input n_3305;
input n_2154;
input n_1825;
input n_1951;
input n_1883;
input n_1906;
input n_2759;
input n_1712;
input n_1387;
input n_3528;
input n_3649;
input n_2262;
input n_2462;
input n_2514;
input n_1532;
input n_2322;
input n_2271;
input n_2625;
input n_18;
input n_3257;
input n_3625;
input n_1027;
input n_971;
input n_1156;
input n_117;
input n_326;
input n_794;
input n_404;
input n_2798;
input n_2331;
input n_2945;
input n_2293;
input n_686;
input n_3989;
input n_2837;
input n_847;
input n_3804;
input n_4051;
input n_1393;
input n_2319;
input n_596;
input n_1775;
input n_2979;
input n_3296;
input n_2028;
input n_1368;
input n_3481;
input n_2762;
input n_558;
input n_3655;
input n_2808;
input n_702;
input n_1276;
input n_3009;
input n_2548;
input n_822;
input n_1412;
input n_2676;
input n_1709;
input n_2679;
input n_3981;
input n_2108;
input n_3640;
input n_728;
input n_266;
input n_1162;
input n_272;
input n_1538;
input n_2930;
input n_1838;
input n_1199;
input n_1847;
input n_1779;
input n_2767;
input n_2777;
input n_2603;
input n_3514;
input n_3116;
input n_352;
input n_1884;
input n_2434;
input n_2660;
input n_53;
input n_3602;
input n_1038;
input n_2967;
input n_520;
input n_1369;
input n_3909;
input n_409;
input n_2611;
input n_1841;
input n_1660;
input n_887;
input n_1905;
input n_2553;
input n_154;
input n_3706;
input n_3207;
input n_2581;
input n_71;
input n_3944;
input n_2195;
input n_2529;
input n_3224;
input n_300;
input n_2698;
input n_3752;
input n_4090;
input n_809;
input n_3923;
input n_870;
input n_931;
input n_599;
input n_1711;
input n_1662;
input n_1891;
input n_1481;
input n_2626;
input n_3441;
input n_3042;
input n_1942;
input n_434;
input n_1978;
input n_1544;
input n_4001;
input n_2510;
input n_3047;
input n_3526;
input n_868;
input n_2454;
input n_639;
input n_2804;
input n_914;
input n_3659;
input n_2120;
input n_411;
input n_414;
input n_2546;
input n_1629;
input n_1293;
input n_2801;
input n_3120;
input n_965;
input n_1876;
input n_1743;
input n_4007;
input n_3790;
input n_4011;
input n_3491;
input n_935;
input n_121;
input n_1175;
input n_817;
input n_2763;
input n_360;
input n_36;
input n_1479;
input n_1810;
input n_2350;
input n_2813;
input n_64;
input n_2825;
input n_1888;
input n_2009;
input n_759;
input n_3643;
input n_3895;
input n_2222;
input n_1892;
input n_3510;
input n_28;
input n_3745;
input n_806;
input n_2990;
input n_1997;
input n_2667;
input n_1766;
input n_3218;
input n_3748;
input n_1477;
input n_3142;
input n_324;
input n_1635;
input n_1963;
input n_2226;
input n_1571;
input n_2891;
input n_3119;
input n_187;
input n_1189;
input n_2690;
input n_4028;
input n_103;
input n_4082;
input n_97;
input n_3370;
input n_11;
input n_2215;
input n_3479;
input n_4085;
input n_7;
input n_1259;
input n_4073;
input n_1690;
input n_3819;
input n_706;
input n_746;
input n_1649;
input n_3150;
input n_747;
input n_2064;
input n_52;
input n_784;
input n_3978;
input n_110;
input n_2449;
input n_3867;
input n_1733;
input n_1244;
input n_3500;
input n_2413;
input n_431;
input n_1194;
input n_1925;
input n_3660;
input n_2297;
input n_1815;
input n_3279;
input n_2621;
input n_615;
input n_851;
input n_1759;
input n_843;
input n_1788;
input n_2177;
input n_2491;
input n_3747;
input n_523;
input n_913;
input n_1537;
input n_705;
input n_3833;
input n_865;
input n_61;
input n_2227;
input n_3775;
input n_678;
input n_2671;
input n_697;
input n_127;
input n_1222;
input n_75;
input n_1679;
input n_2190;
input n_3346;
input n_776;
input n_1798;
input n_2022;
input n_3814;
input n_1790;
input n_2518;
input n_2876;
input n_1415;
input n_367;
input n_2629;
input n_2592;
input n_3416;
input n_452;
input n_525;
input n_3484;
input n_3620;
input n_1260;
input n_1746;
input n_1647;
input n_2181;
input n_2479;
input n_2838;
input n_1829;
input n_1464;
input n_3133;
input n_3513;
input n_649;
input n_547;
input n_2563;
input n_43;
input n_1444;
input n_4030;
input n_1191;
input n_2387;
input n_2992;
input n_1674;
input n_3725;
input n_1833;
input n_116;
input n_3138;
input n_1830;
input n_2517;
input n_2073;
input n_1710;
input n_284;
input n_1128;
input n_2928;
input n_3128;
input n_139;
input n_1734;
input n_3038;
input n_744;
input n_590;
input n_629;
input n_3770;
input n_4014;
input n_2631;
input n_1308;
input n_2871;
input n_2178;
input n_3068;
input n_1767;
input n_3144;
input n_2943;
input n_2913;
input n_2336;
input n_3143;
input n_3168;
input n_254;
input n_1680;
input n_1233;
input n_3469;
input n_2607;
input n_3994;
input n_23;
input n_1615;
input n_1529;
input n_2005;
input n_526;
input n_1916;
input n_3317;
input n_293;
input n_372;
input n_677;
input n_244;
input n_47;
input n_1333;
input n_2469;
input n_1121;
input n_2723;
input n_3355;
input n_314;
input n_368;
input n_433;
input n_604;
input n_2007;
input n_8;
input n_3220;
input n_949;
input n_2539;
input n_3917;
input n_3942;
input n_3263;
input n_100;
input n_2582;
input n_1443;
input n_1008;
input n_3855;
input n_946;
input n_1539;
input n_2736;
input n_1001;
input n_1503;
input n_2054;
input n_3765;
input n_498;
input n_1468;
input n_1559;
input n_3823;
input n_1765;
input n_3455;
input n_1866;
input n_689;
input n_3158;
input n_738;
input n_1624;
input n_3000;
input n_640;
input n_3452;
input n_1510;
input n_252;
input n_624;
input n_1380;
input n_1744;
input n_2623;
input n_1617;
input n_295;
input n_133;
input n_1010;
input n_1994;
input n_1231;
input n_739;
input n_1279;
input n_1406;
input n_3108;
input n_3113;
input n_3111;
input n_2718;
input n_1195;
input n_1837;
input n_1839;
input n_610;
input n_2577;
input n_3760;
input n_4078;
input n_1760;
input n_2875;
input n_936;
input n_568;
input n_1500;
input n_2960;
input n_39;
input n_1090;
input n_2796;
input n_757;
input n_3844;
input n_3280;
input n_2342;
input n_633;
input n_2856;
input n_4054;
input n_439;
input n_3471;
input n_106;
input n_1832;
input n_259;
input n_448;
input n_1851;
input n_758;
input n_999;
input n_3205;
input n_2046;
input n_2848;
input n_2741;
input n_2937;
input n_3666;
input n_3003;
input n_3610;
input n_1933;
input n_3828;
input n_2290;
input n_93;
input n_1656;
input n_3564;
input n_3288;
input n_1158;
input n_3095;
input n_2045;
input n_3369;
input n_3783;
input n_3988;
input n_1509;
input n_1874;
input n_2040;
input n_563;
input n_2060;
input n_3199;
input n_2613;
input n_1987;
input n_2805;
input n_3667;
input n_1145;
input n_878;
input n_524;
input n_3843;
input n_3457;
input n_204;
input n_394;
input n_1678;
input n_1049;
input n_1153;
input n_3856;
input n_2145;
input n_741;
input n_1639;
input n_1306;
input n_3703;
input n_1068;
input n_3030;
input n_3558;
input n_1871;
input n_2580;
input n_3630;
input n_2545;
input n_2787;
input n_3685;
input n_2914;
input n_1964;
input n_2869;
input n_122;
input n_4002;
input n_331;
input n_10;
input n_906;
input n_1163;
input n_3271;
input n_2039;
input n_1207;
input n_919;
input n_908;
input n_4086;
input n_2412;
input n_2406;
input n_3623;
input n_90;
input n_2846;
input n_724;
input n_3753;
input n_1781;
input n_2084;
input n_2925;
input n_3648;
input n_2035;
input n_658;
input n_2061;
input n_3773;
input n_3555;
input n_3579;
input n_3918;
input n_3075;
input n_3173;
input n_2378;
input n_2509;
input n_1740;
input n_3236;
input n_2398;
input n_1362;
input n_3969;
input n_2857;
input n_3932;
input n_1586;
input n_456;
input n_959;
input n_2459;
input n_3031;
input n_535;
input n_152;
input n_3396;
input n_3701;
input n_940;
input n_1445;
input n_9;
input n_3516;
input n_4023;
input n_1492;
input n_2155;
input n_2516;
input n_3797;
input n_1923;
input n_1773;
input n_592;
input n_3243;
input n_1169;
input n_45;
input n_1596;
input n_1692;
input n_2666;
input n_2982;
input n_3385;
input n_1017;
input n_2481;
input n_2947;
input n_3545;
input n_2171;
input n_123;
input n_978;
input n_2768;
input n_2116;
input n_2314;
input n_1434;
input n_1054;
input n_2507;
input n_1474;
input n_1665;
input n_1269;
input n_4019;
input n_2420;
input n_2900;
input n_1095;
input n_3343;
input n_3515;
input n_1828;
input n_1614;
input n_2886;
input n_267;
input n_514;
input n_457;
input n_1079;
input n_1045;
input n_1208;
input n_2093;
input n_2038;
input n_2320;
input n_2339;
input n_2473;
input n_3287;
input n_2137;
input n_3378;
input n_603;
input n_1431;
input n_2583;
input n_484;
input n_1593;
input n_1033;
input n_3767;
input n_442;
input n_3426;
input n_3454;
input n_2299;
input n_131;
input n_2540;
input n_2873;
input n_3820;
input n_636;
input n_3741;
input n_660;
input n_3410;
input n_2087;
input n_1640;
input n_2162;
input n_1732;
input n_1009;
input n_2847;
input n_1148;
input n_2051;
input n_109;
input n_742;
input n_750;
input n_2029;
input n_995;
input n_454;
input n_3221;
input n_2168;
input n_2790;
input n_1609;
input n_374;
input n_3629;
input n_3021;
input n_1989;
input n_3818;
input n_185;
input n_2359;
input n_2941;
input n_3674;
input n_396;
input n_1887;
input n_3502;
input n_2523;
input n_1383;
input n_3098;
input n_1073;
input n_255;
input n_2346;
input n_2457;
input n_662;
input n_459;
input n_2312;
input n_3990;
input n_218;
input n_962;
input n_3475;
input n_1215;
input n_3015;
input n_1171;
input n_1578;
input n_723;
input n_1920;
input n_1065;
input n_1592;
input n_2536;
input n_1336;
input n_2882;
input n_3719;
input n_1721;
input n_1959;
input n_1758;
input n_2338;
input n_3681;
input n_2952;
input n_2737;
input n_1574;
input n_3672;
input n_2399;
input n_3058;
input n_2812;
input n_473;
input n_2048;
input n_3197;
input n_3109;
input n_3607;
input n_2355;
input n_2133;
input n_1921;
input n_2721;
input n_1309;
input n_1878;
input n_1426;
input n_3830;
input n_1043;
input n_2585;
input n_355;
input n_3505;
input n_486;
input n_3002;
input n_1800;
input n_1548;
input n_2725;
input n_614;
input n_337;
input n_1421;
input n_88;
input n_2571;
input n_1286;
input n_3730;
input n_3883;
input n_1177;
input n_3276;
input n_1355;
input n_168;
input n_974;
input n_2565;
input n_727;
input n_3897;
input n_1159;
input n_3845;
input n_957;
input n_3787;
input n_773;
input n_208;
input n_142;
input n_2124;
input n_743;
input n_3001;
input n_2081;
input n_299;
input n_303;
input n_3945;
input n_3149;
input n_296;
input n_613;
input n_1119;
input n_2156;
input n_1240;
input n_2261;
input n_1820;
input n_2729;
input n_3268;
input n_3597;
input n_2418;
input n_3827;
input n_65;
input n_829;
input n_2519;
input n_3354;
input n_2724;
input n_1612;
input n_2179;
input n_1416;
input n_2077;
input n_2897;
input n_3614;
input n_2909;
input n_1724;
input n_2111;
input n_2521;
input n_3301;
input n_361;
input n_3466;
input n_3458;
input n_700;
input n_1237;
input n_573;
input n_69;
input n_1420;
input n_3185;
input n_1132;
input n_3330;
input n_388;
input n_1366;
input n_1300;
input n_3960;
input n_2595;
input n_1127;
input n_3248;
input n_2277;
input n_761;
input n_2477;
input n_3523;
input n_1785;
input n_1568;
input n_2829;
input n_3905;
input n_1006;
input n_3411;
input n_3887;
input n_4087;
input n_2110;
input n_329;
input n_3811;
input n_274;
input n_4093;
input n_1270;
input n_1664;
input n_3200;
input n_1486;
input n_582;
input n_3586;
input n_1332;
input n_3519;
input n_2231;
input n_1390;
input n_2017;
input n_73;
input n_2474;
input n_2879;
input n_2604;
input n_19;
input n_2090;
input n_3374;
input n_3153;
input n_3045;
input n_1870;
input n_309;
input n_30;
input n_512;
input n_2367;
input n_1591;
input n_2033;
input n_4071;
input n_84;
input n_3453;
input n_130;
input n_322;
input n_1682;
input n_1980;
input n_2390;
input n_2628;
input n_1249;
input n_3399;
input n_2896;
input n_652;
input n_1111;
input n_3213;
input n_1365;
input n_4074;
input n_1927;
input n_25;
input n_3065;
input n_2132;
input n_1349;
input n_1093;
input n_288;
input n_2400;
input n_1031;
input n_3645;
input n_263;
input n_609;
input n_1041;
input n_1265;
input n_3223;
input n_1909;
input n_3838;
input n_44;
input n_224;
input n_3077;
input n_3929;
input n_2681;
input n_1562;
input n_383;
input n_3103;
input n_834;
input n_3474;
input n_112;
input n_765;
input n_3675;
input n_2255;
input n_2424;
input n_2272;
input n_893;
input n_3984;
input n_1015;
input n_1140;
input n_891;
input n_1651;
input n_1965;
input n_239;
input n_3387;
input n_630;
input n_1902;
input n_2151;
input n_1941;
input n_55;
input n_2106;
input n_2775;
input n_2716;
input n_3938;
input n_1913;
input n_2878;
input n_504;
input n_1823;
input n_511;
input n_3679;
input n_3779;
input n_874;
input n_2464;
input n_358;
input n_3422;
input n_3888;
input n_1101;
input n_2831;
input n_77;
input n_102;
input n_1106;
input n_1456;
input n_3557;
input n_2230;
input n_3498;
input n_2015;
input n_2365;
input n_1875;
input n_1982;
input n_1304;
input n_2803;
input n_1324;
input n_2851;
input n_3707;
input n_987;
input n_3189;
input n_1846;
input n_3037;
input n_261;
input n_174;
input n_2066;
input n_1885;
input n_1455;
input n_3429;
input n_767;
input n_993;
input n_1903;
input n_2490;
input n_1407;
input n_3849;
input n_3946;
input n_2452;
input n_1551;
input n_3154;
input n_545;
input n_441;
input n_860;
input n_3229;
input n_450;
input n_2849;
input n_1805;
input n_3925;
input n_2176;
input n_2204;
input n_2905;
input n_1816;
input n_3692;
input n_429;
input n_948;
input n_3965;
input n_3566;
input n_1217;
input n_2220;
input n_4059;
input n_2455;
input n_628;
input n_365;
input n_1849;
input n_3788;
input n_4084;
input n_2410;
input n_729;
input n_1131;
input n_1084;
input n_1961;
input n_970;
input n_4037;
input n_1935;
input n_911;
input n_2922;
input n_1430;
input n_83;
input n_3275;
input n_3499;
input n_2645;
input n_2467;
input n_513;
input n_3366;
input n_2727;
input n_1094;
input n_1354;
input n_560;
input n_1534;
input n_340;
input n_2288;
input n_3421;
input n_1351;
input n_2240;
input n_2696;
input n_4063;
input n_1044;
input n_1205;
input n_2436;
input n_346;
input n_1209;
input n_3029;
input n_1552;
input n_2508;
input n_3242;
input n_3592;
input n_3618;
input n_4031;
input n_495;
input n_602;
input n_3525;
input n_574;
input n_2593;
input n_3486;
input n_1435;
input n_879;
input n_3394;
input n_3793;
input n_16;
input n_3683;
input n_2416;
input n_58;
input n_2405;
input n_3642;
input n_623;
input n_3995;
input n_3286;
input n_2088;
input n_405;
input n_2953;
input n_3808;
input n_824;
input n_4036;
input n_359;
input n_1645;
input n_3881;
input n_4041;
input n_2461;
input n_490;
input n_1327;
input n_2858;
input n_2243;
input n_4060;
input n_996;
input n_921;
input n_1684;
input n_233;
input n_2658;
input n_3590;
input n_1717;
input n_572;
input n_366;
input n_2895;
input n_815;
input n_1795;
input n_2128;
input n_2578;
input n_3097;
input n_3483;
input n_128;
input n_1821;
input n_3894;
input n_120;
input n_2929;
input n_3424;
input n_327;
input n_3478;
input n_135;
input n_1381;
input n_2555;
input n_3751;
input n_2662;
input n_2740;
input n_3824;
input n_3890;
input n_1611;
input n_1037;
input n_2368;
input n_3388;
input n_2656;
input n_1080;
input n_2301;
input n_1274;
input n_3583;
input n_2890;
input n_3560;
input n_3059;
input n_3524;
input n_4076;
input n_2554;
input n_3465;
input n_1316;
input n_1708;
input n_2419;
input n_3215;
input n_426;
input n_1438;
input n_3698;
input n_3927;
input n_1082;
input n_1840;
input n_589;
input n_3961;
input n_716;
input n_1630;
input n_2122;
input n_2512;
input n_3589;
input n_562;
input n_1436;
input n_62;
input n_3549;
input n_1691;
input n_952;
input n_2786;
input n_2534;
input n_2092;
input n_3171;
input n_1229;
input n_391;
input n_701;
input n_1437;
input n_1023;
input n_2075;
input n_645;
input n_539;
input n_3658;
input n_3449;
input n_803;
input n_1092;
input n_2694;
input n_238;
input n_1776;
input n_3559;
input n_2198;
input n_2610;
input n_2661;
input n_2572;
input n_2989;
input n_2281;
input n_2131;
input n_2789;
input n_3026;
input n_3993;
input n_2216;
input n_531;
input n_3020;
input n_3677;
input n_1757;
input n_890;
input n_1897;
input n_764;
input n_1919;
input n_1056;
input n_1424;
input n_162;
input n_960;
input n_3462;
input n_3588;
input n_2933;
input n_2308;
input n_3468;
input n_1893;
input n_2910;
input n_222;
input n_3419;
input n_3886;
input n_1290;
input n_1123;
input n_1467;
input n_1047;
input n_2053;
input n_2163;
input n_634;
input n_2328;
input n_199;
input n_1958;
input n_32;
input n_2254;
input n_1252;
input n_348;
input n_3860;
input n_1382;
input n_1029;
input n_925;
input n_3546;
input n_1206;
input n_424;
input n_2647;
input n_3784;
input n_3160;
input n_1311;
input n_2191;
input n_2864;
input n_2969;
input n_3941;
input n_3195;
input n_1519;
input n_256;
input n_950;
input n_3190;
input n_2428;
input n_1553;
input n_3678;
input n_3847;
input n_2664;
input n_1811;
input n_2443;
input n_2624;
input n_3012;
input n_3456;
input n_380;
input n_419;
input n_1346;
input n_3053;
input n_444;
input n_1299;
input n_3244;
input n_2158;
input n_1808;
input n_3893;
input n_3290;
input n_1060;
input n_1141;
input n_316;
input n_2266;
input n_389;
input n_3130;
input n_2465;
input n_2824;
input n_3033;
input n_2650;
input n_3298;
input n_418;
input n_248;
input n_136;
input n_86;
input n_146;
input n_912;
input n_315;
input n_968;
input n_3548;
input n_451;
input n_619;
input n_408;
input n_2440;
input n_1386;
input n_1699;
input n_376;
input n_3334;
input n_967;
input n_1442;
input n_2923;
input n_3665;
input n_3494;
input n_2541;
input n_74;
input n_1139;
input n_2731;
input n_3264;
input n_515;
input n_2333;
input n_57;
input n_351;
input n_3953;
input n_885;
input n_2916;
input n_3166;
input n_397;
input n_1432;
input n_3875;
input n_3976;
input n_1357;
input n_483;
input n_2125;
input n_3771;
input n_3979;
input n_683;
input n_1632;
input n_3110;
input n_2998;
input n_1057;
input n_1051;
input n_1085;
input n_1066;
input n_4003;
input n_3800;
input n_721;
input n_2402;
input n_1157;
input n_3073;
input n_2403;
input n_841;
input n_1050;
input n_22;
input n_802;
input n_1954;
input n_4048;
input n_4026;
input n_2265;
input n_46;
input n_3162;
input n_1608;
input n_983;
input n_1844;
input n_2760;
input n_2792;
input n_3554;
input n_38;
input n_3377;
input n_2870;
input n_3777;
input n_280;
input n_1305;
input n_3749;
input n_3178;
input n_873;
input n_1826;
input n_3962;
input n_3991;
input n_378;
input n_1112;
input n_3134;
input n_2304;
input n_2999;
input n_762;
input n_1283;
input n_1644;
input n_17;
input n_2334;
input n_2637;
input n_3695;
input n_690;
input n_33;
input n_4046;
input n_1974;
input n_2463;
input n_583;
input n_2086;
input n_3537;
input n_2289;
input n_3080;
input n_3051;
input n_302;
input n_4096;
input n_1343;
input n_2701;
input n_2783;
input n_2263;
input n_3362;
input n_2881;
input n_1203;
input n_1631;
input n_3750;
input n_3282;
input n_2472;
input n_821;
input n_3816;
input n_1763;
input n_2341;
input n_3105;
input n_3231;
input n_1966;
input n_3632;
input n_1768;
input n_321;
input n_2294;
input n_1179;
input n_621;
input n_753;
input n_2475;
input n_2733;
input n_455;
input n_1048;
input n_1719;
input n_2993;
input n_3864;
input n_1288;
input n_212;
input n_385;
input n_2785;
input n_2556;
input n_507;
input n_2269;
input n_2732;
input n_3569;
input n_2309;
input n_2415;
input n_2948;
input n_3274;
input n_3041;
input n_3299;
input n_2646;
input n_1560;
input n_3715;
input n_1605;
input n_2236;
input n_330;
input n_1228;
input n_2816;
input n_2123;
input n_3209;
input n_972;
input n_3504;
input n_692;
input n_2037;
input n_2685;
input n_3920;
input n_3040;
input n_1953;
input n_1938;
input n_820;
input n_1200;
input n_2499;
input n_1911;
input n_3616;
input n_2460;
input n_4058;
input n_3568;
input n_3664;
input n_2589;
input n_3203;
input n_1301;
input n_1363;
input n_1668;
input n_3737;
input n_3913;
input n_1185;
input n_991;
input n_2903;
input n_3417;
input n_3482;
input n_3866;
input n_828;
input n_1967;
input n_779;
input n_576;
input n_1143;
input n_1579;
input n_2233;
input n_3717;
input n_4034;
input n_1329;
input n_2743;
input n_2675;
input n_3255;
input n_1312;
input n_1439;
input n_804;
input n_537;
input n_2827;
input n_1688;
input n_3052;
input n_945;
input n_2997;
input n_492;
input n_3743;
input n_3327;
input n_153;
input n_1504;
input n_943;
input n_3326;
input n_3956;
input n_341;
input n_3572;
input n_250;
input n_992;
input n_3067;
input n_1932;
input n_3375;
input n_2755;
input n_4047;
input n_543;
input n_260;
input n_842;
input n_3734;
input n_650;
input n_984;
input n_694;
input n_3237;
input n_2082;
input n_286;
input n_1992;
input n_2429;
input n_1643;
input n_883;
input n_1983;
input n_3167;
input n_4029;
input n_3400;
input n_470;
input n_325;
input n_449;
input n_1594;
input n_132;
input n_1214;
input n_1342;
input n_1400;
input n_3423;
input n_900;
input n_2362;
input n_856;
input n_2609;
input n_3870;
input n_1793;
input n_3382;
input n_1976;
input n_2223;
input n_3044;
input n_3574;
input n_918;
input n_3529;
input n_3854;
input n_942;
input n_2169;
input n_1804;
input n_189;
input n_1147;
input n_1557;
input n_1977;
input n_2153;
input n_2468;
input n_1610;
input n_13;
input n_1077;
input n_1422;
input n_3196;
input n_4095;
input n_3078;
input n_2364;
input n_2533;
input n_540;
input n_3492;
input n_618;
input n_3094;
input n_896;
input n_2310;
input n_2780;
input n_323;
input n_3952;
input n_2287;
input n_2860;
input n_3316;
input n_195;
input n_356;
input n_2291;
input n_3099;
input n_4043;
input n_3704;
input n_2596;
input n_894;
input n_1636;
input n_2056;
input n_3253;
input n_1730;
input n_3601;
input n_3603;
input n_4027;
input n_831;
input n_2280;
input n_2192;
input n_964;
input n_3633;
input n_3363;
input n_1373;
input n_1350;
input n_1511;
input n_1865;
input n_2973;
input n_1470;
input n_1096;
input n_2094;
input n_2670;
input n_234;
input n_1575;
input n_1697;
input n_1735;
input n_833;
input n_2318;
input n_2393;
input n_3689;
input n_2020;
input n_3831;
input n_5;
input n_1646;
input n_2502;
input n_3801;
input n_225;
input n_2504;
input n_1307;
input n_1881;
input n_2974;
input n_988;
input n_2749;
input n_2043;
input n_2901;
input n_1940;
input n_814;
input n_2707;
input n_2751;
input n_2793;
input n_3372;
input n_3451;
input n_192;
input n_2971;
input n_3442;
input n_1549;
input n_1934;
input n_2311;
input n_1201;
input n_1114;
input n_3950;
input n_4000;
input n_655;
input n_3240;
input n_2025;
input n_1616;
input n_3998;
input n_1446;
input n_2285;
input n_3147;
input n_2758;
input n_669;
input n_472;
input n_1458;
input n_1176;
input n_1472;
input n_2298;
input n_2471;
input n_1807;
input n_387;
input n_3869;
input n_1149;
input n_2618;
input n_398;
input n_1671;
input n_635;
input n_2559;
input n_763;
input n_3230;
input n_1020;
input n_1062;
input n_3342;
input n_211;
input n_2303;
input n_1824;
input n_1917;
input n_2295;
input n_1219;
input n_3386;
input n_3931;
input n_3;
input n_3708;
input n_1204;
input n_4010;
input n_2840;
input n_3729;
input n_2810;
input n_2325;
input n_178;
input n_2747;
input n_2446;
input n_3488;
input n_1814;
input n_1035;
input n_2822;
input n_3861;
input n_287;
input n_3780;
input n_555;
input n_783;
input n_1848;
input n_1928;
input n_2126;
input n_2893;
input n_3636;
input n_1188;
input n_2588;
input n_2962;
input n_4004;
input n_1722;
input n_3957;
input n_661;
input n_2441;
input n_3848;
input n_41;
input n_1802;
input n_3083;
input n_2600;
input n_3919;
input n_4079;
input n_3898;
input n_849;
input n_2795;
input n_15;
input n_4091;
input n_336;
input n_584;
input n_681;
input n_1638;
input n_1786;
input n_2981;
input n_50;
input n_430;
input n_2002;
input n_2282;
input n_3608;
input n_510;
input n_2800;
input n_216;
input n_3712;
input n_2371;
input n_2935;
input n_311;
input n_3233;
input n_3829;
input n_3380;
input n_3177;
input n_4053;
input n_830;
input n_2098;
input n_1296;
input n_2627;
input n_3409;
input n_3460;
input n_2352;
input n_3538;
input n_1413;
input n_801;
input n_4040;
input n_2207;
input n_2080;
input n_2377;
input n_2619;
input n_2340;
input n_3085;
input n_2444;
input n_2068;
input n_241;
input n_3552;
input n_875;
input n_357;
input n_1110;
input n_1655;
input n_445;
input n_2641;
input n_3198;
input n_749;
input n_1895;
input n_3123;
input n_3684;
input n_3137;
input n_2574;
input n_1134;
input n_1358;
input n_717;
input n_165;
input n_939;
input n_3697;
input n_482;
input n_2361;
input n_1088;
input n_588;
input n_1173;
input n_789;
input n_3393;
input n_1232;
input n_1603;
input n_734;
input n_638;
input n_2638;
input n_866;
input n_107;
input n_969;
input n_1401;
input n_4018;
input n_4044;
input n_3900;
input n_4062;
input n_3520;
input n_3971;
input n_2492;
input n_1019;
input n_1105;
input n_249;
input n_1998;
input n_304;
input n_3759;
input n_1338;
input n_577;
input n_4005;
input n_2016;
input n_1522;
input n_3872;
input n_2949;
input n_1687;
input n_1637;
input n_2034;
input n_1419;
input n_2711;
input n_3933;
input n_338;
input n_149;
input n_1653;
input n_693;
input n_2270;
input n_1506;
input n_3206;
input n_2653;
input n_3578;
input n_3966;
input n_14;
input n_836;
input n_990;
input n_2867;
input n_3812;
input n_2496;
input n_1886;
input n_1389;
input n_1894;
input n_975;
input n_1908;
input n_1256;
input n_1702;
input n_2259;
input n_2794;
input n_567;
input n_1465;
input n_3145;
input n_3124;
input n_778;
input n_1122;
input n_4068;
input n_151;
input n_3192;
input n_2608;
input n_3877;
input n_306;
input n_3764;
input n_2657;
input n_458;
input n_770;
input n_2995;
input n_1375;
input n_2494;
input n_3547;
input n_2649;
input n_3977;
input n_1102;
input n_3727;
input n_2852;
input n_3774;
input n_4052;
input n_2392;
input n_3459;
input n_3093;
input n_1843;
input n_711;
input n_1499;
input n_3061;
input n_3155;
input n_85;
input n_1187;
input n_3517;
input n_2633;
input n_1441;
input n_3100;
input n_2522;
input n_2435;
input n_1392;
input n_1597;
input n_1929;
input n_2807;
input n_1164;
input n_1659;
input n_1834;
input n_2097;
input n_2313;
input n_2542;
input n_489;
input n_1174;
input n_2431;
input n_3324;
input n_3356;
input n_3758;
input n_2835;
input n_3914;
input n_3911;
input n_2558;
input n_1371;
input n_617;
input n_1303;
input n_2206;
input n_2063;
input n_3803;
input n_3182;
input n_1572;
input n_1968;
input n_3742;
input n_3269;
input n_2564;
input n_2252;
input n_876;
input n_1516;
input n_3736;
input n_1190;
input n_3506;
input n_3896;
input n_1736;
input n_3605;
input n_1685;
input n_3958;
input n_118;
input n_2409;
input n_601;
input n_917;
input n_3450;
input n_1714;
input n_966;
input n_253;
input n_1116;
input n_2000;
input n_1661;
input n_3402;
input n_1212;
input n_2074;
input n_1541;
input n_2576;
input n_3565;
input n_172;
input n_206;
input n_217;
input n_726;
input n_3174;
input n_982;
input n_2575;
input n_2988;
input n_3390;
input n_1573;
input n_1453;
input n_1731;
input n_2217;
input n_3746;
input n_818;
input n_2373;
input n_1970;
input n_861;
input n_1713;
input n_1183;
input n_3398;
input n_2307;
input n_2766;
input n_3817;
input n_1658;
input n_899;
input n_1253;
input n_210;
input n_1737;
input n_2201;
input n_2722;
input n_2117;
input n_2745;
input n_3408;
input n_1904;
input n_2640;
input n_1993;
input n_774;
input n_3835;
input n_1628;
input n_2493;
input n_2205;
input n_3432;
input n_1335;
input n_1514;
input n_1777;
input n_1957;
input n_1059;
input n_1345;
input n_3967;
input n_176;
input n_1133;
input n_1771;
input n_1912;
input n_3401;
input n_1899;
input n_3226;
input n_557;
input n_1410;
input n_1005;
input n_607;
input n_1003;
input n_679;
input n_710;
input n_3090;
input n_2067;
input n_527;
input n_1168;
input n_707;
input n_2219;
input n_2437;
input n_2885;
input n_3762;
input n_3902;
input n_3533;
input n_2877;
input n_3318;
input n_4070;
input n_2148;
input n_937;
input n_2445;
input n_1427;
input n_2779;
input n_3485;
input n_393;
input n_108;
input n_487;
input n_1584;
input n_665;
input n_1726;
input n_1835;
input n_3035;
input n_3654;
input n_66;
input n_1440;
input n_177;
input n_3839;
input n_2164;
input n_421;
input n_1988;
input n_3333;
input n_2115;
input n_1853;
input n_1356;
input n_2845;
input n_1787;
input n_2634;
input n_910;
input n_2232;
input n_3034;
input n_2212;
input n_2602;
input n_1657;
input n_768;
input n_1475;
input n_1302;
input n_1774;
input n_1725;
input n_205;
input n_1136;
input n_1313;
input n_1491;
input n_754;
input n_3972;
input n_2811;
input n_1496;
input n_3348;
input n_179;
input n_1125;
input n_125;
input n_410;
input n_2547;
input n_3014;
input n_3639;
input n_708;
input n_529;
input n_1812;
input n_735;
input n_2501;
input n_3079;
input n_232;
input n_1915;
input n_1109;
input n_126;
input n_895;
input n_2532;
input n_1310;
input n_2605;
input n_3358;
input n_2121;
input n_1803;
input n_202;
input n_3791;
input n_3308;
input n_2665;
input n_427;
input n_1399;
input n_1543;
input n_1991;
input n_1979;
input n_791;
input n_732;
input n_1533;
input n_2224;
input n_193;
input n_3368;
input n_2924;
input n_3467;
input n_808;
input n_2484;
input n_797;
input n_3530;
input n_1025;
input n_1930;
input n_1955;
input n_3731;
input n_2765;
input n_3329;
input n_500;
input n_2994;
input n_1067;
input n_3805;
input n_3825;
input n_2946;
input n_1720;
input n_148;
input n_2830;
input n_2401;
input n_3135;
input n_435;
input n_3657;
input n_2003;
input n_159;
input n_766;
input n_1457;
input n_3928;
input n_541;
input n_2692;
input n_3573;
input n_3148;
input n_538;
input n_2354;
input n_2246;
input n_2008;
input n_1117;
input n_799;
input n_2264;
input n_2754;
input n_687;
input n_3534;
input n_715;
input n_3901;
input n_1742;
input n_1480;
input n_1482;
input n_1213;
input n_2489;
input n_1266;
input n_3970;
input n_3757;
input n_536;
input n_3438;
input n_872;
input n_2012;
input n_594;
input n_3792;
input n_200;
input n_1291;
input n_3974;
input n_3381;
input n_3871;
input n_4094;
input n_3503;
input n_1297;
input n_1753;
input n_2283;
input n_2866;
input n_3278;
input n_1782;
input n_2245;
input n_3561;
input n_1155;
input n_1418;
input n_89;
input n_1972;
input n_1524;
input n_1689;
input n_1485;
input n_2806;
input n_115;
input n_1011;
input n_1184;
input n_2184;
input n_985;
input n_1855;
input n_2425;
input n_2917;
input n_869;
input n_810;
input n_2965;
input n_3536;
input n_3661;
input n_416;
input n_3635;
input n_827;
input n_3217;
input n_3404;
input n_3425;
input n_401;
input n_1703;
input n_3312;
input n_4055;
input n_1352;
input n_2926;
input n_626;
input n_2197;
input n_2199;
input n_3540;
input n_1650;
input n_3670;
input n_1144;
input n_3973;
input n_1137;
input n_1570;
input n_2814;
input n_3046;
input n_3882;
input n_3934;
input n_1170;
input n_305;
input n_2023;
input n_2213;
input n_3826;
input n_3249;
input n_3211;
input n_3285;
input n_2351;
input n_2211;
input n_2095;
input n_3121;
input n_3922;
input n_137;
input n_3846;
input n_676;
input n_294;
input n_318;
input n_2103;
input n_653;
input n_3968;
input n_2160;
input n_642;
input n_3337;
input n_2228;
input n_2527;
input n_1602;
input n_2498;
input n_194;
input n_855;
input n_1178;
input n_1461;
input n_2697;
input n_850;
input n_684;
input n_3074;
input n_124;
input n_3204;
input n_268;
input n_2421;
input n_2286;
input n_2902;
input n_664;
input n_1999;
input n_503;
input n_2372;
input n_2065;
input n_2136;
input n_3673;
input n_2480;
input n_4017;
input n_235;
input n_3768;
input n_1372;
input n_2861;
input n_605;
input n_2630;
input n_1273;
input n_3943;
input n_1822;
input n_3397;
input n_353;
input n_3740;
input n_620;
input n_643;
input n_2363;
input n_2430;
input n_4072;
input n_916;
input n_1081;
input n_2549;
input n_493;
input n_2705;
input n_3005;
input n_2332;
input n_1235;
input n_703;
input n_698;
input n_980;
input n_1115;
input n_2433;
input n_3293;
input n_3129;
input n_1282;
input n_1318;
input n_1783;
input n_780;
input n_2977;
input n_3606;
input n_2601;
input n_3043;
input n_4022;
input n_998;
input n_3802;
input n_2375;
input n_2550;
input n_1454;
input n_3723;
input n_467;
input n_1227;
input n_1531;
input n_840;
input n_1334;
input n_1907;
input n_3600;
input n_501;
input n_823;
input n_245;
input n_2686;
input n_2528;
input n_725;
input n_2344;
input n_3892;
input n_1388;
input n_1417;
input n_1295;
input n_2836;
input n_4035;
input n_2316;
input n_672;
input n_1985;
input n_3055;
input n_1898;
input n_2107;
input n_3294;
input n_3219;
input n_3711;
input n_3315;
input n_581;
input n_2906;
input n_382;
input n_554;
input n_1625;
input n_2130;
input n_3415;
input n_2187;
input n_2284;
input n_898;
input n_2817;
input n_3172;
input n_3139;
input n_2773;
input n_3239;
input n_3292;
input n_2598;
input n_3878;
input n_1762;
input n_1013;
input n_3365;
input n_3476;
input n_3686;
input n_1452;
input n_718;
input n_2687;
input n_265;
input n_3023;
input n_3553;
input n_1120;
input n_719;
input n_443;
input n_1791;
input n_198;
input n_1890;
input n_1747;
input n_714;
input n_2850;
input n_1683;
input n_1817;
input n_909;
input n_1944;
input n_1497;
input n_1530;
input n_4075;
input n_3982;
input n_2654;
input n_997;
input n_3431;
input n_3104;
input n_932;
input n_3169;
input n_3151;
input n_612;
input n_3822;
input n_3131;
input n_2078;
input n_1409;
input n_3850;
input n_788;
input n_1326;
input n_3070;
input n_3284;
input n_4066;
input n_3647;
input n_119;
input n_3176;
input n_2884;
input n_1268;
input n_2996;
input n_559;
input n_825;
input n_2819;
input n_3126;
input n_1981;
input n_508;
input n_2186;
input n_506;
input n_1320;
input n_1663;
input n_737;
input n_1718;
input n_4050;
input n_3700;
input n_3609;
input n_986;
input n_2315;
input n_509;
input n_3228;
input n_1317;
input n_147;
input n_1518;
input n_1715;
input n_2102;
input n_3581;
input n_2562;
input n_1281;
input n_67;
input n_1952;
input n_4077;
input n_1192;
input n_2221;
input n_1024;
input n_3576;
input n_1063;
input n_3720;
input n_1889;
input n_209;
input n_1792;
input n_1564;
input n_1868;
input n_1613;
input n_733;
input n_1489;
input n_1922;
input n_2966;
input n_4049;
input n_1376;
input n_941;
input n_2326;
input n_981;
input n_2560;
input n_3862;
input n_1569;
input n_2188;
input n_68;
input n_3495;
input n_3879;
input n_867;
input n_186;
input n_2348;
input n_2422;
input n_3959;
input n_134;
input n_2239;
input n_587;
input n_2950;
input n_63;
input n_792;
input n_756;
input n_1429;
input n_399;
input n_1238;
input n_2448;
input n_3140;
input n_3852;
input n_548;
input n_3170;
input n_3724;
input n_812;
input n_298;
input n_2104;
input n_2748;
input n_3311;
input n_518;
input n_505;
input n_2057;
input n_3272;
input n_4008;
input n_3011;
input n_1772;
input n_282;
input n_752;
input n_905;
input n_1476;
input n_1108;
input n_2898;
input n_782;
input n_2717;
input n_2818;
input n_1100;
input n_3646;
input n_1861;
input n_2129;
input n_1395;
input n_3345;
input n_862;
input n_3584;
input n_1425;
input n_760;
input n_3858;
input n_1901;
input n_3069;
input n_3756;
input n_1900;
input n_1620;
input n_3032;
input n_381;
input n_3628;
input n_2889;
input n_3691;
input n_220;
input n_390;
input n_1330;
input n_1867;
input n_31;
input n_1945;
input n_2772;
input n_481;
input n_3018;
input n_1675;
input n_3072;
input n_1924;
input n_2573;
input n_3084;
input n_3081;
input n_3313;
input n_1727;
input n_2710;
input n_1554;
input n_2939;
input n_1745;
input n_3924;
input n_2735;
input n_769;
input n_2497;
input n_2006;
input n_3412;
input n_3999;
input n_42;
input n_2844;
input n_1995;
input n_2411;
input n_3807;
input n_2138;
input n_1046;
input n_271;
input n_934;
input n_1618;
input n_2260;
input n_826;
input n_2343;
input n_1813;
input n_2447;
input n_3761;
input n_886;
input n_3439;
input n_2014;
input n_3056;
input n_1221;
input n_2345;
input n_2986;
input n_654;
input n_1172;
input n_167;
input n_2535;
input n_379;
input n_428;
input n_1341;
input n_2726;
input n_570;
input n_2774;
input n_3295;
input n_1641;
input n_1361;
input n_3184;
input n_2382;
input n_1707;
input n_853;
input n_3062;
input n_3161;
input n_377;
input n_2317;
input n_751;
input n_3289;
input n_2799;
input n_2172;
input n_1973;
input n_786;
input n_1083;
input n_1142;
input n_2376;
input n_2488;
input n_1129;
input n_392;
input n_2579;
input n_3477;
input n_3017;
input n_158;
input n_3626;
input n_2476;
input n_704;
input n_787;
input n_1770;
input n_138;
input n_2781;
input n_2456;
input n_3904;
input n_961;
input n_2250;
input n_2678;
input n_1756;
input n_771;
input n_2778;
input n_276;
input n_95;
input n_1716;
input n_2788;
input n_2872;
input n_1225;
input n_2984;
input n_1520;
input n_2451;
input n_169;
input n_2887;
input n_522;
input n_3364;
input n_1287;
input n_1262;
input n_2691;
input n_400;
input n_930;
input n_181;
input n_4092;
input n_3908;
input n_1873;
input n_1411;
input n_3926;
input n_3201;
input n_3054;
input n_221;
input n_622;
input n_1962;
input n_3996;
input n_1577;
input n_2423;
input n_3671;
input n_1087;
input n_3472;
input n_2526;
input n_2854;
input n_386;
input n_994;
input n_1701;
input n_3344;
input n_2194;
input n_848;
input n_1550;
input n_2874;
input n_2764;
input n_2703;
input n_1498;
input n_2167;
input n_3302;
input n_3235;
input n_1223;
input n_1272;
input n_2680;
input n_3391;
input n_104;
input n_682;
input n_1567;
input n_56;
input n_141;
input n_2567;
input n_3949;
input n_3543;
input n_1247;
input n_2709;
input n_3102;
input n_922;
input n_3122;
input n_816;
input n_1648;
input n_4015;
input n_591;
input n_3842;
input n_145;
input n_1536;
input n_3050;
input n_3265;
input n_1857;
input n_4056;
input n_1344;
input n_2041;
input n_313;
input n_631;
input n_3627;
input n_479;
input n_1246;
input n_3840;
input n_1339;
input n_1478;
input n_1797;
input n_432;
input n_1769;
input n_2957;
input n_839;
input n_3551;
input n_3903;
input n_1210;
input n_3518;
input n_2964;
input n_3769;
input n_1364;
input n_2956;
input n_2357;
input n_3733;
input n_2183;
input n_2673;
input n_2742;
input n_3314;
input n_2360;
input n_3254;
input n_328;
input n_140;
input n_2292;
input n_1250;
input n_2173;
input n_3859;
input n_369;
input n_3722;
input n_3865;
input n_1842;
input n_871;
input n_2442;
input n_3309;
input n_3738;
input n_4045;
input n_598;
input n_685;
input n_928;
input n_608;
input n_1367;
input n_78;
input n_1943;
input n_3634;
input n_1460;
input n_772;
input n_2018;
input n_3464;
input n_3260;
input n_1555;
input n_3117;
input n_2834;
input n_3245;
input n_3357;
input n_499;
input n_2531;
input n_1589;
input n_517;
input n_3428;
input n_98;
input n_2961;
input n_402;
input n_413;
input n_1086;
input n_2570;
input n_2702;
input n_796;
input n_1858;
input n_3351;
input n_1619;
input n_3527;
input n_2815;
input n_236;
input n_2119;
input n_1502;
input n_2157;
input n_2552;
input n_3754;
input n_1469;
input n_1012;
input n_1;
input n_1396;
input n_2744;
input n_1348;
input n_2030;
input n_903;
input n_2453;
input n_1525;
input n_1752;
input n_2397;
input n_740;
input n_2883;
input n_3115;
input n_203;
input n_3509;
input n_3352;
input n_384;
input n_2208;
input n_3076;
input n_1404;
input n_80;
input n_3063;
input n_3617;
input n_2912;
input n_1794;
input n_3535;
input n_2182;
input n_35;
input n_1315;
input n_2234;
input n_277;
input n_1061;
input n_3251;
input n_92;
input n_1910;
input n_333;
input n_1298;
input n_3955;
input n_2931;
input n_1652;
input n_2209;
input n_3794;
input n_462;
input n_2050;
input n_2809;
input n_1193;
input n_2797;
input n_1676;
input n_1255;
input n_258;
input n_1113;
input n_3118;
input n_29;
input n_79;
input n_4039;
input n_3227;
input n_3300;
input n_2321;
input n_3511;
input n_1226;
input n_722;
input n_1277;
input n_3680;
input n_2591;
input n_3443;
input n_188;
input n_2146;
input n_844;
input n_201;
input n_3384;
input n_471;
input n_852;
input n_3497;
input n_1487;
input n_40;
input n_1864;
input n_3644;
input n_1028;
input n_1601;
input n_4016;
input n_3336;
input n_3935;
input n_781;
input n_474;
input n_2940;
input n_542;
input n_3435;
input n_3521;
input n_463;
input n_3575;
input n_1546;
input n_595;
input n_502;
input n_3562;
input n_3948;
input n_466;
input n_2612;
input n_420;
input n_1337;
input n_1495;
input n_632;
input n_699;
input n_979;
input n_1515;
input n_2841;
input n_3165;
input n_1627;
input n_2918;
input n_3232;
input n_3322;
input n_3652;
input n_1245;
input n_846;
input n_2427;
input n_2438;
input n_2505;
input n_1673;
input n_465;
input n_2832;
input n_76;
input n_362;
input n_1321;
input n_170;
input n_1975;
input n_27;
input n_2296;
input n_2070;
input n_161;
input n_273;
input n_1937;
input n_585;
input n_2112;
input n_3250;
input n_4083;
input n_1739;
input n_3181;
input n_270;
input n_2958;
input n_616;
input n_2278;
input n_81;
input n_2594;
input n_3114;
input n_3125;
input n_2394;
input n_3234;
input n_1914;
input n_3612;
input n_2954;
input n_2135;
input n_2335;
input n_2904;
input n_3493;
input n_745;
input n_2381;
input n_3303;
input n_1654;
input n_3004;
input n_3323;
input n_3916;
input n_2569;
input n_3112;
input n_2349;
input n_1103;
input n_3921;
input n_4081;
input n_3132;
input n_3556;
input n_648;
input n_1379;
input n_2734;
input n_3874;
input n_312;
input n_2196;
input n_3591;
input n_3951;
input n_3024;
input n_2170;
input n_1076;
input n_2823;
input n_1091;
input n_1408;
input n_3512;
input n_494;
input n_1761;
input n_641;
input n_3238;
input n_3210;
input n_3930;
input n_730;
input n_3175;
input n_3522;
input n_2036;
input n_1325;
input n_3267;
input n_1595;
input n_2161;
input n_354;
input n_575;
input n_480;
input n_425;
input n_795;
input n_2404;
input n_2083;
input n_695;
input n_180;
input n_3281;
input n_656;
input n_3307;
input n_1606;
input n_2503;
input n_1220;
input n_37;
input n_1694;
input n_1540;
input n_3964;
input n_3266;
input n_2485;
input n_3772;
input n_229;
input n_1936;
input n_1956;
input n_437;
input n_1642;
input n_2279;
input n_3373;
input n_2655;
input n_2027;
input n_3884;
input n_60;
input n_403;
input n_453;
input n_2642;
input n_1130;
input n_720;
input n_0;
input n_2500;
input n_2366;
input n_1918;
input n_1526;
input n_863;
input n_3726;
input n_2210;
input n_805;
input n_3247;
input n_3997;
input n_1604;
input n_1275;
input n_2513;
input n_2525;
input n_3091;
input n_2695;
input n_1764;
input n_3480;
input n_2892;
input n_4032;
input n_3057;
input n_3194;
input n_3582;
input n_3066;
input n_113;
input n_712;
input n_2414;
input n_2907;
input n_246;
input n_1583;
input n_2426;
input n_2826;
input n_3577;
input n_3539;
input n_1042;
input n_1402;
input n_2820;
input n_269;
input n_3662;
input n_2049;
input n_2273;
input n_285;
input n_412;
input n_2719;
input n_1493;
input n_657;
input n_644;
input n_1741;
input n_2229;
input n_1160;
input n_1397;
input n_4057;
input n_491;
input n_1258;
input n_1074;
input n_3347;
input n_2004;
input n_3216;
input n_1621;
input n_2708;
input n_3809;
input n_2113;
input n_251;
input n_160;
input n_566;
input n_565;
input n_2586;
input n_3694;
input n_1448;
input n_2225;
input n_3567;
input n_3613;
input n_1507;
input n_1398;
input n_2383;
input n_1879;
input n_597;
input n_1996;
input n_3406;
input n_3604;
input n_3444;
input n_3853;
input n_1181;
input n_1505;
input n_1634;
input n_3939;
input n_1196;
input n_4012;
input n_2019;
input n_651;
input n_1340;
input n_2274;
input n_2972;
input n_334;
input n_811;
input n_1558;
input n_3225;
input n_807;
input n_3321;
input n_2166;
input n_3910;
input n_2938;
input n_3212;
input n_835;
input n_175;
input n_666;
input n_3319;
input n_262;
input n_1433;
input n_3594;
input n_1704;
input n_2256;
input n_3152;
input n_3721;
input n_3335;
input n_99;
input n_1254;
input n_3799;
input n_1026;
input n_3413;
input n_2026;
input n_1969;
input n_1234;
input n_2109;
input n_319;
input n_364;
input n_1138;
input n_927;
input n_20;
input n_1089;
input n_2013;
input n_1990;
input n_2044;
input n_2689;
input n_2920;
input n_3259;
input n_1004;
input n_1186;
input n_1032;
input n_242;
input n_2614;
input n_2511;
input n_1681;
input n_2010;
input n_2991;
input n_3688;
input n_3383;
input n_1018;
input n_2242;
input n_2247;
input n_2752;
input n_2894;
input n_3016;
input n_1693;
input n_3585;
input n_2975;
input n_3473;
input n_438;
input n_2599;
input n_713;
input n_2704;
input n_904;
input n_2839;
input n_3338;
input n_1588;
input n_1622;
input n_2237;
input n_3414;
input n_3463;
input n_3699;
input n_166;
input n_1180;
input n_1827;
input n_3360;
input n_2524;
input n_3873;
input n_1271;
input n_3705;
input n_2802;
input n_533;
input n_1542;
input n_1251;
input n_3693;
input n_4009;
input n_3159;
input n_278;
input n_2728;
input n_3857;
input n_2268;
input n_3778;

output n_16249;

wire n_13115;
wire n_6643;
wire n_6122;
wire n_10564;
wire n_13903;
wire n_7981;
wire n_9936;
wire n_5567;
wire n_4706;
wire n_12148;
wire n_15472;
wire n_14870;
wire n_15741;
wire n_9194;
wire n_15969;
wire n_12407;
wire n_6579;
wire n_15974;
wire n_9325;
wire n_7164;
wire n_10794;
wire n_6546;
wire n_5287;
wire n_12872;
wire n_13683;
wire n_14881;
wire n_15306;
wire n_9655;
wire n_15349;
wire n_14101;
wire n_15948;
wire n_5484;
wire n_10515;
wire n_11207;
wire n_11326;
wire n_5978;
wire n_8174;
wire n_5161;
wire n_15269;
wire n_5776;
wire n_14036;
wire n_13241;
wire n_6551;
wire n_13217;
wire n_16007;
wire n_5512;
wire n_14764;
wire n_10793;
wire n_14635;
wire n_5207;
wire n_12853;
wire n_9044;
wire n_6786;
wire n_12327;
wire n_13927;
wire n_7206;
wire n_7303;
wire n_10552;
wire n_9083;
wire n_12215;
wire n_4963;
wire n_13112;
wire n_15682;
wire n_14631;
wire n_4240;
wire n_4508;
wire n_8363;
wire n_9408;
wire n_13779;
wire n_12975;
wire n_11802;
wire n_7710;
wire n_8383;
wire n_5035;
wire n_5282;
wire n_10885;
wire n_11583;
wire n_11349;
wire n_16000;
wire n_8328;
wire n_13499;
wire n_7461;
wire n_12641;
wire n_9331;
wire n_8060;
wire n_6649;
wire n_14203;
wire n_14939;
wire n_7154;
wire n_8551;
wire n_14264;
wire n_13768;
wire n_8002;
wire n_12924;
wire n_4977;
wire n_15935;
wire n_10108;
wire n_8594;
wire n_6810;
wire n_13386;
wire n_7660;
wire n_14070;
wire n_12071;
wire n_6276;
wire n_11016;
wire n_6072;
wire n_12738;
wire n_4128;
wire n_8976;
wire n_4145;
wire n_8617;
wire n_14144;
wire n_5033;
wire n_10883;
wire n_7686;
wire n_16119;
wire n_4211;
wire n_10117;
wire n_15940;
wire n_16152;
wire n_12139;
wire n_9846;
wire n_12328;
wire n_8603;
wire n_7024;
wire n_12493;
wire n_14762;
wire n_7205;
wire n_9204;
wire n_6742;
wire n_9769;
wire n_11342;
wire n_15734;
wire n_16153;
wire n_9312;
wire n_13493;
wire n_10363;
wire n_16208;
wire n_8319;
wire n_6694;
wire n_9610;
wire n_15411;
wire n_7616;
wire n_4517;
wire n_7486;
wire n_13220;
wire n_15406;
wire n_13822;
wire n_4425;
wire n_4950;
wire n_4988;
wire n_11450;
wire n_14287;
wire n_8244;
wire n_12028;
wire n_9273;
wire n_12357;
wire n_4615;
wire n_6580;
wire n_6090;
wire n_12515;
wire n_7010;
wire n_11678;
wire n_5480;
wire n_6549;
wire n_8105;
wire n_14471;
wire n_6913;
wire n_7867;
wire n_13158;
wire n_10756;
wire n_7315;
wire n_11801;
wire n_14435;
wire n_13516;
wire n_16013;
wire n_11653;
wire n_11737;
wire n_7004;
wire n_8961;
wire n_13415;
wire n_16240;
wire n_4131;
wire n_7772;
wire n_10761;
wire n_11299;
wire n_5402;
wire n_13146;
wire n_5851;
wire n_13889;
wire n_5509;
wire n_13775;
wire n_9773;
wire n_15311;
wire n_8574;
wire n_11089;
wire n_14045;
wire n_11077;
wire n_8864;
wire n_15797;
wire n_12861;
wire n_9173;
wire n_12709;
wire n_7641;
wire n_11296;
wire n_15567;
wire n_5154;
wire n_9363;
wire n_8681;
wire n_7468;
wire n_9796;
wire n_5469;
wire n_6431;
wire n_11800;
wire n_13906;
wire n_14721;
wire n_12012;
wire n_12462;
wire n_5744;
wire n_14714;
wire n_12266;
wire n_9049;
wire n_11947;
wire n_5453;
wire n_14411;
wire n_11917;
wire n_15377;
wire n_14537;
wire n_7861;
wire n_9907;
wire n_4499;
wire n_4927;
wire n_8413;
wire n_9738;
wire n_15543;
wire n_5202;
wire n_5648;
wire n_10745;
wire n_13748;
wire n_14898;
wire n_13178;
wire n_7667;
wire n_13072;
wire n_6931;
wire n_9539;
wire n_14270;
wire n_8114;
wire n_15657;
wire n_9811;
wire n_12970;
wire n_6618;
wire n_13771;
wire n_6408;
wire n_9993;
wire n_9208;
wire n_14729;
wire n_10421;
wire n_7523;
wire n_4311;
wire n_14800;
wire n_8706;
wire n_4691;
wire n_13000;
wire n_5922;
wire n_16182;
wire n_8158;
wire n_11594;
wire n_15727;
wire n_12100;
wire n_14959;
wire n_6698;
wire n_4678;
wire n_15990;
wire n_9500;
wire n_15484;
wire n_16017;
wire n_8104;
wire n_10399;
wire n_5848;
wire n_10420;
wire n_12575;
wire n_11635;
wire n_5406;
wire n_12501;
wire n_6085;
wire n_14408;
wire n_15805;
wire n_12819;
wire n_7421;
wire n_7306;
wire n_11505;
wire n_14403;
wire n_8819;
wire n_15753;
wire n_10535;
wire n_6214;
wire n_7493;
wire n_10360;
wire n_12027;
wire n_9420;
wire n_7804;
wire n_8089;
wire n_12111;
wire n_12075;
wire n_12078;
wire n_13401;
wire n_9557;
wire n_4203;
wire n_13708;
wire n_9382;
wire n_5241;
wire n_12175;
wire n_6939;
wire n_12604;
wire n_7528;
wire n_11615;
wire n_10307;
wire n_14519;
wire n_10781;
wire n_8262;
wire n_8290;
wire n_9206;
wire n_11507;
wire n_7562;
wire n_12626;
wire n_11497;
wire n_5037;
wire n_9388;
wire n_10193;
wire n_14611;
wire n_11541;
wire n_4468;
wire n_5661;
wire n_6991;
wire n_8885;
wire n_5562;
wire n_16192;
wire n_9772;
wire n_10437;
wire n_12142;
wire n_10430;
wire n_8147;
wire n_4976;
wire n_6586;
wire n_11111;
wire n_11354;
wire n_5008;
wire n_10177;
wire n_13782;
wire n_8310;
wire n_11052;
wire n_4811;
wire n_13875;
wire n_5398;
wire n_6096;
wire n_15548;
wire n_6707;
wire n_14170;
wire n_10175;
wire n_5852;
wire n_12767;
wire n_6920;
wire n_13110;
wire n_6868;
wire n_9311;
wire n_12754;
wire n_5144;
wire n_9422;
wire n_14892;
wire n_4758;
wire n_10672;
wire n_9040;
wire n_9795;
wire n_14336;
wire n_15551;
wire n_8380;
wire n_9027;
wire n_15813;
wire n_8962;
wire n_12225;
wire n_7402;
wire n_4255;
wire n_5577;
wire n_10626;
wire n_7592;
wire n_4484;
wire n_15697;
wire n_11316;
wire n_7152;
wire n_14579;
wire n_15312;
wire n_6512;
wire n_9966;
wire n_11272;
wire n_13571;
wire n_13096;
wire n_4237;
wire n_15154;
wire n_8126;
wire n_5689;
wire n_13087;
wire n_13309;
wire n_10392;
wire n_5894;
wire n_12670;
wire n_12152;
wire n_15336;
wire n_7801;
wire n_7992;
wire n_11588;
wire n_11689;
wire n_9161;
wire n_10231;
wire n_7463;
wire n_12101;
wire n_8556;
wire n_10316;
wire n_9369;
wire n_13753;
wire n_13147;
wire n_4901;
wire n_9033;
wire n_13542;
wire n_8305;
wire n_10683;
wire n_6725;
wire n_14109;
wire n_7613;
wire n_9429;
wire n_12576;
wire n_7083;
wire n_4917;
wire n_7086;
wire n_7349;
wire n_14458;
wire n_13610;
wire n_15343;
wire n_10514;
wire n_6464;
wire n_8317;
wire n_10730;
wire n_10958;
wire n_13095;
wire n_10562;
wire n_11273;
wire n_11962;
wire n_14856;
wire n_15008;
wire n_13706;
wire n_8653;
wire n_7647;
wire n_5825;
wire n_7779;
wire n_7712;
wire n_14792;
wire n_11303;
wire n_14711;
wire n_7316;
wire n_6820;
wire n_12224;
wire n_5343;
wire n_9780;
wire n_10252;
wire n_4421;
wire n_10438;
wire n_9824;
wire n_6098;
wire n_12237;
wire n_7019;
wire n_12751;
wire n_13612;
wire n_6686;
wire n_11664;
wire n_10523;
wire n_15481;
wire n_4836;
wire n_11720;
wire n_5062;
wire n_10202;
wire n_11398;
wire n_15106;
wire n_11659;
wire n_4469;
wire n_4414;
wire n_6561;
wire n_6584;
wire n_7452;
wire n_5184;
wire n_7956;
wire n_8939;
wire n_4532;
wire n_12824;
wire n_15823;
wire n_9489;
wire n_8604;
wire n_7323;
wire n_14605;
wire n_14405;
wire n_15932;
wire n_11365;
wire n_13755;
wire n_12269;
wire n_7195;
wire n_6701;
wire n_13243;
wire n_10988;
wire n_7478;
wire n_11836;
wire n_16030;
wire n_6769;
wire n_7683;
wire n_13131;
wire n_6592;
wire n_11150;
wire n_5686;
wire n_12298;
wire n_12019;
wire n_13457;
wire n_5463;
wire n_14263;
wire n_14824;
wire n_5236;
wire n_6062;
wire n_6191;
wire n_7903;
wire n_11003;
wire n_12299;
wire n_9625;
wire n_8440;
wire n_15995;
wire n_10980;
wire n_4405;
wire n_5433;
wire n_10367;
wire n_8525;
wire n_4195;
wire n_8416;
wire n_13734;
wire n_13219;
wire n_4969;
wire n_4504;
wire n_9570;
wire n_12232;
wire n_9368;
wire n_15040;
wire n_15981;
wire n_8064;
wire n_13547;
wire n_5909;
wire n_7575;
wire n_15564;
wire n_8879;
wire n_10664;
wire n_4408;
wire n_13458;
wire n_9115;
wire n_9694;
wire n_9367;
wire n_4531;
wire n_6043;
wire n_15544;
wire n_11520;
wire n_13747;
wire n_12812;
wire n_6271;
wire n_7171;
wire n_4567;
wire n_11099;
wire n_7701;
wire n_4164;
wire n_13223;
wire n_5315;
wire n_4234;
wire n_4130;
wire n_11859;
wire n_13416;
wire n_8931;
wire n_15290;
wire n_5348;
wire n_5055;
wire n_8214;
wire n_9072;
wire n_14973;
wire n_16025;
wire n_6793;
wire n_7873;
wire n_9612;
wire n_16154;
wire n_12777;
wire n_15762;
wire n_9971;
wire n_13620;
wire n_8729;
wire n_14886;
wire n_7127;
wire n_16141;
wire n_5397;
wire n_6550;
wire n_4471;
wire n_5031;
wire n_10575;
wire n_11746;
wire n_5709;
wire n_4444;
wire n_7568;
wire n_10803;
wire n_15331;
wire n_15503;
wire n_6021;
wire n_16179;
wire n_9720;
wire n_5695;
wire n_4983;
wire n_7814;
wire n_9213;
wire n_10187;
wire n_10400;
wire n_14227;
wire n_14345;
wire n_11330;
wire n_14698;
wire n_10778;
wire n_15896;
wire n_5860;
wire n_6926;
wire n_4916;
wire n_11121;
wire n_9607;
wire n_4302;
wire n_7589;
wire n_6928;
wire n_7965;
wire n_13283;
wire n_15911;
wire n_15857;
wire n_5862;
wire n_6304;
wire n_8228;
wire n_8210;
wire n_5189;
wire n_10586;
wire n_6956;
wire n_10040;
wire n_5381;
wire n_13555;
wire n_4786;
wire n_7026;
wire n_4160;
wire n_6782;
wire n_13582;
wire n_5854;
wire n_11911;
wire n_5516;
wire n_15316;
wire n_9554;
wire n_15281;
wire n_9262;
wire n_11599;
wire n_15649;
wire n_12412;
wire n_8387;
wire n_7002;
wire n_12782;
wire n_8898;
wire n_8410;
wire n_14852;
wire n_7141;
wire n_14019;
wire n_10935;
wire n_13809;
wire n_5936;
wire n_6126;
wire n_9761;
wire n_12284;
wire n_12612;
wire n_11102;
wire n_8795;
wire n_9649;
wire n_10164;
wire n_10269;
wire n_11039;
wire n_8501;
wire n_12567;
wire n_15622;
wire n_10401;
wire n_14228;
wire n_15264;
wire n_6027;
wire n_6598;
wire n_9529;
wire n_9254;
wire n_15205;
wire n_15345;
wire n_11535;
wire n_4647;
wire n_6342;
wire n_14854;
wire n_14627;
wire n_6638;
wire n_10651;
wire n_16183;
wire n_7308;
wire n_5254;
wire n_12180;
wire n_15828;
wire n_6900;
wire n_8953;
wire n_14016;
wire n_13295;
wire n_12731;
wire n_13644;
wire n_9726;
wire n_11686;
wire n_8823;
wire n_12153;
wire n_10851;
wire n_7264;
wire n_14046;
wire n_11730;
wire n_12608;
wire n_7457;
wire n_4613;
wire n_12383;
wire n_7718;
wire n_10918;
wire n_4649;
wire n_7617;
wire n_13629;
wire n_14671;
wire n_15041;
wire n_13360;
wire n_9197;
wire n_14265;
wire n_13351;
wire n_6269;
wire n_8843;
wire n_11942;
wire n_14709;
wire n_5615;
wire n_4795;
wire n_12057;
wire n_14098;
wire n_15913;
wire n_5902;
wire n_7768;
wire n_13083;
wire n_5479;
wire n_10964;
wire n_13294;
wire n_14143;
wire n_15165;
wire n_13234;
wire n_16020;
wire n_15632;
wire n_7974;
wire n_13896;
wire n_12902;
wire n_9106;
wire n_6013;
wire n_7357;
wire n_5083;
wire n_8247;
wire n_9564;
wire n_6927;
wire n_15257;
wire n_9627;
wire n_7975;
wire n_10864;
wire n_13380;
wire n_6503;
wire n_5888;
wire n_8172;
wire n_4186;
wire n_8941;
wire n_8940;
wire n_9739;
wire n_7310;
wire n_10598;
wire n_11835;
wire n_12070;
wire n_13021;
wire n_15687;
wire n_16031;
wire n_14797;
wire n_4731;
wire n_11444;
wire n_5698;
wire n_5592;
wire n_7521;
wire n_12430;
wire n_4618;
wire n_7593;
wire n_4742;
wire n_6256;
wire n_7716;
wire n_13971;
wire n_15798;
wire n_4099;
wire n_7406;
wire n_7600;
wire n_11353;
wire n_10223;
wire n_5870;
wire n_13884;
wire n_9812;
wire n_14905;
wire n_4295;
wire n_14415;
wire n_11823;
wire n_9646;
wire n_5303;
wire n_15594;
wire n_13686;
wire n_10451;
wire n_10553;
wire n_12718;
wire n_12393;
wire n_10201;
wire n_12249;
wire n_7076;
wire n_11814;
wire n_12719;
wire n_8780;
wire n_10215;
wire n_11205;
wire n_9465;
wire n_12932;
wire n_14093;
wire n_9928;
wire n_14150;
wire n_4694;
wire n_8456;
wire n_9970;
wire n_13719;
wire n_4533;
wire n_11138;
wire n_14238;
wire n_5081;
wire n_9894;
wire n_10100;
wire n_10278;
wire n_5124;
wire n_10436;
wire n_15425;
wire n_5807;
wire n_5863;
wire n_5943;
wire n_4244;
wire n_4603;
wire n_11048;
wire n_4254;
wire n_15341;
wire n_16203;
wire n_9129;
wire n_14641;
wire n_14842;
wire n_6982;
wire n_14616;
wire n_4697;
wire n_7286;
wire n_7137;
wire n_12625;
wire n_9957;
wire n_10915;
wire n_13172;
wire n_4190;
wire n_9558;
wire n_11292;
wire n_15642;
wire n_13167;
wire n_15185;
wire n_11487;
wire n_11753;
wire n_4810;
wire n_7848;
wire n_6727;
wire n_11782;
wire n_8218;
wire n_10689;
wire n_9267;
wire n_12371;
wire n_7539;
wire n_16231;
wire n_8769;
wire n_7229;
wire n_4391;
wire n_10538;
wire n_8514;
wire n_14628;
wire n_14117;
wire n_13487;
wire n_16232;
wire n_5954;
wire n_11865;
wire n_12258;
wire n_4157;
wire n_4283;
wire n_8368;
wire n_4681;
wire n_12163;
wire n_8334;
wire n_15605;
wire n_15743;
wire n_9918;
wire n_4638;
wire n_8159;
wire n_6097;
wire n_10773;
wire n_11397;
wire n_8639;
wire n_10621;
wire n_5047;
wire n_11600;
wire n_15506;
wire n_14116;
wire n_12516;
wire n_14342;
wire n_16143;
wire n_5346;
wire n_14916;
wire n_5517;
wire n_7125;
wire n_6677;
wire n_7797;
wire n_8216;
wire n_4707;
wire n_14979;
wire n_13887;
wire n_4527;
wire n_14740;
wire n_6624;
wire n_7121;
wire n_5109;
wire n_10924;
wire n_15186;
wire n_11844;
wire n_10874;
wire n_7869;
wire n_6466;
wire n_12871;
wire n_10942;
wire n_12602;
wire n_12295;
wire n_13912;
wire n_14171;
wire n_15307;
wire n_15285;
wire n_14830;
wire n_4156;
wire n_9956;
wire n_15134;
wire n_4848;
wire n_9095;
wire n_9715;
wire n_14975;
wire n_6008;
wire n_15048;
wire n_15338;
wire n_15679;
wire n_12198;
wire n_8337;
wire n_11201;
wire n_14141;
wire n_8257;
wire n_11781;
wire n_10292;
wire n_7983;
wire n_11550;
wire n_12077;
wire n_15404;
wire n_7781;
wire n_8125;
wire n_12166;
wire n_12786;
wire n_13467;
wire n_14677;
wire n_5624;
wire n_14860;
wire n_4918;
wire n_5714;
wire n_16069;
wire n_5806;
wire n_9246;
wire n_13675;
wire n_7624;
wire n_10653;
wire n_9683;
wire n_12117;
wire n_12110;
wire n_11945;
wire n_14716;
wire n_4898;
wire n_12216;
wire n_6221;
wire n_7160;
wire n_8063;
wire n_9931;
wire n_6805;
wire n_12098;
wire n_15229;
wire n_6185;
wire n_5010;
wire n_7762;
wire n_13097;
wire n_13749;
wire n_15064;
wire n_8731;
wire n_14334;
wire n_14683;
wire n_15744;
wire n_12102;
wire n_13009;
wire n_14373;
wire n_14325;
wire n_8950;
wire n_13535;
wire n_14955;
wire n_16075;
wire n_10624;
wire n_15776;
wire n_12802;
wire n_13982;
wire n_6568;
wire n_9011;
wire n_9899;
wire n_5358;
wire n_4528;
wire n_8295;
wire n_13668;
wire n_12570;
wire n_15124;
wire n_13577;
wire n_14836;
wire n_4619;
wire n_4673;
wire n_13034;
wire n_6004;
wire n_6351;
wire n_7552;
wire n_8059;
wire n_14292;
wire n_4822;
wire n_8995;
wire n_8146;
wire n_11502;
wire n_14583;
wire n_6901;
wire n_8082;
wire n_11965;
wire n_13046;
wire n_11997;
wire n_9094;
wire n_5580;
wire n_4299;
wire n_5937;
wire n_14589;
wire n_4801;
wire n_7183;
wire n_13300;
wire n_12456;
wire n_15179;
wire n_11424;
wire n_6411;
wire n_15617;
wire n_8339;
wire n_15898;
wire n_13405;
wire n_11816;
wire n_9195;
wire n_7746;
wire n_13641;
wire n_5435;
wire n_12768;
wire n_10867;
wire n_11361;
wire n_10701;
wire n_14735;
wire n_14233;
wire n_15848;
wire n_11062;
wire n_14068;
wire n_6873;
wire n_14610;
wire n_4279;
wire n_4769;
wire n_15253;
wire n_14584;
wire n_4632;
wire n_10741;
wire n_5373;
wire n_5745;
wire n_15223;
wire n_8032;
wire n_14505;
wire n_7139;
wire n_14655;
wire n_12710;
wire n_12483;
wire n_8640;
wire n_4294;
wire n_9332;
wire n_10016;
wire n_16019;
wire n_10070;
wire n_5279;
wire n_14121;
wire n_4125;
wire n_4232;
wire n_8351;
wire n_4949;
wire n_10190;
wire n_14673;
wire n_11499;
wire n_8196;
wire n_11580;
wire n_15084;
wire n_12128;
wire n_6594;
wire n_5493;
wire n_4790;
wire n_7857;
wire n_9054;
wire n_10812;
wire n_10150;
wire n_15132;
wire n_9460;
wire n_9638;
wire n_12682;
wire n_13028;
wire n_6387;
wire n_14896;
wire n_13613;
wire n_12389;
wire n_7223;
wire n_7890;
wire n_12464;
wire n_4847;
wire n_6179;
wire n_9281;
wire n_7338;
wire n_5321;
wire n_10134;
wire n_11379;
wire n_13700;
wire n_7964;
wire n_13135;
wire n_5096;
wire n_9740;
wire n_16024;
wire n_4365;
wire n_9475;
wire n_8865;
wire n_9661;
wire n_13721;
wire n_13056;
wire n_10861;
wire n_6019;
wire n_12313;
wire n_15672;
wire n_12147;
wire n_11070;
wire n_9190;
wire n_6222;
wire n_7165;
wire n_8110;
wire n_11245;
wire n_10635;
wire n_12874;
wire n_14749;
wire n_6223;
wire n_8475;
wire n_8838;
wire n_4610;
wire n_6435;
wire n_12909;
wire n_9143;
wire n_4489;
wire n_12990;
wire n_14871;
wire n_7235;
wire n_5210;
wire n_6976;
wire n_4967;
wire n_6486;
wire n_8488;
wire n_15547;
wire n_11286;
wire n_16095;
wire n_5657;
wire n_6889;
wire n_6083;
wire n_4992;
wire n_8766;
wire n_15785;
wire n_6844;
wire n_13628;
wire n_7795;
wire n_8969;
wire n_12240;
wire n_11631;
wire n_7404;
wire n_13326;
wire n_9891;
wire n_10555;
wire n_4542;
wire n_6295;
wire n_11147;
wire n_10897;
wire n_9087;
wire n_11700;
wire n_15894;
wire n_15151;
wire n_9804;
wire n_10287;
wire n_8087;
wire n_8119;
wire n_15793;
wire n_15227;
wire n_10135;
wire n_9321;
wire n_7885;
wire n_12468;
wire n_4198;
wire n_5857;
wire n_10983;
wire n_15243;
wire n_16204;
wire n_8173;
wire n_4534;
wire n_4500;
wire n_11833;
wire n_9800;
wire n_7437;
wire n_15242;
wire n_5014;
wire n_11053;
wire n_6241;
wire n_8420;
wire n_15283;
wire n_6087;
wire n_14035;
wire n_8019;
wire n_9186;
wire n_15266;
wire n_15327;
wire n_13307;
wire n_9951;
wire n_6846;
wire n_4597;
wire n_4329;
wire n_9243;
wire n_11335;
wire n_14346;
wire n_14921;
wire n_13509;
wire n_14902;
wire n_15416;
wire n_5756;
wire n_12294;
wire n_11336;
wire n_11247;
wire n_11057;
wire n_6041;
wire n_7822;
wire n_12186;
wire n_15943;
wire n_8851;
wire n_14949;
wire n_6994;
wire n_15069;
wire n_10987;
wire n_15523;
wire n_4257;
wire n_7449;
wire n_11262;
wire n_7329;
wire n_9359;
wire n_5708;
wire n_10402;
wire n_15083;
wire n_15599;
wire n_13238;
wire n_8687;
wire n_6790;
wire n_14813;
wire n_15280;
wire n_12860;
wire n_15357;
wire n_10001;
wire n_13598;
wire n_15801;
wire n_10666;
wire n_7194;
wire n_11363;
wire n_6273;
wire n_14482;
wire n_11783;
wire n_8740;
wire n_11661;
wire n_14450;
wire n_15664;
wire n_11026;
wire n_6807;
wire n_11889;
wire n_15066;
wire n_14806;
wire n_14990;
wire n_5927;
wire n_15433;
wire n_10189;
wire n_12939;
wire n_9879;
wire n_4665;
wire n_8221;
wire n_8468;
wire n_7708;
wire n_7696;
wire n_14708;
wire n_11756;
wire n_13153;
wire n_11232;
wire n_11419;
wire n_13211;
wire n_15570;
wire n_5638;
wire n_9975;
wire n_10997;
wire n_7115;
wire n_9335;
wire n_13763;
wire n_4189;
wire n_5670;
wire n_9171;
wire n_12778;
wire n_8815;
wire n_14994;
wire n_9942;
wire n_11081;
wire n_13304;
wire n_12813;
wire n_13391;
wire n_13711;
wire n_11407;
wire n_5584;
wire n_8952;
wire n_14102;
wire n_11654;
wire n_9247;
wire n_9933;
wire n_5965;
wire n_12907;
wire n_4463;
wire n_7958;
wire n_10209;
wire n_8128;
wire n_11519;
wire n_4687;
wire n_5751;
wire n_13475;
wire n_10434;
wire n_5664;
wire n_12011;
wire n_9441;
wire n_11668;
wire n_11913;
wire n_4670;
wire n_11978;
wire n_15013;
wire n_15718;
wire n_4703;
wire n_15014;
wire n_10829;
wire n_5641;
wire n_8667;
wire n_6218;
wire n_8863;
wire n_7281;
wire n_10233;
wire n_11810;
wire n_8106;
wire n_9362;
wire n_15710;
wire n_10690;
wire n_15723;
wire n_14212;
wire n_10311;
wire n_15639;
wire n_14001;
wire n_6824;
wire n_11198;
wire n_11767;
wire n_8717;
wire n_14712;
wire n_6189;
wire n_11595;
wire n_16201;
wire n_13305;
wire n_9216;
wire n_11168;
wire n_8299;
wire n_5262;
wire n_9200;
wire n_6993;
wire n_6037;
wire n_7245;
wire n_11872;
wire n_13787;
wire n_16187;
wire n_5963;
wire n_5980;
wire n_8892;
wire n_15303;
wire n_11235;
wire n_12007;
wire n_10146;
wire n_4763;
wire n_14445;
wire n_14550;
wire n_9067;
wire n_12712;
wire n_5310;
wire n_9152;
wire n_12846;
wire n_8287;
wire n_11906;
wire n_13837;
wire n_15139;
wire n_14604;
wire n_4594;
wire n_6153;
wire n_15604;
wire n_9074;
wire n_13550;
wire n_7989;
wire n_14528;
wire n_13908;
wire n_15019;
wire n_10790;
wire n_16241;
wire n_5970;
wire n_6418;
wire n_12908;
wire n_6564;
wire n_13461;
wire n_13955;
wire n_15997;
wire n_8657;
wire n_12505;
wire n_12747;
wire n_15150;
wire n_12577;
wire n_4714;
wire n_12426;
wire n_16175;
wire n_5146;
wire n_4776;
wire n_11122;
wire n_9287;
wire n_4102;
wire n_8197;
wire n_9511;
wire n_14500;
wire n_13733;
wire n_15621;
wire n_10052;
wire n_13067;
wire n_8081;
wire n_7192;
wire n_12309;
wire n_13974;
wire n_15158;
wire n_6671;
wire n_10407;
wire n_10449;
wire n_11324;
wire n_12164;
wire n_15803;
wire n_6591;
wire n_6266;
wire n_10950;
wire n_14235;
wire n_14425;
wire n_7161;
wire n_11566;
wire n_14352;
wire n_7580;
wire n_7153;
wire n_9880;
wire n_10072;
wire n_14929;
wire n_9843;
wire n_5213;
wire n_8609;
wire n_11869;
wire n_14609;
wire n_15640;
wire n_5441;
wire n_6517;
wire n_14326;
wire n_11579;
wire n_14196;
wire n_8559;
wire n_7350;
wire n_15938;
wire n_10838;
wire n_5690;
wire n_12140;
wire n_13312;
wire n_10369;
wire n_14075;
wire n_6967;
wire n_5885;
wire n_10920;
wire n_9248;
wire n_6433;
wire n_10321;
wire n_12178;
wire n_7535;
wire n_6893;
wire n_9128;
wire n_13003;
wire n_8452;
wire n_14261;
wire n_10506;
wire n_4443;
wire n_5461;
wire n_11082;
wire n_4507;
wire n_7178;
wire n_13192;
wire n_7480;
wire n_10224;
wire n_7632;
wire n_4575;
wire n_12554;
wire n_10671;
wire n_8771;
wire n_15212;
wire n_8140;
wire n_8476;
wire n_9528;
wire n_12912;
wire n_13213;
wire n_6501;
wire n_8981;
wire n_10157;
wire n_12200;
wire n_11529;
wire n_9507;
wire n_6028;
wire n_14603;
wire n_13557;
wire n_16001;
wire n_14332;
wire n_5629;
wire n_4452;
wire n_4348;
wire n_5634;
wire n_5430;
wire n_9533;
wire n_13890;
wire n_12611;
wire n_13767;
wire n_5362;
wire n_8137;
wire n_6709;
wire n_15630;
wire n_14285;
wire n_4355;
wire n_15924;
wire n_14443;
wire n_12322;
wire n_8469;
wire n_13270;
wire n_10808;
wire n_6798;
wire n_12303;
wire n_12507;
wire n_5702;
wire n_5050;
wire n_16023;
wire n_5063;
wire n_15941;
wire n_5229;
wire n_7844;
wire n_5199;
wire n_11430;
wire n_11882;
wire n_12023;
wire n_14379;
wire n_13802;
wire n_14128;
wire n_14991;
wire n_9665;
wire n_4572;
wire n_8423;
wire n_12171;
wire n_12395;
wire n_12472;
wire n_12815;
wire n_5527;
wire n_6986;
wire n_11146;
wire n_8090;
wire n_5609;
wire n_12239;
wire n_5416;
wire n_10504;
wire n_11279;
wire n_15715;
wire n_4104;
wire n_10975;
wire n_4512;
wire n_13176;
wire n_4377;
wire n_5266;
wire n_7471;
wire n_13443;
wire n_13418;
wire n_9436;
wire n_5355;
wire n_9562;
wire n_6745;
wire n_11516;
wire n_11005;
wire n_8260;
wire n_4521;
wire n_8481;
wire n_13961;
wire n_15261;
wire n_4488;
wire n_5977;
wire n_15342;
wire n_6811;
wire n_15867;
wire n_14811;
wire n_6209;
wire n_6875;
wire n_13799;
wire n_10566;
wire n_15369;
wire n_15745;
wire n_15491;
wire n_14685;
wire n_16215;
wire n_11451;
wire n_4588;
wire n_14146;
wire n_15870;
wire n_15763;
wire n_11980;
wire n_11076;
wire n_7905;
wire n_14877;
wire n_6853;
wire n_4519;
wire n_12121;
wire n_15020;
wire n_5551;
wire n_7594;
wire n_7766;
wire n_7803;
wire n_7340;
wire n_10837;
wire n_6699;
wire n_7747;
wire n_15648;
wire n_6073;
wire n_8205;
wire n_5767;
wire n_8401;
wire n_6324;
wire n_12116;
wire n_8651;
wire n_14260;
wire n_5640;
wire n_10199;
wire n_13020;
wire n_13621;
wire n_8284;
wire n_10688;
wire n_14999;
wire n_12261;
wire n_9255;
wire n_16189;
wire n_15873;
wire n_10039;
wire n_15625;
wire n_8828;
wire n_5655;
wire n_5475;
wire n_11239;
wire n_12259;
wire n_12338;
wire n_14310;
wire n_14608;
wire n_7603;
wire n_6138;
wire n_8510;
wire n_8810;
wire n_13163;
wire n_9034;
wire n_15611;
wire n_15778;
wire n_9203;
wire n_9601;
wire n_13173;
wire n_5692;
wire n_4856;
wire n_7726;
wire n_10443;
wire n_11623;
wire n_12825;
wire n_7494;
wire n_5921;
wire n_12222;
wire n_8024;
wire n_9946;
wire n_14383;
wire n_4400;
wire n_5168;
wire n_10887;
wire n_13253;
wire n_13119;
wire n_9967;
wire n_6477;
wire n_10735;
wire n_10274;
wire n_8739;
wire n_8133;
wire n_8373;
wire n_8919;
wire n_11740;
wire n_14469;
wire n_4778;
wire n_13525;
wire n_10482;
wire n_15478;
wire n_6159;
wire n_11012;
wire n_9647;
wire n_16197;
wire n_6283;
wire n_7396;
wire n_9912;
wire n_14237;
wire n_5322;
wire n_14774;
wire n_11698;
wire n_7116;
wire n_12779;
wire n_14782;
wire n_16018;
wire n_14694;
wire n_7519;
wire n_4352;
wire n_10485;
wire n_6943;
wire n_4441;
wire n_9329;
wire n_6827;
wire n_4761;
wire n_10652;
wire n_12465;
wire n_6173;
wire n_8318;
wire n_13042;
wire n_16170;
wire n_8542;
wire n_11059;
wire n_14592;
wire n_4347;
wire n_8543;
wire n_8846;
wire n_10791;
wire n_6312;
wire n_4593;
wire n_14803;
wire n_14895;
wire n_11236;
wire n_13514;
wire n_14183;
wire n_4727;
wire n_4568;
wire n_12852;
wire n_13994;
wire n_5371;
wire n_12334;
wire n_15502;
wire n_13162;
wire n_6997;
wire n_15044;
wire n_5418;
wire n_15095;
wire n_15910;
wire n_11196;
wire n_11629;
wire n_10411;
wire n_12847;
wire n_7770;
wire n_16037;
wire n_10286;
wire n_14679;
wire n_12511;
wire n_11643;
wire n_7664;
wire n_10913;
wire n_13199;
wire n_15068;
wire n_5316;
wire n_9890;
wire n_13969;
wire n_14736;
wire n_10273;
wire n_15005;
wire n_6300;
wire n_9609;
wire n_9883;
wire n_10172;
wire n_7815;
wire n_16011;
wire n_13209;
wire n_12014;
wire n_9046;
wire n_13407;
wire n_9361;
wire n_8163;
wire n_13980;
wire n_11609;
wire n_6131;
wire n_4893;
wire n_15554;
wire n_5032;
wire n_10806;
wire n_6537;
wire n_13712;
wire n_5933;
wire n_13059;
wire n_15759;
wire n_12305;
wire n_4948;
wire n_13681;
wire n_14864;
wire n_9864;
wire n_13521;
wire n_4406;
wire n_12485;
wire n_7023;
wire n_8972;
wire n_9300;
wire n_12408;
wire n_15749;
wire n_13263;
wire n_12238;
wire n_7428;
wire n_5112;
wire n_10694;
wire n_5386;
wire n_11509;
wire n_6783;
wire n_11351;
wire n_9353;
wire n_4748;
wire n_9766;
wire n_7465;
wire n_13720;
wire n_11271;
wire n_8293;
wire n_5017;
wire n_14421;
wire n_9832;
wire n_16213;
wire n_10754;
wire n_14480;
wire n_4710;
wire n_14663;
wire n_12409;
wire n_13565;
wire n_11307;
wire n_13685;
wire n_5123;
wire n_4607;
wire n_9954;
wire n_4117;
wire n_8737;
wire n_13129;
wire n_14091;
wire n_7961;
wire n_10953;
wire n_15477;
wire n_11761;
wire n_7847;
wire n_9997;
wire n_10703;
wire n_16048;
wire n_11973;
wire n_4487;
wire n_15144;
wire n_5001;
wire n_9334;
wire n_7149;
wire n_8252;
wire n_15052;
wire n_6459;
wire n_9622;
wire n_10847;
wire n_11565;
wire n_14088;
wire n_13446;
wire n_11252;
wire n_15786;
wire n_8450;
wire n_4817;
wire n_7700;
wire n_9284;
wire n_5644;
wire n_14318;
wire n_13865;
wire n_9147;
wire n_8367;
wire n_12454;
wire n_10103;
wire n_8834;
wire n_6869;
wire n_8078;
wire n_10922;
wire n_10413;
wire n_11571;
wire n_4849;
wire n_10738;
wire n_12587;
wire n_4867;
wire n_13197;
wire n_5424;
wire n_15222;
wire n_7914;
wire n_13916;
wire n_10995;
wire n_7967;
wire n_9794;
wire n_11858;
wire n_4728;
wire n_14812;
wire n_13963;
wire n_7117;
wire n_14845;
wire n_9354;
wire n_8471;
wire n_11904;
wire n_15890;
wire n_12324;
wire n_13925;
wire n_4247;
wire n_4933;
wire n_12130;
wire n_6977;
wire n_8474;
wire n_12643;
wire n_7984;
wire n_13448;
wire n_15931;
wire n_10185;
wire n_11131;
wire n_4902;
wire n_11478;
wire n_4518;
wire n_10591;
wire n_11656;
wire n_14426;
wire n_16228;
wire n_12955;
wire n_4409;
wire n_4411;
wire n_11673;
wire n_11821;
wire n_8361;
wire n_15412;
wire n_6313;
wire n_11701;
wire n_10856;
wire n_14348;
wire n_15757;
wire n_13626;
wire n_4336;
wire n_6569;
wire n_4777;
wire n_15356;
wire n_9494;
wire n_16132;
wire n_6555;
wire n_9614;
wire n_11283;
wire n_13616;
wire n_12948;
wire n_14329;
wire n_9551;
wire n_13653;
wire n_6639;
wire n_7516;
wire n_5496;
wire n_13694;
wire n_9154;
wire n_13233;
wire n_10677;
wire n_7596;
wire n_13189;
wire n_16089;
wire n_13640;
wire n_5864;
wire n_6536;
wire n_14211;
wire n_4398;
wire n_8553;
wire n_6490;
wire n_8301;
wire n_15003;
wire n_10610;
wire n_6961;
wire n_13392;
wire n_4954;
wire n_12574;
wire n_12697;
wire n_9437;
wire n_5460;
wire n_7628;
wire n_9276;
wire n_4304;
wire n_6761;
wire n_15760;
wire n_14572;
wire n_9346;
wire n_11229;
wire n_15626;
wire n_5333;
wire n_15724;
wire n_6294;
wire n_14851;
wire n_11636;
wire n_6767;
wire n_8518;
wire n_4431;
wire n_7427;
wire n_4192;
wire n_6802;
wire n_7527;
wire n_13962;
wire n_12162;
wire n_5570;
wire n_6326;
wire n_9514;
wire n_4805;
wire n_11919;
wire n_9402;
wire n_14118;
wire n_10456;
wire n_12634;
wire n_11675;
wire n_10343;
wire n_4885;
wire n_7838;
wire n_8364;
wire n_7786;
wire n_5983;
wire n_9580;
wire n_14134;
wire n_9005;
wire n_5804;
wire n_12236;
wire n_7979;
wire n_6376;
wire n_8621;
wire n_6167;
wire n_15231;
wire n_8993;
wire n_7926;
wire n_4701;
wire n_12632;
wire n_5910;
wire n_7411;
wire n_14545;
wire n_7101;
wire n_12398;
wire n_6730;
wire n_5040;
wire n_6948;
wire n_15415;
wire n_10979;
wire n_13591;
wire n_10487;
wire n_10332;
wire n_9162;
wire n_9921;
wire n_9443;
wire n_6582;
wire n_13479;
wire n_8910;
wire n_7752;
wire n_13631;
wire n_15453;
wire n_9897;
wire n_11570;
wire n_15364;
wire n_10807;
wire n_6996;
wire n_11855;
wire n_9817;
wire n_14930;
wire n_15389;
wire n_11667;
wire n_15166;
wire n_9301;
wire n_6974;
wire n_7731;
wire n_8753;
wire n_15265;
wire n_6765;
wire n_7577;
wire n_8388;
wire n_9401;
wire n_16171;
wire n_8321;
wire n_6921;
wire n_11290;
wire n_13738;
wire n_15739;
wire n_8044;
wire n_15937;
wire n_8091;
wire n_14137;
wire n_8486;
wire n_7845;
wire n_13122;
wire n_10750;
wire n_12292;
wire n_7709;
wire n_9689;
wire n_4631;
wire n_15628;
wire n_11592;
wire n_11466;
wire n_5194;
wire n_15536;
wire n_13346;
wire n_9982;
wire n_6898;
wire n_12056;
wire n_6710;
wire n_13149;
wire n_5717;
wire n_7162;
wire n_6565;
wire n_5464;
wire n_8508;
wire n_12679;
wire n_8261;
wire n_14179;
wire n_15262;
wire n_12811;
wire n_13100;
wire n_14821;
wire n_5886;
wire n_7080;
wire n_16096;
wire n_9886;
wire n_7744;
wire n_13232;
wire n_12897;
wire n_8034;
wire n_8841;
wire n_10970;
wire n_14401;
wire n_7302;
wire n_6533;
wire n_12837;
wire n_4965;
wire n_10264;
wire n_6960;
wire n_8201;
wire n_6426;
wire n_6634;
wire n_7180;
wire n_5610;
wire n_6836;
wire n_5239;
wire n_11983;
wire n_13840;
wire n_15735;
wire n_12605;
wire n_11043;
wire n_4747;
wire n_5197;
wire n_8947;
wire n_15792;
wire n_16233;
wire n_15609;
wire n_9671;
wire n_6972;
wire n_9297;
wire n_8788;
wire n_10472;
wire n_13460;
wire n_13389;
wire n_7111;
wire n_7549;
wire n_4111;
wire n_14180;
wire n_5785;
wire n_4587;
wire n_11415;
wire n_15849;
wire n_13578;
wire n_6344;
wire n_14773;
wire n_5305;
wire n_5994;
wire n_6093;
wire n_4538;
wire n_10499;
wire n_8093;
wire n_11680;
wire n_13870;
wire n_15096;
wire n_6010;
wire n_14958;
wire n_15791;
wire n_15696;
wire n_7247;
wire n_13088;
wire n_11446;
wire n_9225;
wire n_8061;
wire n_6833;
wire n_11972;
wire n_14247;
wire n_5376;
wire n_13862;
wire n_13600;
wire n_11103;
wire n_7481;
wire n_10435;
wire n_12220;
wire n_13843;
wire n_10066;
wire n_13605;
wire n_14707;
wire n_5204;
wire n_7292;
wire n_10341;
wire n_12230;
wire n_15987;
wire n_14511;
wire n_8811;
wire n_12995;
wire n_7150;
wire n_13486;
wire n_14176;
wire n_7687;
wire n_10498;
wire n_10184;
wire n_13599;
wire n_12867;
wire n_9662;
wire n_8507;
wire n_10508;
wire n_9057;
wire n_12497;
wire n_14173;
wire n_14323;
wire n_4150;
wire n_14667;
wire n_4878;
wire n_12406;
wire n_6265;
wire n_8861;
wire n_14544;
wire n_11749;
wire n_14875;
wire n_6821;
wire n_8661;
wire n_15740;
wire n_11417;
wire n_8545;
wire n_12725;
wire n_4985;
wire n_6373;
wire n_6988;
wire n_8755;
wire n_5788;
wire n_11490;
wire n_12401;
wire n_13404;
wire n_8573;
wire n_8191;
wire n_11704;
wire n_7692;
wire n_5897;
wire n_6887;
wire n_10865;
wire n_11343;
wire n_14777;
wire n_15065;
wire n_9809;
wire n_13277;
wire n_12185;
wire n_16041;
wire n_13518;
wire n_14157;
wire n_8683;
wire n_15293;
wire n_10081;
wire n_8836;
wire n_6676;
wire n_7016;
wire n_6347;
wire n_6492;
wire n_13540;
wire n_14366;
wire n_12161;
wire n_15756;
wire n_15676;
wire n_9448;
wire n_16220;
wire n_8136;
wire n_8446;
wire n_9799;
wire n_7742;
wire n_10577;
wire n_9313;
wire n_15085;
wire n_8916;
wire n_14650;
wire n_14657;
wire n_7955;
wire n_5795;
wire n_7072;
wire n_5508;
wire n_10037;
wire n_13370;
wire n_12424;
wire n_5582;
wire n_15844;
wire n_10234;
wire n_14801;
wire n_7374;
wire n_7440;
wire n_9989;
wire n_11766;
wire n_4852;
wire n_7758;
wire n_11639;
wire n_7547;
wire n_14802;
wire n_12114;
wire n_13171;
wire n_11967;
wire n_4869;
wire n_9438;
wire n_13528;
wire n_4700;
wire n_7201;
wire n_13419;
wire n_14087;
wire n_11457;
wire n_4426;
wire n_10832;
wire n_12490;
wire n_10036;
wire n_12571;
wire n_11932;
wire n_15053;
wire n_5746;
wire n_15559;
wire n_5292;
wire n_14656;
wire n_10853;
wire n_12508;
wire n_12582;
wire n_6648;
wire n_7880;
wire n_12052;
wire n_14757;
wire n_4601;
wire n_8075;
wire n_13937;
wire n_14298;
wire n_14623;
wire n_8857;
wire n_11275;
wire n_14253;
wire n_4220;
wire n_8587;
wire n_12337;
wire n_9675;
wire n_10030;
wire n_5630;
wire n_9667;
wire n_10676;
wire n_11819;
wire n_8071;
wire n_13159;
wire n_15766;
wire n_10815;
wire n_12928;
wire n_16064;
wire n_11589;
wire n_11309;
wire n_12927;
wire n_15161;
wire n_15401;
wire n_13347;
wire n_11803;
wire n_7513;
wire n_11067;
wire n_12321;
wire n_4515;
wire n_4351;
wire n_11274;
wire n_5264;
wire n_9537;
wire n_11174;
wire n_7413;
wire n_10833;
wire n_4403;
wire n_11795;
wire n_11770;
wire n_12610;
wire n_7540;
wire n_8646;
wire n_15381;
wire n_4858;
wire n_4509;
wire n_15829;
wire n_9866;
wire n_5504;
wire n_8630;
wire n_7622;
wire n_9602;
wire n_14392;
wire n_15373;
wire n_7005;
wire n_11266;
wire n_11151;
wire n_4223;
wire n_7353;
wire n_6219;
wire n_10071;
wire n_9885;
wire n_15216;
wire n_14115;
wire n_12592;
wire n_15654;
wire n_14992;
wire n_15811;
wire n_12698;
wire n_13343;
wire n_8315;
wire n_14282;
wire n_6965;
wire n_9260;
wire n_13938;
wire n_16063;
wire n_5025;
wire n_8314;
wire n_12048;
wire n_6720;
wire n_14615;
wire n_8149;
wire n_16169;
wire n_6032;
wire n_11413;
wire n_8581;
wire n_15729;
wire n_13932;
wire n_13094;
wire n_7174;
wire n_8565;
wire n_6205;
wire n_6362;
wire n_6402;
wire n_14668;
wire n_14509;
wire n_4644;
wire n_7166;
wire n_4456;
wire n_5060;
wire n_15495;
wire n_7607;
wire n_8209;
wire n_9159;
wire n_5334;
wire n_15973;
wire n_15317;
wire n_4346;
wire n_7816;
wire n_13290;
wire n_9654;
wire n_8560;
wire n_7591;
wire n_15500;
wire n_5775;
wire n_8141;
wire n_14139;
wire n_7830;
wire n_7282;
wire n_6491;
wire n_13198;
wire n_8302;
wire n_10015;
wire n_9306;
wire n_11682;
wire n_7151;
wire n_11652;
wire n_12801;
wire n_6229;
wire n_11091;
wire n_15325;
wire n_11929;
wire n_9978;
wire n_16116;
wire n_5731;
wire n_8612;
wire n_5581;
wire n_7446;
wire n_6668;
wire n_16139;
wire n_10362;
wire n_4235;
wire n_15952;
wire n_7053;
wire n_8724;
wire n_11331;
wire n_11640;
wire n_14702;
wire n_5831;
wire n_10171;
wire n_12552;
wire n_7473;
wire n_4435;
wire n_10183;
wire n_10471;
wire n_14674;
wire n_8070;
wire n_6835;
wire n_13039;
wire n_6419;
wire n_6039;
wire n_12704;
wire n_11237;
wire n_15304;
wire n_11601;
wire n_11741;
wire n_14130;
wire n_14402;
wire n_15839;
wire n_14305;
wire n_5884;
wire n_14400;
wire n_9279;
wire n_8457;
wire n_4764;
wire n_5653;
wire n_8922;
wire n_10095;
wire n_8248;
wire n_7966;
wire n_9509;
wire n_6258;
wire n_10549;
wire n_7070;
wire n_5394;
wire n_15775;
wire n_11721;
wire n_6755;
wire n_9563;
wire n_7276;
wire n_7351;
wire n_12256;
wire n_7942;
wire n_10057;
wire n_4655;
wire n_12477;
wire n_4581;
wire n_12184;
wire n_11093;
wire n_12245;
wire n_6084;
wire n_10301;
wire n_15888;
wire n_4827;
wire n_9496;
wire n_13156;
wire n_15531;
wire n_8411;
wire n_12657;
wire n_12740;
wire n_9644;
wire n_7412;
wire n_7157;
wire n_6436;
wire n_7666;
wire n_12089;
wire n_13957;
wire n_6472;
wire n_14051;
wire n_8527;
wire n_5421;
wire n_11097;
wire n_7211;
wire n_10394;
wire n_10154;
wire n_4399;
wire n_11681;
wire n_6531;
wire n_5309;
wire n_7901;
wire n_8689;
wire n_11522;
wire n_14724;
wire n_9750;
wire n_4782;
wire n_9980;
wire n_13164;
wire n_10818;
wire n_12145;
wire n_8988;
wire n_4363;
wire n_11105;
wire n_12647;
wire n_12377;
wire n_12721;
wire n_4864;
wire n_9251;
wire n_10141;
wire n_15906;
wire n_7368;
wire n_15420;
wire n_13624;
wire n_8549;
wire n_12541;
wire n_12316;
wire n_4335;
wire n_6567;
wire n_5889;
wire n_11849;
wire n_6771;
wire n_11578;
wire n_13484;
wire n_10916;
wire n_10208;
wire n_13714;
wire n_6389;
wire n_10182;
wire n_13655;
wire n_9616;
wire n_15142;
wire n_15037;
wire n_12399;
wire n_8004;
wire n_10929;
wire n_15189;
wire n_8658;
wire n_9959;
wire n_8375;
wire n_10403;
wire n_5764;
wire n_10260;
wire n_6910;
wire n_5428;
wire n_9291;
wire n_9092;
wire n_10261;
wire n_6442;
wire n_12285;
wire n_16180;
wire n_13606;
wire n_6102;
wire n_8908;
wire n_5541;
wire n_4259;
wire n_15067;
wire n_13438;
wire n_16003;
wire n_10384;
wire n_6441;
wire n_15868;
wire n_5543;
wire n_10372;
wire n_9818;
wire n_10237;
wire n_9283;
wire n_5678;
wire n_5935;
wire n_4865;
wire n_11219;
wire n_13498;
wire n_14453;
wire n_4564;
wire n_7677;
wire n_5085;
wire n_8569;
wire n_13661;
wire n_8676;
wire n_10118;
wire n_5950;
wire n_15260;
wire n_12379;
wire n_15413;
wire n_13496;
wire n_7929;
wire n_10028;
wire n_12257;
wire n_10691;
wire n_8399;
wire n_5995;
wire n_12246;
wire n_16060;
wire n_15363;
wire n_11069;
wire n_6162;
wire n_5116;
wire n_4526;
wire n_6331;
wire n_13674;
wire n_14099;
wire n_6006;
wire n_8421;
wire n_4417;
wire n_6109;
wire n_11268;
wire n_6278;
wire n_9304;
wire n_12655;
wire n_13818;
wire n_14855;
wire n_6787;
wire n_10777;
wire n_11066;
wire n_6872;
wire n_6208;
wire n_4899;
wire n_14642;
wire n_15858;
wire n_6632;
wire n_13133;
wire n_9310;
wire n_7754;
wire n_5411;
wire n_14246;
wire n_4798;
wire n_9830;
wire n_9913;
wire n_11728;
wire n_7027;
wire n_8001;
wire n_5671;
wire n_8322;
wire n_12272;
wire n_6990;
wire n_12862;
wire n_8403;
wire n_6349;
wire n_14885;
wire n_13140;
wire n_11796;
wire n_13573;
wire n_7631;
wire n_6830;
wire n_8999;
wire n_12662;
wire n_8754;
wire n_5185;
wire n_7939;
wire n_8675;
wire n_7898;
wire n_10715;
wire n_12136;
wire n_14889;
wire n_6359;
wire n_9375;
wire n_15111;
wire n_16068;
wire n_8596;
wire n_10665;
wire n_10073;
wire n_10291;
wire n_13251;
wire n_14890;
wire n_8858;
wire n_8666;
wire n_11873;
wire n_15579;
wire n_8313;
wire n_7763;
wire n_10296;
wire n_13154;
wire n_7498;
wire n_5076;
wire n_7377;
wire n_11228;
wire n_8555;
wire n_5379;
wire n_15149;
wire n_15769;
wire n_4750;
wire n_12517;
wire n_13796;
wire n_16173;
wire n_6301;
wire n_12031;
wire n_11743;
wire n_14274;
wire n_10512;
wire n_8610;
wire n_13195;
wire n_13314;
wire n_14456;
wire n_13679;
wire n_12993;
wire n_10324;
wire n_13658;
wire n_12663;
wire n_7945;
wire n_5945;
wire n_14850;
wire n_11261;
wire n_13667;
wire n_9323;
wire n_6744;
wire n_4981;
wire n_10765;
wire n_9985;
wire n_12039;
wire n_11023;
wire n_8615;
wire n_11382;
wire n_4835;
wire n_5811;
wire n_4430;
wire n_6439;
wire n_14278;
wire n_10026;
wire n_8677;
wire n_9355;
wire n_8602;
wire n_9714;
wire n_12938;
wire n_7381;
wire n_13772;
wire n_10041;
wire n_5565;
wire n_7948;
wire n_4407;
wire n_8102;
wire n_7291;
wire n_16210;
wire n_9540;
wire n_14840;
wire n_15859;
wire n_4894;
wire n_13033;
wire n_9753;
wire n_5780;
wire n_8460;
wire n_9105;
wire n_13746;
wire n_5643;
wire n_11305;
wire n_10149;
wire n_16088;
wire n_12680;
wire n_13017;
wire n_14530;
wire n_11137;
wire n_11607;
wire n_5846;
wire n_7430;
wire n_9700;
wire n_14234;
wire n_15511;
wire n_12930;
wire n_13914;
wire n_13752;
wire n_4995;
wire n_15093;
wire n_8871;
wire n_10649;
wire n_14360;
wire n_9476;
wire n_12722;
wire n_7870;
wire n_13529;
wire n_9875;
wire n_11265;
wire n_10593;
wire n_12042;
wire n_5524;
wire n_8824;
wire n_14827;
wire n_10597;
wire n_9963;
wire n_6104;
wire n_4446;
wire n_6475;
wire n_8470;
wire n_9582;
wire n_12469;
wire n_16058;
wire n_12172;
wire n_15533;
wire n_11739;
wire n_10817;
wire n_6465;
wire n_10060;
wire n_9574;
wire n_12049;
wire n_6496;
wire n_13229;
wire n_13973;
wire n_11687;
wire n_14160;
wire n_9732;
wire n_11050;
wire n_13070;
wire n_15576;
wire n_14440;
wire n_12666;
wire n_8238;
wire n_9882;
wire n_12205;
wire n_6998;
wire n_10779;
wire n_13177;
wire n_15230;
wire n_6145;
wire n_11789;
wire n_16239;
wire n_8699;
wire n_14946;
wire n_7305;
wire n_13878;
wire n_10242;
wire n_10086;
wire n_16135;
wire n_9992;
wire n_12885;
wire n_14899;
wire n_15204;
wire n_11347;
wire n_15899;
wire n_14166;
wire n_4332;
wire n_4314;
wire n_7980;
wire n_14363;
wire n_11617;
wire n_14952;
wire n_7075;
wire n_7545;
wire n_11581;
wire n_7846;
wire n_10981;
wire n_6076;
wire n_4288;
wire n_14626;
wire n_8438;
wire n_14831;
wire n_6194;
wire n_10673;
wire n_10869;
wire n_7695;
wire n_5066;
wire n_13850;
wire n_12917;
wire n_6092;
wire n_7275;
wire n_15254;
wire n_5401;
wire n_6357;
wire n_5843;
wire n_4241;
wire n_8095;
wire n_12616;
wire n_7537;
wire n_13690;
wire n_14356;
wire n_14429;
wire n_14705;
wire n_10128;
wire n_10746;
wire n_12217;
wire n_12287;
wire n_12950;
wire n_15845;
wire n_7489;
wire n_5106;
wire n_10339;
wire n_15572;
wire n_11559;
wire n_14629;
wire n_5468;
wire n_11867;
wire n_15197;
wire n_4265;
wire n_6335;
wire n_8112;
wire n_12835;
wire n_14727;
wire n_14343;
wire n_5883;
wire n_6985;
wire n_8642;
wire n_5319;
wire n_14996;
wire n_15072;
wire n_13552;
wire n_13432;
wire n_15800;
wire n_7451;
wire n_8624;
wire n_16161;
wire n_6238;
wire n_9090;
wire n_14066;
wire n_15780;
wire n_11989;
wire n_12800;
wire n_13495;
wire n_10684;
wire n_15030;
wire n_10441;
wire n_12177;
wire n_12036;
wire n_9149;
wire n_10590;
wire n_9174;
wire n_12850;
wire n_11175;
wire n_12962;
wire n_6548;
wire n_14755;
wire n_4705;
wire n_5455;
wire n_8894;
wire n_9226;
wire n_6366;
wire n_5706;
wire n_5337;
wire n_9018;
wire n_12336;
wire n_10949;
wire n_7236;
wire n_9835;
wire n_12044;
wire n_15135;
wire n_11727;
wire n_12905;
wire n_7269;
wire n_4604;
wire n_8878;
wire n_15663;
wire n_15706;
wire n_5223;
wire n_10934;
wire n_5962;
wire n_6602;
wire n_5020;
wire n_4419;
wire n_4477;
wire n_14018;
wire n_6620;
wire n_6502;
wire n_15856;
wire n_9702;
wire n_13409;
wire n_7560;
wire n_15348;
wire n_11725;
wire n_15565;
wire n_10279;
wire n_11291;
wire n_15138;
wire n_7326;
wire n_13548;
wire n_7060;
wire n_15643;
wire n_7572;
wire n_15301;
wire n_6885;
wire n_12495;
wire n_13139;
wire n_4217;
wire n_4395;
wire n_8807;
wire n_14207;
wire n_12565;
wire n_9968;
wire n_5074;
wire n_5364;
wire n_9924;
wire n_6529;
wire n_8732;
wire n_8169;
wire n_15174;
wire n_11958;
wire n_15954;
wire n_16207;
wire n_8803;
wire n_9515;
wire n_8017;
wire n_10527;
wire n_13506;
wire n_5895;
wire n_4639;
wire n_14756;
wire n_6951;
wire n_8801;
wire n_12584;
wire n_14258;
wire n_5649;
wire n_5046;
wire n_5166;
wire n_7169;
wire n_12654;
wire n_13255;
wire n_6423;
wire n_9252;
wire n_15017;
wire n_14938;
wire n_15779;
wire n_10785;
wire n_7140;
wire n_7233;
wire n_10228;
wire n_11311;
wire n_12999;
wire n_14084;
wire n_13120;
wire n_5088;
wire n_6558;
wire n_8522;
wire n_5457;
wire n_15123;
wire n_7352;
wire n_15869;
wire n_7986;
wire n_15863;
wire n_9948;
wire n_7134;
wire n_5532;
wire n_12823;
wire n_11528;
wire n_12422;
wire n_6950;
wire n_7246;
wire n_12234;
wire n_6525;
wire n_7650;
wire n_9871;
wire n_11807;
wire n_14907;
wire n_6892;
wire n_6631;
wire n_11705;
wire n_8203;
wire n_15162;
wire n_15653;
wire n_14587;
wire n_15678;
wire n_7663;
wire n_13125;
wire n_15566;
wire n_9423;
wire n_11378;
wire n_11521;
wire n_11998;
wire n_4227;
wire n_4289;
wire n_9660;
wire n_14513;
wire n_9108;
wire n_14472;
wire n_11222;
wire n_15562;
wire n_15015;
wire n_4780;
wire n_14910;
wire n_8680;
wire n_9631;
wire n_10643;
wire n_7056;
wire n_4243;
wire n_14590;
wire n_4982;
wire n_12293;
wire n_16130;
wire n_10427;
wire n_4330;
wire n_6683;
wire n_8727;
wire n_15333;
wire n_10389;
wire n_13069;
wire n_13254;
wire n_16211;
wire n_15658;
wire n_10423;
wire n_6292;
wire n_5544;
wire n_15094;
wire n_9900;
wire n_14042;
wire n_15305;
wire n_11080;
wire n_7729;
wire n_7339;
wire n_5987;
wire n_7740;
wire n_6180;
wire n_5352;
wire n_5824;
wire n_14409;
wire n_4991;
wire n_11533;
wire n_12572;
wire n_5538;
wire n_8138;
wire n_6658;
wire n_10863;
wire n_6264;
wire n_9608;
wire n_9137;
wire n_15344;
wire n_6925;
wire n_8990;
wire n_15616;
wire n_5919;
wire n_10077;
wire n_12988;
wire n_8206;
wire n_9144;
wire n_12512;
wire n_7767;
wire n_11940;
wire n_13736;
wire n_8190;
wire n_6176;
wire n_13727;
wire n_9778;
wire n_16009;
wire n_8622;
wire n_13352;
wire n_15247;
wire n_5410;
wire n_11808;
wire n_13986;
wire n_15035;
wire n_7146;
wire n_8092;
wire n_13953;
wire n_15520;
wire n_10250;
wire n_15819;
wire n_6124;
wire n_7672;
wire n_14251;
wire n_8242;
wire n_4525;
wire n_12118;
wire n_12609;
wire n_14053;
wire n_14494;
wire n_7482;
wire n_12176;
wire n_14503;
wire n_9850;
wire n_14940;
wire n_6864;
wire n_9531;
wire n_13453;
wire n_7893;
wire n_4208;
wire n_8331;
wire n_15921;
wire n_7090;
wire n_15105;
wire n_11549;
wire n_16123;
wire n_7158;
wire n_14174;
wire n_15644;
wire n_7156;
wire n_5742;
wire n_5992;
wire n_8649;
wire n_15438;
wire n_16244;
wire n_8684;
wire n_6494;
wire n_5503;
wire n_8323;
wire n_10828;
wire n_4177;
wire n_12353;
wire n_6199;
wire n_11139;
wire n_8296;
wire n_13846;
wire n_9139;
wire n_11584;
wire n_9430;
wire n_10417;
wire n_5958;
wire n_6614;
wire n_7749;
wire n_15059;
wire n_11695;
wire n_16148;
wire n_7839;
wire n_4264;
wire n_8882;
wire n_10310;
wire n_12053;
wire n_7504;
wire n_10333;
wire n_13316;
wire n_10996;
wire n_13583;
wire n_12795;
wire n_9272;
wire n_10880;
wire n_8708;
wire n_12045;
wire n_7360;
wire n_10810;
wire n_12274;
wire n_7681;
wire n_10636;
wire n_12348;
wire n_8448;
wire n_8076;
wire n_7301;
wire n_9041;
wire n_11360;
wire n_5129;
wire n_11886;
wire n_9643;
wire n_8904;
wire n_7375;
wire n_7102;
wire n_5500;
wire n_8277;
wire n_15883;
wire n_11920;
wire n_4276;
wire n_15215;
wire n_7794;
wire n_11479;
wire n_13388;
wire n_12006;
wire n_7366;
wire n_16196;
wire n_8184;
wire n_13344;
wire n_5219;
wire n_13336;
wire n_14516;
wire n_15851;
wire n_5605;
wire n_9944;
wire n_14103;
wire n_16245;
wire n_5170;
wire n_5654;
wire n_7025;
wire n_8304;
wire n_5320;
wire n_13915;
wire n_14935;
wire n_10258;
wire n_11534;
wire n_6947;
wire n_8586;
wire n_5107;
wire n_9648;
wire n_5999;
wire n_4485;
wire n_9376;
wire n_8557;
wire n_10507;
wire n_16184;
wire n_8636;
wire n_7309;
wire n_13885;
wire n_4626;
wire n_6863;
wire n_9288;
wire n_10835;
wire n_6637;
wire n_15240;
wire n_15507;
wire n_6100;
wire n_13259;
wire n_7860;
wire n_6735;
wire n_14815;
wire n_9521;
wire n_9541;
wire n_13477;
wire n_8212;
wire n_6358;
wire n_4975;
wire n_9759;
wire n_14737;
wire n_12500;
wire n_12781;
wire n_13204;
wire n_16038;
wire n_7911;
wire n_15469;
wire n_13085;
wire n_15455;
wire n_11848;
wire n_8530;
wire n_9278;
wire n_9378;
wire n_11227;
wire n_8665;
wire n_5602;
wire n_9456;
wire n_13778;
wire n_9086;
wire n_7876;
wire n_15532;
wire n_6050;
wire n_11401;
wire n_15329;
wire n_15164;
wire n_14925;
wire n_9711;
wire n_8933;
wire n_14805;
wire n_13206;
wire n_15309;
wire n_7244;
wire n_15709;
wire n_7960;
wire n_5405;
wire n_13462;
wire n_12922;
wire n_14123;
wire n_5253;
wire n_9485;
wire n_4760;
wire n_11375;
wire n_4652;
wire n_4624;
wire n_9555;
wire n_10959;
wire n_7610;
wire n_12842;
wire n_9999;
wire n_11813;
wire n_14353;
wire n_9994;
wire n_10814;
wire n_5903;
wire n_6371;
wire n_8690;
wire n_8538;
wire n_7043;
wire n_12753;
wire n_16248;
wire n_15214;
wire n_10859;
wire n_6171;
wire n_7751;
wire n_8643;
wire n_15366;
wire n_6510;
wire n_15430;
wire n_6468;
wire n_4569;
wire n_9142;
wire n_9613;
wire n_11134;
wire n_4897;
wire n_9440;
wire n_5491;
wire n_8825;
wire n_11716;
wire n_12366;
wire n_7788;
wire n_14548;
wire n_5842;
wire n_6352;
wire n_8300;
wire n_13954;
wire n_10531;
wire n_14419;
wire n_5722;
wire n_7534;
wire n_9462;
wire n_5636;
wire n_7719;
wire n_11357;
wire n_9202;
wire n_7287;
wire n_5065;
wire n_10699;
wire n_12208;
wire n_7032;
wire n_8451;
wire n_11386;
wire n_13383;
wire n_14161;
wire n_4523;
wire n_5492;
wire n_9237;
wire n_10941;
wire n_11448;
wire n_5084;
wire n_10567;
wire n_6850;
wire n_8435;
wire n_5667;
wire n_16120;
wire n_12122;
wire n_14600;
wire n_10770;
wire n_5260;
wire n_11693;
wire n_7119;
wire n_8835;
wire n_4919;
wire n_13728;
wire n_15038;
wire n_10714;
wire n_9788;
wire n_13584;
wire n_15358;
wire n_13722;
wire n_5328;
wire n_14060;
wire n_14936;
wire n_6354;
wire n_5918;
wire n_7634;
wire n_14634;
wire n_16145;
wire n_11755;
wire n_4503;
wire n_6959;
wire n_6909;
wire n_11221;
wire n_7851;
wire n_6332;
wire n_9807;
wire n_14613;
wire n_13642;
wire n_4464;
wire n_13567;
wire n_7006;
wire n_15473;
wire n_15912;
wire n_9573;
wire n_5877;
wire n_8963;
wire n_12351;
wire n_6306;
wire n_7682;
wire n_15659;
wire n_4114;
wire n_14297;
wire n_13618;
wire n_6434;
wire n_12040;
wire n_12443;
wire n_8713;
wire n_6751;
wire n_7068;
wire n_9392;
wire n_12133;
wire n_4556;
wire n_11084;
wire n_13371;
wire n_14573;
wire n_6322;
wire n_14048;
wire n_8668;
wire n_8353;
wire n_13301;
wire n_5454;
wire n_9390;
wire n_13492;
wire n_14376;
wire n_7704;
wire n_10326;
wire n_7773;
wire n_9416;
wire n_14728;
wire n_6667;
wire n_7526;
wire n_13333;
wire n_8817;
wire n_6530;
wire n_9518;
wire n_13329;
wire n_15578;
wire n_12491;
wire n_7376;
wire n_13826;
wire n_6156;
wire n_13966;
wire n_14498;
wire n_5913;
wire n_7268;
wire n_16198;
wire n_7044;
wire n_12452;
wire n_5621;
wire n_13788;
wire n_13437;
wire n_16082;
wire n_8213;
wire n_12233;
wire n_4327;
wire n_8591;
wire n_7973;
wire n_11885;
wire n_4218;
wire n_6429;
wire n_13423;
wire n_10966;
wire n_5165;
wire n_15914;
wire n_7239;
wire n_10047;
wire n_12633;
wire n_5573;
wire n_11253;
wire n_6405;
wire n_11551;
wire n_14761;
wire n_8532;
wire n_11380;
wire n_12936;
wire n_15199;
wire n_12035;
wire n_13928;
wire n_6613;
wire n_4353;
wire n_8043;
wire n_9196;
wire n_11172;
wire n_13947;
wire n_14420;
wire n_15584;
wire n_7969;
wire n_6248;
wire n_14059;
wire n_15462;
wire n_12915;
wire n_7821;
wire n_15854;
wire n_4990;
wire n_6088;
wire n_12275;
wire n_10784;
wire n_5529;
wire n_10248;
wire n_6894;
wire n_12947;
wire n_14678;
wire n_7267;
wire n_4959;
wire n_9589;
wire n_4161;
wire n_5800;
wire n_11539;
wire n_9898;
wire n_14520;
wire n_15224;
wire n_13257;
wire n_9373;
wire n_11976;
wire n_12308;
wire n_13063;
wire n_8606;
wire n_14669;
wire n_4103;
wire n_4466;
wire n_15702;
wire n_6204;
wire n_10351;
wire n_13834;
wire n_13951;
wire n_15236;
wire n_16110;
wire n_7915;
wire n_8121;
wire n_8868;
wire n_10408;
wire n_10921;
wire n_13340;
wire n_7387;
wire n_7431;
wire n_11731;
wire n_7654;
wire n_10551;
wire n_12760;
wire n_10656;
wire n_4844;
wire n_6296;
wire n_11531;
wire n_12318;
wire n_13379;
wire n_15624;
wire n_10313;
wire n_10639;
wire n_15557;
wire n_5257;
wire n_16012;
wire n_9983;
wire n_6290;
wire n_14983;
wire n_6288;
wire n_12700;
wire n_4688;
wire n_14517;
wire n_4765;
wire n_8276;
wire n_8718;
wire n_12364;
wire n_8182;
wire n_14512;
wire n_5645;
wire n_11392;
wire n_15540;
wire n_5180;
wire n_13490;
wire n_11204;
wire n_13025;
wire n_13672;
wire n_13754;
wire n_14785;
wire n_15923;
wire n_12985;
wire n_5779;
wire n_11627;
wire n_13697;
wire n_4388;
wire n_4206;
wire n_12340;
wire n_12478;
wire n_6140;
wire n_9039;
wire n_13744;
wire n_8359;
wire n_7441;
wire n_9849;
wire n_8597;
wire n_4738;
wire n_6211;
wire n_12788;
wire n_8562;
wire n_13470;
wire n_11485;
wire n_8211;
wire n_13998;
wire n_13943;
wire n_9962;
wire n_14814;
wire n_12826;
wire n_8430;
wire n_6307;
wire n_8007;
wire n_10871;
wire n_6164;
wire n_12752;
wire n_15434;
wire n_7394;
wire n_8600;
wire n_8311;
wire n_8943;
wire n_8441;
wire n_12194;
wire n_4434;
wire n_4837;
wire n_10747;
wire n_7022;
wire n_15395;
wire n_9829;
wire n_14772;
wire n_13637;
wire n_15322;
wire n_6860;
wire n_4219;
wire n_10459;
wire n_8978;
wire n_5012;
wire n_10121;
wire n_15558;
wire n_4620;
wire n_11387;
wire n_8198;
wire n_9988;
wire n_14417;
wire n_5697;
wire n_14652;
wire n_14002;
wire n_15596;
wire n_15945;
wire n_7188;
wire n_8526;
wire n_10705;
wire n_13099;
wire n_7573;
wire n_7879;
wire n_4438;
wire n_16242;
wire n_9848;
wire n_7087;
wire n_6147;
wire n_14911;
wire n_10334;
wire n_7985;
wire n_16221;
wire n_12689;
wire n_11691;
wire n_11358;
wire n_9045;
wire n_9466;
wire n_6515;
wire n_15021;
wire n_9348;
wire n_6011;
wire n_8278;
wire n_7722;
wire n_7935;
wire n_8592;
wire n_15783;
wire n_6645;
wire n_11128;
wire n_12271;
wire n_13595;
wire n_14358;
wire n_14006;
wire n_8226;
wire n_15140;
wire n_6984;
wire n_4325;
wire n_12843;
wire n_13780;
wire n_10716;
wire n_12273;
wire n_10235;
wire n_13212;
wire n_15167;
wire n_13701;
wire n_10090;
wire n_13247;
wire n_10153;
wire n_16138;
wire n_14271;
wire n_15681;
wire n_11649;
wire n_10937;
wire n_13922;
wire n_7193;
wire n_10018;
wire n_13278;
wire n_8987;
wire n_13836;
wire n_4133;
wire n_11489;
wire n_6897;
wire n_7256;
wire n_12391;
wire n_4184;
wire n_5203;
wire n_12420;
wire n_14181;
wire n_9071;
wire n_10568;
wire n_9356;
wire n_9464;
wire n_4481;
wire n_12314;
wire n_6460;
wire n_4379;
wire n_7128;
wire n_7595;
wire n_9239;
wire n_10053;
wire n_6183;
wire n_10051;
wire n_11373;
wire n_7522;
wire n_5882;
wire n_13341;
wire n_15388;
wire n_16034;
wire n_9606;
wire n_13856;
wire n_10359;
wire n_7881;
wire n_14416;
wire n_14796;
wire n_14961;
wire n_15619;
wire n_7436;
wire n_4490;
wire n_15726;
wire n_7380;
wire n_7012;
wire n_11216;
wire n_4397;
wire n_12356;
wire n_10998;
wire n_15272;
wire n_7502;
wire n_9492;
wire n_13271;
wire n_8960;
wire n_7335;
wire n_7103;
wire n_13553;
wire n_4820;
wire n_10648;
wire n_10151;
wire n_6246;
wire n_14602;
wire n_14133;
wire n_11194;
wire n_11804;
wire n_8025;
wire n_5094;
wire n_6383;
wire n_9031;
wire n_15612;
wire n_15976;
wire n_11107;
wire n_4938;
wire n_9717;
wire n_11434;
wire n_9516;
wire n_11645;
wire n_12073;
wire n_15732;
wire n_7020;
wire n_8434;
wire n_4179;
wire n_11244;
wire n_12848;
wire n_8175;
wire n_9693;
wire n_9991;
wire n_5336;
wire n_15378;
wire n_12155;
wire n_13356;
wire n_14286;
wire n_9103;
wire n_8850;
wire n_11254;
wire n_14865;
wire n_13693;
wire n_9477;
wire n_15761;
wire n_14277;
wire n_5672;
wire n_4641;
wire n_13673;
wire n_5548;
wire n_10253;
wire n_10822;
wire n_5601;
wire n_7248;
wire n_7662;
wire n_14793;
wire n_8895;
wire n_10589;
wire n_12390;
wire n_12160;
wire n_13501;
wire n_15927;
wire n_11297;
wire n_10349;
wire n_11991;
wire n_5339;
wire n_13376;
wire n_4931;
wire n_6099;
wire n_10946;
wire n_12150;
wire n_5693;
wire n_8046;
wire n_11183;
wire n_11173;
wire n_6904;
wire n_11922;
wire n_16115;
wire n_13897;
wire n_8867;
wire n_15480;
wire n_15651;
wire n_10473;
wire n_8239;
wire n_9599;
wire n_13104;
wire n_4146;
wire n_4360;
wire n_7825;
wire n_8924;
wire n_8183;
wire n_12840;
wire n_9001;
wire n_15339;
wire n_10893;
wire n_13215;
wire n_10218;
wire n_13482;
wire n_16026;
wire n_12964;
wire n_13075;
wire n_5514;
wire n_4404;
wire n_7533;
wire n_5091;
wire n_8578;
wire n_11548;
wire n_9777;
wire n_4787;
wire n_8848;
wire n_10903;
wire n_13562;
wire n_10458;
wire n_11868;
wire n_13445;
wire n_9222;
wire n_10148;
wire n_15198;
wire n_6626;
wire n_6563;
wire n_5486;
wire n_9366;
wire n_6611;
wire n_10775;
wire n_11248;
wire n_10543;
wire n_9449;
wire n_4903;
wire n_15098;
wire n_15669;
wire n_11114;
wire n_11260;
wire n_11901;
wire n_12994;
wire n_5599;
wire n_14771;
wire n_6116;
wire n_16081;
wire n_15834;
wire n_7186;
wire n_10337;
wire n_4356;
wire n_8230;
wire n_9869;
wire n_10478;
wire n_15552;
wire n_12252;
wire n_11981;
wire n_15831;
wire n_6819;
wire n_8725;
wire n_4432;
wire n_13929;
wire n_5251;
wire n_7936;
wire n_13534;
wire n_13680;
wire n_6473;
wire n_12951;
wire n_13750;
wire n_9741;
wire n_13275;
wire n_4291;
wire n_11956;
wire n_10956;
wire n_10637;
wire n_13331;
wire n_13536;
wire n_15996;
wire n_11805;
wire n_15043;
wire n_5403;
wire n_4386;
wire n_12131;
wire n_12280;
wire n_4149;
wire n_8391;
wire n_6310;
wire n_7840;
wire n_10698;
wire n_15728;
wire n_11381;
wire n_14607;
wire n_9397;
wire n_8202;
wire n_11797;
wire n_11775;
wire n_12453;
wire n_10834;
wire n_7429;
wire n_6688;
wire n_12557;
wire n_7906;
wire n_8948;
wire n_8678;
wire n_9754;
wire n_15295;
wire n_10783;
wire n_9179;
wire n_7148;
wire n_15582;
wire n_5782;
wire n_6714;
wire n_7017;
wire n_4637;
wire n_7462;
wire n_7250;
wire n_7658;
wire n_7828;
wire n_8340;
wire n_8905;
wire n_12020;
wire n_13439;
wire n_4935;
wire n_8691;
wire n_13249;
wire n_12051;
wire n_6365;
wire n_16044;
wire n_10619;
wire n_14225;
wire n_4785;
wire n_13502;
wire n_13801;
wire n_5608;
wire n_13468;
wire n_12455;
wire n_11322;
wire n_10136;
wire n_7401;
wire n_13789;
wire n_8812;
wire n_12920;
wire n_14759;
wire n_13403;
wire n_9169;
wire n_6828;
wire n_12785;
wire n_14200;
wire n_11758;
wire n_5298;
wire n_8704;
wire n_6355;
wire n_5596;
wire n_7887;
wire n_11162;
wire n_13996;
wire n_8058;
wire n_4413;
wire n_12559;
wire n_9177;
wire n_10078;
wire n_6777;
wire n_5728;
wire n_11987;
wire n_16162;
wire n_8394;
wire n_9269;
wire n_4493;
wire n_7835;
wire n_10719;
wire n_12614;
wire n_13201;
wire n_14638;
wire n_15326;
wire n_11106;
wire n_9289;
wire n_8181;
wire n_10463;
wire n_12797;
wire n_13737;
wire n_13441;
wire n_14396;
wire n_14687;
wire n_8722;
wire n_10827;
wire n_12429;
wire n_6420;
wire n_6945;
wire n_11218;
wire n_9350;
wire n_7356;
wire n_5726;
wire n_7288;
wire n_7637;
wire n_7124;
wire n_10454;
wire n_11467;
wire n_12384;
wire n_7294;
wire n_12629;
wire n_12668;
wire n_13291;
wire n_12123;
wire n_5290;
wire n_12972;
wire n_14969;
wire n_7018;
wire n_13105;
wire n_10312;
wire n_11374;
wire n_11167;
wire n_13440;
wire n_12146;
wire n_7321;
wire n_9166;
wire n_10663;
wire n_10501;
wire n_5095;
wire n_10265;
wire n_10452;
wire n_15796;
wire n_8707;
wire n_6754;
wire n_10766;
wire n_12435;
wire n_13533;
wire n_11999;
wire n_6583;
wire n_13367;
wire n_6622;
wire n_6936;
wire n_13123;
wire n_8747;
wire n_5324;
wire n_7691;
wire n_15459;
wire n_5928;
wire n_8742;
wire n_10470;
wire n_10563;
wire n_12921;
wire n_16006;
wire n_7108;
wire n_6882;
wire n_15693;
wire n_11455;
wire n_7585;
wire n_13930;
wire n_9125;
wire n_4570;
wire n_7386;
wire n_8552;
wire n_10288;
wire n_5101;
wire n_12581;
wire n_5019;
wire n_5911;
wire n_4296;
wire n_7362;
wire n_7888;
wire n_7417;
wire n_12029;
wire n_12548;
wire n_9641;
wire n_14460;
wire n_9960;
wire n_7187;
wire n_13111;
wire n_11884;
wire n_5589;
wire n_5841;
wire n_13060;
wire n_12727;
wire n_10776;
wire n_11611;
wire n_9785;
wire n_9923;
wire n_8224;
wire n_10771;
wire n_7544;
wire n_11087;
wire n_14556;
wire n_5712;
wire n_11960;
wire n_4606;
wire n_6166;
wire n_8628;
wire n_4774;
wire n_13108;
wire n_11422;
wire n_13948;
wire n_6966;
wire n_13563;
wire n_7542;
wire n_6781;
wire n_9228;
wire n_14828;
wire n_7255;
wire n_15131;
wire n_12227;
wire n_8037;
wire n_8084;
wire n_7120;
wire n_7218;
wire n_12597;
wire n_16056;
wire n_4672;
wire n_7147;
wire n_7221;
wire n_14653;
wire n_15016;
wire n_15601;
wire n_10967;
wire n_4174;
wire n_8289;
wire n_9801;
wire n_14189;
wire n_16021;
wire n_10249;
wire n_11029;
wire n_15057;
wire n_9645;
wire n_4766;
wire n_8045;
wire n_11199;
wire n_15721;
wire n_5633;
wire n_8697;
wire n_13568;
wire n_13396;
wire n_13029;
wire n_13647;
wire n_8077;
wire n_6980;
wire n_4600;
wire n_12674;
wire n_15977;
wire n_5583;
wire n_11826;
wire n_9457;
wire n_15071;
wire n_4460;
wire n_8026;
wire n_11317;
wire n_13652;
wire n_7889;
wire n_6064;
wire n_6110;
wire n_10742;
wire n_6237;
wire n_16083;
wire n_14538;
wire n_7196;
wire n_12913;
wire n_10390;
wire n_9330;
wire n_6341;
wire n_10012;
wire n_9365;
wire n_14861;
wire n_15781;
wire n_6590;
wire n_5501;
wire n_8444;
wire n_9178;
wire n_8654;
wire n_14021;
wire n_10035;
wire n_10753;
wire n_9181;
wire n_12112;
wire n_7923;
wire n_13965;
wire n_14465;
wire n_5377;
wire n_11033;
wire n_6697;
wire n_13168;
wire n_5652;
wire n_6453;
wire n_6135;
wire n_13574;
wire n_14037;
wire n_7559;
wire n_11798;
wire n_15577;
wire n_12346;
wire n_4110;
wire n_11853;
wire n_7081;
wire n_9307;
wire n_15476;
wire n_10795;
wire n_10300;
wire n_10257;
wire n_15752;
wire n_6449;
wire n_7832;
wire n_7968;
wire n_9238;
wire n_12714;
wire n_11079;
wire n_11166;
wire n_13581;
wire n_6141;
wire n_10099;
wire n_8449;
wire n_11217;
wire n_12732;
wire n_13138;
wire n_14481;
wire n_10985;
wire n_15650;
wire n_4349;
wire n_14931;
wire n_8493;
wire n_7584;
wire n_9224;
wire n_10244;
wire n_12400;
wire n_4313;
wire n_6983;
wire n_12671;
wire n_7843;
wire n_13774;
wire n_10377;
wire n_6036;
wire n_11469;
wire n_10984;
wire n_12863;
wire n_12347;
wire n_15188;
wire n_8958;
wire n_10801;
wire n_11898;
wire n_8443;
wire n_4863;
wire n_12041;
wire n_9756;
wire n_7222;
wire n_9624;
wire n_6071;
wire n_8161;
wire n_13435;
wire n_11710;
wire n_6808;
wire n_8734;
wire n_9547;
wire n_11341;
wire n_8271;
wire n_9594;
wire n_9901;
wire n_11619;
wire n_11238;
wire n_9895;
wire n_10878;
wire n_13378;
wire n_6724;
wire n_15460;
wire n_9277;
wire n_11608;
wire n_14169;
wire n_14086;
wire n_12756;
wire n_6571;
wire n_15074;
wire n_7470;
wire n_5100;
wire n_9189;
wire n_15470;
wire n_16059;
wire n_5849;
wire n_8495;
wire n_6251;
wire n_7400;
wire n_14255;
wire n_9548;
wire n_14309;
wire n_12088;
wire n_12218;
wire n_14204;
wire n_6635;
wire n_10000;
wire n_9472;
wire n_13202;
wire n_14738;
wire n_13410;
wire n_11553;
wire n_14432;
wire n_13816;
wire n_5367;
wire n_8994;
wire n_15930;
wire n_8901;
wire n_8056;
wire n_10725;
wire n_12323;
wire n_14767;
wire n_9538;
wire n_7623;
wire n_12387;
wire n_14984;
wire n_10627;
wire n_8954;
wire n_13590;
wire n_15846;
wire n_5616;
wire n_13230;
wire n_7597;
wire n_11996;
wire n_5034;
wire n_6733;
wire n_7071;
wire n_15029;
wire n_8840;
wire n_5988;
wire n_6467;
wire n_6035;
wire n_7859;
wire n_8900;
wire n_13456;
wire n_15194;
wire n_10477;
wire n_14651;
wire n_13321;
wire n_15967;
wire n_12798;
wire n_14306;
wire n_16067;
wire n_11032;
wire n_6522;
wire n_7109;
wire n_11834;
wire n_14057;
wire n_9434;
wire n_10604;
wire n_11110;
wire n_5959;
wire n_9052;
wire n_7645;
wire n_6732;
wire n_13806;
wire n_4807;
wire n_6562;
wire n_16149;
wire n_12780;
wire n_6150;
wire n_9176;
wire n_10461;
wire n_12772;
wire n_10559;
wire n_15314;
wire n_11141;
wire n_8157;
wire n_12539;
wire n_13007;
wire n_8346;
wire n_9697;
wire n_4230;
wire n_15656;
wire n_13651;
wire n_7882;
wire n_13830;
wire n_8827;
wire n_13113;
wire n_8309;
wire n_13196;
wire n_14998;
wire n_8344;
wire n_5917;
wire n_12589;
wire n_9060;
wire n_5754;
wire n_6016;
wire n_12775;
wire n_8096;
wire n_8100;
wire n_8822;
wire n_15670;
wire n_12043;
wire n_9758;
wire n_7212;
wire n_7908;
wire n_15160;
wire n_8222;
wire n_14430;
wire n_10479;
wire n_9876;
wire n_5628;
wire n_10572;
wire n_11971;
wire n_6726;
wire n_8406;
wire n_10277;
wire n_11320;
wire n_14697;
wire n_16091;
wire n_4428;
wire n_5003;
wire n_11028;
wire n_5252;
wire n_7009;
wire n_6554;
wire n_10139;
wire n_10230;
wire n_15847;
wire n_14294;
wire n_6689;
wire n_15708;
wire n_14245;
wire n_12476;
wire n_14858;
wire n_8866;
wire n_13724;
wire n_6143;
wire n_5614;
wire n_8693;
wire n_5134;
wire n_10207;
wire n_12536;
wire n_15597;
wire n_4122;
wire n_11368;
wire n_11144;
wire n_7355;
wire n_7365;
wire n_15286;
wire n_4582;
wire n_7777;
wire n_8794;
wire n_9653;
wire n_6277;
wire n_14993;
wire n_7395;
wire n_4684;
wire n_5981;
wire n_11404;
wire n_12896;
wire n_13373;
wire n_15593;
wire n_6095;
wire n_16079;
wire n_7671;
wire n_10429;
wire n_16222;
wire n_15951;
wire n_8020;
wire n_14241;
wire n_12957;
wire n_13866;
wire n_6247;
wire n_4840;
wire n_10255;
wire n_9257;
wire n_13014;
wire n_15141;
wire n_15235;
wire n_9270;
wire n_6880;
wire n_10901;
wire n_15881;
wire n_10101;
wire n_5720;
wire n_15129;
wire n_14000;
wire n_13022;
wire n_13422;
wire n_5325;
wire n_13633;
wire n_15380;
wire n_5696;
wire n_12549;
wire n_5375;
wire n_4384;
wire n_8736;
wire n_6499;
wire n_12362;
wire n_6837;
wire n_13442;
wire n_14741;
wire n_14972;
wire n_15073;
wire n_4423;
wire n_10063;
wire n_13390;
wire n_12030;
wire n_7393;
wire n_8400;
wire n_6616;
wire n_9686;
wire n_13136;
wire n_13334;
wire n_13408;
wire n_13989;
wire n_14690;
wire n_15288;
wire n_7871;
wire n_14532;
wire n_14859;
wire n_12018;
wire n_10846;
wire n_6946;
wire n_4996;
wire n_8055;
wire n_8333;
wire n_10195;
wire n_11593;
wire n_11847;
wire n_15904;
wire n_9718;
wire n_11773;
wire n_4598;
wire n_14074;
wire n_14944;
wire n_5064;
wire n_9215;
wire n_5759;
wire n_12060;
wire n_4478;
wire n_5753;
wire n_10628;
wire n_8909;
wire n_16033;
wire n_5536;
wire n_15056;
wire n_7484;
wire n_5173;
wire n_11968;
wire n_6305;
wire n_13630;
wire n_14071;
wire n_16053;
wire n_14127;
wire n_6317;
wire n_9762;
wire n_9407;
wire n_10819;
wire n_12315;
wire n_12903;
wire n_4890;
wire n_13269;
wire n_14570;
wire n_5691;
wire n_13103;
wire n_15771;
wire n_15865;
wire n_5794;
wire n_13098;
wire n_11896;
wire n_5027;
wire n_5647;
wire n_7231;
wire n_11897;
wire n_14447;
wire n_13707;
wire n_10368;
wire n_12484;
wire n_14971;
wire n_7272;
wire n_9964;
wire n_4106;
wire n_13031;
wire n_13646;
wire n_5738;
wire n_7649;
wire n_9953;
wire n_10356;
wire n_14154;
wire n_7324;
wire n_5215;
wire n_9153;
wire n_6693;
wire n_8786;
wire n_10931;
wire n_8541;
wire n_11711;
wire n_12673;
wire n_6734;
wire n_12000;
wire n_10173;
wire n_15107;
wire n_9571;
wire n_7135;
wire n_11554;
wire n_7014;
wire n_8263;
wire n_10644;
wire n_8884;
wire n_11159;
wire n_5597;
wire n_4721;
wire n_13062;
wire n_5635;
wire n_13424;
wire n_10323;
wire n_11350;
wire n_6382;
wire n_9019;
wire n_11310;
wire n_13001;
wire n_7328;
wire n_7635;
wire n_6404;
wire n_12063;
wire n_15023;
wire n_10229;
wire n_10693;
wire n_5975;
wire n_9737;
wire n_11688;
wire n_13842;
wire n_10493;
wire n_11125;
wire n_8494;
wire n_10554;
wire n_6379;
wire n_10382;
wire n_11083;
wire n_7703;
wire n_7066;
wire n_4496;
wire n_7358;
wire n_9468;
wire n_10622;
wire n_12449;
wire n_13664;
wire n_11939;
wire n_6235;
wire n_16176;
wire n_13144;
wire n_9870;
wire n_4338;
wire n_7277;
wire n_6504;
wire n_9026;
wire n_13900;
wire n_9710;
wire n_15799;
wire n_7265;
wire n_8638;
wire n_11126;
wire n_15665;
wire n_15958;
wire n_8710;
wire n_10019;
wire n_13512;
wire n_15591;
wire n_6789;
wire n_15719;
wire n_7184;
wire n_11090;
wire n_6440;
wire n_9725;
wire n_11953;
wire n_6417;
wire n_12845;
wire n_14557;
wire n_8177;
wire n_14013;
wire n_15385;
wire n_12062;
wire n_12636;
wire n_14784;
wire n_7491;
wire n_4495;
wire n_4762;
wire n_5942;
wire n_14436;
wire n_15866;
wire n_14524;
wire n_9084;
wire n_7728;
wire n_10488;
wire n_10767;
wire n_7690;
wire n_15360;
wire n_13084;
wire n_15110;
wire n_7219;
wire n_13375;
wire n_7479;
wire n_11040;
wire n_13852;
wire n_11751;
wire n_9419;
wire n_12793;
wire n_13203;
wire n_4141;
wire n_11158;
wire n_14378;
wire n_7270;
wire n_5940;
wire n_8170;
wire n_12367;
wire n_10579;
wire n_14488;
wire n_8893;
wire n_13473;
wire n_14923;
wire n_12317;
wire n_7390;
wire n_15296;
wire n_15586;
wire n_7805;
wire n_10474;
wire n_7807;
wire n_5121;
wire n_9479;
wire n_9820;
wire n_8589;
wire n_4107;
wire n_9973;
wire n_12954;
wire n_12724;
wire n_4667;
wire n_11094;
wire n_8320;
wire n_5555;
wire n_6914;
wire n_7978;
wire n_15155;
wire n_15458;
wire n_12157;
wire n_15379;
wire n_14891;
wire n_11161;
wire n_11182;
wire n_10587;
wire n_15441;
wire n_7182;
wire n_12195;
wire n_4547;
wire n_11839;
wire n_15115;
wire n_11815;
wire n_5784;
wire n_10843;
wire n_12773;
wire n_6272;
wire n_8153;
wire n_7699;
wire n_6484;
wire n_7674;
wire n_12556;
wire n_6236;
wire n_8620;
wire n_10755;
wire n_5576;
wire n_4668;
wire n_8298;
wire n_11614;
wire n_4953;
wire n_5466;
wire n_6958;
wire n_6840;
wire n_13645;
wire n_6871;
wire n_12789;
wire n_10270;
wire n_11590;
wire n_12649;
wire n_8235;
wire n_15201;
wire n_11845;
wire n_5284;
wire n_9294;
wire n_9126;
wire n_8370;
wire n_13773;
wire n_11263;
wire n_11908;
wire n_4997;
wire n_13066;
wire n_15109;
wire n_5308;
wire n_4274;
wire n_13469;
wire n_10573;
wire n_13101;
wire n_6768;
wire n_4759;
wire n_13494;
wire n_13893;
wire n_7951;
wire n_15190;
wire n_10992;
wire n_14490;
wire n_4467;
wire n_7506;
wire n_14210;
wire n_14717;
wire n_12696;
wire n_6717;
wire n_13505;
wire n_11257;
wire n_4735;
wire n_7048;
wire n_11136;
wire n_11142;
wire n_15368;
wire n_10428;
wire n_13569;
wire n_15908;
wire n_12664;
wire n_15885;
wire n_5578;
wire n_8395;
wire n_10989;
wire n_13450;
wire n_11145;
wire n_12206;
wire n_11745;
wire n_13010;
wire n_15081;
wire n_15812;
wire n_14375;
wire n_13181;
wire n_11017;
wire n_4113;
wire n_10805;
wire n_15623;
wire n_8906;
wire n_4686;
wire n_10682;
wire n_5530;
wire n_11414;
wire n_8097;
wire n_10327;
wire n_12940;
wire n_14322;
wire n_6196;
wire n_7416;
wire n_4321;
wire n_4342;
wire n_15608;
wire n_10528;
wire n_5741;
wire n_8570;
wire n_8902;
wire n_12404;
wire n_5991;
wire n_13815;
wire n_10365;
wire n_7330;
wire n_15435;
wire n_15950;
wire n_7928;
wire n_12201;
wire n_5506;
wire n_5243;
wire n_15061;
wire n_9819;
wire n_8477;
wire n_5449;
wire n_10236;
wire n_5221;
wire n_6992;
wire n_10433;
wire n_13725;
wire n_13924;
wire n_4183;
wire n_12312;
wire n_15191;
wire n_4872;
wire n_10625;
wire n_6000;
wire n_16005;
wire n_10303;
wire n_9545;
wire n_4233;
wire n_7283;
wire n_7099;
wire n_11452;
wire n_15270;
wire n_10557;
wire n_4709;
wire n_5038;
wire n_5311;
wire n_6448;
wire n_11323;
wire n_16125;
wire n_13002;
wire n_6655;
wire n_12982;
wire n_7892;
wire n_9165;
wire n_11558;
wire n_14732;
wire n_15256;
wire n_7304;
wire n_10143;
wire n_13018;
wire n_5792;
wire n_13185;
wire n_14872;
wire n_15705;
wire n_14681;
wire n_12002;
wire n_15171;
wire n_6657;
wire n_7756;
wire n_8129;
wire n_13150;
wire n_5575;
wire n_8580;
wire n_11543;
wire n_7990;
wire n_15521;
wire n_4625;
wire n_8122;
wire n_11883;
wire n_10796;
wire n_8259;
wire n_8536;
wire n_7626;
wire n_7474;
wire n_10855;
wire n_8748;
wire n_7612;
wire n_6113;
wire n_16155;
wire n_7789;
wire n_4819;
wire n_9056;
wire n_15826;
wire n_8094;
wire n_9341;
wire n_14164;
wire n_11429;
wire n_14165;
wire n_6242;
wire n_7902;
wire n_7088;
wire n_15027;
wire n_6519;
wire n_10357;
wire n_8572;
wire n_4900;
wire n_10681;
wire n_8120;
wire n_12598;
wire n_6842;
wire n_12942;
wire n_12750;
wire n_13575;
wire n_12729;
wire n_7588;
wire n_12033;
wire n_6206;
wire n_6414;
wire n_11241;
wire n_9172;
wire n_14239;
wire n_12441;
wire n_9145;
wire n_13805;
wire n_6801;
wire n_8099;
wire n_9996;
wire n_11348;
wire n_10059;
wire n_10284;
wire n_7680;
wire n_4930;
wire n_8770;
wire n_5276;
wire n_6308;
wire n_14790;
wire n_7398;
wire n_6906;
wire n_14029;
wire n_5078;
wire n_11169;
wire n_4537;
wire n_11041;
wire n_16039;
wire n_7230;
wire n_8700;
wire n_11160;
wire n_16015;
wire n_9906;
wire n_6629;
wire n_5011;
wire n_10957;
wire n_14250;
wire n_12827;
wire n_11124;
wire n_16028;
wire n_6968;
wire n_9920;
wire n_4282;
wire n_9504;
wire n_6615;
wire n_4180;
wire n_7378;
wire n_15689;
wire n_16206;
wire n_12734;
wire n_12181;
wire n_9482;
wire n_15145;
wire n_5205;
wire n_14032;
wire n_14760;
wire n_16107;
wire n_9138;
wire n_11152;
wire n_9384;
wire n_8637;
wire n_5651;
wire n_6144;
wire n_8757;
wire n_4143;
wire n_4659;
wire n_6188;
wire n_14794;
wire n_5819;
wire n_10147;
wire n_14197;
wire n_4579;
wire n_4616;
wire n_13765;
wire n_8903;
wire n_13709;
wire n_9193;
wire n_15962;
wire n_5998;
wire n_6398;
wire n_11586;
wire n_14660;
wire n_5023;
wire n_12069;
wire n_11990;
wire n_4105;
wire n_5721;
wire n_5673;
wire n_9527;
wire n_14554;
wire n_5351;
wire n_10889;
wire n_12363;
wire n_11019;
wire n_14028;
wire n_15788;
wire n_13170;
wire n_14368;
wire n_14699;
wire n_8585;
wire n_9064;
wire n_14056;
wire n_8982;
wire n_6415;
wire n_10816;
wire n_14374;
wire n_10032;
wire n_13385;
wire n_6857;
wire n_10489;
wire n_15114;
wire n_5476;
wire n_10200;
wire n_12442;
wire n_7842;
wire n_10898;
wire n_12499;
wire n_5856;
wire n_14588;
wire n_8709;
wire n_5446;
wire n_9383;
wire n_10825;
wire n_4895;
wire n_6722;
wire n_9735;
wire n_9943;
wire n_10290;
wire n_6428;
wire n_15853;
wire n_5944;
wire n_7618;
wire n_15569;
wire n_15862;
wire n_12818;
wire n_15078;
wire n_6413;
wire n_7679;
wire n_11132;
wire n_4275;
wire n_13684;
wire n_6361;
wire n_9357;
wire n_11677;
wire n_13608;
wire n_10680;
wire n_12531;
wire n_6231;
wire n_7783;
wire n_4098;
wire n_11036;
wire n_15394;
wire n_14826;
wire n_5684;
wire n_5861;
wire n_11927;
wire n_8108;
wire n_10306;
wire n_5976;
wire n_15445;
wire n_4789;
wire n_11827;
wire n_7862;
wire n_5312;
wire n_10675;
wire n_5850;
wire n_10014;
wire n_16150;
wire n_13454;
wire n_5111;
wire n_16117;
wire n_13829;
wire n_5890;
wire n_15968;
wire n_9986;
wire n_10355;
wire n_13758;
wire n_10830;
wire n_7820;
wire n_7167;
wire n_8692;
wire n_14967;
wire n_7833;
wire n_11118;
wire n_8820;
wire n_12496;
wire n_14750;
wire n_15454;
wire n_7643;
wire n_12460;
wire n_13586;
wire n_8490;
wire n_10380;
wire n_5113;
wire n_4442;
wire n_9491;
wire n_4698;
wire n_12821;
wire n_15028;
wire n_15736;
wire n_14809;
wire n_9922;
wire n_6712;
wire n_5687;
wire n_12479;
wire n_10530;
wire n_13703;
wire n_4779;
wire n_8062;
wire n_8781;
wire n_10999;
wire n_10203;
wire n_4966;
wire n_8000;
wire n_10061;
wire n_13860;
wire n_10899;
wire n_10961;
wire n_8808;
wire n_13359;
wire n_8233;
wire n_15573;
wire n_5839;
wire n_9747;
wire n_11811;
wire n_6953;
wire n_8685;
wire n_4418;
wire n_13877;
wire n_15097;
wire n_9061;
wire n_9168;
wire n_12361;
wire n_11561;
wire n_12345;
wire n_8575;
wire n_8701;
wire n_11690;
wire n_15126;
wire n_11212;
wire n_6303;
wire n_12593;
wire n_6474;
wire n_6182;
wire n_16114;
wire n_11155;
wire n_15118;
wire n_5674;
wire n_8670;
wire n_6573;
wire n_4134;
wire n_13151;
wire n_6053;
wire n_14380;
wire n_7234;
wire n_10425;
wire n_15060;
wire n_8352;
wire n_7993;
wire n_7930;
wire n_5682;
wire n_12984;
wire n_15170;
wire n_16194;
wire n_16094;
wire n_8385;
wire n_14330;
wire n_8875;
wire n_6392;
wire n_8166;
wire n_11433;
wire n_5167;
wire n_9073;
wire n_8934;
wire n_5117;
wire n_11312;
wire n_4913;
wire n_11477;
wire n_15928;
wire n_7999;
wire n_5612;
wire n_14347;
wire n_11988;
wire n_6125;
wire n_7963;
wire n_6599;
wire n_14978;
wire n_15485;
wire n_6685;
wire n_12311;
wire n_12914;
wire n_15213;
wire n_11964;
wire n_12086;
wire n_4251;
wire n_8389;
wire n_9068;
wire n_15289;
wire n_10537;
wire n_4621;
wire n_10158;
wire n_14823;
wire n_6560;
wire n_12787;
wire n_14686;
wire n_10711;
wire n_11933;
wire n_8659;
wire n_8804;
wire n_10043;
wire n_4559;
wire n_12703;
wire n_4368;
wire n_6253;
wire n_12411;
wire n_4740;
wire n_7382;
wire n_8439;
wire n_13337;
wire n_9544;
wire n_14108;
wire n_8814;
wire n_8369;
wire n_13867;
wire n_5301;
wire n_11574;
wire n_7800;
wire n_15575;
wire n_5007;
wire n_7615;
wire n_10930;
wire n_4642;
wire n_9286;
wire n_5898;
wire n_11313;
wire n_14700;
wire n_15633;
wire n_11206;
wire n_12263;
wire n_7298;
wire n_12959;
wire n_10131;
wire n_7581;
wire n_15238;
wire n_6641;
wire n_5214;
wire n_13057;
wire n_13551;
wire n_5563;
wire n_5487;
wire n_6593;
wire n_12461;
wire n_6673;
wire n_10696;
wire n_12893;
wire n_13990;
wire n_8789;
wire n_7172;
wire n_7074;
wire n_10685;
wire n_5497;
wire n_8790;
wire n_11223;
wire n_8234;
wire n_11624;
wire n_4724;
wire n_5832;
wire n_13876;
wire n_13791;
wire n_14438;
wire n_7190;
wire n_11515;
wire n_7112;
wire n_14382;
wire n_13128;
wire n_16217;
wire n_13807;
wire n_13142;
wire n_7678;
wire n_10082;
wire n_15299;
wire n_9265;
wire n_11560;
wire n_15390;
wire n_13678;
wire n_9080;
wire n_13433;
wire n_5526;
wire n_8989;
wire n_10152;
wire n_15063;
wire n_13589;
wire n_12645;
wire n_6367;
wire n_6195;
wire n_4546;
wire n_14192;
wire n_6356;
wire n_8927;
wire n_11055;
wire n_11616;
wire n_9770;
wire n_15824;
wire n_14746;
wire n_9463;
wire n_7001;
wire n_12090;
wire n_13481;
wire n_13743;
wire n_5593;
wire n_5021;
wire n_6514;
wire n_7369;
wire n_5444;
wire n_10580;
wire n_14365;
wire n_7829;
wire n_14131;
wire n_4382;
wire n_9939;
wire n_10159;
wire n_11390;
wire n_8534;
wire n_9911;
wire n_9210;
wire n_6559;
wire n_5211;
wire n_5230;
wire n_10122;
wire n_10302;
wire n_14457;
wire n_7359;
wire n_14398;
wire n_5389;
wire n_15443;
wire n_7144;
wire n_10462;
wire n_4833;
wire n_14244;
wire n_13357;
wire n_8756;
wire n_6841;
wire n_14320;
wire n_11597;
wire n_14918;
wire n_11002;
wire n_13716;
wire n_9691;
wire n_5110;
wire n_16223;
wire n_6653;
wire n_16045;
wire n_12165;
wire n_15970;
wire n_4719;
wire n_4178;
wire n_7450;
wire n_5425;
wire n_13803;
wire n_14455;
wire n_10532;
wire n_8832;
wire n_15583;
wire n_15614;
wire n_5737;
wire n_15178;
wire n_16151;
wire n_9340;
wire n_10350;
wire n_9351;
wire n_8461;
wire n_8042;
wire n_10977;
wire n_11179;
wire n_15128;
wire n_6923;
wire n_6825;
wire n_11708;
wire n_15108;
wire n_10418;
wire n_9950;
wire n_11474;
wire n_15889;
wire n_10336;
wire n_4228;
wire n_4401;
wire n_8021;
wire n_8839;
wire n_12092;
wire n_11369;
wire n_6112;
wire n_6547;
wire n_11738;
wire n_11240;
wire n_14113;
wire n_6198;
wire n_13155;
wire n_7439;
wire n_5560;
wire n_15483;
wire n_12074;
wire n_9155;
wire n_14565;
wire n_11931;
wire n_14231;
wire n_15841;
wire n_10925;
wire n_6399;
wire n_8623;
wire n_15277;
wire n_12109;
wire n_11438;
wire n_8758;
wire n_14508;
wire n_6275;
wire n_5666;
wire n_6575;
wire n_10609;
wire n_13508;
wire n_7924;
wire n_7732;
wire n_6151;
wire n_13058;
wire n_5179;
wire n_7227;
wire n_7040;
wire n_4605;
wire n_15042;
wire n_4877;
wire n_8511;
wire n_7325;
wire n_6469;
wire n_4968;
wire n_6756;
wire n_8595;
wire n_12900;
wire n_8873;
wire n_11376;
wire n_5030;
wire n_13055;
wire n_5961;
wire n_7191;
wire n_7459;
wire n_9201;
wire n_9823;
wire n_11051;
wire n_11812;
wire n_14304;
wire n_9688;
wire n_12330;
wire n_15530;
wire n_7096;
wire n_12519;
wire n_13872;
wire n_13597;
wire n_8455;
wire n_11838;
wire n_12717;
wire n_8280;
wire n_10102;
wire n_4834;
wire n_10908;
wire n_11333;
wire n_9595;
wire n_5272;
wire n_15119;
wire n_9530;
wire n_4158;
wire n_6826;
wire n_9227;
wire n_6015;
wire n_8372;
wire n_8598;
wire n_5361;
wire n_5683;
wire n_10939;
wire n_4171;
wire n_13503;
wire n_11178;
wire n_12595;
wire n_5847;
wire n_7551;
wire n_9400;
wire n_6678;
wire n_11188;
wire n_4562;
wire n_5068;
wire n_9025;
wire n_5740;
wire n_13086;
wire n_8282;
wire n_7750;
wire n_10936;
wire n_11840;
wire n_5015;
wire n_12525;
wire n_7697;
wire n_5729;
wire n_7485;
wire n_11685;
wire n_10955;
wire n_13093;
wire n_10824;
wire n_6748;
wire n_15673;
wire n_12084;
wire n_8616;
wire n_4749;
wire n_10440;
wire n_10630;
wire n_8336;
wire n_4390;
wire n_5302;
wire n_4979;
wire n_11472;
wire n_6752;
wire n_9749;
wire n_14404;
wire n_4804;
wire n_5545;
wire n_6553;
wire n_9285;
wire n_12997;
wire n_11295;
wire n_9972;
wire n_10058;
wire n_7652;
wire n_14533;
wire n_8847;
wire n_7808;
wire n_11171;
wire n_6500;
wire n_4270;
wire n_8135;
wire n_9214;
wire n_13299;
wire n_7051;
wire n_9859;
wire n_11030;
wire n_13394;
wire n_10295;
wire n_5152;
wire n_9003;
wire n_11443;
wire n_9271;
wire n_9258;
wire n_6628;
wire n_13849;
wire n_12661;
wire n_12693;
wire n_6297;
wire n_5905;
wire n_12203;
wire n_6975;
wire n_5409;
wire n_6329;
wire n_7536;
wire n_8979;
wire n_12080;
wire n_8529;
wire n_15514;
wire n_10658;
wire n_5688;
wire n_9763;
wire n_5128;
wire n_10894;
wire n_4566;
wire n_9597;
wire n_6293;
wire n_8417;
wire n_9965;
wire n_9076;
wire n_10912;
wire n_7952;
wire n_4576;
wire n_9393;
wire n_8498;
wire n_7991;
wire n_7676;
wire n_11769;
wire n_16052;
wire n_12486;
wire n_7553;
wire n_6905;
wire n_12623;
wire n_7425;
wire n_13698;
wire n_5798;
wire n_6381;
wire n_6521;
wire n_14701;
wire n_5307;
wire n_12933;
wire n_12489;
wire n_8967;
wire n_8355;
wire n_9736;
wire n_4767;
wire n_13691;
wire n_7998;
wire n_14122;
wire n_4328;
wire n_5986;
wire n_8719;
wire n_16098;
wire n_6581;
wire n_10160;
wire n_10678;
wire n_14372;
wire n_6215;
wire n_7095;
wire n_11794;
wire n_14645;
wire n_15901;
wire n_5415;
wire n_4676;
wire n_10241;
wire n_5770;
wire n_11495;
wire n_14259;
wire n_7064;
wire n_5892;
wire n_8762;
wire n_12480;
wire n_13273;
wire n_4544;
wire n_13265;
wire n_10180;
wire n_8516;
wire n_8880;
wire n_6577;
wire n_6899;
wire n_8784;
wire n_14666;
wire n_12335;
wire n_5676;
wire n_7307;
wire n_6545;
wire n_10631;
wire n_8237;
wire n_5802;
wire n_13372;
wire n_15897;
wire n_10852;
wire n_14546;
wire n_13669;
wire n_9803;
wire n_4429;
wire n_8977;
wire n_13079;
wire n_14371;
wire n_11406;
wire n_8171;
wire n_13121;
wire n_4591;
wire n_10978;
wire n_10500;
wire n_6370;
wire n_9755;
wire n_9805;
wire n_13731;
wire n_15634;
wire n_7210;
wire n_14997;
wire n_4646;
wire n_7899;
wire n_10370;
wire n_15263;
wire n_15836;
wire n_9728;
wire n_5769;
wire n_6065;
wire n_13845;
wire n_15475;
wire n_16051;
wire n_7039;
wire n_9659;
wire n_6987;
wire n_12624;
wire n_14328;
wire n_4563;
wire n_4725;
wire n_9107;
wire n_11428;
wire n_14361;
wire n_4169;
wire n_6190;
wire n_6859;
wire n_5331;
wire n_14311;
wire n_13447;
wire n_12410;
wire n_9917;
wire n_14574;
wire n_14847;
wire n_6309;
wire n_11149;
wire n_9520;
wire n_6623;
wire n_12055;
wire n_12925;
wire n_7723;
wire n_15922;
wire n_12771;
wire n_6527;
wire n_7443;
wire n_16014;
wire n_13262;
wire n_11707;
wire n_10550;
wire n_9583;
wire n_7811;
wire n_12413;
wire n_11086;
wire n_5341;
wire n_4320;
wire n_12182;
wire n_14096;
wire n_15315;
wire n_14943;
wire n_5930;
wire n_13622;
wire n_5814;
wire n_12803;
wire n_4881;
wire n_9036;
wire n_14007;
wire n_15026;
wire n_9522;
wire n_13145;
wire n_16134;
wire n_5979;
wire n_14034;
wire n_5271;
wire n_5089;
wire n_10571;
wire n_7015;
wire n_5263;
wire n_13276;
wire n_14394;
wire n_11772;
wire n_13338;
wire n_14618;
wire n_15806;
wire n_16008;
wire n_12547;
wire n_6929;
wire n_11225;
wire n_11764;
wire n_13904;
wire n_14256;
wire n_12544;
wire n_11339;
wire n_5518;
wire n_10125;
wire n_5637;
wire n_4636;
wire n_12370;
wire n_4584;
wire n_12931;
wire n_14810;
wire n_8279;
wire n_5622;
wire n_13940;
wire n_14054;
wire n_13648;
wire n_14844;
wire n_4711;
wire n_11112;
wire n_9723;
wire n_12986;
wire n_13570;
wire n_7348;
wire n_10254;
wire n_5240;
wire n_5813;
wire n_15589;
wire n_13543;
wire n_5495;
wire n_4680;
wire n_5546;
wire n_8912;
wire n_13873;
wire n_14491;
wire n_9488;
wire n_7143;
wire n_5482;
wire n_7312;
wire n_4191;
wire n_5224;
wire n_4293;
wire n_14267;
wire n_7155;
wire n_8227;
wire n_9231;
wire n_8938;
wire n_15116;
wire n_6865;
wire n_8787;
wire n_16238;
wire n_5393;
wire n_10017;
wire n_6535;
wire n_7213;
wire n_15774;
wire n_14987;
wire n_10866;
wire n_9047;
wire n_10348;
wire n_14846;
wire n_12991;
wire n_4671;
wire n_8270;
wire n_4209;
wire n_5966;
wire n_11072;
wire n_7456;
wire n_8335;
wire n_11359;
wire n_13449;
wire n_13459;
wire n_13781;
wire n_14974;
wire n_10657;
wire n_13899;
wire n_7420;
wire n_5041;
wire n_14223;
wire n_11605;
wire n_15871;
wire n_13395;
wire n_9798;
wire n_14463;
wire n_9681;
wire n_8054;
wire n_9414;
wire n_12419;
wire n_8607;
wire n_5431;
wire n_13760;
wire n_9979;
wire n_9093;
wire n_15677;
wire n_14151;
wire n_11959;
wire n_6482;
wire n_5026;
wire n_15487;
wire n_11830;
wire n_11318;
wire n_10842;
wire n_15428;
wire n_13012;
wire n_15148;
wire n_12865;
wire n_8150;
wire n_9379;
wire n_5059;
wire n_5505;
wire n_7715;
wire n_9486;
wire n_11881;
wire n_6605;
wire n_4250;
wire n_9134;
wire n_5329;
wire n_15210;
wire n_12481;
wire n_4699;
wire n_7007;
wire n_8358;
wire n_9410;
wire n_4127;
wire n_10045;
wire n_14672;
wire n_13594;
wire n_13991;
wire n_15408;
wire n_7909;
wire n_14751;
wire n_15133;
wire n_14307;
wire n_9151;
wire n_12278;
wire n_13102;
wire n_4292;
wire n_14407;
wire n_4577;
wire n_11863;
wire n_14715;
wire n_15595;
wire n_14563;
wire n_13558;
wire n_4854;
wire n_14428;
wire n_8281;
wire n_12562;
wire n_11494;
wire n_9182;
wire n_5908;
wire n_6018;
wire n_12744;
wire n_4202;
wire n_7168;
wire n_11850;
wire n_5212;
wire n_9976;
wire n_7736;
wire n_5000;
wire n_14107;
wire n_8396;
wire n_9591;
wire n_10322;
wire n_13952;
wire n_9838;
wire n_7177;
wire n_5939;
wire n_10033;
wire n_12615;
wire n_13027;
wire n_14478;
wire n_11258;
wire n_9568;
wire n_7780;
wire n_10886;
wire n_15956;
wire n_9261;
wire n_9701;
wire n_7379;
wire n_4165;
wire n_4866;
wire n_7444;
wire n_8223;
wire n_5931;
wire n_11468;
wire n_7435;
wire n_4109;
wire n_5297;
wire n_7813;
wire n_7030;
wire n_8459;
wire n_5420;
wire n_16027;
wire n_6311;
wire n_11192;
wire n_12580;
wire n_11569;
wire n_4412;
wire n_6654;
wire n_6424;
wire n_6816;
wire n_6220;
wire n_9752;
wire n_12769;
wire n_5234;
wire n_6740;
wire n_7122;
wire n_12540;
wire n_5835;
wire n_7049;
wire n_7567;
wire n_6029;
wire n_13607;
wire n_15807;
wire n_13080;
wire n_8379;
wire n_11563;
wire n_15089;
wire n_6879;
wire n_13292;
wire n_5259;
wire n_5440;
wire n_5679;
wire n_5938;
wire n_9079;
wire n_6702;
wire n_4155;
wire n_11846;
wire n_5891;
wire n_14682;
wire n_10383;
wire n_13377;
wire n_4144;
wire n_5724;
wire n_10064;
wire n_10876;
wire n_5774;
wire n_8793;
wire n_11852;
wire n_6452;
wire n_15637;
wire n_4374;
wire n_12619;
wire n_14527;
wire n_8975;
wire n_14020;
wire n_6791;
wire n_11679;
wire n_9170;
wire n_8792;
wire n_5131;
wire n_7280;
wire n_8671;
wire n_8489;
wire n_6915;
wire n_7110;
wire n_7511;
wire n_10831;
wire n_6856;
wire n_7941;
wire n_7791;
wire n_9385;
wire n_11186;
wire n_11870;
wire n_12960;
wire n_13519;
wire n_8484;
wire n_8454;
wire n_11492;
wire n_13984;
wire n_10536;
wire n_10238;
wire n_7232;
wire n_8759;
wire n_12268;
wire n_11544;
wire n_4548;
wire n_7345;
wire n_5923;
wire n_8703;
wire n_11233;
wire n_12656;
wire n_15193;
wire n_5790;
wire n_12678;
wire n_14521;
wire n_10206;
wire n_14726;
wire n_4989;
wire n_14924;
wire n_4622;
wire n_4315;
wire n_12880;
wire n_9670;
wire n_12876;
wire n_6364;
wire n_6451;
wire n_13107;
wire n_12711;
wire n_13511;
wire n_6552;
wire n_14205;
wire n_15667;
wire n_15168;
wire n_10786;
wire n_8325;
wire n_13523;
wire n_6328;
wire n_5140;
wire n_9598;
wire n_4816;
wire n_8382;
wire n_7827;
wire n_8971;
wire n_15815;
wire n_6363;
wire n_11646;
wire n_10602;
wire n_10620;
wire n_13699;
wire n_14049;
wire n_16049;
wire n_13420;
wire n_7159;
wire n_8127;
wire n_11878;
wire n_10079;
wire n_10188;
wire n_8721;
wire n_9391;
wire n_15751;
wire n_12458;
wire n_6132;
wire n_6578;
wire n_8889;
wire n_6406;
wire n_10319;
wire n_5598;
wire n_13643;
wire n_13603;
wire n_11900;
wire n_9470;
wire n_12132;
wire n_14434;
wire n_15429;
wire n_5306;
wire n_6978;
wire n_12104;
wire n_12037;
wire n_9328;
wire n_12467;
wire n_4483;
wire n_12870;
wire n_5342;
wire n_9245;
wire n_16156;
wire n_10739;
wire n_12911;
wire n_8232;
wire n_4358;
wire n_7477;
wire n_5147;
wire n_6918;
wire n_12386;
wire n_7363;
wire n_4793;
wire n_9833;
wire n_11837;
wire n_10213;
wire n_6612;
wire n_15588;
wire n_10107;
wire n_8664;
wire n_5677;
wire n_4168;
wire n_10872;
wire n_5997;
wire n_9455;
wire n_12651;
wire n_5511;
wire n_7863;
wire n_9719;
wire n_5680;
wire n_4806;
wire n_4350;
wire n_7295;
wire n_8633;
wire n_9744;
wire n_8842;
wire n_15900;
wire n_5533;
wire n_5838;
wire n_6058;
wire n_11871;
wire n_8956;
wire n_5280;
wire n_10969;
wire n_6375;
wire n_6479;
wire n_14507;
wire n_6866;
wire n_12563;
wire n_7831;
wire n_13825;
wire n_11674;
wire n_12621;
wire n_5235;
wire n_15234;
wire n_13798;
wire n_14564;
wire n_12331;
wire n_12304;
wire n_9698;
wire n_12339;
wire n_6170;
wire n_12270;
wire n_14599;
wire n_15049;
wire n_9124;
wire n_10669;
wire n_10718;
wire n_9695;
wire n_4187;
wire n_4166;
wire n_6447;
wire n_6263;
wire n_7093;
wire n_9497;
wire n_5206;
wire n_10895;
wire n_8641;
wire n_15903;
wire n_8479;
wire n_11610;
wire n_15983;
wire n_11187;
wire n_12210;
wire n_7466;
wire n_14525;
wire n_16246;
wire n_14058;
wire n_15249;
wire n_15255;
wire n_5419;
wire n_6130;
wire n_12858;
wire n_14153;
wire n_15101;
wire n_12382;
wire n_11280;
wire n_10757;
wire n_7651;
wire n_4937;
wire n_13324;
wire n_10513;
wire n_15018;
wire n_5103;
wire n_11148;
wire n_8179;
wire n_15825;
wire n_5803;
wire n_13286;
wire n_4258;
wire n_14272;
wire n_6014;
wire n_4498;
wire n_11396;
wire n_8973;
wire n_6935;
wire n_14953;
wire n_10194;
wire n_9775;
wire n_7530;
wire n_5285;
wire n_11426;
wire n_14980;
wire n_9038;
wire n_8308;
wire n_15537;
wire n_4936;
wire n_13406;
wire n_5387;
wire n_9630;
wire n_13071;
wire n_10692;
wire n_16164;
wire n_8378;
wire n_8733;
wire n_12107;
wire n_14337;
wire n_8809;
wire n_14427;
wire n_4770;
wire n_5985;
wire n_14439;
wire n_11723;
wire n_11009;
wire n_4907;
wire n_9652;
wire n_10021;
wire n_5058;
wire n_12381;
wire n_6907;
wire n_11706;
wire n_13284;
wire n_8500;
wire n_12653;
wire n_6158;
wire n_7661;
wire n_10782;
wire n_9709;
wire n_6541;
wire n_6119;
wire n_8447;
wire n_14202;
wire n_5018;
wire n_11949;
wire n_5896;
wire n_4861;
wire n_13303;
wire n_15004;
wire n_10457;
wire n_9324;
wire n_13311;
wire n_9934;
wire n_13364;
wire n_13813;
wire n_11957;
wire n_5192;
wire n_8548;
wire n_11538;
wire n_5141;
wire n_14743;
wire n_5133;
wire n_8412;
wire n_6226;
wire n_4712;
wire n_11264;
wire n_12774;
wire n_11211;
wire n_11880;
wire n_9668;
wire n_14340;
wire n_7145;
wire n_10385;
wire n_15526;
wire n_11377;
wire n_12064;
wire n_9877;
wire n_4310;
wire n_12503;
wire n_9657;
wire n_10111;
wire n_11302;
wire n_6338;
wire n_12425;
wire n_14319;
wire n_14922;
wire n_15181;
wire n_11921;
wire n_13358;
wire n_5159;
wire n_15248;
wire n_9352;
wire n_15917;
wire n_9395;
wire n_12807;
wire n_14621;
wire n_15211;
wire n_8425;
wire n_10809;
wire n_9349;
wire n_4674;
wire n_4908;
wire n_14734;
wire n_8241;
wire n_7823;
wire n_15268;
wire n_9209;
wire n_7467;
wire n_5097;
wire n_14555;
wire n_10113;
wire n_15010;
wire n_11267;
wire n_10990;
wire n_7932;
wire n_11626;
wire n_14957;
wire n_15308;
wire n_5730;
wire n_7550;
wire n_11694;
wire n_13811;
wire n_14014;
wire n_4159;
wire n_16109;
wire n_11618;
wire n_9969;
wire n_9937;
wire n_15754;
wire n_5816;
wire n_7541;
wire n_10545;
wire n_12715;
wire n_4862;
wire n_7241;
wire n_7717;
wire n_14945;
wire n_5300;
wire n_10595;
wire n_10973;
wire n_13883;
wire n_11011;
wire n_13814;
wire n_12015;
wire n_12968;
wire n_9618;
wire n_10732;
wire n_14257;
wire n_10009;
wire n_11776;
wire n_4850;
wire n_6625;
wire n_11165;
wire n_4813;
wire n_4912;
wire n_12135;
wire n_7464;
wire n_9082;
wire n_11366;
wire n_6302;
wire n_14279;
wire n_9424;
wire n_8274;
wire n_9453;
wire n_15239;
wire n_5748;
wire n_13757;
wire n_6759;
wire n_16199;
wire n_5525;
wire n_9637;
wire n_8152;
wire n_6706;
wire n_10526;
wire n_8550;
wire n_6139;
wire n_14190;
wire n_4256;
wire n_14185;
wire n_8264;
wire n_7434;
wire n_7636;
wire n_6999;
wire n_7054;
wire n_12817;
wire n_13832;
wire n_4224;
wire n_6403;
wire n_6483;
wire n_9183;
wire n_8829;
wire n_9205;
wire n_14630;
wire n_13935;
wire n_12869;
wire n_9009;
wire n_13325;
wire n_15764;
wire n_13841;
wire n_6228;
wire n_11315;
wire n_5650;
wire n_14104;
wire n_14344;
wire n_10044;
wire n_16181;
wire n_13207;
wire n_12059;
wire n_14188;
wire n_15482;
wire n_16219;
wire n_12586;
wire n_11098;
wire n_5400;
wire n_13043;
wire n_4415;
wire n_5552;
wire n_7299;
wire n_10221;
wire n_4702;
wire n_13281;
wire n_6888;
wire n_8266;
wire n_13960;
wire n_15086;
wire n_14069;
wire n_8515;
wire n_10109;
wire n_10169;
wire n_4252;
wire n_13556;
wire n_4457;
wire n_8648;
wire n_15707;
wire n_6063;
wire n_10329;
wire n_10928;
wire n_9030;
wire n_9024;
wire n_9523;
wire n_15875;
wire n_9377;
wire n_10891;
wire n_8946;
wire n_15099;
wire n_16074;
wire n_10839;
wire n_11875;
wire n_6800;
wire n_5139;
wire n_13260;
wire n_9716;
wire n_6922;
wire n_9380;
wire n_14543;
wire n_6890;
wire n_5481;
wire n_14474;
wire n_8744;
wire n_9000;
wire n_9679;
wire n_9116;
wire n_9742;
wire n_9016;
wire n_7503;
wire n_6070;
wire n_13979;
wire n_13308;
wire n_9006;
wire n_12514;
wire n_13381;
wire n_11524;
wire n_10091;
wire n_6651;
wire n_5821;
wire n_7091;
wire n_7296;
wire n_7273;
wire n_6647;
wire n_4491;
wire n_5733;
wire n_14704;
wire n_10029;
wire n_9690;
wire n_8765;
wire n_15183;
wire n_4132;
wire n_13483;
wire n_14675;
wire n_5871;
wire n_9852;
wire n_7543;
wire n_4261;
wire n_13400;
wire n_10600;
wire n_15424;
wire n_9914;
wire n_11056;
wire n_11514;
wire n_12438;
wire n_6184;
wire n_14268;
wire n_16157;
wire n_4886;
wire n_11774;
wire n_8627;
wire n_7507;
wire n_9451;
wire n_10849;
wire n_15456;
wire n_5043;
wire n_15466;
wire n_11108;
wire n_9760;
wire n_7555;
wire n_15509;
wire n_13910;
wire n_15874;
wire n_5707;
wire n_13907;
wire n_10947;
wire n_13369;
wire n_10272;
wire n_12099;
wire n_9035;
wire n_12009;
wire n_12806;
wire n_4371;
wire n_5836;
wire n_9211;
wire n_15077;
wire n_5281;
wire n_14873;
wire n_6716;
wire n_16043;
wire n_6422;
wire n_12887;
wire n_12776;
wire n_4473;
wire n_12898;
wire n_4268;
wire n_9677;
wire n_13464;
wire n_5048;
wire n_11954;
wire n_14965;
wire n_5521;
wire n_12191;
wire n_7578;
wire n_5028;
wire n_13611;
wire n_4480;
wire n_7475;
wire n_4194;
wire n_8195;
wire n_9070;
wire n_5585;
wire n_6397;
wire n_12578;
wire n_4824;
wire n_4120;
wire n_14012;
wire n_4427;
wire n_11864;
wire n_14221;
wire n_14232;
wire n_7033;
wire n_9881;
wire n_6121;
wire n_16010;
wire n_9669;
wire n_7531;
wire n_4142;
wire n_9958;
wire n_9858;
wire n_8462;
wire n_5561;
wire n_9981;
wire n_10391;
wire n_4260;
wire n_8377;
wire n_11157;
wire n_14390;
wire n_4163;
wire n_4439;
wire n_12509;
wire n_13345;
wire n_12235;
wire n_6981;
wire n_15647;
wire n_4372;
wire n_14932;
wire n_15666;
wire n_9588;
wire n_6954;
wire n_11733;
wire n_5799;
wire n_5073;
wire n_5024;
wire n_12471;
wire n_13632;
wire n_13756;
wire n_15208;
wire n_12365;
wire n_5875;
wire n_8428;
wire n_8103;
wire n_13417;
wire n_4262;
wire n_14350;
wire n_9021;
wire n_13130;
wire n_6646;
wire n_8936;
wire n_8414;
wire n_8362;
wire n_15529;
wire n_12083;
wire n_15251;
wire n_9682;
wire n_10137;
wire n_10344;
wire n_7131;
wire n_4720;
wire n_7769;
wire n_10882;
wire n_11540;
wire n_11861;
wire n_15397;
wire n_6903;
wire n_9050;
wire n_11724;
wire n_9303;
wire n_14775;
wire n_12065;
wire n_9495;
wire n_13970;
wire n_15156;
wire n_15971;
wire n_12167;
wire n_11220;
wire n_14220;
wire n_4685;
wire n_6101;
wire n_9415;
wire n_5968;
wire n_14451;
wire n_10196;
wire n_8491;
wire n_9058;
wire n_4334;
wire n_6941;
wire n_9845;
wire n_8831;
wire n_4511;
wire n_5812;
wire n_14100;
wire n_6148;
wire n_15704;
wire n_5515;
wire n_8324;
wire n_11459;
wire n_11355;
wire n_6106;
wire n_9822;
wire n_12087;
wire n_6604;
wire n_14510;
wire n_12243;
wire n_7418;
wire n_12267;
wire n_5250;
wire n_12569;
wire n_4757;
wire n_7688;
wire n_10518;
wire n_11101;
wire n_9640;
wire n_11899;
wire n_8348;
wire n_5607;
wire n_14313;
wire n_15842;
wire n_4175;
wire n_8288;
wire n_10613;
wire n_15688;
wire n_10583;
wire n_14719;
wire n_4648;
wire n_14452;
wire n_15447;
wire n_11481;
wire n_14308;
wire n_16046;
wire n_11712;
wire n_11612;
wire n_8269;
wire n_5006;
wire n_14288;
wire n_7806;
wire n_10335;
wire n_10085;
wire n_10840;
wire n_6566;
wire n_14833;
wire n_13152;
wire n_12599;
wire n_8625;
wire n_5734;
wire n_6081;
wire n_8458;
wire n_4892;
wire n_8806;
wire n_13857;
wire n_7204;
wire n_16071;
wire n_10560;
wire n_8180;
wire n_16160;
wire n_4173;
wire n_8601;
wire n_8499;
wire n_4970;
wire n_9062;
wire n_13315;
wire n_14606;
wire n_13180;
wire n_14097;
wire n_5404;
wire n_4108;
wire n_4486;
wire n_8306;
wire n_15510;
wire n_12375;
wire n_12091;
wire n_9722;
wire n_12513;
wire n_6047;
wire n_14788;
wire n_8167;
wire n_5438;
wire n_10486;
wire n_9791;
wire n_12307;
wire n_16086;
wire n_9229;
wire n_11603;
wire n_11890;
wire n_4627;
wire n_8613;
wire n_9603;
wire n_11790;
wire n_8913;
wire n_11060;
wire n_7354;
wire n_7448;
wire n_15550;
wire n_8800;
wire n_16047;
wire n_6244;
wire n_13474;
wire n_13224;
wire n_16212;
wire n_12684;
wire n_8768;
wire n_6861;
wire n_13702;
wire n_9099;
wire n_10919;
wire n_13797;
wire n_14388;
wire n_12288;
wire n_9309;
wire n_12418;
wire n_13853;
wire n_7852;
wire n_13762;
wire n_15957;
wire n_10952;
wire n_5725;
wire n_12566;
wire n_7925;
wire n_12415;
wire n_13037;
wire n_9432;
wire n_16054;
wire n_9454;
wire n_4249;
wire n_7571;
wire n_15351;
wire n_11744;
wire n_13919;
wire n_14466;
wire n_9065;
wire n_11650;
wire n_5163;
wire n_11518;
wire n_7748;
wire n_5768;
wire n_12949;
wire n_4961;
wire n_7556;
wire n_14061;
wire n_7640;
wire n_8187;
wire n_10352;
wire n_14962;
wire n_15365;
wire n_8881;
wire n_9704;
wire n_4718;
wire n_15615;
wire n_11663;
wire n_5190;
wire n_7422;
wire n_7920;
wire n_8433;
wire n_9837;
wire n_10991;
wire n_4317;
wire n_4855;
wire n_9431;
wire n_10167;
wire n_12681;
wire n_12859;
wire n_14413;
wire n_9160;
wire n_10911;
wire n_4154;
wire n_9433;
wire n_14050;
wire n_15587;
wire n_6588;
wire n_9256;
wire n_10442;
wire n_12829;
wire n_13593;
wire n_11282;
wire n_14912;
wire n_9706;
wire n_12448;
wire n_13044;
wire n_7900;
wire n_7050;
wire n_9808;
wire n_9915;
wire n_13723;
wire n_10534;
wire n_14156;
wire n_5685;
wire n_4420;
wire n_11726;
wire n_13188;
wire n_5773;
wire n_7136;
wire n_10465;
wire n_10406;
wire n_12188;
wire n_12943;
wire n_8316;
wire n_7318;
wire n_13923;
wire n_12149;
wire n_6055;
wire n_5138;
wire n_12783;
wire n_8397;
wire n_9184;
wire n_15136;
wire n_5374;
wire n_10373;
wire n_13472;
wire n_9133;
wire n_6108;
wire n_8115;
wire n_12129;
wire n_12631;
wire n_6165;
wire n_14387;
wire n_10965;
wire n_6621;
wire n_13148;
wire n_7175;
wire n_5349;
wire n_15645;
wire n_4973;
wire n_7810;
wire n_9109;
wire n_4640;
wire n_13964;
wire n_10517;
wire n_6323;
wire n_12588;
wire n_12652;
wire n_8523;
wire n_9207;
wire n_11458;
wire n_4396;
wire n_13485;
wire n_5127;
wire n_6587;
wire n_4367;
wire n_16214;
wire n_6480;
wire n_13531;
wire n_13355;
wire n_13368;
wire n_7733;
wire n_6731;
wire n_5485;
wire n_13160;
wire n_10484;
wire n_5766;
wire n_11255;
wire n_6597;
wire n_5216;
wire n_13676;
wire n_16004;
wire n_10561;
wire n_13183;
wire n_9673;
wire n_13601;
wire n_15282;
wire n_8891;
wire n_12523;
wire n_7817;
wire n_8294;
wire n_11856;
wire n_14312;
wire n_6933;
wire n_4387;
wire n_7878;
wire n_8338;
wire n_15176;
wire n_15972;
wire n_4951;
wire n_12579;
wire n_9010;
wire n_14904;
wire n_8915;
wire n_4453;
wire n_4170;
wire n_6881;
wire n_11442;
wire n_13052;
wire n_7289;
wire n_14754;
wire n_5805;
wire n_7665;
wire n_8131;
wire n_11747;
wire n_9552;
wire n_7855;
wire n_11008;
wire n_10371;
wire n_11243;
wire n_12675;
wire n_9841;
wire n_13006;
wire n_12174;
wire n_9230;
wire n_14947;
wire n_14659;
wire n_7764;
wire n_4308;
wire n_15747;
wire n_12113;
wire n_12831;
wire n_15516;
wire n_10198;
wire n_8027;
wire n_6216;
wire n_10096;
wire n_10582;
wire n_11425;
wire n_10638;
wire n_8162;
wire n_6817;
wire n_7170;
wire n_7314;
wire n_9132;
wire n_11992;
wire n_6949;
wire n_6509;
wire n_14198;
wire n_15882;
wire n_5175;
wire n_7260;
wire n_8855;
wire n_10483;
wire n_11657;
wire n_4152;
wire n_13820;
wire n_12470;
wire n_14039;
wire n_8546;
wire n_9878;
wire n_11536;
wire n_11717;
wire n_9069;
wire n_8966;
wire n_12154;
wire n_15323;
wire n_8487;
wire n_7263;
wire n_8844;
wire n_14995;
wire n_5948;
wire n_4392;
wire n_4660;
wire n_5611;
wire n_10662;
wire n_13471;
wire n_15817;
wire n_6911;
wire n_9674;
wire n_11512;
wire n_11327;
wire n_8533;
wire n_4281;
wire n_4661;
wire n_12799;
wire n_15555;
wire n_4200;
wire n_13114;
wire n_15002;
wire n_8869;
wire n_5900;
wire n_15860;
wire n_4962;
wire n_14956;
wire n_15731;
wire n_15684;
wire n_9786;
wire n_13976;
wire n_6327;
wire n_8584;
wire n_13200;
wire n_11140;
wire n_8932;
wire n_14862;
wire n_9063;
wire n_8998;
wire n_6607;
wire n_15833;
wire n_9188;
wire n_9467;
wire n_15652;
wire n_9372;
wire n_10960;
wire n_11078;
wire n_4958;
wire n_9743;
wire n_4271;
wire n_7850;
wire n_7509;
wire n_11620;
wire n_7209;
wire n_5171;
wire n_15592;
wire n_12617;
wire n_6401;
wire n_5554;
wire n_6227;
wire n_12919;
wire n_8480;
wire n_9926;
wire n_7240;
wire n_10094;
wire n_12095;
wire n_14620;
wire n_10749;
wire n_11907;
wire n_14291;
wire n_15933;
wire n_4921;
wire n_14092;
wire n_12432;
wire n_12796;
wire n_8911;
wire n_11352;
wire n_5427;
wire n_15876;
wire n_5639;
wire n_14293;
wire n_7725;
wire n_8398;
wire n_4361;
wire n_10585;
wire n_15039;
wire n_5417;
wire n_8772;
wire n_12279;
wire n_4614;
wire n_12008;
wire n_9480;
wire n_8307;
wire n_14005;
wire n_14884;
wire n_10896;
wire n_8767;
wire n_15273;
wire n_9113;
wire n_13764;
wire n_9158;
wire n_12156;
wire n_11851;
wire n_4945;
wire n_14441;
wire n_4922;
wire n_4732;
wire n_7609;
wire n_14688;
wire n_15827;
wire n_13264;
wire n_8010;
wire n_7278;
wire n_11986;
wire n_12637;
wire n_15878;
wire n_15965;
wire n_12301;
wire n_9263;
wire n_8347;
wire n_11734;
wire n_7630;
wire n_11517;
wire n_11022;
wire n_14468;
wire n_11831;
wire n_14766;
wire n_10162;
wire n_12302;
wire n_8466;
wire n_6416;
wire n_5488;
wire n_4693;
wire n_12190;
wire n_14222;
wire n_15054;
wire n_9632;
wire n_10353;
wire n_8813;
wire n_8354;
wire n_4326;
wire n_8204;
wire n_6695;
wire n_14067;
wire n_7741;
wire n_5447;
wire n_5383;
wire n_4744;
wire n_14598;
wire n_6127;
wire n_7565;
wire n_11259;
wire n_14446;
wire n_11197;
wire n_9282;
wire n_4305;
wire n_14747;
wire n_14909;
wire n_15635;
wire n_5781;
wire n_15403;
wire n_7883;
wire n_6600;
wire n_10933;
wire n_12192;
wire n_7410;
wire n_12010;
wire n_12977;
wire n_4213;
wire n_10546;
wire n_7097;
wire n_12864;
wire n_13227;
wire n_13869;
wire n_9503;
wire n_6421;
wire n_10724;
wire n_5747;
wire n_7414;
wire n_15486;
wire n_11427;
wire n_10660;
wire n_13348;
wire n_13166;
wire n_7495;
wire n_9782;
wire n_5969;
wire n_13350;
wire n_9114;
wire n_8312;
wire n_9855;
wire n_4929;
wire n_15400;
wire n_8040;
wire n_14242;
wire n_11153;
wire n_9347;
wire n_4964;
wire n_13615;
wire n_9469;
wire n_9680;
wire n_9746;
wire n_10923;
wire n_6079;
wire n_4802;
wire n_6192;
wire n_9633;
wire n_12746;
wire n_15452;
wire n_10836;
wire n_13266;
wire n_6458;
wire n_10884;
wire n_4139;
wire n_13319;
wire n_13623;
wire n_15062;
wire n_15698;
wire n_6746;
wire n_8132;
wire n_12436;
wire n_7586;
wire n_10780;
wire n_9501;
wire n_12528;
wire n_7720;
wire n_6719;
wire n_13544;
wire n_12792;
wire n_15556;
wire n_14586;
wire n_5437;
wire n_9148;
wire n_15417;
wire n_15959;
wire n_13530;
wire n_11475;
wire n_5826;
wire n_7659;
wire n_12973;
wire n_14095;
wire n_11385;
wire n_14191;
wire n_6506;
wire n_14289;
wire n_4583;
wire n_6287;
wire n_13092;
wire n_6662;
wire n_8650;
wire n_12923;
wire n_10870;
wire n_12916;
wire n_16202;
wire n_9585;
wire n_10267;
wire n_13888;
wire n_8974;
wire n_10379;
wire n_4210;
wire n_5245;
wire n_14561;
wire n_7189;
wire n_8688;
wire n_4666;
wire n_10821;
wire n_10740;
wire n_16108;
wire n_8983;
wire n_10558;
wire n_6851;
wire n_8116;
wire n_12144;
wire n_9338;
wire n_12716;
wire n_6687;
wire n_10297;
wire n_6884;
wire n_8356;
wire n_8013;
wire n_9075;
wire n_13981;
wire n_14614;
wire n_4540;
wire n_6780;
wire n_6513;
wire n_12463;
wire n_12524;
wire n_16216;
wire n_4891;
wire n_8519;
wire n_14484;
wire n_7841;
wire n_15399;
wire n_10497;
wire n_6619;
wire n_10354;
wire n_11456;
wire n_8193;
wire n_15620;
wire n_14536;
wire n_5603;
wire n_10888;
wire n_6804;
wire n_9370;
wire n_15717;
wire n_11647;
wire n_12392;
wire n_13205;
wire n_13421;
wire n_12173;
wire n_9409;
wire n_14140;
wire n_5716;
wire n_10138;
wire n_4940;
wire n_6516;
wire n_10358;
wire n_5208;
wire n_7490;
wire n_7792;
wire n_10578;
wire n_15902;
wire n_6924;
wire n_4590;
wire n_13745;
wire n_7492;
wire n_12168;
wire n_12349;
wire n_13349;
wire n_10948;
wire n_5606;
wire n_13730;
wire n_15087;
wire n_4830;
wire n_12665;
wire n_5231;
wire n_8329;
wire n_5237;
wire n_7809;
wire n_11736;
wire n_14339;
wire n_14804;
wire n_4664;
wire n_9626;
wire n_14501;
wire n_16073;
wire n_8154;
wire n_15007;
wire n_12067;
wire n_5456;
wire n_12546;
wire n_7073;
wire n_13489;
wire n_14825;
wire n_11393;
wire n_10007;
wire n_5093;
wire n_10904;
wire n_10386;
wire n_6040;
wire n_4946;
wire n_15125;
wire n_15479;
wire n_9961;
wire n_13488;
wire n_15542;
wire n_14718;
wire n_5727;
wire n_4906;
wire n_9098;
wire n_4663;
wire n_5390;
wire n_7114;
wire n_5347;
wire n_11325;
wire n_14612;
wire n_9861;
wire n_6788;
wire n_13638;
wire n_15686;
wire n_14869;
wire n_16190;
wire n_4883;
wire n_11660;
wire n_4162;
wire n_10448;
wire n_14985;
wire n_5115;
wire n_12963;
wire n_14110;
wire n_6393;
wire n_9536;
wire n_8566;
wire n_12282;
wire n_8086;
wire n_14316;
wire n_12620;
wire n_8746;
wire n_11411;
wire n_6249;
wire n_14506;
wire n_4297;
wire n_5833;
wire n_6849;
wire n_13268;
wire n_12431;
wire n_9593;
wire n_15613;
wire n_9017;
wire n_5407;
wire n_14595;
wire n_11281;
wire n_15218;
wire n_11841;
wire n_4608;
wire n_11658;
wire n_5232;
wire n_14765;
wire n_9703;
wire n_14215;
wire n_15437;
wire n_7271;
wire n_12830;
wire n_15991;
wire n_11025;
wire n_6572;
wire n_12213;
wire n_4172;
wire n_4791;
wire n_6739;
wire n_11372;
wire n_4536;
wire n_10450;
wire n_13117;
wire n_13510;
wire n_12397;
wire n_14781;
wire n_14920;
wire n_13665;
wire n_5967;
wire n_5149;
wire n_7569;
wire n_5151;
wire n_7003;
wire n_9565;
wire n_7897;
wire n_4773;
wire n_14954;
wire n_7962;
wire n_8942;
wire n_5345;
wire n_5357;
wire n_4497;
wire n_6666;
wire n_13179;
wire n_13429;
wire n_10320;
wire n_4611;
wire n_14835;
wire n_8113;
wire n_6812;
wire n_4755;
wire n_15284;
wire n_5982;
wire n_4960;
wire n_10308;
wire n_14216;
wire n_8652;
wire n_16032;
wire n_13993;
wire n_4658;
wire n_5135;
wire n_15711;
wire n_16092;
wire n_15701;
wire n_7419;
wire n_15025;
wire n_11545;
wire n_12974;
wire n_14078;
wire n_13717;
wire n_5827;
wire n_9337;
wire n_5494;
wire n_11465;
wire n_4362;
wire n_14314;
wire n_15298;
wire n_15409;
wire n_4306;
wire n_6200;
wire n_11437;
wire n_15602;
wire n_10304;
wire n_16243;
wire n_11436;
wire n_7784;
wire n_13804;
wire n_4422;
wire n_10902;
wire n_8714;
wire n_6123;
wire n_10607;
wire n_6934;
wire n_7500;
wire n_7094;
wire n_11463;
wire n_14152;
wire n_10605;
wire n_11394;
wire n_6082;
wire n_10668;
wire n_8944;
wire n_12487;
wire n_13660;
wire n_13861;
wire n_9232;
wire n_12385;
wire n_15471;
wire n_9320;
wire n_10713;
wire n_4555;
wire n_11191;
wire n_14937;
wire n_9167;
wire n_10464;
wire n_5136;
wire n_15451;
wire n_7864;
wire n_5228;
wire n_14580;
wire n_10596;
wire n_14654;
wire n_10034;
wire n_11068;
wire n_15130;
wire n_7129;
wire n_5758;
wire n_5323;
wire n_13081;
wire n_7790;
wire n_14249;
wire n_4215;
wire n_6952;
wire n_4280;
wire n_7062;
wire n_10875;
wire n_15287;
wire n_16166;
wire n_12735;
wire n_9526;
wire n_8107;
wire n_5471;
wire n_7642;
wire n_5434;
wire n_12475;
wire n_15375;
wire n_14300;
wire n_15461;
wire n_9077;
wire n_5941;
wire n_15993;
wire n_16186;
wire n_7045;
wire n_12646;
wire n_5879;
wire n_11277;
wire n_15340;
wire n_11665;
wire n_15880;
wire n_15195;
wire n_5558;
wire n_11061;
wire n_13777;
wire n_9692;
wire n_13444;
wire n_13800;
wire n_14022;
wire n_5350;
wire n_13267;
wire n_15737;
wire n_13959;
wire n_9141;
wire n_11483;
wire n_5338;
wire n_7238;
wire n_12733;
wire n_7126;
wire n_9745;
wire n_5669;
wire n_9787;
wire n_8674;
wire n_11073;
wire n_14105;
wire n_12944;
wire n_13362;
wire n_14637;
wire n_15120;
wire n_7931;
wire n_10309;
wire n_12061;
wire n_12265;
wire n_13190;
wire n_12380;
wire n_15546;
wire n_8482;
wire n_11462;
wire n_8992;
wire n_14703;
wire n_13032;
wire n_6979;
wire n_11224;
wire n_10024;
wire n_9892;
wire n_6203;
wire n_7405;
wire n_10762;
wire n_7739;
wire n_16227;
wire n_13790;
wire n_10490;
wire n_14357;
wire n_8761;
wire n_7207;
wire n_9078;
wire n_8899;
wire n_11127;
wire n_7934;
wire n_9015;
wire n_7454;
wire n_14283;
wire n_9012;
wire n_4599;
wire n_12794;
wire n_5830;
wire n_6796;
wire n_4812;
wire n_9233;
wire n_12890;
wire n_14492;
wire n_9217;
wire n_13576;
wire n_14644;
wire n_5760;
wire n_6368;
wire n_15457;
wire n_6556;
wire n_4628;
wire n_11632;
wire n_15893;
wire n_10974;
wire n_9435;
wire n_5668;
wire n_5878;
wire n_4873;
wire n_8926;
wire n_5588;
wire n_4657;
wire n_11692;
wire n_11762;
wire n_14662;
wire n_5765;
wire n_11843;
wire n_14341;
wire n_14470;
wire n_9389;
wire n_11344;
wire n_4458;
wire n_11403;
wire n_6596;
wire n_12926;
wire n_15794;
wire n_4121;
wire n_5090;
wire n_14159;
wire n_6870;
wire n_10520;
wire n_7639;
wire n_13666;
wire n_12247;
wire n_12881;
wire n_5613;
wire n_4476;
wire n_10914;
wire n_10129;
wire n_4756;
wire n_4307;
wire n_5104;
wire n_5042;
wire n_4860;
wire n_4359;
wire n_13710;
wire n_11510;
wire n_10084;
wire n_14082;
wire n_7251;
wire n_15966;
wire n_16193;
wire n_10519;
wire n_7776;
wire n_12966;
wire n_6080;
wire n_10318;
wire n_13785;
wire n_7059;
wire n_13287;
wire n_14665;
wire n_8561;
wire n_10877;
wire n_8255;
wire n_7035;
wire n_10468;
wire n_14752;
wire n_5571;
wire n_11854;
wire n_12894;
wire n_8029;
wire n_10906;
wire n_4573;
wire n_6713;
wire n_4118;
wire n_5289;
wire n_14632;
wire n_5513;
wire n_6747;
wire n_12276;
wire n_6281;
wire n_13588;
wire n_15925;
wire n_4803;
wire n_5972;
wire n_10289;
wire n_14496;
wire n_9381;
wire n_13261;
wire n_13634;
wire n_9873;
wire n_15738;
wire n_11925;
wire n_12594;
wire n_10905;
wire n_5916;
wire n_5984;
wire n_7029;
wire n_7317;
wire n_13030;
wire n_14043;
wire n_15855;
wire n_9575;
wire n_5145;
wire n_12529;
wire n_14636;
wire n_11817;
wire n_15887;
wire n_6094;
wire n_15036;
wire n_6444;
wire n_11961;
wire n_12001;
wire n_5132;
wire n_15879;
wire n_5191;
wire n_10298;
wire n_12433;
wire n_6333;
wire n_10940;
wire n_6262;
wire n_16103;
wire n_12765;
wire n_13704;
wire n_5869;
wire n_8130;
wire n_5925;
wire n_9023;
wire n_12097;
wire n_6240;
wire n_10723;
wire n_5359;
wire n_13627;
wire n_6412;
wire n_9412;
wire n_7782;
wire n_5293;
wire n_7220;
wire n_10293;
wire n_11824;
wire n_15427;
wire n_4316;
wire n_15228;
wire n_10361;
wire n_7438;
wire n_11269;
wire n_11270;
wire n_9955;
wire n_10161;
wire n_10432;
wire n_15192;
wire n_7515;
wire n_11532;
wire n_7574;
wire n_12402;
wire n_12728;
wire n_6684;
wire n_4524;
wire n_4843;
wire n_8921;
wire n_13191;
wire n_13766;
wire n_13784;
wire n_10640;
wire n_11546;
wire n_7065;
wire n_10271;
wire n_11314;
wire n_5510;
wire n_6046;
wire n_15359;
wire n_7894;
wire n_9418;
wire n_7868;
wire n_6973;
wire n_9733;
wire n_14963;
wire n_5363;
wire n_7285;
wire n_8286;
wire n_5200;
wire n_9502;
wire n_5659;
wire n_5618;
wire n_15045;
wire n_6325;
wire n_15802;
wire n_13374;
wire n_9765;
wire n_9029;
wire n_11130;
wire n_10163;
wire n_13824;
wire n_6737;
wire n_12262;
wire n_6454;
wire n_4253;
wire n_5356;
wire n_6721;
wire n_8178;
wire n_14175;
wire n_5369;
wire n_11935;
wire n_13452;
wire n_5258;
wire n_12708;
wire n_5255;
wire n_14423;
wire n_15202;
wire n_15919;
wire n_13656;
wire n_10576;
wire n_9623;
wire n_11822;
wire n_10424;
wire n_12805;
wire n_7008;
wire n_11035;
wire n_8925;
wire n_10404;
wire n_14138;
wire n_15318;
wire n_15986;
wire n_8432;
wire n_16040;
wire n_6111;
wire n_16163;
wire n_10130;
wire n_12901;
wire n_7505;
wire n_8047;
wire n_6260;
wire n_7501;
wire n_10214;
wire n_12971;
wire n_15636;
wire n_5080;
wire n_11389;
wire n_6665;
wire n_9783;
wire n_7566;
wire n_7937;
wire n_12658;
wire n_7055;
wire n_14568;
wire n_14562;
wire n_8268;
wire n_11501;
wire n_12372;
wire n_12564;
wire n_8053;
wire n_13141;
wire n_11015;
wire n_5858;
wire n_5817;
wire n_10317;
wire n_6690;
wire n_9840;
wire n_5723;
wire n_10491;
wire n_5295;
wire n_6137;
wire n_10712;
wire n_4679;
wire n_4115;
wire n_6201;
wire n_9909;
wire n_10192;
wire n_7113;
wire n_12204;
wire n_14684;
wire n_4998;
wire n_15055;
wire n_10453;
wire n_11034;
wire n_15852;
wire n_8735;
wire n_11895;
wire n_15291;
wire n_7872;
wire n_12543;
wire n_13895;
wire n_10219;
wire n_15541;
wire n_15722;
wire n_5627;
wire n_12888;
wire n_13854;
wire n_4167;
wire n_14062;
wire n_8845;
wire n_7242;
wire n_5155;
wire n_16235;
wire n_14467;
wire n_6461;
wire n_12013;
wire n_8830;
wire n_11662;
wire n_5016;
wire n_14706;
wire n_7954;
wire n_6212;
wire n_15703;
wire n_6908;
wire n_7819;
wire n_6570;
wire n_14362;
wire n_12741;
wire n_8022;
wire n_9532;
wire n_8415;
wire n_9112;
wire n_6498;
wire n_10062;
wire n_4730;
wire n_7228;
wire n_9561;
wire n_6692;
wire n_8547;
wire n_14553;
wire n_10788;
wire n_11500;
wire n_15092;
wire n_6074;
wire n_10910;
wire n_7561;
wire n_6380;
wire n_10892;
wire n_10216;
wire n_9091;
wire n_14377;
wire n_5996;
wire n_8386;
wire n_8426;
wire n_9326;
wire n_8672;
wire n_11977;
wire n_10049;
wire n_5327;
wire n_7994;
wire n_9180;
wire n_10431;
wire n_11215;
wire n_8540;
wire n_6045;
wire n_9932;
wire n_15274;
wire n_15421;
wire n_4713;
wire n_5137;
wire n_6505;
wire n_13705;
wire n_14535;
wire n_15767;
wire n_16097;
wire n_14776;
wire n_9220;
wire n_9834;
wire n_15814;
wire n_7415;
wire n_13726;
wire n_9474;
wire n_14770;
wire n_14551;
wire n_7793;
wire n_5796;
wire n_7702;
wire n_9542;
wire n_11530;
wire n_7598;
wire n_14406;
wire n_15001;
wire n_6320;
wire n_6489;
wire n_6068;
wire n_15000;
wire n_14449;
wire n_12889;
wire n_14290;
wire n_15765;
wire n_14919;
wire n_8192;
wire n_5791;
wire n_8791;
wire n_9458;
wire n_10608;
wire n_15535;
wire n_4204;
wire n_9642;
wire n_14768;
wire n_5098;
wire n_6877;
wire n_6772;
wire n_6823;
wire n_9020;
wire n_9910;
wire n_6806;
wire n_7426;
wire n_11014;
wire n_15355;
wire n_5906;
wire n_8350;
wire n_11439;
wire n_14744;
wire n_16036;
wire n_12526;
wire n_9100;
wire n_11119;
wire n_11752;
wire n_14081;
wire n_14410;
wire n_4743;
wire n_8816;
wire n_7957;
wire n_14549;
wire n_8712;
wire n_8048;
wire n_6831;
wire n_15058;
wire n_16172;
wire n_10395;
wire n_4924;
wire n_12255;
wire n_9781;
wire n_13881;
wire n_8663;
wire n_15861;
wire n_7217;
wire n_4859;
wire n_9940;
wire n_12068;
wire n_10802;
wire n_6284;
wire n_7058;
wire n_6157;
wire n_4654;
wire n_5423;
wire n_7497;
wire n_8503;
wire n_6785;
wire n_8254;
wire n_6374;
wire n_8959;
wire n_13280;
wire n_9117;
wire n_6930;
wire n_12784;
wire n_9198;
wire n_6017;
wire n_4733;
wire n_11729;
wire n_8506;
wire n_4272;
wire n_11289;
wire n_11699;
wire n_7735;
wire n_8265;
wire n_8465;
wire n_8049;
wire n_12277;
wire n_4269;
wire n_4695;
wire n_6838;
wire n_11902;
wire n_12212;
wire n_12126;
wire n_5736;
wire n_6937;
wire n_12686;
wire n_15716;
wire n_6443;
wire n_13328;
wire n_6105;
wire n_10080;
wire n_16236;
wire n_7558;
wire n_13554;
wire n_12344;
wire n_12250;
wire n_8937;
wire n_12961;
wire n_14142;
wire n_5069;
wire n_7442;
wire n_10574;
wire n_8272;
wire n_5700;
wire n_6543;
wire n_9249;
wire n_15527;
wire n_11628;
wire n_10594;
wire n_11784;
wire n_12193;
wire n_9398;
wire n_5099;
wire n_16144;
wire n_15748;
wire n_11622;
wire n_14033;
wire n_4704;
wire n_14269;
wire n_4551;
wire n_11763;
wire n_13393;
wire n_5052;
wire n_6091;
wire n_11606;
wire n_12749;
wire n_4957;
wire n_6674;
wire n_15821;
wire n_10155;
wire n_14585;
wire n_6034;
wire n_15683;
wire n_15964;
wire n_15032;
wire n_7499;
wire n_9751;
wire n_14866;
wire n_13134;
wire n_5579;
wire n_8381;
wire n_13399;
wire n_7085;
wire n_13413;
wire n_12079;
wire n_4781;
wire n_9579;
wire n_11006;
wire n_10879;
wire n_6652;
wire n_7098;
wire n_5004;
wire n_6762;
wire n_15090;
wire n_7341;
wire n_7895;
wire n_13602;
wire n_4424;
wire n_11321;
wire n_13250;
wire n_15980;
wire n_8366;
wire n_10792;
wire n_16137;
wire n_8101;
wire n_7611;
wire n_9925;
wire n_10655;
wire n_14065;
wire n_7391;
wire n_14713;
wire n_10890;
wire n_12187;
wire n_12093;
wire n_5837;
wire n_14539;
wire n_15963;
wire n_4436;
wire n_6895;
wire n_7646;
wire n_4450;
wire n_8384;
wire n_13035;
wire n_9889;
wire n_5642;
wire n_14299;
wire n_12705;
wire n_7224;
wire n_5880;
wire n_8728;
wire n_6169;
wire n_11133;
wire n_4746;
wire n_12241;
wire n_14114;
wire n_12211;
wire n_15082;
wire n_7524;
wire n_5713;
wire n_6005;
wire n_15100;
wire n_10212;
wire n_8023;
wire n_13770;
wire n_13975;
wire n_8052;
wire n_11001;
wire n_7627;
wire n_9998;
wire n_11143;
wire n_10654;
wire n_9729;
wire n_5118;
wire n_5105;
wire n_14112;
wire n_15367;
wire n_13833;
wire n_13886;
wire n_15402;
wire n_15934;
wire n_4459;
wire n_11757;
wire n_13169;
wire n_8614;
wire n_16124;
wire n_5793;
wire n_5591;
wire n_13237;
wire n_7856;
wire n_16055;
wire n_9081;
wire n_7496;
wire n_12446;
wire n_12640;
wire n_15302;
wire n_12699;
wire n_9784;
wire n_13354;
wire n_13696;
wire n_15250;
wire n_5623;
wire n_12856;
wire n_14834;
wire n_16106;
wire n_10005;
wire n_10544;
wire n_10217;
wire n_12231;
wire n_5681;
wire n_4853;
wire n_11421;
wire n_11780;
wire n_12745;
wire n_14798;
wire n_9856;
wire n_15474;
wire n_15768;
wire n_9101;
wire n_7399;
wire n_12841;
wire n_15955;
wire n_6213;
wire n_8656;
wire n_10393;
wire n_6118;
wire n_5256;
wire n_11793;
wire n_12527;
wire n_7605;
wire n_14386;
wire n_11400;
wire n_5220;
wire n_12814;
wire n_5732;
wire n_8897;
wire n_9696;
wire n_12545;
wire n_5178;
wire n_11621;
wire n_15436;
wire n_6814;
wire n_4520;
wire n_13913;
wire n_7342;
wire n_12354;
wire n_8014;
wire n_9825;
wire n_13783;
wire n_15493;
wire n_16078;
wire n_5507;
wire n_10093;
wire n_8564;
wire n_11969;
wire n_14926;
wire n_7472;
wire n_7214;
wire n_12685;
wire n_5077;
wire n_10850;
wire n_12886;
wire n_13297;
wire n_8371;
wire n_10945;
wire n_5872;
wire n_13564;
wire n_14601;
wire n_15984;
wire n_11791;
wire n_7408;
wire n_8231;
wire n_9250;
wire n_6115;
wire n_4502;
wire n_9572;
wire n_10541;
wire n_6858;
wire n_12196;
wire n_10375;
wire n_11948;
wire n_11910;
wire n_8558;
wire n_5735;
wire n_4851;
wire n_9483;
wire n_10275;
wire n_9816;
wire n_12119;
wire n_9253;
wire n_15080;
wire n_8164;
wire n_7254;
wire n_6944;
wire n_7384;
wire n_9136;
wire n_14280;
wire n_7837;
wire n_8357;
wire n_10726;
wire n_9426;
wire n_8870;
wire n_9831;
wire n_4571;
wire n_13434;
wire n_14017;
wire n_14395;
wire n_8143;
wire n_11064;
wire n_14187;
wire n_6430;
wire n_14027;
wire n_6193;
wire n_10614;
wire n_8422;
wire n_6462;
wire n_5314;
wire n_12094;
wire n_15916;
wire n_12096;
wire n_9896;
wire n_9650;
wire n_13657;
wire n_12730;
wire n_10002;
wire n_5049;
wire n_6757;
wire n_6822;
wire n_14639;
wire n_4205;
wire n_5953;
wire n_7599;
wire n_16218;
wire n_5277;
wire n_4723;
wire n_5176;
wire n_11974;
wire n_12202;
wire n_6779;
wire n_6518;
wire n_9767;
wire n_15258;
wire n_16085;
wire n_6797;
wire n_11367;
wire n_14094;
wire n_4454;
wire n_7938;
wire n_8253;
wire n_4229;
wire n_14730;
wire n_5952;
wire n_15207;
wire n_4739;
wire n_12534;
wire n_13692;
wire n_5820;
wire n_5483;
wire n_12120;
wire n_9028;
wire n_9055;
wire n_5718;
wire n_10251;
wire n_14722;
wire n_11562;
wire n_11866;
wire n_13585;
wire n_6916;
wire n_5150;
wire n_11383;
wire n_12854;
wire n_8563;
wire n_15988;
wire n_9949;
wire n_4838;
wire n_16168;
wire n_5075;
wire n_11655;
wire n_12553;
wire n_7812;
wire n_12816;
wire n_14906;
wire n_4879;
wire n_5051;
wire n_14486;
wire n_11552;
wire n_14807;
wire n_9684;
wire n_15418;
wire n_6152;
wire n_10010;
wire n_9724;
wire n_13430;
wire n_4221;
wire n_8243;
wire n_10226;
wire n_11117;
wire n_8236;
wire n_14964;
wire n_11046;
wire n_8292;
wire n_14640;
wire n_14901;
wire n_11547;
wire n_12676;
wire n_13327;
wire n_4181;
wire n_14412;
wire n_14391;
wire n_5777;
wire n_7949;
wire n_8611;
wire n_7046;
wire n_12720;
wire n_4225;
wire n_10475;
wire n_13365;
wire n_10020;
wire n_9826;
wire n_5142;
wire n_14195;
wire n_10467;
wire n_4153;
wire n_5156;
wire n_13118;
wire n_5926;
wire n_8011;
wire n_15271;
wire n_9839;
wire n_15816;
wire n_14431;
wire n_4300;
wire n_9399;
wire n_4783;
wire n_12535;
wire n_14254;
wire n_13279;
wire n_15497;
wire n_12283;
wire n_12506;
wire n_14044;
wire n_6589;
wire n_7579;
wire n_4530;
wire n_15393;
wire n_4267;
wire n_8139;
wire n_12046;
wire n_8123;
wire n_15104;
wire n_7173;
wire n_10720;
wire n_7917;
wire n_5951;
wire n_7092;
wire n_10907;
wire n_6197;
wire n_6971;
wire n_9938;
wire n_8424;
wire n_9776;
wire n_8859;
wire n_13844;
wire n_14462;
wire n_11256;
wire n_7460;
wire n_9658;
wire n_15773;
wire n_11914;
wire n_9605;
wire n_12124;
wire n_11934;
wire n_14731;
wire n_15638;
wire n_10868;
wire n_11047;
wire n_9013;
wire n_14004;
wire n_8730;
wire n_9417;
wire n_14841;
wire n_13945;
wire n_8156;
wire n_9290;
wire n_9212;
wire n_13431;
wire n_15446;
wire n_13342;
wire n_9721;
wire n_14913;
wire n_14789;
wire n_12189;
wire n_10615;
wire n_7698;
wire n_12884;
wire n_13187;
wire n_7886;
wire n_6154;
wire n_7344;
wire n_14504;
wire n_6020;
wire n_15884;
wire n_13082;
wire n_9586;
wire n_7904;
wire n_12310;
wire n_11004;
wire n_4182;
wire n_10751;
wire n_12683;
wire n_13821;
wire n_11287;
wire n_5701;
wire n_4825;
wire n_10706;
wire n_4440;
wire n_10774;
wire n_11208;
wire n_4549;
wire n_12108;
wire n_12502;
wire n_15267;
wire n_9104;
wire n_7079;
wire n_10225;
wire n_11963;
wire n_10570;
wire n_9293;
wire n_15517;
wire n_11860;
wire n_13298;
wire n_5120;
wire n_8645;
wire n_10744;
wire n_11625;
wire n_5470;
wire n_16174;
wire n_4565;
wire n_7675;
wire n_10416;
wire n_4303;
wire n_4574;
wire n_14933;
wire n_7774;
wire n_5797;
wire n_7922;
wire n_8189;
wire n_8618;
wire n_6696;
wire n_11181;
wire n_11787;
wire n_14024;
wire n_4839;
wire n_5222;
wire n_13810;
wire n_8285;
wire n_5743;
wire n_10396;
wire n_9919;
wire n_8826;
wire n_6210;
wire n_10123;
wire n_5772;
wire n_12899;
wire n_14252;
wire n_8715;
wire n_12761;
wire n_14522;
wire n_8782;
wire n_6964;
wire n_14399;
wire n_10083;
wire n_5801;
wire n_6117;
wire n_14331;
wire n_4231;
wire n_15561;
wire n_8117;
wire n_12918;
wire n_11825;
wire n_6202;
wire n_7279;
wire n_7670;
wire n_11364;
wire n_4923;
wire n_12713;
wire n_15585;
wire n_14126;
wire n_12522;
wire n_12822;
wire n_9445;
wire n_14148;
wire n_4097;
wire n_14031;
wire n_6681;
wire n_13539;
wire n_5971;
wire n_11420;
wire n_12223;
wire n_13532;
wire n_15892;
wire n_11470;
wire n_4461;
wire n_13089;
wire n_5392;
wire n_8497;
wire n_12082;
wire n_9930;
wire n_6661;
wire n_8018;
wire n_6640;
wire n_12151;
wire n_15755;
wire n_13335;
wire n_7940;
wire n_14493;
wire n_11230;
wire n_12757;
wire n_7371;
wire n_10731;
wire n_6962;
wire n_4101;
wire n_13411;
wire n_11074;
wire n_10347;
wire n_11063;
wire n_15468;
wire n_6455;
wire n_7721;
wire n_9727;
wire n_4273;
wire n_15034;
wire n_7606;
wire n_5443;
wire n_12025;
wire n_5600;
wire n_4939;
wire n_15895;
wire n_5169;
wire n_6963;
wire n_10926;
wire n_6644;
wire n_13848;
wire n_13879;
wire n_14534;
wire n_4389;
wire n_6896;
wire n_14475;
wire n_12183;
wire n_14633;
wire n_4448;
wire n_11669;
wire n_10734;
wire n_6832;
wire n_8798;
wire n_7836;
wire n_16128;
wire n_16224;
wire n_12143;
wire n_6160;
wire n_14473;
wire n_7564;
wire n_11493;
wire n_12158;
wire n_7884;
wire n_8673;
wire n_10281;
wire n_6718;
wire n_9685;
wire n_11486;
wire n_8502;
wire n_6542;
wire n_10126;
wire n_10759;
wire n_13293;
wire n_11786;
wire n_10650;
wire n_14083;
wire n_11777;
wire n_6031;
wire n_5568;
wire n_5502;
wire n_9421;
wire n_8577;
wire n_11722;
wire n_14487;
wire n_7653;
wire n_15835;
wire n_10445;
wire n_10092;
wire n_15241;
wire n_5656;
wire n_8531;
wire n_8635;
wire n_6763;
wire n_4831;
wire n_5974;
wire n_9567;
wire n_6280;
wire n_9298;
wire n_11941;
wire n_10116;
wire n_6438;
wire n_13614;
wire n_10048;
wire n_9059;
wire n_12937;
wire n_15372;
wire n_8485;
wire n_13285;
wire n_6316;
wire n_7383;
wire n_4319;
wire n_5474;
wire n_13596;
wire n_8872;
wire n_8752;
wire n_13609;
wire n_9396;
wire n_4596;
wire n_6758;
wire n_5413;
wire n_12459;
wire n_13715;
wire n_13398;
wire n_7976;
wire n_9234;
wire n_9425;
wire n_12648;
wire n_10364;
wire n_5412;
wire n_9620;
wire n_6069;
wire n_10963;
wire n_5752;
wire n_10191;
wire n_6874;
wire n_13330;
wire n_4726;
wire n_16127;
wire n_13235;
wire n_4751;
wire n_15319;
wire n_4222;
wire n_8341;
wire n_13412;
wire n_13995;
wire n_14867;
wire n_12638;
wire n_8521;
wire n_6030;
wire n_11209;
wire n_8199;
wire n_12976;
wire n_13091;
wire n_13306;
wire n_13561;
wire n_6077;
wire n_8005;
wire n_11718;
wire n_4119;
wire n_7743;
wire n_4298;
wire n_16122;
wire n_5201;
wire n_6299;
wire n_9280;
wire n_9517;
wire n_4474;
wire n_6386;
wire n_9639;
wire n_9192;
wire n_14089;
wire n_12762;
wire n_9102;
wire n_5217;
wire n_10003;
wire n_10025;
wire n_8016;
wire n_10156;
wire n_8669;
wire n_5957;
wire n_15603;
wire n_12066;
wire n_11234;
wire n_16101;
wire n_12021;
wire n_14822;
wire n_8283;
wire n_13016;
wire n_13048;
wire n_10502;
wire n_7655;
wire n_5490;
wire n_16102;
wire n_5029;
wire n_8291;
wire n_4214;
wire n_8176;
wire n_10674;
wire n_15337;
wire n_5158;
wire n_4884;
wire n_14942;
wire n_6708;
wire n_7737;
wire n_10179;
wire n_14076;
wire n_7433;
wire n_11000;
wire n_12447;
wire n_13939;
wire n_11702;
wire n_4366;
wire n_10466;
wire n_12667;
wire n_15782;
wire n_12221;
wire n_7347;
wire n_8145;
wire n_9487;
wire n_10268;
wire n_4580;
wire n_13560;
wire n_6792;
wire n_14389;
wire n_12906;
wire n_15392;
wire n_7633;
wire n_12851;
wire n_6177;
wire n_5912;
wire n_11431;
wire n_10679;
wire n_12691;
wire n_7798;
wire n_10492;
wire n_11177;
wire n_12980;
wire n_4129;
wire n_4871;
wire n_12416;
wire n_13436;
wire n_4999;
wire n_13023;
wire n_13985;
wire n_11454;
wire n_6033;
wire n_9221;
wire n_12989;
wire n_11418;
wire n_5557;
wire n_7397;
wire n_12739;
wire n_7389;
wire n_13074;
wire n_12791;
wire n_5472;
wire n_7602;
wire n_13920;
wire n_13795;
wire n_14483;
wire n_4112;
wire n_8069;
wire n_6002;
wire n_14696;
wire n_14571;
wire n_14753;
wire n_4337;
wire n_5711;
wire n_4138;
wire n_7554;
wire n_14903;
wire n_5396;
wire n_7693;
wire n_14052;
wire n_5335;
wire n_8888;
wire n_12650;
wire n_12319;
wire n_15661;
wire n_15391;
wire n_6557;
wire n_7300;
wire n_15515;
wire n_9566;
wire n_12692;
wire n_12403;
wire n_14908;
wire n_15522;
wire n_9578;
wire n_8483;
wire n_15534;
wire n_14820;
wire n_8797;
wire n_5960;
wire n_8605;
wire n_8041;
wire n_4236;
wire n_9868;
wire n_13451;
wire n_14778;
wire n_5002;
wire n_15225;
wire n_11750;
wire n_14124;
wire n_14442;
wire n_15386;
wire n_11572;
wire n_7532;
wire n_11049;
wire n_11038;
wire n_9292;
wire n_10460;
wire n_13363;
wire n_5143;
wire n_7724;
wire n_4238;
wire n_12669;
wire n_15492;
wire n_15508;
wire n_11491;
wire n_14838;
wire n_6142;
wire n_6917;
wire n_7510;
wire n_11109;
wire n_5859;
wire n_10968;
wire n_8760;
wire n_4734;
wire n_8928;
wire n_10004;
wire n_11894;
wire n_10729;
wire n_13689;
wire n_8374;
wire n_14276;
wire n_8917;
wire n_6163;
wire n_4635;
wire n_10811;
wire n_14540;
wire n_7118;
wire n_8006;
wire n_11806;
wire n_9884;
wire n_11504;
wire n_6285;
wire n_6778;
wire n_7946;
wire n_8723;
wire n_9857;
wire n_12127;
wire n_11637;
wire n_14622;
wire n_6025;
wire n_13769;
wire n_8957;
wire n_12058;
wire n_7257;
wire n_4242;
wire n_11799;
wire n_10944;
wire n_11788;
wire n_13537;
wire n_15809;
wire n_6862;
wire n_6319;
wire n_7067;
wire n_4984;
wire n_13143;
wire n_13808;
wire n_10140;
wire n_14226;
wire n_12868;
wire n_12642;
wire n_10013;
wire n_14106;
wire n_12600;
wire n_7933;
wire n_5283;
wire n_8409;
wire n_9815;
wire n_9110;
wire n_7669;
wire n_5268;
wire n_10110;
wire n_13909;
wire n_6318;
wire n_10133;
wire n_14531;
wire n_14720;
wire n_8215;
wire n_11453;
wire n_16234;
wire n_11184;
wire n_8220;
wire n_9471;
wire n_9048;
wire n_4561;
wire n_7927;
wire n_11356;
wire n_6089;
wire n_8629;
wire n_13045;
wire n_5122;
wire n_7910;
wire n_12005;
wire n_11955;
wire n_13426;
wire n_14596;
wire n_6315;
wire n_10592;
wire n_14887;
wire n_7970;
wire n_14172;
wire n_15518;
wire n_4955;
wire n_15985;
wire n_10476;
wire n_8407;
wire n_5556;
wire n_5462;
wire n_16100;
wire n_4501;
wire n_15153;
wire n_14147;
wire n_12953;
wire n_14593;
wire n_13507;
wire n_15159;
wire n_11488;
wire n_13040;
wire n_15432;
wire n_12369;
wire n_9394;
wire n_8991;
wire n_12300;
wire n_5840;
wire n_13015;
wire n_14934;
wire n_6343;
wire n_10186;
wire n_11938;
wire n_15505;
wire n_14988;
wire n_11946;
wire n_9191;
wire n_11918;
wire n_9004;
wire n_12832;
wire n_13839;
wire n_6049;
wire n_6919;
wire n_7423;
wire n_7865;
wire n_6052;
wire n_11412;
wire n_13522;
wire n_10700;
wire n_5330;
wire n_4197;
wire n_15690;
wire n_4829;
wire n_15746;
wire n_7069;
wire n_12290;
wire n_13208;
wire n_6886;
wire n_13761;
wire n_14219;
wire n_12169;
wire n_8783;
wire n_6912;
wire n_8326;
wire n_10496;
wire n_11249;
wire n_13538;
wire n_10521;
wire n_12838;
wire n_5914;
wire n_14523;
wire n_11464;
wire n_12325;
wire n_15465;
wire n_8504;
wire n_10695;
wire n_14763;
wire n_8445;
wire n_11950;
wire n_13847;
wire n_11648;
wire n_8250;
wire n_10994;
wire n_11576;
wire n_4715;
wire n_5039;
wire n_9118;
wire n_13950;
wire n_6061;
wire n_4369;
wire n_14025;
wire n_15006;
wire n_12969;
wire n_13214;
wire n_5378;
wire n_10758;
wire n_13559;
wire n_8408;
wire n_4543;
wire n_10120;
wire n_11410;
wire n_15499;
wire n_4941;
wire n_11251;
wire n_7252;
wire n_5542;
wire n_15450;
wire n_4394;
wire n_9051;
wire n_16159;
wire n_7133;
wire n_6883;
wire n_10345;
wire n_13065;
wire n_5519;
wire n_12809;
wire n_9908;
wire n_12748;
wire n_13639;
wire n_6009;
wire n_7061;
wire n_8155;
wire n_5278;
wire n_8818;
wire n_11641;
wire n_11633;
wire n_12264;
wire n_7518;
wire n_9123;
wire n_12352;
wire n_5586;
wire n_13221;
wire n_15297;
wire n_10232;
wire n_6378;
wire n_8660;
wire n_5187;
wire n_4944;
wire n_13619;
wire n_15581;
wire n_12054;
wire n_5675;
wire n_14055;
wire n_4135;
wire n_8275;
wire n_9327;
wire n_6601;
wire n_5771;
wire n_7216;
wire n_6407;
wire n_15488;
wire n_11555;
wire n_9687;
wire n_14552;
wire n_8297;
wire n_9828;
wire n_6749;
wire n_13921;
wire n_11984;
wire n_14355;
wire n_6839;
wire n_10533;
wire n_13053;
wire n_14448;
wire n_9519;
wire n_10611;
wire n_7711;
wire n_15431;
wire n_13635;
wire n_12368;
wire n_10089;
wire n_15206;
wire n_12137;
wire n_15538;
wire n_4263;
wire n_11651;
wire n_14038;
wire n_7705;
wire n_10455;
wire n_6051;
wire n_4716;
wire n_8590;
wire n_15259;
wire n_12538;
wire n_4942;
wire n_6217;
wire n_13671;
wire n_6680;
wire n_5844;
wire n_12016;
wire n_15610;
wire n_7972;
wire n_15075;
wire n_6532;
wire n_13517;
wire n_15837;
wire n_6155;
wire n_4745;
wire n_6446;
wire n_8072;
wire n_12644;
wire n_6738;
wire n_6250;
wire n_7614;
wire n_7458;
wire n_7854;
wire n_12017;
wire n_7707;
wire n_10632;
wire n_13428;
wire n_11672;
wire n_16016;
wire n_11696;
wire n_8050;
wire n_6736;
wire n_5344;
wire n_15398;
wire n_6526;
wire n_8142;
wire n_10820;
wire n_14914;
wire n_10601;
wire n_13455;
wire n_6339;
wire n_4629;
wire n_14594;
wire n_12197;
wire n_5225;
wire n_8151;
wire n_6350;
wire n_7013;
wire n_12892;
wire n_5662;
wire n_4857;
wire n_16061;
wire n_14213;
wire n_9802;
wire n_9315;
wire n_9296;
wire n_8599;
wire n_10447;
wire n_12373;
wire n_12660;
wire n_14393;
wire n_4226;
wire n_4741;
wire n_10022;
wire n_14526;
wire n_15278;
wire n_4752;
wire n_5265;
wire n_14184;
wire n_11567;
wire n_10305;
wire n_14769;
wire n_12855;
wire n_15777;
wire n_14795;
wire n_4376;
wire n_10031;
wire n_12877;
wire n_5705;
wire n_4753;
wire n_12350;
wire n_14691;
wire n_15730;
wire n_14576;
wire n_15944;
wire n_13137;
wire n_10798;
wire n_12388;
wire n_4552;
wire n_7656;
wire n_11202;
wire n_10760;
wire n_6845;
wire n_9405;
wire n_14647;
wire n_12891;
wire n_9302;
wire n_7105;
wire n_12836;
wire n_5196;
wire n_13892;
wire n_5181;
wire n_13636;
wire n_16057;
wire n_11779;
wire n_11888;
wire n_10166;
wire n_14317;
wire n_15024;
wire n_6829;
wire n_11684;
wire n_11879;
wire n_5574;
wire n_15843;
wire n_11054;
wire n_5126;
wire n_6508;
wire n_9842;
wire n_9977;
wire n_9887;
wire n_15820;
wire n_14893;
wire n_15370;
wire n_5553;
wire n_4176;
wire n_7570;
wire n_8246;
wire n_11116;
wire n_15220;
wire n_9524;
wire n_11129;
wire n_7771;
wire n_4385;
wire n_13742;
wire n_7052;
wire n_5009;
wire n_7262;
wire n_5368;
wire n_9322;
wire n_11937;
wire n_10098;
wire n_15079;
wire n_10510;
wire n_13934;
wire n_13905;
wire n_10848;
wire n_10042;
wire n_8057;
wire n_9122;
wire n_8349;
wire n_5626;
wire n_9333;
wire n_13240;
wire n_16131;
wire n_15947;
wire n_8743;
wire n_6603;
wire n_6114;
wire n_14073;
wire n_16136;
wire n_9590;
wire n_13515;
wire n_6576;
wire n_15915;
wire n_7943;
wire n_4333;
wire n_7364;
wire n_8473;
wire n_10993;
wire n_13838;
wire n_10342;
wire n_7208;
wire n_12286;
wire n_6245;
wire n_15353;
wire n_12992;
wire n_14132;
wire n_10439;
wire n_11923;
wire n_12844;
wire n_14284;
wire n_5499;
wire n_6703;
wire n_4788;
wire n_4375;
wire n_4717;
wire n_4986;
wire n_5604;
wire n_13868;
wire n_9676;
wire n_10444;
wire n_15103;
wire n_7714;
wire n_9902;
wire n_10054;
wire n_12759;
wire n_8535;
wire n_10728;
wire n_4815;
wire n_9621;
wire n_13175;
wire n_7202;
wire n_9140;
wire n_4246;
wire n_9604;
wire n_7011;
wire n_4609;
wire n_13759;
wire n_7621;
wire n_8068;
wire n_5291;
wire n_10565;
wire n_10540;
wire n_14444;
wire n_12935;
wire n_16230;
wire n_9821;
wire n_11943;
wire n_14158;
wire n_10748;
wire n_5876;
wire n_10178;
wire n_11995;
wire n_15294;
wire n_11058;
wire n_6970;
wire n_11842;
wire n_12076;
wire n_12790;
wire n_12979;
wire n_5114;
wire n_6409;
wire n_6704;
wire n_16191;
wire n_6876;
wire n_12659;
wire n_7778;
wire n_4357;
wire n_9343;
wire n_15563;
wire n_7028;
wire n_12532;
wire n_4462;
wire n_4472;
wire n_7313;
wire n_7320;
wire n_6255;
wire n_14437;
wire n_7343;
wire n_5288;
wire n_5540;
wire n_5699;
wire n_11473;
wire n_7525;
wire n_13735;
wire n_7875;
wire n_16065;
wire n_5810;
wire n_11568;
wire n_14384;
wire n_16113;
wire n_13258;
wire n_15784;
wire n_15891;
wire n_4151;
wire n_4148;
wire n_13617;
wire n_12702;
wire n_16077;
wire n_6938;
wire n_12050;
wire n_4373;
wire n_12138;
wire n_5762;
wire n_13713;
wire n_4934;
wire n_5218;
wire n_8785;
wire n_9952;
wire n_12473;
wire n_13013;
wire n_14577;
wire n_15175;
wire n_10686;
wire n_15975;
wire n_8327;
wire n_12606;
wire n_9219;
wire n_7337;
wire n_6989;
wire n_8512;
wire n_13625;
wire n_4630;
wire n_5408;
wire n_10971;
wire n_4643;
wire n_6427;
wire n_4331;
wire n_15810;
wire n_13051;
wire n_13054;
wire n_4475;
wire n_7753;
wire n_10076;
wire n_4846;
wire n_11924;
wire n_4344;
wire n_15410;
wire n_12374;
wire n_8168;
wire n_14837;
wire n_16099;
wire n_14266;
wire n_14064;
wire n_8392;
wire n_7038;
wire n_12967;
wire n_15440;
wire n_14745;
wire n_4683;
wire n_15383;
wire n_5366;
wire n_10132;
wire n_10282;
wire n_13649;
wire n_9872;
wire n_16080;
wire n_15354;
wire n_12956;
wire n_6360;
wire n_11203;
wire n_13026;
wire n_9553;
wire n_10900;
wire n_6146;
wire n_10616;
wire n_9447;
wire n_6270;
wire n_11585;
wire n_9150;
wire n_5477;
wire n_9592;
wire n_5451;
wire n_9984;
wire n_12695;
wire n_14111;
wire n_11416;
wire n_4696;
wire n_11526;
wire n_11742;
wire n_13476;
wire n_13855;
wire n_12179;
wire n_8419;
wire n_11809;
wire n_15187;
wire n_5086;
wire n_9814;
wire n_10858;
wire n_12038;
wire n_5901;
wire n_6353;
wire n_14359;
wire n_10769;
wire n_15513;
wire n_9446;
wire n_4905;
wire n_14689;
wire n_15088;
wire n_10211;
wire n_10023;
wire n_15335;
wire n_11877;
wire n_4876;
wire n_15384;
wire n_6345;
wire n_12105;
wire n_9461;
wire n_10772;
wire n_9793;
wire n_6691;
wire n_8997;
wire n_14324;
wire n_4278;
wire n_15939;
wire n_13184;
wire n_15641;
wire n_4623;
wire n_4910;
wire n_12360;
wire n_15330;
wire n_15361;
wire n_12297;
wire n_4410;
wire n_12952;
wire n_9874;
wire n_15838;
wire n_7392;
wire n_5053;
wire n_7912;
wire n_8245;
wire n_14567;
wire n_6239;
wire n_4553;
wire n_6803;
wire n_10446;
wire n_11735;
wire n_14981;
wire n_7919;
wire n_15050;
wire n_6340;
wire n_7583;
wire n_14281;
wire n_4809;
wire n_14876;
wire n_8109;
wire n_5226;
wire n_7657;
wire n_14129;
wire n_15936;
wire n_7995;
wire n_11405;
wire n_15382;
wire n_5867;
wire n_6048;
wire n_8985;
wire n_13318;
wire n_14733;
wire n_5079;
wire n_5590;
wire n_10331;
wire n_12103;
wire n_6773;
wire n_9403;
wire n_5632;
wire n_14515;
wire n_8390;
wire n_15252;
wire n_11480;
wire n_11874;
wire n_4841;
wire n_12115;
wire n_6336;
wire n_8463;
wire n_14120;
wire n_7041;
wire n_15324;
wire n_7802;
wire n_15489;
wire n_4911;
wire n_4842;
wire n_14243;
wire n_4340;
wire n_7370;
wire n_13366;
wire n_10181;
wire n_10074;
wire n_9731;
wire n_5660;
wire n_11104;
wire n_13677;
wire n_4645;
wire n_7557;
wire n_11862;
wire n_11952;
wire n_14529;
wire n_6174;
wire n_4920;
wire n_12828;
wire n_4972;
wire n_13322;
wire n_6023;
wire n_6776;
wire n_14894;
wire n_13078;
wire n_5426;
wire n_15496;
wire n_9947;
wire n_15758;
wire n_6463;
wire n_15423;
wire n_13387;
wire n_14370;
wire n_7896;
wire n_13226;
wire n_9699;
wire n_6372;
wire n_10962;
wire n_11037;
wire n_9305;
wire n_10481;
wire n_14624;
wire n_7176;
wire n_12003;
wire n_14194;
wire n_14868;
wire n_15770;
wire n_10220;
wire n_13917;
wire n_10381;
wire n_15237;
wire n_8517;
wire n_12332;
wire n_5625;
wire n_5778;
wire n_6396;
wire n_10642;
wire n_9218;
wire n_13317;
wire n_11556;
wire n_6669;
wire n_9096;
wire n_10634;
wire n_13480;
wire n_10170;
wire n_10142;
wire n_10569;
wire n_12326;
wire n_15449;
wire n_14489;
wire n_15830;
wire n_5531;
wire n_15321;
wire n_9534;
wire n_7826;
wire n_5429;
wire n_11044;
wire n_5818;
wire n_5646;
wire n_6940;
wire n_4557;
wire n_5248;
wire n_11042;
wire n_12141;
wire n_4451;
wire n_6394;
wire n_9164;
wire n_9546;
wire n_12622;
wire n_11226;
wire n_5448;
wire n_7590;
wire n_5432;
wire n_14977;
wire n_16126;
wire n_13732;
wire n_15804;
wire n_9358;
wire n_11985;
wire n_5160;
wire n_11328;
wire n_13545;
wire n_8208;
wire n_15117;
wire n_6995;
wire n_7185;
wire n_10127;
wire n_14214;
wire n_11525;
wire n_9730;
wire n_6254;
wire n_6161;
wire n_13246;
wire n_9066;
wire n_16209;
wire n_10800;
wire n_11020;
wire n_9185;
wire n_15233;
wire n_9318;
wire n_10374;
wire n_7987;
wire n_8134;
wire n_14367;
wire n_4324;
wire n_4821;
wire n_10328;
wire n_8631;
wire n_14542;
wire n_5445;
wire n_8694;
wire n_11892;
wire n_8965;
wire n_8647;
wire n_13288;
wire n_11013;
wire n_12343;
wire n_7332;
wire n_6660;
wire n_15396;
wire n_4771;
wire n_5719;
wire n_15422;
wire n_7225;
wire n_10529;
wire n_12396;
wire n_13823;
wire n_6128;
wire n_7037;
wire n_15350;
wire n_11820;
wire n_14900;
wire n_11587;
wire n_14863;
wire n_4814;
wire n_12081;
wire n_13157;
wire n_10314;
wire n_14966;
wire n_15982;
wire n_15646;
wire n_5749;
wire n_11697;
wire n_12296;
wire n_8427;
wire n_9339;
wire n_5332;
wire n_13038;
wire n_9596;
wire n_5108;
wire n_7409;
wire n_4692;
wire n_10006;
wire n_10667;
wire n_7258;
wire n_7432;
wire n_9156;
wire n_11441;
wire n_11242;
wire n_11916;
wire n_15209;
wire n_14591;
wire n_15818;
wire n_11435;
wire n_12804;
wire n_13999;
wire n_11471;
wire n_6334;
wire n_10346;
wire n_13236;
wire n_8984;
wire n_6848;
wire n_14502;
wire n_10539;
wire n_8345;
wire n_15590;
wire n_10414;
wire n_6321;
wire n_7765;
wire n_4708;
wire n_9708;
wire n_9268;
wire n_8764;
wire n_6794;
wire n_10340;
wire n_4826;
wire n_13310;
wire n_10245;
wire n_14479;
wire n_11644;
wire n_7761;
wire n_7197;
wire n_12466;
wire n_12701;
wire n_5489;
wire n_15560;
wire n_12106;
wire n_6400;
wire n_12560;
wire n_4589;
wire n_9097;
wire n_5057;
wire n_10280;
wire n_15909;
wire n_12895;
wire n_16066;
wire n_11432;
wire n_4578;
wire n_12342;
wire n_6705;
wire n_7775;
wire n_9636;
wire n_10256;
wire n_14559;
wire n_14676;
wire n_7619;
wire n_12125;
wire n_5436;
wire n_5907;
wire n_11120;
wire n_5072;
wire n_11391;
wire n_11164;
wire n_6044;
wire n_11527;
wire n_5286;
wire n_8083;
wire n_8853;
wire n_11371;
wire n_6495;
wire n_5013;
wire n_10917;
wire n_7403;
wire n_13933;
wire n_6902;
wire n_6470;
wire n_14619;
wire n_9473;
wire n_10727;
wire n_11591;
wire n_10145;
wire n_12341;
wire n_9560;
wire n_5569;
wire n_8038;
wire n_10938;
wire n_15631;
wire n_15525;
wire n_9175;
wire n_8711;
wire n_10976;
wire n_5439;
wire n_8229;
wire n_8949;
wire n_14248;
wire n_14928;
wire n_10612;
wire n_5619;
wire n_4147;
wire n_15127;
wire n_6481;
wire n_9810;
wire n_14079;
wire n_4925;
wire n_7548;
wire n_9244;
wire n_14878;
wire n_15444;
wire n_9584;
wire n_12047;
wire n_6534;
wire n_11460;
wire n_15112;
wire n_13289;
wire n_4974;
wire n_8567;
wire n_10797;
wire n_13320;
wire n_9439;
wire n_11915;
wire n_14224;
wire n_13210;
wire n_14015;
wire n_4932;
wire n_4510;
wire n_8655;
wire n_9235;
wire n_6181;
wire n_8705;
wire n_6728;
wire n_11642;
wire n_15313;
wire n_9043;
wire n_9768;
wire n_11306;
wire n_14566;
wire n_13549;
wire n_5119;
wire n_9037;
wire n_15334;
wire n_12434;
wire n_5715;
wire n_9085;
wire n_8085;
wire n_14874;
wire n_8777;
wire n_6133;
wire n_11891;
wire n_14951;
wire n_8852;
wire n_9264;
wire n_6528;
wire n_10114;
wire n_7604;
wire n_7407;
wire n_14499;
wire n_8185;
wire n_12998;
wire n_13427;
wire n_10845;
wire n_4447;
wire n_8513;
wire n_15942;
wire n_6670;
wire n_12248;
wire n_14155;
wire n_16226;
wire n_6774;
wire n_8365;
wire n_11007;
wire n_14229;
wire n_4285;
wire n_5887;
wire n_4651;
wire n_6741;
wire n_7424;
wire n_11557;
wire n_12405;
wire n_6038;
wire n_4818;
wire n_15320;
wire n_7727;
wire n_4514;
wire n_4800;
wire n_10599;
wire n_11231;
wire n_9550;
wire n_9836;
wire n_13228;
wire n_6282;
wire n_13244;
wire n_9929;
wire n_12134;
wire n_15877;
wire n_8035;
wire n_8505;
wire n_11399;
wire n_11092;
wire n_4433;
wire n_11163;
wire n_8874;
wire n_11542;
wire n_10008;
wire n_16195;
wire n_6700;
wire n_15362;
wire n_15742;
wire n_7334;
wire n_8098;
wire n_7684;
wire n_7755;
wire n_10623;
wire n_4341;
wire n_9187;
wire n_13880;
wire n_11276;
wire n_4312;
wire n_10511;
wire n_12770;
wire n_5932;
wire n_13011;
wire n_14418;
wire n_15629;
wire n_6178;
wire n_11575;
wire n_10503;
wire n_6234;
wire n_15226;
wire n_15180;
wire n_14880;
wire n_11732;
wire n_6012;
wire n_4633;
wire n_14518;
wire n_9406;
wire n_10857;
wire n_9342;
wire n_13323;
wire n_4277;
wire n_13222;
wire n_13604;
wire n_14119;
wire n_14321;
wire n_15146;
wire n_15279;
wire n_7787;
wire n_14808;
wire n_15750;
wire n_4140;
wire n_8067;
wire n_12421;
wire n_5092;
wire n_10708;
wire n_14136;
wire n_13106;
wire n_14950;
wire n_15961;
wire n_7849;
wire n_12550;
wire n_5186;
wire n_13126;
wire n_15772;
wire n_11045;
wire n_7367;
wire n_8619;
wire n_9851;
wire n_9559;
wire n_11993;
wire n_14818;
wire n_15448;
wire n_11508;
wire n_12755;
wire n_8679;
wire n_9806;
wire n_8644;
wire n_12306;
wire n_12965;
wire n_11982;
wire n_10516;
wire n_4662;
wire n_6715;
wire n_11395;
wire n_5828;
wire n_11634;
wire n_7200;
wire n_13068;
wire n_9860;
wire n_4882;
wire n_4993;
wire n_11887;
wire n_11301;
wire n_15031;
wire n_7582;
wire n_4832;
wire n_4207;
wire n_4545;
wire n_13402;
wire n_6337;
wire n_13997;
wire n_4868;
wire n_8923;
wire n_8970;
wire n_10119;
wire n_8332;
wire n_14302;
wire n_10548;
wire n_11010;
wire n_11408;
wire n_15182;
wire n_8632;
wire n_14829;
wire n_6770;
wire n_7745;
wire n_6743;
wire n_8876;
wire n_10733;
wire n_10547;
wire n_11670;
wire n_13218;
wire n_14011;
wire n_5238;
wire n_10067;
wire n_14646;
wire n_13958;
wire n_13239;
wire n_8856;
wire n_12603;
wire n_14230;
wire n_11604;
wire n_15907;
wire n_9240;
wire n_4595;
wire n_7877;
wire n_11506;
wire n_11666;
wire n_8945;
wire n_11503;
wire n_8918;
wire n_14433;
wire n_16140;
wire n_7799;
wire n_16022;
wire n_6682;
wire n_5054;
wire n_7673;
wire n_11857;
wire n_15886;
wire n_5631;
wire n_8028;
wire n_6539;
wire n_16035;
wire n_7243;
wire n_7179;
wire n_9345;
wire n_5399;
wire n_6314;
wire n_6617;
wire n_10222;
wire n_11193;
wire n_13983;
wire n_11293;
wire n_12439;
wire n_5694;
wire n_4650;
wire n_4888;
wire n_8774;
wire n_7274;
wire n_5326;
wire n_12072;
wire n_14199;
wire n_15920;
wire n_8779;
wire n_13949;
wire n_8968;
wire n_13941;
wire n_4874;
wire n_7608;
wire n_8404;
wire n_4669;
wire n_13090;
wire n_6595;
wire n_4339;
wire n_12558;
wire n_12244;
wire n_12199;
wire n_11214;
wire n_5459;
wire n_7738;
wire n_13851;
wire n_14209;
wire n_14986;
wire n_9223;
wire n_9499;
wire n_10647;
wire n_14177;
wire n_14495;
wire n_11362;
wire n_11288;
wire n_11409;
wire n_15091;
wire n_5528;
wire n_13036;
wire n_11027;
wire n_12996;
wire n_5391;
wire n_12873;
wire n_8073;
wire n_4541;
wire n_7785;
wire n_5422;
wire n_13225;
wire n_16129;
wire n_6385;
wire n_14485;
wire n_6289;
wire n_12591;
wire n_5267;
wire n_4494;
wire n_10581;
wire n_13587;
wire n_5523;
wire n_16205;
wire n_4796;
wire n_7373;
wire n_9576;
wire n_9120;
wire n_14832;
wire n_14917;
wire n_10097;
wire n_10405;
wire n_15009;
wire n_6186;
wire n_4799;
wire n_5153;
wire n_12726;
wire n_9651;
wire n_12833;
wire n_14206;
wire n_6257;
wire n_14240;
wire n_12690;
wire n_11031;
wire n_14080;
wire n_13076;
wire n_15787;
wire n_9386;
wire n_11285;
wire n_10813;
wire n_6852;
wire n_6346;
wire n_11346;
wire n_12618;
wire n_16087;
wire n_4775;
wire n_9779;
wire n_5044;
wire n_5809;
wire n_12414;
wire n_11513;
wire n_16142;
wire n_5365;
wire n_14888;
wire n_7587;
wire n_13729;
wire n_5045;
wire n_4381;
wire n_4266;
wire n_11250;
wire n_7874;
wire n_11340;
wire n_5354;
wire n_15992;
wire n_4455;
wire n_6274;
wire n_14381;
wire n_14739;
wire n_7372;
wire n_7760;
wire n_10588;
wire n_15699;
wire n_4248;
wire n_9635;
wire n_5915;
wire n_6818;
wire n_9444;
wire n_10943;
wire n_11190;
wire n_7226;
wire n_5452;
wire n_8930;
wire n_4754;
wire n_13992;
wire n_7057;
wire n_12736;
wire n_7685;
wire n_8031;
wire n_11818;
wire n_8750;
wire n_14193;
wire n_15840;
wire n_14649;
wire n_4554;
wire n_5595;
wire n_6609;
wire n_6815;
wire n_6753;
wire n_4845;
wire n_9364;
wire n_9581;
wire n_9512;
wire n_9317;
wire n_14625;
wire n_14661;
wire n_14968;
wire n_8593;
wire n_14047;
wire n_13592;
wire n_4585;
wire n_7730;
wire n_14262;
wire n_14723;
wire n_13165;
wire n_8509;
wire n_9314;
wire n_9459;
wire n_8405;
wire n_13659;
wire n_14558;
wire n_9549;
wire n_11564;
wire n_10641;
wire n_7913;
wire n_4383;
wire n_11719;
wire n_8492;
wire n_6764;
wire n_14569;
wire n_5535;
wire n_15795;
wire n_9275;
wire n_13670;
wire n_15245;
wire n_15598;
wire n_15102;
wire n_10210;
wire n_5370;
wire n_11944;
wire n_13967;
wire n_7706;
wire n_7891;
wire n_6391;
wire n_13248;
wire n_16093;
wire n_11785;
wire n_8088;
wire n_5372;
wire n_5299;
wire n_5594;
wire n_4301;
wire n_11754;
wire n_4586;
wire n_14369;
wire n_14301;
wire n_9865;
wire n_6471;
wire n_11075;
wire n_15960;
wire n_11511;
wire n_12981;
wire n_13061;
wire n_13546;
wire n_6627;
wire n_10027;
wire n_5761;
wire n_10263;
wire n_10722;
wire n_14422;
wire n_13005;
wire n_13978;
wire n_11771;
wire n_4784;
wire n_7203;
wire n_8429;
wire n_8854;
wire n_9757;
wire n_15121;
wire n_7512;
wire n_5550;
wire n_12333;
wire n_11912;
wire n_15405;
wire n_5082;
wire n_9656;
wire n_15442;
wire n_10426;
wire n_11284;
wire n_5209;
wire n_7215;
wire n_15033;
wire n_10246;
wire n_6636;
wire n_13500;
wire n_4199;
wire n_13004;
wire n_10617;
wire n_5929;
wire n_16146;
wire n_10909;
wire n_15347;
wire n_5559;
wire n_12694;
wire n_13972;
wire n_14295;
wire n_5478;
wire n_11298;
wire n_15733;
wire n_7388;
wire n_16225;
wire n_7694;
wire n_6243;
wire n_6488;
wire n_4286;
wire n_9629;
wire n_13864;
wire n_11185;
wire n_5102;
wire n_11498;
wire n_6022;
wire n_8686;
wire n_6457;
wire n_10299;
wire n_4470;
wire n_12904;
wire n_7982;
wire n_13874;
wire n_11384;
wire n_10763;
wire n_10494;
wire n_13520;
wire n_8773;
wire n_10743;
wire n_8225;
wire n_8583;
wire n_4188;
wire n_6867;
wire n_8887;
wire n_9556;
wire n_15494;
wire n_5868;
wire n_6230;
wire n_6538;
wire n_15524;
wire n_12810;
wire n_15989;
wire n_9259;
wire n_9995;
wire n_14680;
wire n_15946;
wire n_12820;
wire n_6633;
wire n_9371;
wire n_8080;
wire n_11496;
wire n_6187;
wire n_15662;
wire n_6172;
wire n_13274;
wire n_10050;
wire n_13827;
wire n_5275;
wire n_14927;
wire n_15196;
wire n_10702;
wire n_4689;
wire n_13572;
wire n_14236;
wire n_5071;
wire n_7311;
wire n_15606;
wire n_5989;
wire n_8964;
wire n_11768;
wire n_15051;
wire n_12085;
wire n_14748;
wire n_9008;
wire n_6574;
wire n_11683;
wire n_11388;
wire n_13786;
wire n_8929;
wire n_8539;
wire n_6395;
wire n_4402;
wire n_9484;
wire n_15660;
wire n_8745;
wire n_4239;
wire n_6854;
wire n_7996;
wire n_6233;
wire n_4550;
wire n_6456;
wire n_8776;
wire n_8588;
wire n_8554;
wire n_9319;
wire n_15568;
wire n_11748;
wire n_7488;
wire n_5227;
wire n_13463;
wire n_9442;
wire n_14351;
wire n_10165;
wire n_14385;
wire n_7198;
wire n_4201;
wire n_10366;
wire n_12207;
wire n_8802;
wire n_13242;
wire n_13194;
wire n_9587;
wire n_6784;
wire n_14915;
wire n_6168;
wire n_16076;
wire n_13871;
wire n_14168;
wire n_9904;
wire n_9157;
wire n_8431;
wire n_8453;
wire n_6766;
wire n_5242;
wire n_8955;
wire n_12510;
wire n_8634;
wire n_14575;
wire n_4123;
wire n_6330;
wire n_15978;
wire n_5520;
wire n_8896;
wire n_14695;
wire n_4479;
wire n_7950;
wire n_7249;
wire n_13741;
wire n_9713;
wire n_11210;
wire n_9452;
wire n_10104;
wire n_16111;
wire n_15539;
wire n_14186;
wire n_5947;
wire n_7336;
wire n_4416;
wire n_8837;
wire n_7031;
wire n_4539;
wire n_8907;
wire n_6799;
wire n_10115;
wire n_14514;
wire n_14853;
wire n_13654;
wire n_8015;
wire n_14149;
wire n_10397;
wire n_14454;
wire n_9974;
wire n_13245;
wire n_15221;
wire n_10398;
wire n_5920;
wire n_6672;
wire n_13193;
wire n_6149;
wire n_8256;
wire n_13739;
wire n_14578;
wire n_10065;
wire n_11156;
wire n_12628;
wire n_10087;
wire n_14003;
wire n_7142;
wire n_11598;
wire n_13977;
wire n_5808;
wire n_15692;
wire n_6054;
wire n_7089;
wire n_11176;
wire n_12687;
wire n_4682;
wire n_7916;
wire n_12260;
wire n_6450;
wire n_5353;
wire n_5294;
wire n_12445;
wire n_13776;
wire n_8074;
wire n_12878;
wire n_14023;
wire n_4978;
wire n_4690;
wire n_10174;
wire n_12281;
wire n_10266;
wire n_12879;
wire n_16050;
wire n_10509;
wire n_12355;
wire n_4437;
wire n_5458;
wire n_5617;
wire n_4736;
wire n_7042;
wire n_8778;
wire n_8039;
wire n_10415;
wire n_5244;
wire n_6523;
wire n_13127;
wire n_5382;
wire n_14581;
wire n_8065;
wire n_6107;
wire n_9634;
wire n_12601;
wire n_12004;
wire n_11893;
wire n_11828;
wire n_6775;
wire n_5274;
wire n_10873;
wire n_12291;
wire n_8194;
wire n_4284;
wire n_14125;
wire n_11582;
wire n_8207;
wire n_13109;
wire n_10106;
wire n_12474;
wire n_13414;
wire n_9241;
wire n_6232;
wire n_13688;
wire n_6445;
wire n_10422;
wire n_10736;
wire n_7181;
wire n_6134;
wire n_5384;
wire n_9903;
wire n_15712;
wire n_8582;
wire n_10378;
wire n_6056;
wire n_8537;
wire n_6932;
wire n_13425;
wire n_7036;
wire n_4513;
wire n_9615;
wire n_8951;
wire n_7759;
wire n_9600;
wire n_11095;
wire n_7818;
wire n_11180;
wire n_9748;
wire n_9945;
wire n_5125;
wire n_12024;
wire n_9927;
wire n_15574;
wire n_5587;
wire n_6855;
wire n_14072;
wire n_11876;
wire n_5789;
wire n_8217;
wire n_10046;
wire n_15157;
wire n_13182;
wire n_14787;
wire n_16237;
wire n_13911;
wire n_16165;
wire n_5787;
wire n_6585;
wire n_6369;
wire n_5056;
wire n_10954;
wire n_10388;
wire n_14883;
wire n_8437;
wire n_5249;
wire n_8849;
wire n_7447;
wire n_10659;
wire n_13124;
wire n_13956;
wire n_14617;
wire n_7944;
wire n_5198;
wire n_11709;
wire n_5360;
wire n_10804;
wire n_7455;
wire n_5829;
wire n_5233;
wire n_4887;
wire n_4617;
wire n_9295;
wire n_5269;
wire n_13819;
wire n_11602;
wire n_11304;
wire n_6252;
wire n_12934;
wire n_5866;
wire n_6493;
wire n_14843;
wire n_8568;
wire n_10239;
wire n_12723;
wire n_7947;
wire n_12428;
wire n_10841;
wire n_12857;
wire n_13566;
wire n_14315;
wire n_9916;
wire n_4904;
wire n_8980;
wire n_13682;
wire n_5899;
wire n_11630;
wire n_13339;
wire n_7629;
wire n_13478;
wire n_8051;
wire n_4792;
wire n_7104;
wire n_8716;
wire n_11461;
wire n_9844;
wire n_15376;
wire n_7601;
wire n_4980;
wire n_11135;
wire n_15467;
wire n_15790;
wire n_12520;
wire n_14303;
wire n_11994;
wire n_15998;
wire n_12457;
wire n_12743;
wire n_6026;
wire n_15177;
wire n_4290;
wire n_7757;
wire n_8030;
wire n_5247;
wire n_9316;
wire n_9663;
wire n_13918;
wire n_15714;
wire n_10168;
wire n_13526;
wire n_5865;
wire n_13019;
wire n_14335;
wire n_10075;
wire n_15275;
wire n_6544;
wire n_5317;
wire n_14848;
wire n_14989;
wire n_10068;
wire n_11596;
wire n_10276;
wire n_15332;
wire n_12533;
wire n_8749;
wire n_11024;
wire n_7138;
wire n_7290;
wire n_14424;
wire n_8544;
wire n_13077;
wire n_15419;
wire n_13524;
wire n_8249;
wire n_12555;
wire n_9628;
wire n_14560;
wire n_6679;
wire n_8496;
wire n_9789;
wire n_14273;
wire n_13296;
wire n_13891;
wire n_4956;
wire n_14090;
wire n_5380;
wire n_5924;
wire n_12839;
wire n_7625;
wire n_5822;
wire n_10495;
wire n_9299;
wire n_6259;
wire n_12251;
wire n_4947;
wire n_7284;
wire n_11246;
wire n_14693;
wire n_11715;
wire n_4656;
wire n_12983;
wire n_12766;
wire n_6390;
wire n_12573;
wire n_12945;
wire n_11970;
wire n_15047;
wire n_4729;
wire n_14839;
wire n_5786;
wire n_4987;
wire n_13466;
wire n_5182;
wire n_4971;
wire n_11113;
wire n_12451;
wire n_7971;
wire n_15310;
wire n_12542;
wire n_12376;
wire n_9022;
wire n_10927;
wire n_6630;
wire n_15463;
wire n_13116;
wire n_12585;
wire n_10704;
wire n_5658;
wire n_16133;
wire n_11613;
wire n_5388;
wire n_13256;
wire n_13968;
wire n_4823;
wire n_13942;
wire n_9427;
wire n_4875;
wire n_13231;
wire n_6279;
wire n_8698;
wire n_8695;
wire n_9344;
wire n_14461;
wire n_12530;
wire n_13718;
wire n_8751;
wire n_15618;
wire n_15671;
wire n_15789;
wire n_15979;
wire n_10603;
wire n_12875;
wire n_11085;
wire n_15864;
wire n_6813;
wire n_9764;
wire n_15720;
wire n_12808;
wire n_5564;
wire n_11294;
wire n_13024;
wire n_8273;
wire n_14897;
wire n_11021;
wire n_15918;
wire n_14041;
wire n_14817;
wire n_15675;
wire n_9242;
wire n_9498;
wire n_8442;
wire n_14799;
wire n_7106;
wire n_8472;
wire n_9535;
wire n_6042;
wire n_7644;
wire n_12494;
wire n_6057;
wire n_4137;
wire n_7529;
wire n_8986;
wire n_10011;
wire n_11905;
wire n_6675;
wire n_12488;
wire n_4529;
wire n_4323;
wire n_12229;
wire n_13740;
wire n_6476;
wire n_8200;
wire n_14397;
wire n_10055;
wire n_7907;
wire n_13064;
wire n_10982;
wire n_8188;
wire n_11926;
wire n_12219;
wire n_8528;
wire n_11951;
wire n_13041;
wire n_14879;
wire n_6207;
wire n_5539;
wire n_10764;
wire n_16177;
wire n_14333;
wire n_6268;
wire n_6878;
wire n_6286;
wire n_9088;
wire n_15490;
wire n_12630;
wire n_6524;
wire n_10787;
wire n_5036;
wire n_12910;
wire n_5547;
wire n_4772;
wire n_6225;
wire n_4322;
wire n_8920;
wire n_8267;
wire n_12758;
wire n_13302;
wire n_10972;
wire n_7297;
wire n_6291;
wire n_5893;
wire n_4354;
wire n_4653;
wire n_12883;
wire n_16042;
wire n_9734;
wire n_9505;
wire n_9664;
wire n_12672;
wire n_7199;
wire n_14167;
wire n_5273;
wire n_10262;
wire n_10826;
wire n_8360;
wire n_13828;
wire n_4677;
wire n_8036;
wire n_9510;
wire n_5261;
wire n_16121;
wire n_11423;
wire n_6520;
wire n_14162;
wire n_7853;
wire n_7648;
wire n_9413;
wire n_9888;
wire n_14085;
wire n_8393;
wire n_11484;
wire n_8821;
wire n_11760;
wire n_9863;
wire n_12946;
wire n_13397;
wire n_10881;
wire n_8160;
wire n_9199;
wire n_11370;
wire n_5193;
wire n_10707;
wire n_9014;
wire n_10204;
wire n_9411;
wire n_12394;
wire n_12613;
wire n_12706;
wire n_4909;
wire n_11909;
wire n_13882;
wire n_9336;
wire n_9360;
wire n_10556;
wire n_9543;
wire n_15374;
wire n_6024;
wire n_7866;
wire n_5022;
wire n_13252;
wire n_14783;
wire n_5005;
wire n_13174;
wire n_7487;
wire n_15553;
wire n_10717;
wire n_6425;
wire n_13931;
wire n_5993;
wire n_13541;
wire n_12978;
wire n_14201;
wire n_14710;
wire n_12253;
wire n_7638;
wire n_8833;
wire n_14296;
wire n_5703;
wire n_15169;
wire n_8240;
wire n_12450;
wire n_14857;
wire n_4634;
wire n_7988;
wire n_13579;
wire n_9404;
wire n_14643;
wire n_8579;
wire n_5534;
wire n_6432;
wire n_14354;
wire n_9678;
wire n_16104;
wire n_12444;
wire n_8258;
wire n_9854;
wire n_7259;
wire n_11071;
wire n_11979;
wire n_15414;
wire n_13050;
wire n_8626;
wire n_13384;
wire n_12289;
wire n_6955;
wire n_6540;
wire n_9481;
wire n_5174;
wire n_10862;
wire n_4952;
wire n_12583;
wire n_15872;
wire n_5157;
wire n_13936;
wire n_4380;
wire n_9672;
wire n_14009;
wire n_9893;
wire n_4126;
wire n_7237;
wire n_8935;
wire n_11928;
wire n_5087;
wire n_12590;
wire n_12596;
wire n_6388;
wire n_4506;
wire n_10240;
wire n_5904;
wire n_9478;
wire n_13465;
wire n_4880;
wire n_11792;
wire n_9266;
wire n_9813;
wire n_12551;
wire n_14026;
wire n_6760;
wire n_13817;
wire n_8009;
wire n_11329;
wire n_15700;
wire n_4896;
wire n_15929;
wire n_5620;
wire n_5061;
wire n_5750;
wire n_5572;
wire n_7063;
wire n_10338;
wire n_10205;
wire n_12034;
wire n_14275;
wire n_11573;
wire n_11703;
wire n_9042;
wire n_4943;
wire n_11671;
wire n_8012;
wire n_11445;
wire n_14692;
wire n_7576;
wire n_9506;
wire n_8608;
wire n_13946;
wire n_15655;
wire n_8008;
wire n_12498;
wire n_10285;
wire n_14040;
wire n_6795;
wire n_14464;
wire n_5881;
wire n_8079;
wire n_6664;
wire n_15695;
wire n_16090;
wire n_12228;
wire n_5815;
wire n_12378;
wire n_11832;
wire n_6261;
wire n_15953;
wire n_4193;
wire n_5873;
wire n_13926;
wire n_9666;
wire n_10112;
wire n_15200;
wire n_14163;
wire n_6487;
wire n_9146;
wire n_4737;
wire n_7734;
wire n_6729;
wire n_15046;
wire n_10056;
wire n_9862;
wire n_5755;
wire n_10283;
wire n_9274;
wire n_15407;
wire n_15680;
wire n_8702;
wire n_5949;
wire n_10469;
wire n_15999;
wire n_13944;
wire n_5195;
wire n_7483;
wire n_4136;
wire n_15926;
wire n_6608;
wire n_15498;
wire n_14145;
wire n_7858;
wire n_9619;
wire n_12742;
wire n_15172;
wire n_7385;
wire n_4393;
wire n_11088;
wire n_12423;
wire n_10618;
wire n_13902;
wire n_8576;
wire n_9508;
wire n_4535;
wire n_10105;
wire n_7668;
wire n_13008;
wire n_8662;
wire n_15694;
wire n_4522;
wire n_6663;
wire n_4794;
wire n_13504;
wire n_5955;
wire n_7476;
wire n_15022;
wire n_7327;
wire n_5763;
wire n_6656;
wire n_8436;
wire n_11154;
wire n_13491;
wire n_9987;
wire n_8124;
wire n_8148;
wire n_14135;
wire n_12518;
wire n_15519;
wire n_8033;
wire n_6843;
wire n_12764;
wire n_7953;
wire n_8343;
wire n_5246;
wire n_5964;
wire n_11065;
wire n_13812;
wire n_12417;
wire n_8118;
wire n_14182;
wire n_13751;
wire n_15850;
wire n_12209;
wire n_15143;
wire n_12882;
wire n_7266;
wire n_5164;
wire n_11449;
wire n_4196;
wire n_6969;
wire n_11447;
wire n_8741;
wire n_12427;
wire n_13894;
wire n_14217;
wire n_4592;
wire n_4675;
wire n_5665;
wire n_6485;
wire n_5340;
wire n_14882;
wire n_5498;
wire n_7100;
wire n_15173;
wire n_15012;
wire n_4370;
wire n_14541;
wire n_5783;
wire n_11123;
wire n_8478;
wire n_5183;
wire n_11319;
wire n_11676;
wire n_6075;
wire n_7082;
wire n_9569;
wire n_15439;
wire n_6120;
wire n_6659;
wire n_13513;
wire n_6750;
wire n_15685;
wire n_15808;
wire n_11018;
wire n_5549;
wire n_9935;
wire n_14477;
wire n_9707;
wire n_13663;
wire n_14664;
wire n_8376;
wire n_9827;
wire n_7689;
wire n_13858;
wire n_4889;
wire n_15674;
wire n_7132;
wire n_11537;
wire n_8763;
wire n_13361;
wire n_5442;
wire n_13792;
wire n_5739;
wire n_7824;
wire n_8996;
wire n_12707;
wire n_15832;
wire n_15949;
wire n_16112;
wire n_13161;
wire n_9007;
wire n_4828;
wire n_9797;
wire n_13132;
wire n_6003;
wire n_16167;
wire n_5385;
wire n_8726;
wire n_13662;
wire n_8799;
wire n_4558;
wire n_7796;
wire n_10670;
wire n_9053;
wire n_6478;
wire n_6066;
wire n_15607;
wire n_15232;
wire n_9450;
wire n_13272;
wire n_15512;
wire n_12437;
wire n_7034;
wire n_6086;
wire n_9121;
wire n_6650;
wire n_4722;
wire n_6224;
wire n_10789;
wire n_14725;
wire n_10387;
wire n_8303;
wire n_8796;
wire n_4768;
wire n_12941;
wire n_10661;
wire n_13859;
wire n_11638;
wire n_14476;
wire n_4100;
wire n_10088;
wire n_12026;
wire n_10629;
wire n_15246;
wire n_14208;
wire n_13898;
wire n_7084;
wire n_5845;
wire n_9617;
wire n_9089;
wire n_8883;
wire n_7293;
wire n_10505;
wire n_8251;
wire n_10247;
wire n_9236;
wire n_5990;
wire n_6175;
wire n_10860;
wire n_15464;
wire n_15387;
wire n_6060;
wire n_7253;
wire n_6891;
wire n_5663;
wire n_12537;
wire n_14547;
wire n_9493;
wire n_8860;
wire n_14364;
wire n_8003;
wire n_6410;
wire n_12607;
wire n_5973;
wire n_4465;
wire n_15184;
wire n_12958;
wire n_12849;
wire n_16185;
wire n_14849;
wire n_15822;
wire n_5537;
wire n_5304;
wire n_8524;
wire n_13835;
wire n_13863;
wire n_6059;
wire n_15713;
wire n_16200;
wire n_5130;
wire n_12329;
wire n_13650;
wire n_8914;
wire n_10524;
wire n_7520;
wire n_12032;
wire n_12159;
wire n_5162;
wire n_4808;
wire n_8520;
wire n_9490;
wire n_12737;
wire n_6103;
wire n_6809;
wire n_10376;
wire n_4482;
wire n_15328;
wire n_11213;
wire n_10986;
wire n_12504;
wire n_12987;
wire n_14780;
wire n_6267;
wire n_8165;
wire n_15163;
wire n_11523;
wire n_9525;
wire n_9127;
wire n_9119;
wire n_12521;
wire n_5855;
wire n_11903;
wire n_9002;
wire n_10069;
wire n_10697;
wire n_15300;
wire n_11100;
wire n_13695;
wire n_12866;
wire n_14030;
wire n_8330;
wire n_12226;
wire n_8682;
wire n_5757;
wire n_6437;
wire n_7331;
wire n_6610;
wire n_7918;
wire n_12170;
wire n_11440;
wire n_10259;
wire n_8467;
wire n_13216;
wire n_8775;
wire n_8886;
wire n_10844;
wire n_15371;
wire n_12482;
wire n_4926;
wire n_11476;
wire n_8696;
wire n_16002;
wire n_4116;
wire n_14742;
wire n_6957;
wire n_14658;
wire n_15600;
wire n_5704;
wire n_7514;
wire n_11966;
wire n_10330;
wire n_15571;
wire n_7163;
wire n_7620;
wire n_11115;
wire n_16105;
wire n_9867;
wire n_5473;
wire n_15113;
wire n_11765;
wire n_4612;
wire n_5946;
wire n_10197;
wire n_6711;
wire n_14648;
wire n_15501;
wire n_8464;
wire n_12440;
wire n_4287;
wire n_15580;
wire n_13313;
wire n_7445;
wire n_10584;
wire n_6847;
wire n_9131;
wire n_9790;
wire n_10522;
wire n_5177;
wire n_15011;
wire n_11200;
wire n_16072;
wire n_10752;
wire n_16188;
wire n_15152;
wire n_11332;
wire n_15426;
wire n_7123;
wire n_6384;
wire n_10854;
wire n_16118;
wire n_15244;
wire n_15122;
wire n_4516;
wire n_11189;
wire n_12834;
wire n_10768;
wire n_14791;
wire n_8720;
wire n_14779;
wire n_4505;
wire n_7959;
wire n_10542;
wire n_9611;
wire n_15203;
wire n_15352;
wire n_7563;
wire n_15217;
wire n_6298;
wire n_11170;
wire n_11337;
wire n_13987;
wire n_9032;
wire n_14218;
wire n_14982;
wire n_9428;
wire n_9990;
wire n_16062;
wire n_7361;
wire n_12929;
wire n_11278;
wire n_16029;
wire n_4602;
wire n_8186;
wire n_5172;
wire n_4449;
wire n_9705;
wire n_8890;
wire n_13497;
wire n_7322;
wire n_8219;
wire n_5710;
wire n_7453;
wire n_6067;
wire n_9774;
wire n_5070;
wire n_14941;
wire n_12022;
wire n_15725;
wire n_6377;
wire n_12358;
wire n_13793;
wire n_12242;
wire n_4445;
wire n_14010;
wire n_5566;
wire n_10419;
wire n_5414;
wire n_8738;
wire n_16084;
wire n_13186;
wire n_4870;
wire n_10645;
wire n_11713;
wire n_15691;
wire n_12214;
wire n_13282;
wire n_13988;
wire n_6348;
wire n_7713;
wire n_10412;
wire n_4915;
wire n_15545;
wire n_6129;
wire n_5296;
wire n_5450;
wire n_15147;
wire n_11195;
wire n_6834;
wire n_10124;
wire n_11975;
wire n_5313;
wire n_12254;
wire n_13073;
wire n_13580;
wire n_14178;
wire n_14816;
wire n_12320;
wire n_9374;
wire n_14960;
wire n_4914;
wire n_10737;
wire n_9792;
wire n_6136;
wire n_7261;
wire n_6723;
wire n_5834;
wire n_14008;
wire n_8066;
wire n_5874;
wire n_14459;
wire n_16229;
wire n_7977;
wire n_14582;
wire n_14970;
wire n_10294;
wire n_14063;
wire n_10687;
wire n_12763;
wire n_11402;
wire n_14597;
wire n_14976;
wire n_8342;
wire n_13527;
wire n_7508;
wire n_9771;
wire n_10480;
wire n_15549;
wire n_9712;
wire n_7021;
wire n_13831;
wire n_12627;
wire n_5270;
wire n_11345;
wire n_5956;
wire n_7834;
wire n_14670;
wire n_4345;
wire n_16147;
wire n_14349;
wire n_5188;
wire n_9905;
wire n_8571;
wire n_6078;
wire n_7000;
wire n_9163;
wire n_9308;
wire n_10243;
wire n_15627;
wire n_4318;
wire n_10038;
wire n_10721;
wire n_15905;
wire n_7921;
wire n_8877;
wire n_4185;
wire n_16178;
wire n_8862;
wire n_16247;
wire n_10144;
wire n_8402;
wire n_10410;
wire n_4797;
wire n_7130;
wire n_10823;
wire n_15070;
wire n_10176;
wire n_11714;
wire n_5823;
wire n_13687;
wire n_5465;
wire n_9387;
wire n_7538;
wire n_11778;
wire n_12492;
wire n_13794;
wire n_7517;
wire n_14948;
wire n_5853;
wire n_15504;
wire n_14758;
wire n_10799;
wire n_15994;
wire n_10315;
wire n_7077;
wire n_11300;
wire n_12561;
wire n_14497;
wire n_4343;
wire n_13382;
wire n_11338;
wire n_4212;
wire n_12359;
wire n_15528;
wire n_6642;
wire n_4124;
wire n_11577;
wire n_15276;
wire n_5467;
wire n_5522;
wire n_4492;
wire n_7346;
wire n_10525;
wire n_11930;
wire n_5148;
wire n_4994;
wire n_13353;
wire n_15076;
wire n_7333;
wire n_4245;
wire n_4364;
wire n_4928;
wire n_11334;
wire n_4378;
wire n_16158;
wire n_7546;
wire n_4216;
wire n_9847;
wire n_12688;
wire n_5934;
wire n_6942;
wire n_8418;
wire n_10932;
wire n_10227;
wire n_11096;
wire n_9577;
wire n_10951;
wire n_4309;
wire n_9111;
wire n_8805;
wire n_10646;
wire n_6511;
wire n_15219;
wire n_12635;
wire n_6507;
wire n_12677;
wire n_14338;
wire n_9513;
wire n_12568;
wire n_11482;
wire n_14819;
wire n_9853;
wire n_11759;
wire n_10710;
wire n_15137;
wire n_7319;
wire n_7997;
wire n_12639;
wire n_6497;
wire n_6001;
wire n_6007;
wire n_9130;
wire n_10409;
wire n_9941;
wire n_9135;
wire n_14414;
wire n_6606;
wire n_4560;
wire n_10709;
wire n_10633;
wire n_5318;
wire n_11829;
wire n_5395;
wire n_14327;
wire n_13901;
wire n_15346;
wire n_7078;
wire n_15292;
wire n_7047;
wire n_8144;
wire n_5067;
wire n_7107;
wire n_10606;
wire n_13047;
wire n_14077;
wire n_16070;
wire n_13049;
wire n_11936;
wire n_10325;
wire n_7469;
wire n_15668;
wire n_13332;
wire n_14786;
wire n_8111;
wire n_11308;

INVx1_ASAP7_75t_L g4097 ( 
.A(n_488),
.Y(n_4097)
);

INVx1_ASAP7_75t_L g4098 ( 
.A(n_2595),
.Y(n_4098)
);

CKINVDCx5p33_ASAP7_75t_R g4099 ( 
.A(n_922),
.Y(n_4099)
);

CKINVDCx20_ASAP7_75t_R g4100 ( 
.A(n_1340),
.Y(n_4100)
);

BUFx6f_ASAP7_75t_L g4101 ( 
.A(n_3906),
.Y(n_4101)
);

CKINVDCx5p33_ASAP7_75t_R g4102 ( 
.A(n_3773),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_3115),
.Y(n_4103)
);

CKINVDCx5p33_ASAP7_75t_R g4104 ( 
.A(n_3898),
.Y(n_4104)
);

CKINVDCx5p33_ASAP7_75t_R g4105 ( 
.A(n_2510),
.Y(n_4105)
);

CKINVDCx5p33_ASAP7_75t_R g4106 ( 
.A(n_2568),
.Y(n_4106)
);

INVx2_ASAP7_75t_L g4107 ( 
.A(n_12),
.Y(n_4107)
);

CKINVDCx20_ASAP7_75t_R g4108 ( 
.A(n_2756),
.Y(n_4108)
);

BUFx6f_ASAP7_75t_L g4109 ( 
.A(n_1808),
.Y(n_4109)
);

CKINVDCx5p33_ASAP7_75t_R g4110 ( 
.A(n_3891),
.Y(n_4110)
);

CKINVDCx5p33_ASAP7_75t_R g4111 ( 
.A(n_3421),
.Y(n_4111)
);

CKINVDCx5p33_ASAP7_75t_R g4112 ( 
.A(n_4050),
.Y(n_4112)
);

CKINVDCx5p33_ASAP7_75t_R g4113 ( 
.A(n_3693),
.Y(n_4113)
);

INVx1_ASAP7_75t_L g4114 ( 
.A(n_4027),
.Y(n_4114)
);

CKINVDCx16_ASAP7_75t_R g4115 ( 
.A(n_3183),
.Y(n_4115)
);

BUFx3_ASAP7_75t_L g4116 ( 
.A(n_2558),
.Y(n_4116)
);

INVx1_ASAP7_75t_L g4117 ( 
.A(n_1835),
.Y(n_4117)
);

CKINVDCx5p33_ASAP7_75t_R g4118 ( 
.A(n_2042),
.Y(n_4118)
);

BUFx2_ASAP7_75t_L g4119 ( 
.A(n_3348),
.Y(n_4119)
);

CKINVDCx20_ASAP7_75t_R g4120 ( 
.A(n_1989),
.Y(n_4120)
);

INVx1_ASAP7_75t_L g4121 ( 
.A(n_651),
.Y(n_4121)
);

INVx1_ASAP7_75t_L g4122 ( 
.A(n_3466),
.Y(n_4122)
);

INVx1_ASAP7_75t_L g4123 ( 
.A(n_3623),
.Y(n_4123)
);

CKINVDCx5p33_ASAP7_75t_R g4124 ( 
.A(n_3992),
.Y(n_4124)
);

CKINVDCx5p33_ASAP7_75t_R g4125 ( 
.A(n_1485),
.Y(n_4125)
);

BUFx8_ASAP7_75t_SL g4126 ( 
.A(n_3597),
.Y(n_4126)
);

INVx1_ASAP7_75t_L g4127 ( 
.A(n_2493),
.Y(n_4127)
);

INVx1_ASAP7_75t_L g4128 ( 
.A(n_3019),
.Y(n_4128)
);

INVx1_ASAP7_75t_L g4129 ( 
.A(n_1357),
.Y(n_4129)
);

INVx1_ASAP7_75t_L g4130 ( 
.A(n_256),
.Y(n_4130)
);

CKINVDCx5p33_ASAP7_75t_R g4131 ( 
.A(n_1403),
.Y(n_4131)
);

CKINVDCx14_ASAP7_75t_R g4132 ( 
.A(n_3661),
.Y(n_4132)
);

BUFx3_ASAP7_75t_L g4133 ( 
.A(n_1674),
.Y(n_4133)
);

INVx1_ASAP7_75t_L g4134 ( 
.A(n_2982),
.Y(n_4134)
);

INVx1_ASAP7_75t_L g4135 ( 
.A(n_4009),
.Y(n_4135)
);

INVx1_ASAP7_75t_L g4136 ( 
.A(n_1173),
.Y(n_4136)
);

CKINVDCx5p33_ASAP7_75t_R g4137 ( 
.A(n_3976),
.Y(n_4137)
);

INVx1_ASAP7_75t_L g4138 ( 
.A(n_3926),
.Y(n_4138)
);

CKINVDCx5p33_ASAP7_75t_R g4139 ( 
.A(n_3818),
.Y(n_4139)
);

INVx1_ASAP7_75t_L g4140 ( 
.A(n_3371),
.Y(n_4140)
);

CKINVDCx5p33_ASAP7_75t_R g4141 ( 
.A(n_720),
.Y(n_4141)
);

CKINVDCx5p33_ASAP7_75t_R g4142 ( 
.A(n_3935),
.Y(n_4142)
);

CKINVDCx5p33_ASAP7_75t_R g4143 ( 
.A(n_2253),
.Y(n_4143)
);

CKINVDCx5p33_ASAP7_75t_R g4144 ( 
.A(n_2028),
.Y(n_4144)
);

CKINVDCx5p33_ASAP7_75t_R g4145 ( 
.A(n_1491),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_3423),
.Y(n_4146)
);

INVx1_ASAP7_75t_SL g4147 ( 
.A(n_1685),
.Y(n_4147)
);

CKINVDCx5p33_ASAP7_75t_R g4148 ( 
.A(n_2686),
.Y(n_4148)
);

CKINVDCx5p33_ASAP7_75t_R g4149 ( 
.A(n_3894),
.Y(n_4149)
);

CKINVDCx20_ASAP7_75t_R g4150 ( 
.A(n_2579),
.Y(n_4150)
);

CKINVDCx20_ASAP7_75t_R g4151 ( 
.A(n_2767),
.Y(n_4151)
);

INVx1_ASAP7_75t_L g4152 ( 
.A(n_3328),
.Y(n_4152)
);

CKINVDCx5p33_ASAP7_75t_R g4153 ( 
.A(n_2296),
.Y(n_4153)
);

CKINVDCx5p33_ASAP7_75t_R g4154 ( 
.A(n_2260),
.Y(n_4154)
);

CKINVDCx5p33_ASAP7_75t_R g4155 ( 
.A(n_2851),
.Y(n_4155)
);

CKINVDCx5p33_ASAP7_75t_R g4156 ( 
.A(n_3535),
.Y(n_4156)
);

CKINVDCx5p33_ASAP7_75t_R g4157 ( 
.A(n_636),
.Y(n_4157)
);

BUFx3_ASAP7_75t_L g4158 ( 
.A(n_3893),
.Y(n_4158)
);

INVx1_ASAP7_75t_L g4159 ( 
.A(n_3687),
.Y(n_4159)
);

CKINVDCx5p33_ASAP7_75t_R g4160 ( 
.A(n_3995),
.Y(n_4160)
);

INVx2_ASAP7_75t_L g4161 ( 
.A(n_3636),
.Y(n_4161)
);

CKINVDCx5p33_ASAP7_75t_R g4162 ( 
.A(n_1593),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_73),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_3993),
.Y(n_4164)
);

BUFx2_ASAP7_75t_SL g4165 ( 
.A(n_1808),
.Y(n_4165)
);

INVx1_ASAP7_75t_L g4166 ( 
.A(n_3430),
.Y(n_4166)
);

CKINVDCx16_ASAP7_75t_R g4167 ( 
.A(n_3590),
.Y(n_4167)
);

CKINVDCx5p33_ASAP7_75t_R g4168 ( 
.A(n_2010),
.Y(n_4168)
);

CKINVDCx5p33_ASAP7_75t_R g4169 ( 
.A(n_1409),
.Y(n_4169)
);

CKINVDCx5p33_ASAP7_75t_R g4170 ( 
.A(n_1096),
.Y(n_4170)
);

BUFx5_ASAP7_75t_L g4171 ( 
.A(n_3907),
.Y(n_4171)
);

INVx1_ASAP7_75t_L g4172 ( 
.A(n_3727),
.Y(n_4172)
);

INVx2_ASAP7_75t_L g4173 ( 
.A(n_2125),
.Y(n_4173)
);

HB1xp67_ASAP7_75t_L g4174 ( 
.A(n_4033),
.Y(n_4174)
);

INVx2_ASAP7_75t_L g4175 ( 
.A(n_4021),
.Y(n_4175)
);

CKINVDCx5p33_ASAP7_75t_R g4176 ( 
.A(n_734),
.Y(n_4176)
);

CKINVDCx20_ASAP7_75t_R g4177 ( 
.A(n_2892),
.Y(n_4177)
);

CKINVDCx5p33_ASAP7_75t_R g4178 ( 
.A(n_4058),
.Y(n_4178)
);

INVx1_ASAP7_75t_SL g4179 ( 
.A(n_1440),
.Y(n_4179)
);

CKINVDCx5p33_ASAP7_75t_R g4180 ( 
.A(n_3483),
.Y(n_4180)
);

BUFx6f_ASAP7_75t_L g4181 ( 
.A(n_2334),
.Y(n_4181)
);

INVx1_ASAP7_75t_L g4182 ( 
.A(n_4016),
.Y(n_4182)
);

CKINVDCx5p33_ASAP7_75t_R g4183 ( 
.A(n_2696),
.Y(n_4183)
);

INVxp67_ASAP7_75t_SL g4184 ( 
.A(n_3472),
.Y(n_4184)
);

INVx1_ASAP7_75t_L g4185 ( 
.A(n_3640),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_2276),
.Y(n_4186)
);

CKINVDCx5p33_ASAP7_75t_R g4187 ( 
.A(n_1158),
.Y(n_4187)
);

HB1xp67_ASAP7_75t_L g4188 ( 
.A(n_3897),
.Y(n_4188)
);

INVx2_ASAP7_75t_L g4189 ( 
.A(n_1041),
.Y(n_4189)
);

CKINVDCx5p33_ASAP7_75t_R g4190 ( 
.A(n_3203),
.Y(n_4190)
);

INVx2_ASAP7_75t_SL g4191 ( 
.A(n_3525),
.Y(n_4191)
);

CKINVDCx5p33_ASAP7_75t_R g4192 ( 
.A(n_1988),
.Y(n_4192)
);

CKINVDCx5p33_ASAP7_75t_R g4193 ( 
.A(n_2673),
.Y(n_4193)
);

CKINVDCx5p33_ASAP7_75t_R g4194 ( 
.A(n_3611),
.Y(n_4194)
);

INVx1_ASAP7_75t_L g4195 ( 
.A(n_2565),
.Y(n_4195)
);

INVx2_ASAP7_75t_L g4196 ( 
.A(n_2135),
.Y(n_4196)
);

CKINVDCx5p33_ASAP7_75t_R g4197 ( 
.A(n_476),
.Y(n_4197)
);

BUFx6f_ASAP7_75t_L g4198 ( 
.A(n_3299),
.Y(n_4198)
);

BUFx6f_ASAP7_75t_L g4199 ( 
.A(n_3244),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_3031),
.Y(n_4200)
);

INVx1_ASAP7_75t_L g4201 ( 
.A(n_1950),
.Y(n_4201)
);

INVx1_ASAP7_75t_L g4202 ( 
.A(n_4014),
.Y(n_4202)
);

CKINVDCx5p33_ASAP7_75t_R g4203 ( 
.A(n_1976),
.Y(n_4203)
);

CKINVDCx5p33_ASAP7_75t_R g4204 ( 
.A(n_3991),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_905),
.Y(n_4205)
);

CKINVDCx16_ASAP7_75t_R g4206 ( 
.A(n_3617),
.Y(n_4206)
);

CKINVDCx5p33_ASAP7_75t_R g4207 ( 
.A(n_3940),
.Y(n_4207)
);

CKINVDCx5p33_ASAP7_75t_R g4208 ( 
.A(n_916),
.Y(n_4208)
);

CKINVDCx20_ASAP7_75t_R g4209 ( 
.A(n_2558),
.Y(n_4209)
);

INVx1_ASAP7_75t_L g4210 ( 
.A(n_619),
.Y(n_4210)
);

CKINVDCx5p33_ASAP7_75t_R g4211 ( 
.A(n_3599),
.Y(n_4211)
);

INVx2_ASAP7_75t_SL g4212 ( 
.A(n_3435),
.Y(n_4212)
);

INVx1_ASAP7_75t_L g4213 ( 
.A(n_172),
.Y(n_4213)
);

INVx1_ASAP7_75t_L g4214 ( 
.A(n_849),
.Y(n_4214)
);

CKINVDCx5p33_ASAP7_75t_R g4215 ( 
.A(n_2019),
.Y(n_4215)
);

CKINVDCx5p33_ASAP7_75t_R g4216 ( 
.A(n_2485),
.Y(n_4216)
);

INVx1_ASAP7_75t_L g4217 ( 
.A(n_3590),
.Y(n_4217)
);

CKINVDCx5p33_ASAP7_75t_R g4218 ( 
.A(n_1918),
.Y(n_4218)
);

CKINVDCx5p33_ASAP7_75t_R g4219 ( 
.A(n_4026),
.Y(n_4219)
);

CKINVDCx5p33_ASAP7_75t_R g4220 ( 
.A(n_555),
.Y(n_4220)
);

BUFx5_ASAP7_75t_L g4221 ( 
.A(n_3318),
.Y(n_4221)
);

CKINVDCx5p33_ASAP7_75t_R g4222 ( 
.A(n_821),
.Y(n_4222)
);

CKINVDCx5p33_ASAP7_75t_R g4223 ( 
.A(n_2746),
.Y(n_4223)
);

CKINVDCx5p33_ASAP7_75t_R g4224 ( 
.A(n_1266),
.Y(n_4224)
);

CKINVDCx5p33_ASAP7_75t_R g4225 ( 
.A(n_702),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_1371),
.Y(n_4226)
);

BUFx8_ASAP7_75t_SL g4227 ( 
.A(n_553),
.Y(n_4227)
);

CKINVDCx5p33_ASAP7_75t_R g4228 ( 
.A(n_3854),
.Y(n_4228)
);

INVx2_ASAP7_75t_SL g4229 ( 
.A(n_3032),
.Y(n_4229)
);

CKINVDCx5p33_ASAP7_75t_R g4230 ( 
.A(n_2373),
.Y(n_4230)
);

CKINVDCx5p33_ASAP7_75t_R g4231 ( 
.A(n_3725),
.Y(n_4231)
);

CKINVDCx5p33_ASAP7_75t_R g4232 ( 
.A(n_2672),
.Y(n_4232)
);

BUFx2_ASAP7_75t_L g4233 ( 
.A(n_4023),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_2128),
.Y(n_4234)
);

CKINVDCx5p33_ASAP7_75t_R g4235 ( 
.A(n_164),
.Y(n_4235)
);

CKINVDCx5p33_ASAP7_75t_R g4236 ( 
.A(n_1992),
.Y(n_4236)
);

BUFx6f_ASAP7_75t_L g4237 ( 
.A(n_749),
.Y(n_4237)
);

CKINVDCx5p33_ASAP7_75t_R g4238 ( 
.A(n_1056),
.Y(n_4238)
);

CKINVDCx5p33_ASAP7_75t_R g4239 ( 
.A(n_3031),
.Y(n_4239)
);

CKINVDCx5p33_ASAP7_75t_R g4240 ( 
.A(n_2754),
.Y(n_4240)
);

BUFx3_ASAP7_75t_L g4241 ( 
.A(n_1878),
.Y(n_4241)
);

CKINVDCx5p33_ASAP7_75t_R g4242 ( 
.A(n_3599),
.Y(n_4242)
);

CKINVDCx5p33_ASAP7_75t_R g4243 ( 
.A(n_230),
.Y(n_4243)
);

CKINVDCx5p33_ASAP7_75t_R g4244 ( 
.A(n_54),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_2377),
.Y(n_4245)
);

CKINVDCx5p33_ASAP7_75t_R g4246 ( 
.A(n_4024),
.Y(n_4246)
);

CKINVDCx5p33_ASAP7_75t_R g4247 ( 
.A(n_1579),
.Y(n_4247)
);

CKINVDCx5p33_ASAP7_75t_R g4248 ( 
.A(n_1827),
.Y(n_4248)
);

CKINVDCx20_ASAP7_75t_R g4249 ( 
.A(n_378),
.Y(n_4249)
);

BUFx6f_ASAP7_75t_L g4250 ( 
.A(n_1937),
.Y(n_4250)
);

BUFx6f_ASAP7_75t_L g4251 ( 
.A(n_1587),
.Y(n_4251)
);

INVx1_ASAP7_75t_L g4252 ( 
.A(n_356),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_3363),
.Y(n_4253)
);

BUFx10_ASAP7_75t_L g4254 ( 
.A(n_1007),
.Y(n_4254)
);

CKINVDCx5p33_ASAP7_75t_R g4255 ( 
.A(n_340),
.Y(n_4255)
);

INVx3_ASAP7_75t_L g4256 ( 
.A(n_2851),
.Y(n_4256)
);

CKINVDCx20_ASAP7_75t_R g4257 ( 
.A(n_1098),
.Y(n_4257)
);

BUFx3_ASAP7_75t_L g4258 ( 
.A(n_3217),
.Y(n_4258)
);

CKINVDCx5p33_ASAP7_75t_R g4259 ( 
.A(n_3792),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_1045),
.Y(n_4260)
);

CKINVDCx5p33_ASAP7_75t_R g4261 ( 
.A(n_3373),
.Y(n_4261)
);

CKINVDCx5p33_ASAP7_75t_R g4262 ( 
.A(n_663),
.Y(n_4262)
);

CKINVDCx5p33_ASAP7_75t_R g4263 ( 
.A(n_47),
.Y(n_4263)
);

CKINVDCx5p33_ASAP7_75t_R g4264 ( 
.A(n_3866),
.Y(n_4264)
);

CKINVDCx5p33_ASAP7_75t_R g4265 ( 
.A(n_298),
.Y(n_4265)
);

INVx1_ASAP7_75t_L g4266 ( 
.A(n_205),
.Y(n_4266)
);

INVx1_ASAP7_75t_L g4267 ( 
.A(n_843),
.Y(n_4267)
);

CKINVDCx5p33_ASAP7_75t_R g4268 ( 
.A(n_1024),
.Y(n_4268)
);

HB1xp67_ASAP7_75t_L g4269 ( 
.A(n_2209),
.Y(n_4269)
);

INVxp67_ASAP7_75t_L g4270 ( 
.A(n_1088),
.Y(n_4270)
);

CKINVDCx5p33_ASAP7_75t_R g4271 ( 
.A(n_382),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_1726),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_3856),
.Y(n_4273)
);

INVx1_ASAP7_75t_L g4274 ( 
.A(n_3732),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_3416),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_448),
.Y(n_4276)
);

BUFx2_ASAP7_75t_L g4277 ( 
.A(n_3361),
.Y(n_4277)
);

INVx2_ASAP7_75t_L g4278 ( 
.A(n_365),
.Y(n_4278)
);

CKINVDCx5p33_ASAP7_75t_R g4279 ( 
.A(n_1581),
.Y(n_4279)
);

CKINVDCx20_ASAP7_75t_R g4280 ( 
.A(n_1437),
.Y(n_4280)
);

CKINVDCx5p33_ASAP7_75t_R g4281 ( 
.A(n_7),
.Y(n_4281)
);

INVx2_ASAP7_75t_L g4282 ( 
.A(n_557),
.Y(n_4282)
);

CKINVDCx16_ASAP7_75t_R g4283 ( 
.A(n_2339),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_207),
.Y(n_4284)
);

CKINVDCx5p33_ASAP7_75t_R g4285 ( 
.A(n_501),
.Y(n_4285)
);

INVx1_ASAP7_75t_L g4286 ( 
.A(n_674),
.Y(n_4286)
);

BUFx10_ASAP7_75t_L g4287 ( 
.A(n_3942),
.Y(n_4287)
);

INVx1_ASAP7_75t_L g4288 ( 
.A(n_4020),
.Y(n_4288)
);

INVx1_ASAP7_75t_L g4289 ( 
.A(n_1217),
.Y(n_4289)
);

CKINVDCx5p33_ASAP7_75t_R g4290 ( 
.A(n_491),
.Y(n_4290)
);

INVx2_ASAP7_75t_SL g4291 ( 
.A(n_2382),
.Y(n_4291)
);

BUFx3_ASAP7_75t_L g4292 ( 
.A(n_3825),
.Y(n_4292)
);

CKINVDCx5p33_ASAP7_75t_R g4293 ( 
.A(n_2175),
.Y(n_4293)
);

CKINVDCx5p33_ASAP7_75t_R g4294 ( 
.A(n_1744),
.Y(n_4294)
);

CKINVDCx5p33_ASAP7_75t_R g4295 ( 
.A(n_1853),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_910),
.Y(n_4296)
);

BUFx2_ASAP7_75t_L g4297 ( 
.A(n_3418),
.Y(n_4297)
);

CKINVDCx5p33_ASAP7_75t_R g4298 ( 
.A(n_2198),
.Y(n_4298)
);

BUFx6f_ASAP7_75t_L g4299 ( 
.A(n_1324),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_152),
.Y(n_4300)
);

BUFx2_ASAP7_75t_L g4301 ( 
.A(n_93),
.Y(n_4301)
);

CKINVDCx5p33_ASAP7_75t_R g4302 ( 
.A(n_3998),
.Y(n_4302)
);

CKINVDCx5p33_ASAP7_75t_R g4303 ( 
.A(n_750),
.Y(n_4303)
);

BUFx3_ASAP7_75t_L g4304 ( 
.A(n_2981),
.Y(n_4304)
);

CKINVDCx5p33_ASAP7_75t_R g4305 ( 
.A(n_1441),
.Y(n_4305)
);

CKINVDCx5p33_ASAP7_75t_R g4306 ( 
.A(n_3624),
.Y(n_4306)
);

CKINVDCx5p33_ASAP7_75t_R g4307 ( 
.A(n_2219),
.Y(n_4307)
);

INVx2_ASAP7_75t_L g4308 ( 
.A(n_3952),
.Y(n_4308)
);

CKINVDCx5p33_ASAP7_75t_R g4309 ( 
.A(n_2794),
.Y(n_4309)
);

CKINVDCx5p33_ASAP7_75t_R g4310 ( 
.A(n_2969),
.Y(n_4310)
);

INVx1_ASAP7_75t_L g4311 ( 
.A(n_479),
.Y(n_4311)
);

INVx2_ASAP7_75t_SL g4312 ( 
.A(n_1862),
.Y(n_4312)
);

CKINVDCx20_ASAP7_75t_R g4313 ( 
.A(n_253),
.Y(n_4313)
);

INVx1_ASAP7_75t_L g4314 ( 
.A(n_3861),
.Y(n_4314)
);

INVx1_ASAP7_75t_L g4315 ( 
.A(n_1343),
.Y(n_4315)
);

CKINVDCx5p33_ASAP7_75t_R g4316 ( 
.A(n_666),
.Y(n_4316)
);

INVxp67_ASAP7_75t_SL g4317 ( 
.A(n_3623),
.Y(n_4317)
);

BUFx10_ASAP7_75t_L g4318 ( 
.A(n_210),
.Y(n_4318)
);

INVx1_ASAP7_75t_SL g4319 ( 
.A(n_2853),
.Y(n_4319)
);

CKINVDCx20_ASAP7_75t_R g4320 ( 
.A(n_3806),
.Y(n_4320)
);

CKINVDCx5p33_ASAP7_75t_R g4321 ( 
.A(n_2578),
.Y(n_4321)
);

CKINVDCx5p33_ASAP7_75t_R g4322 ( 
.A(n_994),
.Y(n_4322)
);

CKINVDCx5p33_ASAP7_75t_R g4323 ( 
.A(n_1632),
.Y(n_4323)
);

CKINVDCx5p33_ASAP7_75t_R g4324 ( 
.A(n_3519),
.Y(n_4324)
);

INVx1_ASAP7_75t_L g4325 ( 
.A(n_3969),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_27),
.Y(n_4326)
);

CKINVDCx5p33_ASAP7_75t_R g4327 ( 
.A(n_2532),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_487),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_3436),
.Y(n_4329)
);

INVx1_ASAP7_75t_SL g4330 ( 
.A(n_1457),
.Y(n_4330)
);

INVx1_ASAP7_75t_L g4331 ( 
.A(n_2228),
.Y(n_4331)
);

CKINVDCx5p33_ASAP7_75t_R g4332 ( 
.A(n_1784),
.Y(n_4332)
);

CKINVDCx5p33_ASAP7_75t_R g4333 ( 
.A(n_3930),
.Y(n_4333)
);

INVx1_ASAP7_75t_L g4334 ( 
.A(n_2288),
.Y(n_4334)
);

CKINVDCx5p33_ASAP7_75t_R g4335 ( 
.A(n_2774),
.Y(n_4335)
);

INVx1_ASAP7_75t_SL g4336 ( 
.A(n_1889),
.Y(n_4336)
);

BUFx3_ASAP7_75t_L g4337 ( 
.A(n_2759),
.Y(n_4337)
);

INVxp67_ASAP7_75t_L g4338 ( 
.A(n_1598),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_1029),
.Y(n_4339)
);

CKINVDCx5p33_ASAP7_75t_R g4340 ( 
.A(n_1647),
.Y(n_4340)
);

INVx1_ASAP7_75t_L g4341 ( 
.A(n_2393),
.Y(n_4341)
);

INVx1_ASAP7_75t_L g4342 ( 
.A(n_4037),
.Y(n_4342)
);

CKINVDCx5p33_ASAP7_75t_R g4343 ( 
.A(n_788),
.Y(n_4343)
);

INVx1_ASAP7_75t_L g4344 ( 
.A(n_3903),
.Y(n_4344)
);

CKINVDCx5p33_ASAP7_75t_R g4345 ( 
.A(n_174),
.Y(n_4345)
);

INVx2_ASAP7_75t_L g4346 ( 
.A(n_4072),
.Y(n_4346)
);

BUFx6f_ASAP7_75t_L g4347 ( 
.A(n_3963),
.Y(n_4347)
);

CKINVDCx20_ASAP7_75t_R g4348 ( 
.A(n_1735),
.Y(n_4348)
);

CKINVDCx5p33_ASAP7_75t_R g4349 ( 
.A(n_3934),
.Y(n_4349)
);

INVx1_ASAP7_75t_L g4350 ( 
.A(n_2534),
.Y(n_4350)
);

CKINVDCx5p33_ASAP7_75t_R g4351 ( 
.A(n_2516),
.Y(n_4351)
);

CKINVDCx5p33_ASAP7_75t_R g4352 ( 
.A(n_3396),
.Y(n_4352)
);

CKINVDCx5p33_ASAP7_75t_R g4353 ( 
.A(n_1792),
.Y(n_4353)
);

CKINVDCx5p33_ASAP7_75t_R g4354 ( 
.A(n_1239),
.Y(n_4354)
);

CKINVDCx5p33_ASAP7_75t_R g4355 ( 
.A(n_3165),
.Y(n_4355)
);

CKINVDCx5p33_ASAP7_75t_R g4356 ( 
.A(n_1096),
.Y(n_4356)
);

INVx1_ASAP7_75t_SL g4357 ( 
.A(n_1410),
.Y(n_4357)
);

CKINVDCx5p33_ASAP7_75t_R g4358 ( 
.A(n_553),
.Y(n_4358)
);

INVx1_ASAP7_75t_SL g4359 ( 
.A(n_3477),
.Y(n_4359)
);

CKINVDCx5p33_ASAP7_75t_R g4360 ( 
.A(n_3569),
.Y(n_4360)
);

CKINVDCx5p33_ASAP7_75t_R g4361 ( 
.A(n_3498),
.Y(n_4361)
);

INVxp67_ASAP7_75t_SL g4362 ( 
.A(n_3570),
.Y(n_4362)
);

INVx1_ASAP7_75t_L g4363 ( 
.A(n_1980),
.Y(n_4363)
);

CKINVDCx5p33_ASAP7_75t_R g4364 ( 
.A(n_3939),
.Y(n_4364)
);

CKINVDCx5p33_ASAP7_75t_R g4365 ( 
.A(n_2683),
.Y(n_4365)
);

BUFx6f_ASAP7_75t_L g4366 ( 
.A(n_629),
.Y(n_4366)
);

INVx1_ASAP7_75t_L g4367 ( 
.A(n_891),
.Y(n_4367)
);

CKINVDCx5p33_ASAP7_75t_R g4368 ( 
.A(n_3969),
.Y(n_4368)
);

CKINVDCx5p33_ASAP7_75t_R g4369 ( 
.A(n_1628),
.Y(n_4369)
);

CKINVDCx5p33_ASAP7_75t_R g4370 ( 
.A(n_181),
.Y(n_4370)
);

CKINVDCx20_ASAP7_75t_R g4371 ( 
.A(n_656),
.Y(n_4371)
);

CKINVDCx5p33_ASAP7_75t_R g4372 ( 
.A(n_3680),
.Y(n_4372)
);

CKINVDCx5p33_ASAP7_75t_R g4373 ( 
.A(n_1619),
.Y(n_4373)
);

CKINVDCx5p33_ASAP7_75t_R g4374 ( 
.A(n_945),
.Y(n_4374)
);

INVx1_ASAP7_75t_L g4375 ( 
.A(n_1581),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_4025),
.Y(n_4376)
);

CKINVDCx5p33_ASAP7_75t_R g4377 ( 
.A(n_936),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_2534),
.Y(n_4378)
);

CKINVDCx5p33_ASAP7_75t_R g4379 ( 
.A(n_964),
.Y(n_4379)
);

CKINVDCx20_ASAP7_75t_R g4380 ( 
.A(n_1932),
.Y(n_4380)
);

CKINVDCx5p33_ASAP7_75t_R g4381 ( 
.A(n_1727),
.Y(n_4381)
);

BUFx3_ASAP7_75t_L g4382 ( 
.A(n_1736),
.Y(n_4382)
);

CKINVDCx5p33_ASAP7_75t_R g4383 ( 
.A(n_3327),
.Y(n_4383)
);

CKINVDCx5p33_ASAP7_75t_R g4384 ( 
.A(n_484),
.Y(n_4384)
);

CKINVDCx5p33_ASAP7_75t_R g4385 ( 
.A(n_3728),
.Y(n_4385)
);

BUFx2_ASAP7_75t_SL g4386 ( 
.A(n_2899),
.Y(n_4386)
);

CKINVDCx5p33_ASAP7_75t_R g4387 ( 
.A(n_1560),
.Y(n_4387)
);

CKINVDCx5p33_ASAP7_75t_R g4388 ( 
.A(n_490),
.Y(n_4388)
);

BUFx2_ASAP7_75t_L g4389 ( 
.A(n_3226),
.Y(n_4389)
);

CKINVDCx5p33_ASAP7_75t_R g4390 ( 
.A(n_2022),
.Y(n_4390)
);

CKINVDCx5p33_ASAP7_75t_R g4391 ( 
.A(n_321),
.Y(n_4391)
);

CKINVDCx5p33_ASAP7_75t_R g4392 ( 
.A(n_380),
.Y(n_4392)
);

INVx1_ASAP7_75t_L g4393 ( 
.A(n_868),
.Y(n_4393)
);

BUFx6f_ASAP7_75t_L g4394 ( 
.A(n_1207),
.Y(n_4394)
);

INVx1_ASAP7_75t_L g4395 ( 
.A(n_4013),
.Y(n_4395)
);

INVx2_ASAP7_75t_L g4396 ( 
.A(n_3116),
.Y(n_4396)
);

BUFx3_ASAP7_75t_L g4397 ( 
.A(n_274),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_3046),
.Y(n_4398)
);

CKINVDCx5p33_ASAP7_75t_R g4399 ( 
.A(n_479),
.Y(n_4399)
);

INVx1_ASAP7_75t_L g4400 ( 
.A(n_711),
.Y(n_4400)
);

CKINVDCx5p33_ASAP7_75t_R g4401 ( 
.A(n_3382),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_3719),
.Y(n_4402)
);

CKINVDCx20_ASAP7_75t_R g4403 ( 
.A(n_4028),
.Y(n_4403)
);

INVx2_ASAP7_75t_L g4404 ( 
.A(n_1305),
.Y(n_4404)
);

CKINVDCx5p33_ASAP7_75t_R g4405 ( 
.A(n_515),
.Y(n_4405)
);

CKINVDCx20_ASAP7_75t_R g4406 ( 
.A(n_2232),
.Y(n_4406)
);

CKINVDCx5p33_ASAP7_75t_R g4407 ( 
.A(n_3924),
.Y(n_4407)
);

CKINVDCx5p33_ASAP7_75t_R g4408 ( 
.A(n_1035),
.Y(n_4408)
);

INVx1_ASAP7_75t_SL g4409 ( 
.A(n_2219),
.Y(n_4409)
);

CKINVDCx5p33_ASAP7_75t_R g4410 ( 
.A(n_122),
.Y(n_4410)
);

CKINVDCx5p33_ASAP7_75t_R g4411 ( 
.A(n_3247),
.Y(n_4411)
);

INVx1_ASAP7_75t_L g4412 ( 
.A(n_658),
.Y(n_4412)
);

INVx1_ASAP7_75t_L g4413 ( 
.A(n_24),
.Y(n_4413)
);

CKINVDCx5p33_ASAP7_75t_R g4414 ( 
.A(n_2765),
.Y(n_4414)
);

CKINVDCx5p33_ASAP7_75t_R g4415 ( 
.A(n_2715),
.Y(n_4415)
);

INVx1_ASAP7_75t_L g4416 ( 
.A(n_4095),
.Y(n_4416)
);

INVx2_ASAP7_75t_L g4417 ( 
.A(n_379),
.Y(n_4417)
);

INVx1_ASAP7_75t_L g4418 ( 
.A(n_2734),
.Y(n_4418)
);

CKINVDCx5p33_ASAP7_75t_R g4419 ( 
.A(n_1356),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_639),
.Y(n_4420)
);

INVx1_ASAP7_75t_L g4421 ( 
.A(n_613),
.Y(n_4421)
);

CKINVDCx5p33_ASAP7_75t_R g4422 ( 
.A(n_3543),
.Y(n_4422)
);

INVx1_ASAP7_75t_L g4423 ( 
.A(n_3238),
.Y(n_4423)
);

INVx2_ASAP7_75t_SL g4424 ( 
.A(n_2618),
.Y(n_4424)
);

BUFx3_ASAP7_75t_L g4425 ( 
.A(n_210),
.Y(n_4425)
);

CKINVDCx5p33_ASAP7_75t_R g4426 ( 
.A(n_1145),
.Y(n_4426)
);

CKINVDCx5p33_ASAP7_75t_R g4427 ( 
.A(n_2224),
.Y(n_4427)
);

INVx4_ASAP7_75t_R g4428 ( 
.A(n_320),
.Y(n_4428)
);

BUFx2_ASAP7_75t_L g4429 ( 
.A(n_3927),
.Y(n_4429)
);

CKINVDCx5p33_ASAP7_75t_R g4430 ( 
.A(n_1151),
.Y(n_4430)
);

INVx3_ASAP7_75t_L g4431 ( 
.A(n_1561),
.Y(n_4431)
);

INVx2_ASAP7_75t_L g4432 ( 
.A(n_3412),
.Y(n_4432)
);

CKINVDCx5p33_ASAP7_75t_R g4433 ( 
.A(n_3273),
.Y(n_4433)
);

INVx1_ASAP7_75t_L g4434 ( 
.A(n_1006),
.Y(n_4434)
);

INVx1_ASAP7_75t_L g4435 ( 
.A(n_1489),
.Y(n_4435)
);

INVx1_ASAP7_75t_L g4436 ( 
.A(n_1189),
.Y(n_4436)
);

CKINVDCx5p33_ASAP7_75t_R g4437 ( 
.A(n_3132),
.Y(n_4437)
);

INVx1_ASAP7_75t_L g4438 ( 
.A(n_868),
.Y(n_4438)
);

INVx2_ASAP7_75t_L g4439 ( 
.A(n_818),
.Y(n_4439)
);

CKINVDCx5p33_ASAP7_75t_R g4440 ( 
.A(n_3598),
.Y(n_4440)
);

CKINVDCx5p33_ASAP7_75t_R g4441 ( 
.A(n_3262),
.Y(n_4441)
);

CKINVDCx5p33_ASAP7_75t_R g4442 ( 
.A(n_1692),
.Y(n_4442)
);

INVx2_ASAP7_75t_SL g4443 ( 
.A(n_58),
.Y(n_4443)
);

INVx1_ASAP7_75t_L g4444 ( 
.A(n_580),
.Y(n_4444)
);

CKINVDCx20_ASAP7_75t_R g4445 ( 
.A(n_3443),
.Y(n_4445)
);

CKINVDCx5p33_ASAP7_75t_R g4446 ( 
.A(n_3958),
.Y(n_4446)
);

CKINVDCx5p33_ASAP7_75t_R g4447 ( 
.A(n_1526),
.Y(n_4447)
);

CKINVDCx5p33_ASAP7_75t_R g4448 ( 
.A(n_1276),
.Y(n_4448)
);

CKINVDCx5p33_ASAP7_75t_R g4449 ( 
.A(n_640),
.Y(n_4449)
);

INVx1_ASAP7_75t_L g4450 ( 
.A(n_3298),
.Y(n_4450)
);

BUFx3_ASAP7_75t_L g4451 ( 
.A(n_3217),
.Y(n_4451)
);

INVx1_ASAP7_75t_L g4452 ( 
.A(n_1313),
.Y(n_4452)
);

BUFx6f_ASAP7_75t_L g4453 ( 
.A(n_4029),
.Y(n_4453)
);

CKINVDCx5p33_ASAP7_75t_R g4454 ( 
.A(n_1557),
.Y(n_4454)
);

CKINVDCx5p33_ASAP7_75t_R g4455 ( 
.A(n_3207),
.Y(n_4455)
);

CKINVDCx5p33_ASAP7_75t_R g4456 ( 
.A(n_3932),
.Y(n_4456)
);

INVx1_ASAP7_75t_L g4457 ( 
.A(n_4037),
.Y(n_4457)
);

INVx1_ASAP7_75t_L g4458 ( 
.A(n_537),
.Y(n_4458)
);

INVx1_ASAP7_75t_L g4459 ( 
.A(n_3770),
.Y(n_4459)
);

INVx1_ASAP7_75t_L g4460 ( 
.A(n_1227),
.Y(n_4460)
);

CKINVDCx5p33_ASAP7_75t_R g4461 ( 
.A(n_3396),
.Y(n_4461)
);

CKINVDCx5p33_ASAP7_75t_R g4462 ( 
.A(n_85),
.Y(n_4462)
);

INVx2_ASAP7_75t_L g4463 ( 
.A(n_2040),
.Y(n_4463)
);

INVx1_ASAP7_75t_L g4464 ( 
.A(n_1095),
.Y(n_4464)
);

CKINVDCx5p33_ASAP7_75t_R g4465 ( 
.A(n_2962),
.Y(n_4465)
);

BUFx2_ASAP7_75t_L g4466 ( 
.A(n_516),
.Y(n_4466)
);

CKINVDCx5p33_ASAP7_75t_R g4467 ( 
.A(n_933),
.Y(n_4467)
);

BUFx3_ASAP7_75t_L g4468 ( 
.A(n_153),
.Y(n_4468)
);

HB1xp67_ASAP7_75t_L g4469 ( 
.A(n_3984),
.Y(n_4469)
);

INVx1_ASAP7_75t_L g4470 ( 
.A(n_4010),
.Y(n_4470)
);

CKINVDCx5p33_ASAP7_75t_R g4471 ( 
.A(n_3770),
.Y(n_4471)
);

INVx1_ASAP7_75t_L g4472 ( 
.A(n_3971),
.Y(n_4472)
);

CKINVDCx5p33_ASAP7_75t_R g4473 ( 
.A(n_2650),
.Y(n_4473)
);

INVx1_ASAP7_75t_L g4474 ( 
.A(n_1310),
.Y(n_4474)
);

CKINVDCx5p33_ASAP7_75t_R g4475 ( 
.A(n_990),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_3914),
.Y(n_4476)
);

INVx1_ASAP7_75t_L g4477 ( 
.A(n_3073),
.Y(n_4477)
);

CKINVDCx14_ASAP7_75t_R g4478 ( 
.A(n_3155),
.Y(n_4478)
);

CKINVDCx5p33_ASAP7_75t_R g4479 ( 
.A(n_3420),
.Y(n_4479)
);

BUFx3_ASAP7_75t_L g4480 ( 
.A(n_2597),
.Y(n_4480)
);

CKINVDCx5p33_ASAP7_75t_R g4481 ( 
.A(n_2880),
.Y(n_4481)
);

CKINVDCx5p33_ASAP7_75t_R g4482 ( 
.A(n_3847),
.Y(n_4482)
);

CKINVDCx16_ASAP7_75t_R g4483 ( 
.A(n_1095),
.Y(n_4483)
);

CKINVDCx5p33_ASAP7_75t_R g4484 ( 
.A(n_1706),
.Y(n_4484)
);

BUFx5_ASAP7_75t_L g4485 ( 
.A(n_2261),
.Y(n_4485)
);

CKINVDCx5p33_ASAP7_75t_R g4486 ( 
.A(n_3341),
.Y(n_4486)
);

INVx1_ASAP7_75t_L g4487 ( 
.A(n_3978),
.Y(n_4487)
);

BUFx5_ASAP7_75t_L g4488 ( 
.A(n_3024),
.Y(n_4488)
);

INVx2_ASAP7_75t_L g4489 ( 
.A(n_1543),
.Y(n_4489)
);

BUFx6f_ASAP7_75t_L g4490 ( 
.A(n_3415),
.Y(n_4490)
);

INVx1_ASAP7_75t_L g4491 ( 
.A(n_1712),
.Y(n_4491)
);

INVx1_ASAP7_75t_L g4492 ( 
.A(n_343),
.Y(n_4492)
);

CKINVDCx5p33_ASAP7_75t_R g4493 ( 
.A(n_1541),
.Y(n_4493)
);

INVx2_ASAP7_75t_SL g4494 ( 
.A(n_3973),
.Y(n_4494)
);

BUFx2_ASAP7_75t_L g4495 ( 
.A(n_1021),
.Y(n_4495)
);

CKINVDCx20_ASAP7_75t_R g4496 ( 
.A(n_3736),
.Y(n_4496)
);

CKINVDCx5p33_ASAP7_75t_R g4497 ( 
.A(n_3560),
.Y(n_4497)
);

CKINVDCx20_ASAP7_75t_R g4498 ( 
.A(n_574),
.Y(n_4498)
);

BUFx2_ASAP7_75t_SL g4499 ( 
.A(n_2742),
.Y(n_4499)
);

INVxp67_ASAP7_75t_L g4500 ( 
.A(n_1687),
.Y(n_4500)
);

INVx1_ASAP7_75t_SL g4501 ( 
.A(n_2359),
.Y(n_4501)
);

CKINVDCx5p33_ASAP7_75t_R g4502 ( 
.A(n_10),
.Y(n_4502)
);

CKINVDCx20_ASAP7_75t_R g4503 ( 
.A(n_3721),
.Y(n_4503)
);

CKINVDCx5p33_ASAP7_75t_R g4504 ( 
.A(n_3858),
.Y(n_4504)
);

CKINVDCx5p33_ASAP7_75t_R g4505 ( 
.A(n_1381),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_343),
.Y(n_4506)
);

CKINVDCx5p33_ASAP7_75t_R g4507 ( 
.A(n_3922),
.Y(n_4507)
);

CKINVDCx5p33_ASAP7_75t_R g4508 ( 
.A(n_851),
.Y(n_4508)
);

INVx1_ASAP7_75t_L g4509 ( 
.A(n_3002),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_3574),
.Y(n_4510)
);

CKINVDCx20_ASAP7_75t_R g4511 ( 
.A(n_3147),
.Y(n_4511)
);

CKINVDCx5p33_ASAP7_75t_R g4512 ( 
.A(n_1309),
.Y(n_4512)
);

INVx1_ASAP7_75t_L g4513 ( 
.A(n_2846),
.Y(n_4513)
);

CKINVDCx5p33_ASAP7_75t_R g4514 ( 
.A(n_3257),
.Y(n_4514)
);

CKINVDCx5p33_ASAP7_75t_R g4515 ( 
.A(n_2311),
.Y(n_4515)
);

CKINVDCx5p33_ASAP7_75t_R g4516 ( 
.A(n_1381),
.Y(n_4516)
);

CKINVDCx5p33_ASAP7_75t_R g4517 ( 
.A(n_1645),
.Y(n_4517)
);

BUFx3_ASAP7_75t_L g4518 ( 
.A(n_1345),
.Y(n_4518)
);

CKINVDCx5p33_ASAP7_75t_R g4519 ( 
.A(n_3535),
.Y(n_4519)
);

CKINVDCx5p33_ASAP7_75t_R g4520 ( 
.A(n_2551),
.Y(n_4520)
);

INVx1_ASAP7_75t_L g4521 ( 
.A(n_2634),
.Y(n_4521)
);

BUFx8_ASAP7_75t_SL g4522 ( 
.A(n_3751),
.Y(n_4522)
);

CKINVDCx5p33_ASAP7_75t_R g4523 ( 
.A(n_4000),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_4035),
.Y(n_4524)
);

CKINVDCx5p33_ASAP7_75t_R g4525 ( 
.A(n_818),
.Y(n_4525)
);

CKINVDCx5p33_ASAP7_75t_R g4526 ( 
.A(n_2939),
.Y(n_4526)
);

CKINVDCx5p33_ASAP7_75t_R g4527 ( 
.A(n_174),
.Y(n_4527)
);

INVx1_ASAP7_75t_L g4528 ( 
.A(n_3733),
.Y(n_4528)
);

INVx1_ASAP7_75t_L g4529 ( 
.A(n_3947),
.Y(n_4529)
);

CKINVDCx5p33_ASAP7_75t_R g4530 ( 
.A(n_3763),
.Y(n_4530)
);

CKINVDCx5p33_ASAP7_75t_R g4531 ( 
.A(n_2944),
.Y(n_4531)
);

BUFx3_ASAP7_75t_L g4532 ( 
.A(n_1492),
.Y(n_4532)
);

CKINVDCx5p33_ASAP7_75t_R g4533 ( 
.A(n_3568),
.Y(n_4533)
);

INVx2_ASAP7_75t_L g4534 ( 
.A(n_917),
.Y(n_4534)
);

CKINVDCx5p33_ASAP7_75t_R g4535 ( 
.A(n_3743),
.Y(n_4535)
);

CKINVDCx5p33_ASAP7_75t_R g4536 ( 
.A(n_1584),
.Y(n_4536)
);

CKINVDCx5p33_ASAP7_75t_R g4537 ( 
.A(n_2847),
.Y(n_4537)
);

CKINVDCx5p33_ASAP7_75t_R g4538 ( 
.A(n_3955),
.Y(n_4538)
);

INVx1_ASAP7_75t_L g4539 ( 
.A(n_3921),
.Y(n_4539)
);

CKINVDCx20_ASAP7_75t_R g4540 ( 
.A(n_1262),
.Y(n_4540)
);

INVx2_ASAP7_75t_L g4541 ( 
.A(n_3809),
.Y(n_4541)
);

INVx1_ASAP7_75t_L g4542 ( 
.A(n_1525),
.Y(n_4542)
);

CKINVDCx5p33_ASAP7_75t_R g4543 ( 
.A(n_112),
.Y(n_4543)
);

INVx2_ASAP7_75t_L g4544 ( 
.A(n_3057),
.Y(n_4544)
);

CKINVDCx5p33_ASAP7_75t_R g4545 ( 
.A(n_3766),
.Y(n_4545)
);

CKINVDCx5p33_ASAP7_75t_R g4546 ( 
.A(n_202),
.Y(n_4546)
);

CKINVDCx5p33_ASAP7_75t_R g4547 ( 
.A(n_3141),
.Y(n_4547)
);

INVx2_ASAP7_75t_L g4548 ( 
.A(n_1313),
.Y(n_4548)
);

CKINVDCx5p33_ASAP7_75t_R g4549 ( 
.A(n_3064),
.Y(n_4549)
);

INVx2_ASAP7_75t_L g4550 ( 
.A(n_1276),
.Y(n_4550)
);

INVx1_ASAP7_75t_L g4551 ( 
.A(n_119),
.Y(n_4551)
);

BUFx6f_ASAP7_75t_L g4552 ( 
.A(n_2338),
.Y(n_4552)
);

INVxp67_ASAP7_75t_L g4553 ( 
.A(n_3268),
.Y(n_4553)
);

CKINVDCx20_ASAP7_75t_R g4554 ( 
.A(n_3859),
.Y(n_4554)
);

CKINVDCx5p33_ASAP7_75t_R g4555 ( 
.A(n_4072),
.Y(n_4555)
);

INVx1_ASAP7_75t_L g4556 ( 
.A(n_1986),
.Y(n_4556)
);

INVx1_ASAP7_75t_L g4557 ( 
.A(n_244),
.Y(n_4557)
);

CKINVDCx5p33_ASAP7_75t_R g4558 ( 
.A(n_3959),
.Y(n_4558)
);

CKINVDCx16_ASAP7_75t_R g4559 ( 
.A(n_1543),
.Y(n_4559)
);

BUFx10_ASAP7_75t_L g4560 ( 
.A(n_2429),
.Y(n_4560)
);

BUFx3_ASAP7_75t_L g4561 ( 
.A(n_103),
.Y(n_4561)
);

CKINVDCx5p33_ASAP7_75t_R g4562 ( 
.A(n_349),
.Y(n_4562)
);

CKINVDCx5p33_ASAP7_75t_R g4563 ( 
.A(n_1914),
.Y(n_4563)
);

INVx1_ASAP7_75t_L g4564 ( 
.A(n_2788),
.Y(n_4564)
);

CKINVDCx5p33_ASAP7_75t_R g4565 ( 
.A(n_3975),
.Y(n_4565)
);

INVx1_ASAP7_75t_L g4566 ( 
.A(n_3414),
.Y(n_4566)
);

CKINVDCx20_ASAP7_75t_R g4567 ( 
.A(n_1887),
.Y(n_4567)
);

CKINVDCx5p33_ASAP7_75t_R g4568 ( 
.A(n_1147),
.Y(n_4568)
);

CKINVDCx5p33_ASAP7_75t_R g4569 ( 
.A(n_3886),
.Y(n_4569)
);

INVx1_ASAP7_75t_SL g4570 ( 
.A(n_2248),
.Y(n_4570)
);

BUFx8_ASAP7_75t_SL g4571 ( 
.A(n_3493),
.Y(n_4571)
);

CKINVDCx5p33_ASAP7_75t_R g4572 ( 
.A(n_315),
.Y(n_4572)
);

INVx1_ASAP7_75t_L g4573 ( 
.A(n_1275),
.Y(n_4573)
);

INVx1_ASAP7_75t_L g4574 ( 
.A(n_3370),
.Y(n_4574)
);

INVx1_ASAP7_75t_L g4575 ( 
.A(n_529),
.Y(n_4575)
);

CKINVDCx5p33_ASAP7_75t_R g4576 ( 
.A(n_1379),
.Y(n_4576)
);

CKINVDCx5p33_ASAP7_75t_R g4577 ( 
.A(n_599),
.Y(n_4577)
);

HB1xp67_ASAP7_75t_L g4578 ( 
.A(n_1922),
.Y(n_4578)
);

CKINVDCx20_ASAP7_75t_R g4579 ( 
.A(n_451),
.Y(n_4579)
);

INVx2_ASAP7_75t_L g4580 ( 
.A(n_1919),
.Y(n_4580)
);

CKINVDCx20_ASAP7_75t_R g4581 ( 
.A(n_1836),
.Y(n_4581)
);

INVx1_ASAP7_75t_L g4582 ( 
.A(n_1151),
.Y(n_4582)
);

INVx1_ASAP7_75t_L g4583 ( 
.A(n_1144),
.Y(n_4583)
);

BUFx10_ASAP7_75t_L g4584 ( 
.A(n_2029),
.Y(n_4584)
);

CKINVDCx5p33_ASAP7_75t_R g4585 ( 
.A(n_2924),
.Y(n_4585)
);

INVx1_ASAP7_75t_L g4586 ( 
.A(n_3975),
.Y(n_4586)
);

CKINVDCx5p33_ASAP7_75t_R g4587 ( 
.A(n_1104),
.Y(n_4587)
);

HB1xp67_ASAP7_75t_SL g4588 ( 
.A(n_690),
.Y(n_4588)
);

CKINVDCx5p33_ASAP7_75t_R g4589 ( 
.A(n_1487),
.Y(n_4589)
);

CKINVDCx20_ASAP7_75t_R g4590 ( 
.A(n_1513),
.Y(n_4590)
);

CKINVDCx5p33_ASAP7_75t_R g4591 ( 
.A(n_1010),
.Y(n_4591)
);

CKINVDCx5p33_ASAP7_75t_R g4592 ( 
.A(n_2507),
.Y(n_4592)
);

BUFx10_ASAP7_75t_L g4593 ( 
.A(n_314),
.Y(n_4593)
);

CKINVDCx5p33_ASAP7_75t_R g4594 ( 
.A(n_650),
.Y(n_4594)
);

CKINVDCx5p33_ASAP7_75t_R g4595 ( 
.A(n_3310),
.Y(n_4595)
);

CKINVDCx5p33_ASAP7_75t_R g4596 ( 
.A(n_95),
.Y(n_4596)
);

INVx1_ASAP7_75t_L g4597 ( 
.A(n_2091),
.Y(n_4597)
);

INVx1_ASAP7_75t_L g4598 ( 
.A(n_3511),
.Y(n_4598)
);

INVx1_ASAP7_75t_L g4599 ( 
.A(n_3726),
.Y(n_4599)
);

CKINVDCx5p33_ASAP7_75t_R g4600 ( 
.A(n_2564),
.Y(n_4600)
);

CKINVDCx20_ASAP7_75t_R g4601 ( 
.A(n_3872),
.Y(n_4601)
);

CKINVDCx5p33_ASAP7_75t_R g4602 ( 
.A(n_1013),
.Y(n_4602)
);

INVx2_ASAP7_75t_L g4603 ( 
.A(n_1085),
.Y(n_4603)
);

CKINVDCx5p33_ASAP7_75t_R g4604 ( 
.A(n_1138),
.Y(n_4604)
);

BUFx10_ASAP7_75t_L g4605 ( 
.A(n_2300),
.Y(n_4605)
);

INVx1_ASAP7_75t_L g4606 ( 
.A(n_3188),
.Y(n_4606)
);

CKINVDCx5p33_ASAP7_75t_R g4607 ( 
.A(n_679),
.Y(n_4607)
);

CKINVDCx5p33_ASAP7_75t_R g4608 ( 
.A(n_306),
.Y(n_4608)
);

INVx1_ASAP7_75t_SL g4609 ( 
.A(n_3099),
.Y(n_4609)
);

CKINVDCx5p33_ASAP7_75t_R g4610 ( 
.A(n_1341),
.Y(n_4610)
);

BUFx5_ASAP7_75t_L g4611 ( 
.A(n_595),
.Y(n_4611)
);

CKINVDCx5p33_ASAP7_75t_R g4612 ( 
.A(n_3394),
.Y(n_4612)
);

CKINVDCx14_ASAP7_75t_R g4613 ( 
.A(n_3435),
.Y(n_4613)
);

CKINVDCx20_ASAP7_75t_R g4614 ( 
.A(n_2723),
.Y(n_4614)
);

CKINVDCx20_ASAP7_75t_R g4615 ( 
.A(n_369),
.Y(n_4615)
);

CKINVDCx5p33_ASAP7_75t_R g4616 ( 
.A(n_3750),
.Y(n_4616)
);

CKINVDCx20_ASAP7_75t_R g4617 ( 
.A(n_1958),
.Y(n_4617)
);

CKINVDCx5p33_ASAP7_75t_R g4618 ( 
.A(n_3764),
.Y(n_4618)
);

INVx1_ASAP7_75t_L g4619 ( 
.A(n_1212),
.Y(n_4619)
);

INVx1_ASAP7_75t_L g4620 ( 
.A(n_2254),
.Y(n_4620)
);

INVx1_ASAP7_75t_L g4621 ( 
.A(n_2733),
.Y(n_4621)
);

CKINVDCx5p33_ASAP7_75t_R g4622 ( 
.A(n_2577),
.Y(n_4622)
);

CKINVDCx20_ASAP7_75t_R g4623 ( 
.A(n_1223),
.Y(n_4623)
);

CKINVDCx5p33_ASAP7_75t_R g4624 ( 
.A(n_3957),
.Y(n_4624)
);

BUFx6f_ASAP7_75t_L g4625 ( 
.A(n_43),
.Y(n_4625)
);

INVx1_ASAP7_75t_L g4626 ( 
.A(n_1528),
.Y(n_4626)
);

CKINVDCx5p33_ASAP7_75t_R g4627 ( 
.A(n_3323),
.Y(n_4627)
);

CKINVDCx5p33_ASAP7_75t_R g4628 ( 
.A(n_3983),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_2252),
.Y(n_4629)
);

CKINVDCx5p33_ASAP7_75t_R g4630 ( 
.A(n_724),
.Y(n_4630)
);

INVx1_ASAP7_75t_L g4631 ( 
.A(n_3869),
.Y(n_4631)
);

BUFx3_ASAP7_75t_L g4632 ( 
.A(n_648),
.Y(n_4632)
);

INVx1_ASAP7_75t_L g4633 ( 
.A(n_1744),
.Y(n_4633)
);

CKINVDCx5p33_ASAP7_75t_R g4634 ( 
.A(n_1636),
.Y(n_4634)
);

CKINVDCx5p33_ASAP7_75t_R g4635 ( 
.A(n_3290),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_3028),
.Y(n_4636)
);

CKINVDCx5p33_ASAP7_75t_R g4637 ( 
.A(n_3721),
.Y(n_4637)
);

INVx1_ASAP7_75t_L g4638 ( 
.A(n_2174),
.Y(n_4638)
);

CKINVDCx5p33_ASAP7_75t_R g4639 ( 
.A(n_727),
.Y(n_4639)
);

INVx1_ASAP7_75t_L g4640 ( 
.A(n_3834),
.Y(n_4640)
);

CKINVDCx20_ASAP7_75t_R g4641 ( 
.A(n_2826),
.Y(n_4641)
);

CKINVDCx5p33_ASAP7_75t_R g4642 ( 
.A(n_3862),
.Y(n_4642)
);

INVx1_ASAP7_75t_L g4643 ( 
.A(n_53),
.Y(n_4643)
);

CKINVDCx5p33_ASAP7_75t_R g4644 ( 
.A(n_3108),
.Y(n_4644)
);

CKINVDCx5p33_ASAP7_75t_R g4645 ( 
.A(n_3703),
.Y(n_4645)
);

CKINVDCx5p33_ASAP7_75t_R g4646 ( 
.A(n_901),
.Y(n_4646)
);

CKINVDCx5p33_ASAP7_75t_R g4647 ( 
.A(n_2456),
.Y(n_4647)
);

CKINVDCx5p33_ASAP7_75t_R g4648 ( 
.A(n_1812),
.Y(n_4648)
);

CKINVDCx5p33_ASAP7_75t_R g4649 ( 
.A(n_3378),
.Y(n_4649)
);

BUFx10_ASAP7_75t_L g4650 ( 
.A(n_3280),
.Y(n_4650)
);

INVx1_ASAP7_75t_L g4651 ( 
.A(n_1970),
.Y(n_4651)
);

INVx1_ASAP7_75t_L g4652 ( 
.A(n_2167),
.Y(n_4652)
);

CKINVDCx5p33_ASAP7_75t_R g4653 ( 
.A(n_3896),
.Y(n_4653)
);

INVx2_ASAP7_75t_L g4654 ( 
.A(n_391),
.Y(n_4654)
);

CKINVDCx5p33_ASAP7_75t_R g4655 ( 
.A(n_1292),
.Y(n_4655)
);

CKINVDCx5p33_ASAP7_75t_R g4656 ( 
.A(n_2087),
.Y(n_4656)
);

INVx1_ASAP7_75t_L g4657 ( 
.A(n_3956),
.Y(n_4657)
);

CKINVDCx5p33_ASAP7_75t_R g4658 ( 
.A(n_3443),
.Y(n_4658)
);

CKINVDCx5p33_ASAP7_75t_R g4659 ( 
.A(n_3080),
.Y(n_4659)
);

CKINVDCx5p33_ASAP7_75t_R g4660 ( 
.A(n_1907),
.Y(n_4660)
);

CKINVDCx5p33_ASAP7_75t_R g4661 ( 
.A(n_3324),
.Y(n_4661)
);

CKINVDCx5p33_ASAP7_75t_R g4662 ( 
.A(n_2021),
.Y(n_4662)
);

INVx1_ASAP7_75t_L g4663 ( 
.A(n_3029),
.Y(n_4663)
);

INVx1_ASAP7_75t_L g4664 ( 
.A(n_3467),
.Y(n_4664)
);

INVx1_ASAP7_75t_L g4665 ( 
.A(n_2635),
.Y(n_4665)
);

BUFx6f_ASAP7_75t_L g4666 ( 
.A(n_1649),
.Y(n_4666)
);

BUFx2_ASAP7_75t_L g4667 ( 
.A(n_3341),
.Y(n_4667)
);

CKINVDCx5p33_ASAP7_75t_R g4668 ( 
.A(n_29),
.Y(n_4668)
);

INVx1_ASAP7_75t_L g4669 ( 
.A(n_3967),
.Y(n_4669)
);

INVx1_ASAP7_75t_L g4670 ( 
.A(n_3751),
.Y(n_4670)
);

BUFx6f_ASAP7_75t_L g4671 ( 
.A(n_3033),
.Y(n_4671)
);

INVx1_ASAP7_75t_L g4672 ( 
.A(n_2146),
.Y(n_4672)
);

CKINVDCx5p33_ASAP7_75t_R g4673 ( 
.A(n_2944),
.Y(n_4673)
);

INVx1_ASAP7_75t_SL g4674 ( 
.A(n_3962),
.Y(n_4674)
);

INVx1_ASAP7_75t_L g4675 ( 
.A(n_2325),
.Y(n_4675)
);

INVx1_ASAP7_75t_L g4676 ( 
.A(n_2378),
.Y(n_4676)
);

BUFx3_ASAP7_75t_L g4677 ( 
.A(n_1911),
.Y(n_4677)
);

INVx1_ASAP7_75t_L g4678 ( 
.A(n_3399),
.Y(n_4678)
);

CKINVDCx5p33_ASAP7_75t_R g4679 ( 
.A(n_721),
.Y(n_4679)
);

CKINVDCx5p33_ASAP7_75t_R g4680 ( 
.A(n_2972),
.Y(n_4680)
);

CKINVDCx5p33_ASAP7_75t_R g4681 ( 
.A(n_524),
.Y(n_4681)
);

CKINVDCx16_ASAP7_75t_R g4682 ( 
.A(n_1254),
.Y(n_4682)
);

CKINVDCx5p33_ASAP7_75t_R g4683 ( 
.A(n_88),
.Y(n_4683)
);

INVx1_ASAP7_75t_L g4684 ( 
.A(n_3996),
.Y(n_4684)
);

INVx1_ASAP7_75t_L g4685 ( 
.A(n_1239),
.Y(n_4685)
);

CKINVDCx5p33_ASAP7_75t_R g4686 ( 
.A(n_2480),
.Y(n_4686)
);

INVx1_ASAP7_75t_SL g4687 ( 
.A(n_2088),
.Y(n_4687)
);

INVx1_ASAP7_75t_L g4688 ( 
.A(n_2695),
.Y(n_4688)
);

INVx1_ASAP7_75t_L g4689 ( 
.A(n_3496),
.Y(n_4689)
);

CKINVDCx16_ASAP7_75t_R g4690 ( 
.A(n_1444),
.Y(n_4690)
);

CKINVDCx5p33_ASAP7_75t_R g4691 ( 
.A(n_2136),
.Y(n_4691)
);

BUFx2_ASAP7_75t_L g4692 ( 
.A(n_1359),
.Y(n_4692)
);

CKINVDCx5p33_ASAP7_75t_R g4693 ( 
.A(n_2984),
.Y(n_4693)
);

CKINVDCx5p33_ASAP7_75t_R g4694 ( 
.A(n_515),
.Y(n_4694)
);

CKINVDCx5p33_ASAP7_75t_R g4695 ( 
.A(n_572),
.Y(n_4695)
);

BUFx3_ASAP7_75t_L g4696 ( 
.A(n_1420),
.Y(n_4696)
);

INVx1_ASAP7_75t_L g4697 ( 
.A(n_3916),
.Y(n_4697)
);

INVx1_ASAP7_75t_L g4698 ( 
.A(n_3137),
.Y(n_4698)
);

INVxp33_ASAP7_75t_SL g4699 ( 
.A(n_2546),
.Y(n_4699)
);

INVx2_ASAP7_75t_SL g4700 ( 
.A(n_3925),
.Y(n_4700)
);

CKINVDCx5p33_ASAP7_75t_R g4701 ( 
.A(n_3119),
.Y(n_4701)
);

CKINVDCx5p33_ASAP7_75t_R g4702 ( 
.A(n_134),
.Y(n_4702)
);

INVx1_ASAP7_75t_L g4703 ( 
.A(n_1812),
.Y(n_4703)
);

INVx1_ASAP7_75t_L g4704 ( 
.A(n_4088),
.Y(n_4704)
);

INVx1_ASAP7_75t_SL g4705 ( 
.A(n_2062),
.Y(n_4705)
);

INVx1_ASAP7_75t_L g4706 ( 
.A(n_508),
.Y(n_4706)
);

CKINVDCx5p33_ASAP7_75t_R g4707 ( 
.A(n_3907),
.Y(n_4707)
);

INVx1_ASAP7_75t_L g4708 ( 
.A(n_3961),
.Y(n_4708)
);

CKINVDCx5p33_ASAP7_75t_R g4709 ( 
.A(n_1703),
.Y(n_4709)
);

HB1xp67_ASAP7_75t_L g4710 ( 
.A(n_221),
.Y(n_4710)
);

CKINVDCx5p33_ASAP7_75t_R g4711 ( 
.A(n_877),
.Y(n_4711)
);

CKINVDCx20_ASAP7_75t_R g4712 ( 
.A(n_1833),
.Y(n_4712)
);

CKINVDCx5p33_ASAP7_75t_R g4713 ( 
.A(n_3515),
.Y(n_4713)
);

BUFx10_ASAP7_75t_L g4714 ( 
.A(n_3912),
.Y(n_4714)
);

INVx1_ASAP7_75t_L g4715 ( 
.A(n_99),
.Y(n_4715)
);

CKINVDCx5p33_ASAP7_75t_R g4716 ( 
.A(n_2507),
.Y(n_4716)
);

INVx1_ASAP7_75t_L g4717 ( 
.A(n_3777),
.Y(n_4717)
);

CKINVDCx5p33_ASAP7_75t_R g4718 ( 
.A(n_3931),
.Y(n_4718)
);

CKINVDCx5p33_ASAP7_75t_R g4719 ( 
.A(n_958),
.Y(n_4719)
);

CKINVDCx5p33_ASAP7_75t_R g4720 ( 
.A(n_1041),
.Y(n_4720)
);

CKINVDCx5p33_ASAP7_75t_R g4721 ( 
.A(n_3816),
.Y(n_4721)
);

CKINVDCx5p33_ASAP7_75t_R g4722 ( 
.A(n_3979),
.Y(n_4722)
);

BUFx3_ASAP7_75t_L g4723 ( 
.A(n_1031),
.Y(n_4723)
);

INVx2_ASAP7_75t_L g4724 ( 
.A(n_1663),
.Y(n_4724)
);

CKINVDCx5p33_ASAP7_75t_R g4725 ( 
.A(n_749),
.Y(n_4725)
);

CKINVDCx5p33_ASAP7_75t_R g4726 ( 
.A(n_29),
.Y(n_4726)
);

CKINVDCx5p33_ASAP7_75t_R g4727 ( 
.A(n_1853),
.Y(n_4727)
);

CKINVDCx5p33_ASAP7_75t_R g4728 ( 
.A(n_451),
.Y(n_4728)
);

CKINVDCx20_ASAP7_75t_R g4729 ( 
.A(n_2397),
.Y(n_4729)
);

INVx1_ASAP7_75t_L g4730 ( 
.A(n_2854),
.Y(n_4730)
);

CKINVDCx5p33_ASAP7_75t_R g4731 ( 
.A(n_1546),
.Y(n_4731)
);

CKINVDCx5p33_ASAP7_75t_R g4732 ( 
.A(n_248),
.Y(n_4732)
);

CKINVDCx5p33_ASAP7_75t_R g4733 ( 
.A(n_3878),
.Y(n_4733)
);

CKINVDCx20_ASAP7_75t_R g4734 ( 
.A(n_3913),
.Y(n_4734)
);

CKINVDCx20_ASAP7_75t_R g4735 ( 
.A(n_2592),
.Y(n_4735)
);

INVx1_ASAP7_75t_SL g4736 ( 
.A(n_980),
.Y(n_4736)
);

INVx1_ASAP7_75t_L g4737 ( 
.A(n_3851),
.Y(n_4737)
);

INVx2_ASAP7_75t_L g4738 ( 
.A(n_3988),
.Y(n_4738)
);

CKINVDCx5p33_ASAP7_75t_R g4739 ( 
.A(n_3860),
.Y(n_4739)
);

INVx1_ASAP7_75t_L g4740 ( 
.A(n_498),
.Y(n_4740)
);

INVx1_ASAP7_75t_L g4741 ( 
.A(n_2669),
.Y(n_4741)
);

INVx2_ASAP7_75t_L g4742 ( 
.A(n_3944),
.Y(n_4742)
);

HB1xp67_ASAP7_75t_L g4743 ( 
.A(n_2657),
.Y(n_4743)
);

INVx2_ASAP7_75t_SL g4744 ( 
.A(n_3855),
.Y(n_4744)
);

INVx1_ASAP7_75t_L g4745 ( 
.A(n_2015),
.Y(n_4745)
);

BUFx6f_ASAP7_75t_L g4746 ( 
.A(n_3604),
.Y(n_4746)
);

INVx1_ASAP7_75t_L g4747 ( 
.A(n_743),
.Y(n_4747)
);

BUFx2_ASAP7_75t_L g4748 ( 
.A(n_3265),
.Y(n_4748)
);

INVx1_ASAP7_75t_L g4749 ( 
.A(n_4044),
.Y(n_4749)
);

INVx2_ASAP7_75t_L g4750 ( 
.A(n_3353),
.Y(n_4750)
);

INVx1_ASAP7_75t_SL g4751 ( 
.A(n_3529),
.Y(n_4751)
);

BUFx3_ASAP7_75t_L g4752 ( 
.A(n_362),
.Y(n_4752)
);

INVx2_ASAP7_75t_L g4753 ( 
.A(n_3214),
.Y(n_4753)
);

BUFx3_ASAP7_75t_L g4754 ( 
.A(n_72),
.Y(n_4754)
);

CKINVDCx5p33_ASAP7_75t_R g4755 ( 
.A(n_2351),
.Y(n_4755)
);

CKINVDCx5p33_ASAP7_75t_R g4756 ( 
.A(n_2527),
.Y(n_4756)
);

INVx2_ASAP7_75t_SL g4757 ( 
.A(n_3198),
.Y(n_4757)
);

CKINVDCx5p33_ASAP7_75t_R g4758 ( 
.A(n_588),
.Y(n_4758)
);

CKINVDCx5p33_ASAP7_75t_R g4759 ( 
.A(n_2364),
.Y(n_4759)
);

CKINVDCx5p33_ASAP7_75t_R g4760 ( 
.A(n_2591),
.Y(n_4760)
);

CKINVDCx5p33_ASAP7_75t_R g4761 ( 
.A(n_1920),
.Y(n_4761)
);

INVx1_ASAP7_75t_L g4762 ( 
.A(n_4011),
.Y(n_4762)
);

INVx1_ASAP7_75t_L g4763 ( 
.A(n_4038),
.Y(n_4763)
);

CKINVDCx5p33_ASAP7_75t_R g4764 ( 
.A(n_2761),
.Y(n_4764)
);

INVx1_ASAP7_75t_L g4765 ( 
.A(n_3180),
.Y(n_4765)
);

INVx1_ASAP7_75t_L g4766 ( 
.A(n_2123),
.Y(n_4766)
);

INVx1_ASAP7_75t_L g4767 ( 
.A(n_3507),
.Y(n_4767)
);

CKINVDCx5p33_ASAP7_75t_R g4768 ( 
.A(n_3853),
.Y(n_4768)
);

CKINVDCx5p33_ASAP7_75t_R g4769 ( 
.A(n_1923),
.Y(n_4769)
);

CKINVDCx5p33_ASAP7_75t_R g4770 ( 
.A(n_4007),
.Y(n_4770)
);

INVxp67_ASAP7_75t_L g4771 ( 
.A(n_2683),
.Y(n_4771)
);

CKINVDCx5p33_ASAP7_75t_R g4772 ( 
.A(n_799),
.Y(n_4772)
);

INVx1_ASAP7_75t_L g4773 ( 
.A(n_67),
.Y(n_4773)
);

CKINVDCx5p33_ASAP7_75t_R g4774 ( 
.A(n_3868),
.Y(n_4774)
);

INVx1_ASAP7_75t_L g4775 ( 
.A(n_1520),
.Y(n_4775)
);

INVx1_ASAP7_75t_L g4776 ( 
.A(n_1075),
.Y(n_4776)
);

INVx1_ASAP7_75t_L g4777 ( 
.A(n_2783),
.Y(n_4777)
);

INVxp67_ASAP7_75t_L g4778 ( 
.A(n_3025),
.Y(n_4778)
);

CKINVDCx5p33_ASAP7_75t_R g4779 ( 
.A(n_1535),
.Y(n_4779)
);

BUFx10_ASAP7_75t_L g4780 ( 
.A(n_1348),
.Y(n_4780)
);

INVx1_ASAP7_75t_SL g4781 ( 
.A(n_4043),
.Y(n_4781)
);

INVx1_ASAP7_75t_L g4782 ( 
.A(n_1094),
.Y(n_4782)
);

CKINVDCx5p33_ASAP7_75t_R g4783 ( 
.A(n_153),
.Y(n_4783)
);

CKINVDCx5p33_ASAP7_75t_R g4784 ( 
.A(n_3539),
.Y(n_4784)
);

INVx1_ASAP7_75t_L g4785 ( 
.A(n_3527),
.Y(n_4785)
);

INVx1_ASAP7_75t_L g4786 ( 
.A(n_4091),
.Y(n_4786)
);

INVx1_ASAP7_75t_L g4787 ( 
.A(n_700),
.Y(n_4787)
);

INVx2_ASAP7_75t_SL g4788 ( 
.A(n_3110),
.Y(n_4788)
);

CKINVDCx20_ASAP7_75t_R g4789 ( 
.A(n_3793),
.Y(n_4789)
);

CKINVDCx5p33_ASAP7_75t_R g4790 ( 
.A(n_222),
.Y(n_4790)
);

BUFx3_ASAP7_75t_L g4791 ( 
.A(n_1301),
.Y(n_4791)
);

BUFx6f_ASAP7_75t_L g4792 ( 
.A(n_1323),
.Y(n_4792)
);

CKINVDCx20_ASAP7_75t_R g4793 ( 
.A(n_2025),
.Y(n_4793)
);

CKINVDCx5p33_ASAP7_75t_R g4794 ( 
.A(n_3812),
.Y(n_4794)
);

INVx2_ASAP7_75t_SL g4795 ( 
.A(n_3877),
.Y(n_4795)
);

INVx2_ASAP7_75t_L g4796 ( 
.A(n_1132),
.Y(n_4796)
);

INVx1_ASAP7_75t_L g4797 ( 
.A(n_1742),
.Y(n_4797)
);

CKINVDCx16_ASAP7_75t_R g4798 ( 
.A(n_2253),
.Y(n_4798)
);

BUFx6f_ASAP7_75t_L g4799 ( 
.A(n_1166),
.Y(n_4799)
);

CKINVDCx5p33_ASAP7_75t_R g4800 ( 
.A(n_1685),
.Y(n_4800)
);

CKINVDCx5p33_ASAP7_75t_R g4801 ( 
.A(n_3974),
.Y(n_4801)
);

INVx2_ASAP7_75t_L g4802 ( 
.A(n_3980),
.Y(n_4802)
);

CKINVDCx5p33_ASAP7_75t_R g4803 ( 
.A(n_2465),
.Y(n_4803)
);

CKINVDCx5p33_ASAP7_75t_R g4804 ( 
.A(n_1690),
.Y(n_4804)
);

INVx1_ASAP7_75t_L g4805 ( 
.A(n_496),
.Y(n_4805)
);

BUFx6f_ASAP7_75t_L g4806 ( 
.A(n_3912),
.Y(n_4806)
);

CKINVDCx5p33_ASAP7_75t_R g4807 ( 
.A(n_1921),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4018),
.Y(n_4808)
);

CKINVDCx20_ASAP7_75t_R g4809 ( 
.A(n_1377),
.Y(n_4809)
);

CKINVDCx5p33_ASAP7_75t_R g4810 ( 
.A(n_3250),
.Y(n_4810)
);

CKINVDCx5p33_ASAP7_75t_R g4811 ( 
.A(n_3631),
.Y(n_4811)
);

CKINVDCx20_ASAP7_75t_R g4812 ( 
.A(n_1819),
.Y(n_4812)
);

INVx2_ASAP7_75t_L g4813 ( 
.A(n_3917),
.Y(n_4813)
);

CKINVDCx20_ASAP7_75t_R g4814 ( 
.A(n_185),
.Y(n_4814)
);

BUFx3_ASAP7_75t_L g4815 ( 
.A(n_1516),
.Y(n_4815)
);

CKINVDCx5p33_ASAP7_75t_R g4816 ( 
.A(n_2283),
.Y(n_4816)
);

CKINVDCx5p33_ASAP7_75t_R g4817 ( 
.A(n_951),
.Y(n_4817)
);

BUFx3_ASAP7_75t_L g4818 ( 
.A(n_3881),
.Y(n_4818)
);

CKINVDCx20_ASAP7_75t_R g4819 ( 
.A(n_1497),
.Y(n_4819)
);

CKINVDCx5p33_ASAP7_75t_R g4820 ( 
.A(n_1815),
.Y(n_4820)
);

INVx1_ASAP7_75t_L g4821 ( 
.A(n_3105),
.Y(n_4821)
);

INVxp67_ASAP7_75t_L g4822 ( 
.A(n_2393),
.Y(n_4822)
);

CKINVDCx5p33_ASAP7_75t_R g4823 ( 
.A(n_3997),
.Y(n_4823)
);

CKINVDCx5p33_ASAP7_75t_R g4824 ( 
.A(n_2170),
.Y(n_4824)
);

CKINVDCx5p33_ASAP7_75t_R g4825 ( 
.A(n_419),
.Y(n_4825)
);

CKINVDCx5p33_ASAP7_75t_R g4826 ( 
.A(n_3500),
.Y(n_4826)
);

CKINVDCx5p33_ASAP7_75t_R g4827 ( 
.A(n_2132),
.Y(n_4827)
);

CKINVDCx20_ASAP7_75t_R g4828 ( 
.A(n_985),
.Y(n_4828)
);

BUFx3_ASAP7_75t_L g4829 ( 
.A(n_805),
.Y(n_4829)
);

CKINVDCx5p33_ASAP7_75t_R g4830 ( 
.A(n_3911),
.Y(n_4830)
);

INVx2_ASAP7_75t_L g4831 ( 
.A(n_2982),
.Y(n_4831)
);

CKINVDCx5p33_ASAP7_75t_R g4832 ( 
.A(n_2235),
.Y(n_4832)
);

CKINVDCx16_ASAP7_75t_R g4833 ( 
.A(n_4006),
.Y(n_4833)
);

CKINVDCx5p33_ASAP7_75t_R g4834 ( 
.A(n_2626),
.Y(n_4834)
);

CKINVDCx5p33_ASAP7_75t_R g4835 ( 
.A(n_3593),
.Y(n_4835)
);

BUFx5_ASAP7_75t_L g4836 ( 
.A(n_3880),
.Y(n_4836)
);

INVx1_ASAP7_75t_L g4837 ( 
.A(n_1397),
.Y(n_4837)
);

CKINVDCx5p33_ASAP7_75t_R g4838 ( 
.A(n_3745),
.Y(n_4838)
);

INVx2_ASAP7_75t_SL g4839 ( 
.A(n_3538),
.Y(n_4839)
);

INVx2_ASAP7_75t_L g4840 ( 
.A(n_387),
.Y(n_4840)
);

INVx1_ASAP7_75t_L g4841 ( 
.A(n_2456),
.Y(n_4841)
);

INVx1_ASAP7_75t_L g4842 ( 
.A(n_3471),
.Y(n_4842)
);

INVx1_ASAP7_75t_SL g4843 ( 
.A(n_2543),
.Y(n_4843)
);

CKINVDCx5p33_ASAP7_75t_R g4844 ( 
.A(n_2825),
.Y(n_4844)
);

INVx1_ASAP7_75t_L g4845 ( 
.A(n_3887),
.Y(n_4845)
);

INVx1_ASAP7_75t_SL g4846 ( 
.A(n_3667),
.Y(n_4846)
);

CKINVDCx5p33_ASAP7_75t_R g4847 ( 
.A(n_272),
.Y(n_4847)
);

CKINVDCx20_ASAP7_75t_R g4848 ( 
.A(n_1836),
.Y(n_4848)
);

INVx1_ASAP7_75t_L g4849 ( 
.A(n_151),
.Y(n_4849)
);

CKINVDCx20_ASAP7_75t_R g4850 ( 
.A(n_1425),
.Y(n_4850)
);

CKINVDCx5p33_ASAP7_75t_R g4851 ( 
.A(n_4017),
.Y(n_4851)
);

CKINVDCx5p33_ASAP7_75t_R g4852 ( 
.A(n_3070),
.Y(n_4852)
);

INVx2_ASAP7_75t_SL g4853 ( 
.A(n_2929),
.Y(n_4853)
);

BUFx6f_ASAP7_75t_L g4854 ( 
.A(n_4045),
.Y(n_4854)
);

CKINVDCx5p33_ASAP7_75t_R g4855 ( 
.A(n_3603),
.Y(n_4855)
);

CKINVDCx16_ASAP7_75t_R g4856 ( 
.A(n_3908),
.Y(n_4856)
);

CKINVDCx5p33_ASAP7_75t_R g4857 ( 
.A(n_3994),
.Y(n_4857)
);

CKINVDCx5p33_ASAP7_75t_R g4858 ( 
.A(n_1495),
.Y(n_4858)
);

CKINVDCx5p33_ASAP7_75t_R g4859 ( 
.A(n_1571),
.Y(n_4859)
);

CKINVDCx5p33_ASAP7_75t_R g4860 ( 
.A(n_3427),
.Y(n_4860)
);

CKINVDCx5p33_ASAP7_75t_R g4861 ( 
.A(n_3075),
.Y(n_4861)
);

BUFx3_ASAP7_75t_L g4862 ( 
.A(n_652),
.Y(n_4862)
);

CKINVDCx5p33_ASAP7_75t_R g4863 ( 
.A(n_2093),
.Y(n_4863)
);

CKINVDCx5p33_ASAP7_75t_R g4864 ( 
.A(n_1554),
.Y(n_4864)
);

INVx2_ASAP7_75t_L g4865 ( 
.A(n_91),
.Y(n_4865)
);

BUFx3_ASAP7_75t_L g4866 ( 
.A(n_3011),
.Y(n_4866)
);

INVx1_ASAP7_75t_L g4867 ( 
.A(n_696),
.Y(n_4867)
);

INVx1_ASAP7_75t_L g4868 ( 
.A(n_838),
.Y(n_4868)
);

CKINVDCx5p33_ASAP7_75t_R g4869 ( 
.A(n_2663),
.Y(n_4869)
);

CKINVDCx5p33_ASAP7_75t_R g4870 ( 
.A(n_4053),
.Y(n_4870)
);

BUFx3_ASAP7_75t_L g4871 ( 
.A(n_4001),
.Y(n_4871)
);

CKINVDCx5p33_ASAP7_75t_R g4872 ( 
.A(n_1187),
.Y(n_4872)
);

CKINVDCx20_ASAP7_75t_R g4873 ( 
.A(n_3792),
.Y(n_4873)
);

INVx1_ASAP7_75t_L g4874 ( 
.A(n_1930),
.Y(n_4874)
);

CKINVDCx5p33_ASAP7_75t_R g4875 ( 
.A(n_3985),
.Y(n_4875)
);

INVx1_ASAP7_75t_L g4876 ( 
.A(n_3291),
.Y(n_4876)
);

CKINVDCx5p33_ASAP7_75t_R g4877 ( 
.A(n_258),
.Y(n_4877)
);

BUFx6f_ASAP7_75t_L g4878 ( 
.A(n_3268),
.Y(n_4878)
);

INVx1_ASAP7_75t_L g4879 ( 
.A(n_150),
.Y(n_4879)
);

CKINVDCx5p33_ASAP7_75t_R g4880 ( 
.A(n_3954),
.Y(n_4880)
);

INVx2_ASAP7_75t_L g4881 ( 
.A(n_3196),
.Y(n_4881)
);

CKINVDCx5p33_ASAP7_75t_R g4882 ( 
.A(n_3897),
.Y(n_4882)
);

CKINVDCx5p33_ASAP7_75t_R g4883 ( 
.A(n_265),
.Y(n_4883)
);

CKINVDCx5p33_ASAP7_75t_R g4884 ( 
.A(n_2981),
.Y(n_4884)
);

CKINVDCx5p33_ASAP7_75t_R g4885 ( 
.A(n_1668),
.Y(n_4885)
);

CKINVDCx5p33_ASAP7_75t_R g4886 ( 
.A(n_353),
.Y(n_4886)
);

CKINVDCx5p33_ASAP7_75t_R g4887 ( 
.A(n_2389),
.Y(n_4887)
);

BUFx3_ASAP7_75t_L g4888 ( 
.A(n_856),
.Y(n_4888)
);

CKINVDCx5p33_ASAP7_75t_R g4889 ( 
.A(n_2649),
.Y(n_4889)
);

CKINVDCx5p33_ASAP7_75t_R g4890 ( 
.A(n_932),
.Y(n_4890)
);

BUFx5_ASAP7_75t_L g4891 ( 
.A(n_2445),
.Y(n_4891)
);

CKINVDCx16_ASAP7_75t_R g4892 ( 
.A(n_4042),
.Y(n_4892)
);

CKINVDCx5p33_ASAP7_75t_R g4893 ( 
.A(n_3789),
.Y(n_4893)
);

BUFx6f_ASAP7_75t_L g4894 ( 
.A(n_1694),
.Y(n_4894)
);

BUFx3_ASAP7_75t_L g4895 ( 
.A(n_4071),
.Y(n_4895)
);

CKINVDCx5p33_ASAP7_75t_R g4896 ( 
.A(n_4022),
.Y(n_4896)
);

CKINVDCx5p33_ASAP7_75t_R g4897 ( 
.A(n_678),
.Y(n_4897)
);

CKINVDCx5p33_ASAP7_75t_R g4898 ( 
.A(n_2340),
.Y(n_4898)
);

CKINVDCx5p33_ASAP7_75t_R g4899 ( 
.A(n_4021),
.Y(n_4899)
);

CKINVDCx5p33_ASAP7_75t_R g4900 ( 
.A(n_946),
.Y(n_4900)
);

CKINVDCx5p33_ASAP7_75t_R g4901 ( 
.A(n_3933),
.Y(n_4901)
);

CKINVDCx5p33_ASAP7_75t_R g4902 ( 
.A(n_2684),
.Y(n_4902)
);

CKINVDCx5p33_ASAP7_75t_R g4903 ( 
.A(n_1657),
.Y(n_4903)
);

BUFx3_ASAP7_75t_L g4904 ( 
.A(n_354),
.Y(n_4904)
);

CKINVDCx5p33_ASAP7_75t_R g4905 ( 
.A(n_3945),
.Y(n_4905)
);

CKINVDCx20_ASAP7_75t_R g4906 ( 
.A(n_2200),
.Y(n_4906)
);

INVx1_ASAP7_75t_L g4907 ( 
.A(n_3867),
.Y(n_4907)
);

HB1xp67_ASAP7_75t_L g4908 ( 
.A(n_1913),
.Y(n_4908)
);

INVx1_ASAP7_75t_L g4909 ( 
.A(n_599),
.Y(n_4909)
);

INVx1_ASAP7_75t_L g4910 ( 
.A(n_200),
.Y(n_4910)
);

CKINVDCx5p33_ASAP7_75t_R g4911 ( 
.A(n_118),
.Y(n_4911)
);

CKINVDCx5p33_ASAP7_75t_R g4912 ( 
.A(n_1203),
.Y(n_4912)
);

INVx1_ASAP7_75t_L g4913 ( 
.A(n_2691),
.Y(n_4913)
);

INVx1_ASAP7_75t_L g4914 ( 
.A(n_970),
.Y(n_4914)
);

CKINVDCx5p33_ASAP7_75t_R g4915 ( 
.A(n_3981),
.Y(n_4915)
);

CKINVDCx5p33_ASAP7_75t_R g4916 ( 
.A(n_2881),
.Y(n_4916)
);

CKINVDCx20_ASAP7_75t_R g4917 ( 
.A(n_245),
.Y(n_4917)
);

CKINVDCx5p33_ASAP7_75t_R g4918 ( 
.A(n_846),
.Y(n_4918)
);

CKINVDCx5p33_ASAP7_75t_R g4919 ( 
.A(n_2374),
.Y(n_4919)
);

CKINVDCx5p33_ASAP7_75t_R g4920 ( 
.A(n_3982),
.Y(n_4920)
);

CKINVDCx5p33_ASAP7_75t_R g4921 ( 
.A(n_1774),
.Y(n_4921)
);

BUFx5_ASAP7_75t_L g4922 ( 
.A(n_2282),
.Y(n_4922)
);

CKINVDCx5p33_ASAP7_75t_R g4923 ( 
.A(n_3194),
.Y(n_4923)
);

INVx2_ASAP7_75t_L g4924 ( 
.A(n_766),
.Y(n_4924)
);

INVx2_ASAP7_75t_SL g4925 ( 
.A(n_3923),
.Y(n_4925)
);

CKINVDCx5p33_ASAP7_75t_R g4926 ( 
.A(n_3979),
.Y(n_4926)
);

CKINVDCx5p33_ASAP7_75t_R g4927 ( 
.A(n_3244),
.Y(n_4927)
);

INVx1_ASAP7_75t_L g4928 ( 
.A(n_3826),
.Y(n_4928)
);

INVx2_ASAP7_75t_SL g4929 ( 
.A(n_686),
.Y(n_4929)
);

CKINVDCx5p33_ASAP7_75t_R g4930 ( 
.A(n_873),
.Y(n_4930)
);

INVxp67_ASAP7_75t_L g4931 ( 
.A(n_3905),
.Y(n_4931)
);

CKINVDCx16_ASAP7_75t_R g4932 ( 
.A(n_3282),
.Y(n_4932)
);

INVx2_ASAP7_75t_L g4933 ( 
.A(n_2415),
.Y(n_4933)
);

CKINVDCx20_ASAP7_75t_R g4934 ( 
.A(n_2011),
.Y(n_4934)
);

CKINVDCx5p33_ASAP7_75t_R g4935 ( 
.A(n_2955),
.Y(n_4935)
);

INVx1_ASAP7_75t_L g4936 ( 
.A(n_3903),
.Y(n_4936)
);

INVx1_ASAP7_75t_L g4937 ( 
.A(n_3604),
.Y(n_4937)
);

CKINVDCx5p33_ASAP7_75t_R g4938 ( 
.A(n_2957),
.Y(n_4938)
);

CKINVDCx5p33_ASAP7_75t_R g4939 ( 
.A(n_3908),
.Y(n_4939)
);

CKINVDCx5p33_ASAP7_75t_R g4940 ( 
.A(n_3430),
.Y(n_4940)
);

BUFx10_ASAP7_75t_L g4941 ( 
.A(n_1673),
.Y(n_4941)
);

BUFx6f_ASAP7_75t_L g4942 ( 
.A(n_90),
.Y(n_4942)
);

INVx1_ASAP7_75t_L g4943 ( 
.A(n_27),
.Y(n_4943)
);

CKINVDCx5p33_ASAP7_75t_R g4944 ( 
.A(n_794),
.Y(n_4944)
);

CKINVDCx5p33_ASAP7_75t_R g4945 ( 
.A(n_1307),
.Y(n_4945)
);

CKINVDCx5p33_ASAP7_75t_R g4946 ( 
.A(n_1656),
.Y(n_4946)
);

CKINVDCx5p33_ASAP7_75t_R g4947 ( 
.A(n_3900),
.Y(n_4947)
);

INVx1_ASAP7_75t_L g4948 ( 
.A(n_977),
.Y(n_4948)
);

INVx2_ASAP7_75t_L g4949 ( 
.A(n_1901),
.Y(n_4949)
);

INVx1_ASAP7_75t_L g4950 ( 
.A(n_97),
.Y(n_4950)
);

CKINVDCx5p33_ASAP7_75t_R g4951 ( 
.A(n_1341),
.Y(n_4951)
);

INVx1_ASAP7_75t_L g4952 ( 
.A(n_3685),
.Y(n_4952)
);

CKINVDCx5p33_ASAP7_75t_R g4953 ( 
.A(n_3970),
.Y(n_4953)
);

CKINVDCx5p33_ASAP7_75t_R g4954 ( 
.A(n_4036),
.Y(n_4954)
);

CKINVDCx5p33_ASAP7_75t_R g4955 ( 
.A(n_29),
.Y(n_4955)
);

CKINVDCx5p33_ASAP7_75t_R g4956 ( 
.A(n_757),
.Y(n_4956)
);

CKINVDCx20_ASAP7_75t_R g4957 ( 
.A(n_3480),
.Y(n_4957)
);

CKINVDCx5p33_ASAP7_75t_R g4958 ( 
.A(n_3216),
.Y(n_4958)
);

INVxp67_ASAP7_75t_L g4959 ( 
.A(n_596),
.Y(n_4959)
);

CKINVDCx14_ASAP7_75t_R g4960 ( 
.A(n_1363),
.Y(n_4960)
);

INVx1_ASAP7_75t_L g4961 ( 
.A(n_3990),
.Y(n_4961)
);

INVx1_ASAP7_75t_L g4962 ( 
.A(n_1116),
.Y(n_4962)
);

CKINVDCx5p33_ASAP7_75t_R g4963 ( 
.A(n_3873),
.Y(n_4963)
);

CKINVDCx5p33_ASAP7_75t_R g4964 ( 
.A(n_590),
.Y(n_4964)
);

CKINVDCx5p33_ASAP7_75t_R g4965 ( 
.A(n_803),
.Y(n_4965)
);

INVx1_ASAP7_75t_L g4966 ( 
.A(n_2186),
.Y(n_4966)
);

INVx1_ASAP7_75t_SL g4967 ( 
.A(n_3729),
.Y(n_4967)
);

CKINVDCx5p33_ASAP7_75t_R g4968 ( 
.A(n_3007),
.Y(n_4968)
);

CKINVDCx20_ASAP7_75t_R g4969 ( 
.A(n_1412),
.Y(n_4969)
);

CKINVDCx5p33_ASAP7_75t_R g4970 ( 
.A(n_4018),
.Y(n_4970)
);

CKINVDCx5p33_ASAP7_75t_R g4971 ( 
.A(n_3837),
.Y(n_4971)
);

INVx1_ASAP7_75t_SL g4972 ( 
.A(n_2020),
.Y(n_4972)
);

CKINVDCx5p33_ASAP7_75t_R g4973 ( 
.A(n_345),
.Y(n_4973)
);

BUFx10_ASAP7_75t_L g4974 ( 
.A(n_177),
.Y(n_4974)
);

CKINVDCx20_ASAP7_75t_R g4975 ( 
.A(n_3989),
.Y(n_4975)
);

CKINVDCx16_ASAP7_75t_R g4976 ( 
.A(n_2665),
.Y(n_4976)
);

CKINVDCx5p33_ASAP7_75t_R g4977 ( 
.A(n_3218),
.Y(n_4977)
);

CKINVDCx5p33_ASAP7_75t_R g4978 ( 
.A(n_3546),
.Y(n_4978)
);

INVx1_ASAP7_75t_L g4979 ( 
.A(n_3852),
.Y(n_4979)
);

CKINVDCx5p33_ASAP7_75t_R g4980 ( 
.A(n_2051),
.Y(n_4980)
);

CKINVDCx20_ASAP7_75t_R g4981 ( 
.A(n_371),
.Y(n_4981)
);

INVx1_ASAP7_75t_L g4982 ( 
.A(n_3960),
.Y(n_4982)
);

INVx1_ASAP7_75t_L g4983 ( 
.A(n_3086),
.Y(n_4983)
);

INVx1_ASAP7_75t_L g4984 ( 
.A(n_3690),
.Y(n_4984)
);

INVx1_ASAP7_75t_L g4985 ( 
.A(n_3291),
.Y(n_4985)
);

CKINVDCx5p33_ASAP7_75t_R g4986 ( 
.A(n_834),
.Y(n_4986)
);

INVx1_ASAP7_75t_L g4987 ( 
.A(n_1227),
.Y(n_4987)
);

CKINVDCx5p33_ASAP7_75t_R g4988 ( 
.A(n_2068),
.Y(n_4988)
);

INVx1_ASAP7_75t_L g4989 ( 
.A(n_40),
.Y(n_4989)
);

INVx1_ASAP7_75t_L g4990 ( 
.A(n_2934),
.Y(n_4990)
);

CKINVDCx5p33_ASAP7_75t_R g4991 ( 
.A(n_3045),
.Y(n_4991)
);

INVx1_ASAP7_75t_L g4992 ( 
.A(n_3550),
.Y(n_4992)
);

BUFx3_ASAP7_75t_L g4993 ( 
.A(n_9),
.Y(n_4993)
);

BUFx10_ASAP7_75t_L g4994 ( 
.A(n_3940),
.Y(n_4994)
);

CKINVDCx5p33_ASAP7_75t_R g4995 ( 
.A(n_69),
.Y(n_4995)
);

INVx1_ASAP7_75t_L g4996 ( 
.A(n_3977),
.Y(n_4996)
);

CKINVDCx5p33_ASAP7_75t_R g4997 ( 
.A(n_200),
.Y(n_4997)
);

INVx1_ASAP7_75t_L g4998 ( 
.A(n_3888),
.Y(n_4998)
);

BUFx10_ASAP7_75t_L g4999 ( 
.A(n_3638),
.Y(n_4999)
);

CKINVDCx5p33_ASAP7_75t_R g5000 ( 
.A(n_4078),
.Y(n_5000)
);

INVx1_ASAP7_75t_SL g5001 ( 
.A(n_1601),
.Y(n_5001)
);

CKINVDCx5p33_ASAP7_75t_R g5002 ( 
.A(n_3762),
.Y(n_5002)
);

CKINVDCx5p33_ASAP7_75t_R g5003 ( 
.A(n_3188),
.Y(n_5003)
);

INVx1_ASAP7_75t_L g5004 ( 
.A(n_3909),
.Y(n_5004)
);

INVx1_ASAP7_75t_SL g5005 ( 
.A(n_4080),
.Y(n_5005)
);

CKINVDCx5p33_ASAP7_75t_R g5006 ( 
.A(n_3964),
.Y(n_5006)
);

CKINVDCx5p33_ASAP7_75t_R g5007 ( 
.A(n_470),
.Y(n_5007)
);

CKINVDCx5p33_ASAP7_75t_R g5008 ( 
.A(n_3941),
.Y(n_5008)
);

CKINVDCx5p33_ASAP7_75t_R g5009 ( 
.A(n_3269),
.Y(n_5009)
);

CKINVDCx14_ASAP7_75t_R g5010 ( 
.A(n_3352),
.Y(n_5010)
);

CKINVDCx5p33_ASAP7_75t_R g5011 ( 
.A(n_1100),
.Y(n_5011)
);

BUFx10_ASAP7_75t_L g5012 ( 
.A(n_3253),
.Y(n_5012)
);

INVx1_ASAP7_75t_SL g5013 ( 
.A(n_1893),
.Y(n_5013)
);

BUFx6f_ASAP7_75t_L g5014 ( 
.A(n_2066),
.Y(n_5014)
);

INVx2_ASAP7_75t_L g5015 ( 
.A(n_161),
.Y(n_5015)
);

CKINVDCx5p33_ASAP7_75t_R g5016 ( 
.A(n_3361),
.Y(n_5016)
);

CKINVDCx20_ASAP7_75t_R g5017 ( 
.A(n_1108),
.Y(n_5017)
);

INVx1_ASAP7_75t_L g5018 ( 
.A(n_3462),
.Y(n_5018)
);

BUFx2_ASAP7_75t_L g5019 ( 
.A(n_2368),
.Y(n_5019)
);

CKINVDCx5p33_ASAP7_75t_R g5020 ( 
.A(n_2678),
.Y(n_5020)
);

CKINVDCx5p33_ASAP7_75t_R g5021 ( 
.A(n_2474),
.Y(n_5021)
);

CKINVDCx20_ASAP7_75t_R g5022 ( 
.A(n_2799),
.Y(n_5022)
);

BUFx10_ASAP7_75t_L g5023 ( 
.A(n_2579),
.Y(n_5023)
);

INVx2_ASAP7_75t_SL g5024 ( 
.A(n_3879),
.Y(n_5024)
);

INVx1_ASAP7_75t_L g5025 ( 
.A(n_2307),
.Y(n_5025)
);

INVx1_ASAP7_75t_L g5026 ( 
.A(n_1688),
.Y(n_5026)
);

CKINVDCx5p33_ASAP7_75t_R g5027 ( 
.A(n_3359),
.Y(n_5027)
);

CKINVDCx5p33_ASAP7_75t_R g5028 ( 
.A(n_2409),
.Y(n_5028)
);

INVx2_ASAP7_75t_L g5029 ( 
.A(n_2272),
.Y(n_5029)
);

CKINVDCx5p33_ASAP7_75t_R g5030 ( 
.A(n_270),
.Y(n_5030)
);

BUFx6f_ASAP7_75t_L g5031 ( 
.A(n_2225),
.Y(n_5031)
);

BUFx2_ASAP7_75t_L g5032 ( 
.A(n_160),
.Y(n_5032)
);

CKINVDCx20_ASAP7_75t_R g5033 ( 
.A(n_4044),
.Y(n_5033)
);

CKINVDCx5p33_ASAP7_75t_R g5034 ( 
.A(n_1085),
.Y(n_5034)
);

CKINVDCx5p33_ASAP7_75t_R g5035 ( 
.A(n_2388),
.Y(n_5035)
);

CKINVDCx5p33_ASAP7_75t_R g5036 ( 
.A(n_2109),
.Y(n_5036)
);

CKINVDCx5p33_ASAP7_75t_R g5037 ( 
.A(n_3901),
.Y(n_5037)
);

CKINVDCx5p33_ASAP7_75t_R g5038 ( 
.A(n_3210),
.Y(n_5038)
);

CKINVDCx5p33_ASAP7_75t_R g5039 ( 
.A(n_3987),
.Y(n_5039)
);

CKINVDCx5p33_ASAP7_75t_R g5040 ( 
.A(n_1657),
.Y(n_5040)
);

INVx1_ASAP7_75t_L g5041 ( 
.A(n_1957),
.Y(n_5041)
);

CKINVDCx16_ASAP7_75t_R g5042 ( 
.A(n_3043),
.Y(n_5042)
);

INVx1_ASAP7_75t_L g5043 ( 
.A(n_1868),
.Y(n_5043)
);

CKINVDCx5p33_ASAP7_75t_R g5044 ( 
.A(n_2037),
.Y(n_5044)
);

INVx1_ASAP7_75t_L g5045 ( 
.A(n_40),
.Y(n_5045)
);

CKINVDCx5p33_ASAP7_75t_R g5046 ( 
.A(n_3885),
.Y(n_5046)
);

INVx1_ASAP7_75t_L g5047 ( 
.A(n_1571),
.Y(n_5047)
);

INVx1_ASAP7_75t_L g5048 ( 
.A(n_523),
.Y(n_5048)
);

CKINVDCx5p33_ASAP7_75t_R g5049 ( 
.A(n_3655),
.Y(n_5049)
);

CKINVDCx20_ASAP7_75t_R g5050 ( 
.A(n_3449),
.Y(n_5050)
);

CKINVDCx5p33_ASAP7_75t_R g5051 ( 
.A(n_1760),
.Y(n_5051)
);

INVx1_ASAP7_75t_L g5052 ( 
.A(n_4032),
.Y(n_5052)
);

BUFx6f_ASAP7_75t_L g5053 ( 
.A(n_3064),
.Y(n_5053)
);

INVx1_ASAP7_75t_L g5054 ( 
.A(n_2538),
.Y(n_5054)
);

CKINVDCx5p33_ASAP7_75t_R g5055 ( 
.A(n_1186),
.Y(n_5055)
);

CKINVDCx5p33_ASAP7_75t_R g5056 ( 
.A(n_1793),
.Y(n_5056)
);

INVx1_ASAP7_75t_L g5057 ( 
.A(n_3701),
.Y(n_5057)
);

CKINVDCx5p33_ASAP7_75t_R g5058 ( 
.A(n_3682),
.Y(n_5058)
);

CKINVDCx5p33_ASAP7_75t_R g5059 ( 
.A(n_750),
.Y(n_5059)
);

CKINVDCx5p33_ASAP7_75t_R g5060 ( 
.A(n_1570),
.Y(n_5060)
);

CKINVDCx5p33_ASAP7_75t_R g5061 ( 
.A(n_2806),
.Y(n_5061)
);

INVx1_ASAP7_75t_L g5062 ( 
.A(n_1630),
.Y(n_5062)
);

INVx2_ASAP7_75t_L g5063 ( 
.A(n_1749),
.Y(n_5063)
);

CKINVDCx5p33_ASAP7_75t_R g5064 ( 
.A(n_1804),
.Y(n_5064)
);

CKINVDCx5p33_ASAP7_75t_R g5065 ( 
.A(n_3918),
.Y(n_5065)
);

INVx2_ASAP7_75t_L g5066 ( 
.A(n_1893),
.Y(n_5066)
);

CKINVDCx16_ASAP7_75t_R g5067 ( 
.A(n_1913),
.Y(n_5067)
);

INVx1_ASAP7_75t_L g5068 ( 
.A(n_3328),
.Y(n_5068)
);

INVx1_ASAP7_75t_L g5069 ( 
.A(n_3006),
.Y(n_5069)
);

BUFx10_ASAP7_75t_L g5070 ( 
.A(n_1105),
.Y(n_5070)
);

CKINVDCx16_ASAP7_75t_R g5071 ( 
.A(n_812),
.Y(n_5071)
);

CKINVDCx5p33_ASAP7_75t_R g5072 ( 
.A(n_949),
.Y(n_5072)
);

INVx1_ASAP7_75t_L g5073 ( 
.A(n_2831),
.Y(n_5073)
);

INVx1_ASAP7_75t_SL g5074 ( 
.A(n_959),
.Y(n_5074)
);

CKINVDCx5p33_ASAP7_75t_R g5075 ( 
.A(n_1094),
.Y(n_5075)
);

CKINVDCx5p33_ASAP7_75t_R g5076 ( 
.A(n_3943),
.Y(n_5076)
);

INVx1_ASAP7_75t_L g5077 ( 
.A(n_496),
.Y(n_5077)
);

CKINVDCx5p33_ASAP7_75t_R g5078 ( 
.A(n_3315),
.Y(n_5078)
);

CKINVDCx5p33_ASAP7_75t_R g5079 ( 
.A(n_2910),
.Y(n_5079)
);

CKINVDCx5p33_ASAP7_75t_R g5080 ( 
.A(n_3207),
.Y(n_5080)
);

CKINVDCx5p33_ASAP7_75t_R g5081 ( 
.A(n_1524),
.Y(n_5081)
);

CKINVDCx5p33_ASAP7_75t_R g5082 ( 
.A(n_3939),
.Y(n_5082)
);

INVx2_ASAP7_75t_SL g5083 ( 
.A(n_1459),
.Y(n_5083)
);

INVx1_ASAP7_75t_L g5084 ( 
.A(n_4030),
.Y(n_5084)
);

CKINVDCx5p33_ASAP7_75t_R g5085 ( 
.A(n_2549),
.Y(n_5085)
);

CKINVDCx5p33_ASAP7_75t_R g5086 ( 
.A(n_1182),
.Y(n_5086)
);

BUFx6f_ASAP7_75t_L g5087 ( 
.A(n_3948),
.Y(n_5087)
);

INVx1_ASAP7_75t_L g5088 ( 
.A(n_118),
.Y(n_5088)
);

CKINVDCx20_ASAP7_75t_R g5089 ( 
.A(n_900),
.Y(n_5089)
);

INVx1_ASAP7_75t_L g5090 ( 
.A(n_444),
.Y(n_5090)
);

INVx1_ASAP7_75t_L g5091 ( 
.A(n_3662),
.Y(n_5091)
);

CKINVDCx5p33_ASAP7_75t_R g5092 ( 
.A(n_354),
.Y(n_5092)
);

INVx1_ASAP7_75t_L g5093 ( 
.A(n_1916),
.Y(n_5093)
);

BUFx6f_ASAP7_75t_L g5094 ( 
.A(n_1028),
.Y(n_5094)
);

INVx1_ASAP7_75t_L g5095 ( 
.A(n_3274),
.Y(n_5095)
);

INVx1_ASAP7_75t_L g5096 ( 
.A(n_725),
.Y(n_5096)
);

INVx1_ASAP7_75t_L g5097 ( 
.A(n_3541),
.Y(n_5097)
);

BUFx10_ASAP7_75t_L g5098 ( 
.A(n_87),
.Y(n_5098)
);

CKINVDCx5p33_ASAP7_75t_R g5099 ( 
.A(n_3937),
.Y(n_5099)
);

CKINVDCx5p33_ASAP7_75t_R g5100 ( 
.A(n_628),
.Y(n_5100)
);

BUFx2_ASAP7_75t_L g5101 ( 
.A(n_3686),
.Y(n_5101)
);

CKINVDCx5p33_ASAP7_75t_R g5102 ( 
.A(n_3946),
.Y(n_5102)
);

CKINVDCx20_ASAP7_75t_R g5103 ( 
.A(n_3906),
.Y(n_5103)
);

INVx1_ASAP7_75t_L g5104 ( 
.A(n_3724),
.Y(n_5104)
);

INVx1_ASAP7_75t_L g5105 ( 
.A(n_1417),
.Y(n_5105)
);

INVx1_ASAP7_75t_L g5106 ( 
.A(n_1396),
.Y(n_5106)
);

CKINVDCx5p33_ASAP7_75t_R g5107 ( 
.A(n_638),
.Y(n_5107)
);

INVx1_ASAP7_75t_SL g5108 ( 
.A(n_1683),
.Y(n_5108)
);

CKINVDCx5p33_ASAP7_75t_R g5109 ( 
.A(n_447),
.Y(n_5109)
);

INVx1_ASAP7_75t_L g5110 ( 
.A(n_2422),
.Y(n_5110)
);

INVx1_ASAP7_75t_L g5111 ( 
.A(n_2248),
.Y(n_5111)
);

INVx1_ASAP7_75t_L g5112 ( 
.A(n_2179),
.Y(n_5112)
);

CKINVDCx5p33_ASAP7_75t_R g5113 ( 
.A(n_438),
.Y(n_5113)
);

CKINVDCx5p33_ASAP7_75t_R g5114 ( 
.A(n_4041),
.Y(n_5114)
);

HB1xp67_ASAP7_75t_L g5115 ( 
.A(n_1907),
.Y(n_5115)
);

BUFx10_ASAP7_75t_L g5116 ( 
.A(n_2720),
.Y(n_5116)
);

CKINVDCx5p33_ASAP7_75t_R g5117 ( 
.A(n_3061),
.Y(n_5117)
);

INVx1_ASAP7_75t_L g5118 ( 
.A(n_530),
.Y(n_5118)
);

INVx1_ASAP7_75t_L g5119 ( 
.A(n_3106),
.Y(n_5119)
);

BUFx6f_ASAP7_75t_L g5120 ( 
.A(n_404),
.Y(n_5120)
);

BUFx6f_ASAP7_75t_L g5121 ( 
.A(n_1102),
.Y(n_5121)
);

CKINVDCx5p33_ASAP7_75t_R g5122 ( 
.A(n_3997),
.Y(n_5122)
);

BUFx10_ASAP7_75t_L g5123 ( 
.A(n_1116),
.Y(n_5123)
);

CKINVDCx5p33_ASAP7_75t_R g5124 ( 
.A(n_3642),
.Y(n_5124)
);

CKINVDCx5p33_ASAP7_75t_R g5125 ( 
.A(n_4008),
.Y(n_5125)
);

CKINVDCx5p33_ASAP7_75t_R g5126 ( 
.A(n_185),
.Y(n_5126)
);

INVx1_ASAP7_75t_L g5127 ( 
.A(n_2616),
.Y(n_5127)
);

CKINVDCx5p33_ASAP7_75t_R g5128 ( 
.A(n_1800),
.Y(n_5128)
);

CKINVDCx5p33_ASAP7_75t_R g5129 ( 
.A(n_2962),
.Y(n_5129)
);

CKINVDCx5p33_ASAP7_75t_R g5130 ( 
.A(n_3090),
.Y(n_5130)
);

INVx1_ASAP7_75t_L g5131 ( 
.A(n_209),
.Y(n_5131)
);

BUFx3_ASAP7_75t_L g5132 ( 
.A(n_1740),
.Y(n_5132)
);

INVx1_ASAP7_75t_L g5133 ( 
.A(n_3775),
.Y(n_5133)
);

INVx1_ASAP7_75t_L g5134 ( 
.A(n_3245),
.Y(n_5134)
);

INVx1_ASAP7_75t_L g5135 ( 
.A(n_1506),
.Y(n_5135)
);

CKINVDCx5p33_ASAP7_75t_R g5136 ( 
.A(n_2160),
.Y(n_5136)
);

CKINVDCx5p33_ASAP7_75t_R g5137 ( 
.A(n_3640),
.Y(n_5137)
);

INVx1_ASAP7_75t_L g5138 ( 
.A(n_1720),
.Y(n_5138)
);

INVx1_ASAP7_75t_L g5139 ( 
.A(n_426),
.Y(n_5139)
);

CKINVDCx5p33_ASAP7_75t_R g5140 ( 
.A(n_2078),
.Y(n_5140)
);

CKINVDCx5p33_ASAP7_75t_R g5141 ( 
.A(n_107),
.Y(n_5141)
);

CKINVDCx5p33_ASAP7_75t_R g5142 ( 
.A(n_1408),
.Y(n_5142)
);

HB1xp67_ASAP7_75t_SL g5143 ( 
.A(n_1921),
.Y(n_5143)
);

CKINVDCx20_ASAP7_75t_R g5144 ( 
.A(n_2870),
.Y(n_5144)
);

CKINVDCx5p33_ASAP7_75t_R g5145 ( 
.A(n_3949),
.Y(n_5145)
);

CKINVDCx5p33_ASAP7_75t_R g5146 ( 
.A(n_2591),
.Y(n_5146)
);

CKINVDCx5p33_ASAP7_75t_R g5147 ( 
.A(n_1780),
.Y(n_5147)
);

CKINVDCx5p33_ASAP7_75t_R g5148 ( 
.A(n_79),
.Y(n_5148)
);

CKINVDCx20_ASAP7_75t_R g5149 ( 
.A(n_3418),
.Y(n_5149)
);

CKINVDCx20_ASAP7_75t_R g5150 ( 
.A(n_1067),
.Y(n_5150)
);

CKINVDCx5p33_ASAP7_75t_R g5151 ( 
.A(n_3864),
.Y(n_5151)
);

HB1xp67_ASAP7_75t_L g5152 ( 
.A(n_447),
.Y(n_5152)
);

CKINVDCx5p33_ASAP7_75t_R g5153 ( 
.A(n_1740),
.Y(n_5153)
);

CKINVDCx5p33_ASAP7_75t_R g5154 ( 
.A(n_500),
.Y(n_5154)
);

CKINVDCx5p33_ASAP7_75t_R g5155 ( 
.A(n_549),
.Y(n_5155)
);

CKINVDCx5p33_ASAP7_75t_R g5156 ( 
.A(n_3061),
.Y(n_5156)
);

CKINVDCx5p33_ASAP7_75t_R g5157 ( 
.A(n_2272),
.Y(n_5157)
);

CKINVDCx5p33_ASAP7_75t_R g5158 ( 
.A(n_2783),
.Y(n_5158)
);

INVxp67_ASAP7_75t_SL g5159 ( 
.A(n_2658),
.Y(n_5159)
);

CKINVDCx5p33_ASAP7_75t_R g5160 ( 
.A(n_1665),
.Y(n_5160)
);

INVx1_ASAP7_75t_L g5161 ( 
.A(n_3870),
.Y(n_5161)
);

INVx1_ASAP7_75t_L g5162 ( 
.A(n_3988),
.Y(n_5162)
);

INVx1_ASAP7_75t_L g5163 ( 
.A(n_90),
.Y(n_5163)
);

BUFx10_ASAP7_75t_L g5164 ( 
.A(n_3715),
.Y(n_5164)
);

INVx2_ASAP7_75t_L g5165 ( 
.A(n_3986),
.Y(n_5165)
);

CKINVDCx5p33_ASAP7_75t_R g5166 ( 
.A(n_1245),
.Y(n_5166)
);

CKINVDCx5p33_ASAP7_75t_R g5167 ( 
.A(n_2668),
.Y(n_5167)
);

CKINVDCx5p33_ASAP7_75t_R g5168 ( 
.A(n_1988),
.Y(n_5168)
);

BUFx6f_ASAP7_75t_L g5169 ( 
.A(n_2145),
.Y(n_5169)
);

CKINVDCx5p33_ASAP7_75t_R g5170 ( 
.A(n_3736),
.Y(n_5170)
);

CKINVDCx20_ASAP7_75t_R g5171 ( 
.A(n_2093),
.Y(n_5171)
);

INVx1_ASAP7_75t_L g5172 ( 
.A(n_3365),
.Y(n_5172)
);

CKINVDCx5p33_ASAP7_75t_R g5173 ( 
.A(n_1375),
.Y(n_5173)
);

CKINVDCx5p33_ASAP7_75t_R g5174 ( 
.A(n_829),
.Y(n_5174)
);

CKINVDCx5p33_ASAP7_75t_R g5175 ( 
.A(n_1309),
.Y(n_5175)
);

INVx1_ASAP7_75t_SL g5176 ( 
.A(n_411),
.Y(n_5176)
);

CKINVDCx5p33_ASAP7_75t_R g5177 ( 
.A(n_1469),
.Y(n_5177)
);

INVx1_ASAP7_75t_L g5178 ( 
.A(n_3298),
.Y(n_5178)
);

CKINVDCx5p33_ASAP7_75t_R g5179 ( 
.A(n_1794),
.Y(n_5179)
);

INVx1_ASAP7_75t_L g5180 ( 
.A(n_2345),
.Y(n_5180)
);

CKINVDCx5p33_ASAP7_75t_R g5181 ( 
.A(n_471),
.Y(n_5181)
);

CKINVDCx5p33_ASAP7_75t_R g5182 ( 
.A(n_2232),
.Y(n_5182)
);

CKINVDCx5p33_ASAP7_75t_R g5183 ( 
.A(n_4005),
.Y(n_5183)
);

INVx1_ASAP7_75t_SL g5184 ( 
.A(n_442),
.Y(n_5184)
);

INVx1_ASAP7_75t_L g5185 ( 
.A(n_3178),
.Y(n_5185)
);

INVx1_ASAP7_75t_L g5186 ( 
.A(n_2428),
.Y(n_5186)
);

CKINVDCx16_ASAP7_75t_R g5187 ( 
.A(n_630),
.Y(n_5187)
);

CKINVDCx20_ASAP7_75t_R g5188 ( 
.A(n_791),
.Y(n_5188)
);

INVx1_ASAP7_75t_L g5189 ( 
.A(n_4002),
.Y(n_5189)
);

BUFx6f_ASAP7_75t_L g5190 ( 
.A(n_3911),
.Y(n_5190)
);

CKINVDCx5p33_ASAP7_75t_R g5191 ( 
.A(n_539),
.Y(n_5191)
);

CKINVDCx20_ASAP7_75t_R g5192 ( 
.A(n_3553),
.Y(n_5192)
);

CKINVDCx5p33_ASAP7_75t_R g5193 ( 
.A(n_2842),
.Y(n_5193)
);

CKINVDCx5p33_ASAP7_75t_R g5194 ( 
.A(n_1601),
.Y(n_5194)
);

CKINVDCx5p33_ASAP7_75t_R g5195 ( 
.A(n_3116),
.Y(n_5195)
);

BUFx10_ASAP7_75t_L g5196 ( 
.A(n_467),
.Y(n_5196)
);

CKINVDCx5p33_ASAP7_75t_R g5197 ( 
.A(n_319),
.Y(n_5197)
);

CKINVDCx5p33_ASAP7_75t_R g5198 ( 
.A(n_4055),
.Y(n_5198)
);

CKINVDCx14_ASAP7_75t_R g5199 ( 
.A(n_1418),
.Y(n_5199)
);

CKINVDCx5p33_ASAP7_75t_R g5200 ( 
.A(n_2991),
.Y(n_5200)
);

CKINVDCx20_ASAP7_75t_R g5201 ( 
.A(n_248),
.Y(n_5201)
);

CKINVDCx5p33_ASAP7_75t_R g5202 ( 
.A(n_4077),
.Y(n_5202)
);

CKINVDCx5p33_ASAP7_75t_R g5203 ( 
.A(n_2360),
.Y(n_5203)
);

CKINVDCx5p33_ASAP7_75t_R g5204 ( 
.A(n_3335),
.Y(n_5204)
);

INVx1_ASAP7_75t_L g5205 ( 
.A(n_143),
.Y(n_5205)
);

CKINVDCx5p33_ASAP7_75t_R g5206 ( 
.A(n_2103),
.Y(n_5206)
);

CKINVDCx5p33_ASAP7_75t_R g5207 ( 
.A(n_3007),
.Y(n_5207)
);

CKINVDCx5p33_ASAP7_75t_R g5208 ( 
.A(n_1051),
.Y(n_5208)
);

INVx1_ASAP7_75t_L g5209 ( 
.A(n_951),
.Y(n_5209)
);

INVx1_ASAP7_75t_L g5210 ( 
.A(n_1493),
.Y(n_5210)
);

CKINVDCx5p33_ASAP7_75t_R g5211 ( 
.A(n_4088),
.Y(n_5211)
);

INVx2_ASAP7_75t_L g5212 ( 
.A(n_725),
.Y(n_5212)
);

CKINVDCx5p33_ASAP7_75t_R g5213 ( 
.A(n_607),
.Y(n_5213)
);

BUFx2_ASAP7_75t_L g5214 ( 
.A(n_2056),
.Y(n_5214)
);

CKINVDCx5p33_ASAP7_75t_R g5215 ( 
.A(n_889),
.Y(n_5215)
);

CKINVDCx20_ASAP7_75t_R g5216 ( 
.A(n_3540),
.Y(n_5216)
);

INVx1_ASAP7_75t_L g5217 ( 
.A(n_1971),
.Y(n_5217)
);

INVx1_ASAP7_75t_L g5218 ( 
.A(n_1420),
.Y(n_5218)
);

CKINVDCx5p33_ASAP7_75t_R g5219 ( 
.A(n_3824),
.Y(n_5219)
);

INVx1_ASAP7_75t_L g5220 ( 
.A(n_3551),
.Y(n_5220)
);

BUFx2_ASAP7_75t_L g5221 ( 
.A(n_3627),
.Y(n_5221)
);

INVx1_ASAP7_75t_L g5222 ( 
.A(n_573),
.Y(n_5222)
);

INVx1_ASAP7_75t_L g5223 ( 
.A(n_3707),
.Y(n_5223)
);

INVx1_ASAP7_75t_SL g5224 ( 
.A(n_1680),
.Y(n_5224)
);

BUFx8_ASAP7_75t_SL g5225 ( 
.A(n_2823),
.Y(n_5225)
);

INVx2_ASAP7_75t_L g5226 ( 
.A(n_519),
.Y(n_5226)
);

INVx1_ASAP7_75t_L g5227 ( 
.A(n_2552),
.Y(n_5227)
);

CKINVDCx5p33_ASAP7_75t_R g5228 ( 
.A(n_1),
.Y(n_5228)
);

BUFx6f_ASAP7_75t_L g5229 ( 
.A(n_3863),
.Y(n_5229)
);

CKINVDCx5p33_ASAP7_75t_R g5230 ( 
.A(n_1847),
.Y(n_5230)
);

INVx1_ASAP7_75t_SL g5231 ( 
.A(n_2207),
.Y(n_5231)
);

CKINVDCx5p33_ASAP7_75t_R g5232 ( 
.A(n_346),
.Y(n_5232)
);

CKINVDCx20_ASAP7_75t_R g5233 ( 
.A(n_3764),
.Y(n_5233)
);

CKINVDCx20_ASAP7_75t_R g5234 ( 
.A(n_1453),
.Y(n_5234)
);

CKINVDCx5p33_ASAP7_75t_R g5235 ( 
.A(n_137),
.Y(n_5235)
);

CKINVDCx20_ASAP7_75t_R g5236 ( 
.A(n_1322),
.Y(n_5236)
);

INVx2_ASAP7_75t_SL g5237 ( 
.A(n_1550),
.Y(n_5237)
);

CKINVDCx14_ASAP7_75t_R g5238 ( 
.A(n_3933),
.Y(n_5238)
);

CKINVDCx20_ASAP7_75t_R g5239 ( 
.A(n_1589),
.Y(n_5239)
);

INVx1_ASAP7_75t_L g5240 ( 
.A(n_1569),
.Y(n_5240)
);

CKINVDCx5p33_ASAP7_75t_R g5241 ( 
.A(n_2789),
.Y(n_5241)
);

CKINVDCx5p33_ASAP7_75t_R g5242 ( 
.A(n_2392),
.Y(n_5242)
);

BUFx3_ASAP7_75t_L g5243 ( 
.A(n_570),
.Y(n_5243)
);

BUFx6f_ASAP7_75t_L g5244 ( 
.A(n_3904),
.Y(n_5244)
);

INVx1_ASAP7_75t_L g5245 ( 
.A(n_3367),
.Y(n_5245)
);

CKINVDCx5p33_ASAP7_75t_R g5246 ( 
.A(n_4040),
.Y(n_5246)
);

CKINVDCx5p33_ASAP7_75t_R g5247 ( 
.A(n_2953),
.Y(n_5247)
);

CKINVDCx20_ASAP7_75t_R g5248 ( 
.A(n_3929),
.Y(n_5248)
);

INVx1_ASAP7_75t_L g5249 ( 
.A(n_1008),
.Y(n_5249)
);

INVx1_ASAP7_75t_L g5250 ( 
.A(n_3966),
.Y(n_5250)
);

CKINVDCx5p33_ASAP7_75t_R g5251 ( 
.A(n_3524),
.Y(n_5251)
);

CKINVDCx5p33_ASAP7_75t_R g5252 ( 
.A(n_1049),
.Y(n_5252)
);

INVx1_ASAP7_75t_L g5253 ( 
.A(n_1800),
.Y(n_5253)
);

INVx1_ASAP7_75t_SL g5254 ( 
.A(n_4004),
.Y(n_5254)
);

INVx1_ASAP7_75t_L g5255 ( 
.A(n_2197),
.Y(n_5255)
);

CKINVDCx5p33_ASAP7_75t_R g5256 ( 
.A(n_1199),
.Y(n_5256)
);

INVx2_ASAP7_75t_L g5257 ( 
.A(n_3999),
.Y(n_5257)
);

CKINVDCx5p33_ASAP7_75t_R g5258 ( 
.A(n_1816),
.Y(n_5258)
);

CKINVDCx5p33_ASAP7_75t_R g5259 ( 
.A(n_1157),
.Y(n_5259)
);

INVx1_ASAP7_75t_L g5260 ( 
.A(n_1119),
.Y(n_5260)
);

INVx1_ASAP7_75t_L g5261 ( 
.A(n_1516),
.Y(n_5261)
);

CKINVDCx5p33_ASAP7_75t_R g5262 ( 
.A(n_651),
.Y(n_5262)
);

CKINVDCx5p33_ASAP7_75t_R g5263 ( 
.A(n_1795),
.Y(n_5263)
);

CKINVDCx5p33_ASAP7_75t_R g5264 ( 
.A(n_3290),
.Y(n_5264)
);

CKINVDCx5p33_ASAP7_75t_R g5265 ( 
.A(n_4015),
.Y(n_5265)
);

CKINVDCx5p33_ASAP7_75t_R g5266 ( 
.A(n_2071),
.Y(n_5266)
);

INVx1_ASAP7_75t_L g5267 ( 
.A(n_623),
.Y(n_5267)
);

CKINVDCx20_ASAP7_75t_R g5268 ( 
.A(n_3899),
.Y(n_5268)
);

CKINVDCx5p33_ASAP7_75t_R g5269 ( 
.A(n_3883),
.Y(n_5269)
);

INVx1_ASAP7_75t_L g5270 ( 
.A(n_3919),
.Y(n_5270)
);

CKINVDCx5p33_ASAP7_75t_R g5271 ( 
.A(n_215),
.Y(n_5271)
);

INVx1_ASAP7_75t_L g5272 ( 
.A(n_2161),
.Y(n_5272)
);

INVx1_ASAP7_75t_L g5273 ( 
.A(n_3857),
.Y(n_5273)
);

CKINVDCx5p33_ASAP7_75t_R g5274 ( 
.A(n_1280),
.Y(n_5274)
);

INVx1_ASAP7_75t_L g5275 ( 
.A(n_4019),
.Y(n_5275)
);

CKINVDCx5p33_ASAP7_75t_R g5276 ( 
.A(n_3871),
.Y(n_5276)
);

CKINVDCx5p33_ASAP7_75t_R g5277 ( 
.A(n_3631),
.Y(n_5277)
);

INVx1_ASAP7_75t_L g5278 ( 
.A(n_2926),
.Y(n_5278)
);

INVx1_ASAP7_75t_L g5279 ( 
.A(n_1868),
.Y(n_5279)
);

CKINVDCx5p33_ASAP7_75t_R g5280 ( 
.A(n_1346),
.Y(n_5280)
);

BUFx3_ASAP7_75t_L g5281 ( 
.A(n_2357),
.Y(n_5281)
);

CKINVDCx5p33_ASAP7_75t_R g5282 ( 
.A(n_3587),
.Y(n_5282)
);

CKINVDCx5p33_ASAP7_75t_R g5283 ( 
.A(n_3220),
.Y(n_5283)
);

INVx1_ASAP7_75t_L g5284 ( 
.A(n_3265),
.Y(n_5284)
);

CKINVDCx5p33_ASAP7_75t_R g5285 ( 
.A(n_3797),
.Y(n_5285)
);

BUFx10_ASAP7_75t_L g5286 ( 
.A(n_2423),
.Y(n_5286)
);

INVx1_ASAP7_75t_L g5287 ( 
.A(n_2779),
.Y(n_5287)
);

CKINVDCx5p33_ASAP7_75t_R g5288 ( 
.A(n_4023),
.Y(n_5288)
);

CKINVDCx5p33_ASAP7_75t_R g5289 ( 
.A(n_2684),
.Y(n_5289)
);

BUFx10_ASAP7_75t_L g5290 ( 
.A(n_834),
.Y(n_5290)
);

INVx1_ASAP7_75t_L g5291 ( 
.A(n_1174),
.Y(n_5291)
);

CKINVDCx5p33_ASAP7_75t_R g5292 ( 
.A(n_855),
.Y(n_5292)
);

INVx1_ASAP7_75t_L g5293 ( 
.A(n_3889),
.Y(n_5293)
);

CKINVDCx5p33_ASAP7_75t_R g5294 ( 
.A(n_2007),
.Y(n_5294)
);

BUFx6f_ASAP7_75t_L g5295 ( 
.A(n_1863),
.Y(n_5295)
);

INVx1_ASAP7_75t_SL g5296 ( 
.A(n_3895),
.Y(n_5296)
);

BUFx2_ASAP7_75t_L g5297 ( 
.A(n_1437),
.Y(n_5297)
);

CKINVDCx5p33_ASAP7_75t_R g5298 ( 
.A(n_4062),
.Y(n_5298)
);

CKINVDCx5p33_ASAP7_75t_R g5299 ( 
.A(n_2654),
.Y(n_5299)
);

CKINVDCx5p33_ASAP7_75t_R g5300 ( 
.A(n_396),
.Y(n_5300)
);

BUFx2_ASAP7_75t_L g5301 ( 
.A(n_1720),
.Y(n_5301)
);

CKINVDCx5p33_ASAP7_75t_R g5302 ( 
.A(n_1568),
.Y(n_5302)
);

BUFx2_ASAP7_75t_L g5303 ( 
.A(n_3323),
.Y(n_5303)
);

CKINVDCx5p33_ASAP7_75t_R g5304 ( 
.A(n_2159),
.Y(n_5304)
);

CKINVDCx5p33_ASAP7_75t_R g5305 ( 
.A(n_150),
.Y(n_5305)
);

BUFx6f_ASAP7_75t_L g5306 ( 
.A(n_3254),
.Y(n_5306)
);

HB1xp67_ASAP7_75t_L g5307 ( 
.A(n_2748),
.Y(n_5307)
);

INVx1_ASAP7_75t_L g5308 ( 
.A(n_2374),
.Y(n_5308)
);

INVx1_ASAP7_75t_L g5309 ( 
.A(n_1121),
.Y(n_5309)
);

CKINVDCx5p33_ASAP7_75t_R g5310 ( 
.A(n_1895),
.Y(n_5310)
);

CKINVDCx5p33_ASAP7_75t_R g5311 ( 
.A(n_3680),
.Y(n_5311)
);

CKINVDCx5p33_ASAP7_75t_R g5312 ( 
.A(n_2786),
.Y(n_5312)
);

INVx1_ASAP7_75t_L g5313 ( 
.A(n_1234),
.Y(n_5313)
);

CKINVDCx5p33_ASAP7_75t_R g5314 ( 
.A(n_1950),
.Y(n_5314)
);

CKINVDCx5p33_ASAP7_75t_R g5315 ( 
.A(n_189),
.Y(n_5315)
);

INVx1_ASAP7_75t_L g5316 ( 
.A(n_1272),
.Y(n_5316)
);

CKINVDCx5p33_ASAP7_75t_R g5317 ( 
.A(n_2279),
.Y(n_5317)
);

CKINVDCx5p33_ASAP7_75t_R g5318 ( 
.A(n_3127),
.Y(n_5318)
);

CKINVDCx5p33_ASAP7_75t_R g5319 ( 
.A(n_3882),
.Y(n_5319)
);

CKINVDCx5p33_ASAP7_75t_R g5320 ( 
.A(n_243),
.Y(n_5320)
);

INVx1_ASAP7_75t_L g5321 ( 
.A(n_820),
.Y(n_5321)
);

CKINVDCx5p33_ASAP7_75t_R g5322 ( 
.A(n_3547),
.Y(n_5322)
);

CKINVDCx5p33_ASAP7_75t_R g5323 ( 
.A(n_470),
.Y(n_5323)
);

INVx2_ASAP7_75t_L g5324 ( 
.A(n_3884),
.Y(n_5324)
);

BUFx10_ASAP7_75t_L g5325 ( 
.A(n_2868),
.Y(n_5325)
);

CKINVDCx5p33_ASAP7_75t_R g5326 ( 
.A(n_2240),
.Y(n_5326)
);

INVx1_ASAP7_75t_L g5327 ( 
.A(n_900),
.Y(n_5327)
);

INVx1_ASAP7_75t_L g5328 ( 
.A(n_2096),
.Y(n_5328)
);

INVx2_ASAP7_75t_L g5329 ( 
.A(n_1965),
.Y(n_5329)
);

CKINVDCx5p33_ASAP7_75t_R g5330 ( 
.A(n_1167),
.Y(n_5330)
);

CKINVDCx5p33_ASAP7_75t_R g5331 ( 
.A(n_3704),
.Y(n_5331)
);

BUFx8_ASAP7_75t_SL g5332 ( 
.A(n_1940),
.Y(n_5332)
);

INVx1_ASAP7_75t_L g5333 ( 
.A(n_96),
.Y(n_5333)
);

CKINVDCx5p33_ASAP7_75t_R g5334 ( 
.A(n_3984),
.Y(n_5334)
);

CKINVDCx5p33_ASAP7_75t_R g5335 ( 
.A(n_377),
.Y(n_5335)
);

CKINVDCx5p33_ASAP7_75t_R g5336 ( 
.A(n_3812),
.Y(n_5336)
);

BUFx10_ASAP7_75t_L g5337 ( 
.A(n_3398),
.Y(n_5337)
);

CKINVDCx5p33_ASAP7_75t_R g5338 ( 
.A(n_135),
.Y(n_5338)
);

INVx1_ASAP7_75t_L g5339 ( 
.A(n_199),
.Y(n_5339)
);

CKINVDCx5p33_ASAP7_75t_R g5340 ( 
.A(n_3479),
.Y(n_5340)
);

INVxp67_ASAP7_75t_L g5341 ( 
.A(n_3775),
.Y(n_5341)
);

INVx1_ASAP7_75t_L g5342 ( 
.A(n_1856),
.Y(n_5342)
);

CKINVDCx5p33_ASAP7_75t_R g5343 ( 
.A(n_3910),
.Y(n_5343)
);

CKINVDCx5p33_ASAP7_75t_R g5344 ( 
.A(n_686),
.Y(n_5344)
);

HB1xp67_ASAP7_75t_L g5345 ( 
.A(n_3024),
.Y(n_5345)
);

INVx1_ASAP7_75t_L g5346 ( 
.A(n_1662),
.Y(n_5346)
);

CKINVDCx5p33_ASAP7_75t_R g5347 ( 
.A(n_4046),
.Y(n_5347)
);

INVx2_ASAP7_75t_L g5348 ( 
.A(n_3968),
.Y(n_5348)
);

CKINVDCx5p33_ASAP7_75t_R g5349 ( 
.A(n_2257),
.Y(n_5349)
);

CKINVDCx5p33_ASAP7_75t_R g5350 ( 
.A(n_2777),
.Y(n_5350)
);

CKINVDCx5p33_ASAP7_75t_R g5351 ( 
.A(n_2978),
.Y(n_5351)
);

CKINVDCx16_ASAP7_75t_R g5352 ( 
.A(n_2560),
.Y(n_5352)
);

INVx1_ASAP7_75t_L g5353 ( 
.A(n_4095),
.Y(n_5353)
);

CKINVDCx5p33_ASAP7_75t_R g5354 ( 
.A(n_1023),
.Y(n_5354)
);

CKINVDCx5p33_ASAP7_75t_R g5355 ( 
.A(n_3634),
.Y(n_5355)
);

INVx1_ASAP7_75t_L g5356 ( 
.A(n_923),
.Y(n_5356)
);

INVx1_ASAP7_75t_L g5357 ( 
.A(n_3876),
.Y(n_5357)
);

CKINVDCx5p33_ASAP7_75t_R g5358 ( 
.A(n_2477),
.Y(n_5358)
);

CKINVDCx5p33_ASAP7_75t_R g5359 ( 
.A(n_4030),
.Y(n_5359)
);

CKINVDCx5p33_ASAP7_75t_R g5360 ( 
.A(n_2147),
.Y(n_5360)
);

INVx1_ASAP7_75t_L g5361 ( 
.A(n_356),
.Y(n_5361)
);

CKINVDCx5p33_ASAP7_75t_R g5362 ( 
.A(n_577),
.Y(n_5362)
);

CKINVDCx5p33_ASAP7_75t_R g5363 ( 
.A(n_2069),
.Y(n_5363)
);

CKINVDCx5p33_ASAP7_75t_R g5364 ( 
.A(n_286),
.Y(n_5364)
);

CKINVDCx5p33_ASAP7_75t_R g5365 ( 
.A(n_4031),
.Y(n_5365)
);

INVx1_ASAP7_75t_L g5366 ( 
.A(n_3952),
.Y(n_5366)
);

CKINVDCx20_ASAP7_75t_R g5367 ( 
.A(n_1338),
.Y(n_5367)
);

BUFx6f_ASAP7_75t_L g5368 ( 
.A(n_3826),
.Y(n_5368)
);

INVx1_ASAP7_75t_SL g5369 ( 
.A(n_2383),
.Y(n_5369)
);

CKINVDCx5p33_ASAP7_75t_R g5370 ( 
.A(n_2392),
.Y(n_5370)
);

HB1xp67_ASAP7_75t_L g5371 ( 
.A(n_495),
.Y(n_5371)
);

CKINVDCx20_ASAP7_75t_R g5372 ( 
.A(n_3902),
.Y(n_5372)
);

CKINVDCx5p33_ASAP7_75t_R g5373 ( 
.A(n_3354),
.Y(n_5373)
);

INVx1_ASAP7_75t_SL g5374 ( 
.A(n_3738),
.Y(n_5374)
);

INVx1_ASAP7_75t_L g5375 ( 
.A(n_2309),
.Y(n_5375)
);

INVx2_ASAP7_75t_L g5376 ( 
.A(n_3002),
.Y(n_5376)
);

CKINVDCx5p33_ASAP7_75t_R g5377 ( 
.A(n_3890),
.Y(n_5377)
);

CKINVDCx5p33_ASAP7_75t_R g5378 ( 
.A(n_3153),
.Y(n_5378)
);

CKINVDCx5p33_ASAP7_75t_R g5379 ( 
.A(n_2384),
.Y(n_5379)
);

CKINVDCx5p33_ASAP7_75t_R g5380 ( 
.A(n_3734),
.Y(n_5380)
);

INVx1_ASAP7_75t_L g5381 ( 
.A(n_3971),
.Y(n_5381)
);

CKINVDCx5p33_ASAP7_75t_R g5382 ( 
.A(n_2042),
.Y(n_5382)
);

CKINVDCx5p33_ASAP7_75t_R g5383 ( 
.A(n_936),
.Y(n_5383)
);

INVx1_ASAP7_75t_L g5384 ( 
.A(n_2877),
.Y(n_5384)
);

CKINVDCx5p33_ASAP7_75t_R g5385 ( 
.A(n_2638),
.Y(n_5385)
);

INVx1_ASAP7_75t_L g5386 ( 
.A(n_3746),
.Y(n_5386)
);

CKINVDCx5p33_ASAP7_75t_R g5387 ( 
.A(n_1738),
.Y(n_5387)
);

CKINVDCx5p33_ASAP7_75t_R g5388 ( 
.A(n_1376),
.Y(n_5388)
);

INVx1_ASAP7_75t_L g5389 ( 
.A(n_866),
.Y(n_5389)
);

CKINVDCx5p33_ASAP7_75t_R g5390 ( 
.A(n_623),
.Y(n_5390)
);

CKINVDCx5p33_ASAP7_75t_R g5391 ( 
.A(n_972),
.Y(n_5391)
);

BUFx6f_ASAP7_75t_L g5392 ( 
.A(n_2342),
.Y(n_5392)
);

CKINVDCx5p33_ASAP7_75t_R g5393 ( 
.A(n_2652),
.Y(n_5393)
);

INVx2_ASAP7_75t_L g5394 ( 
.A(n_4039),
.Y(n_5394)
);

CKINVDCx20_ASAP7_75t_R g5395 ( 
.A(n_3208),
.Y(n_5395)
);

INVx2_ASAP7_75t_SL g5396 ( 
.A(n_2875),
.Y(n_5396)
);

CKINVDCx5p33_ASAP7_75t_R g5397 ( 
.A(n_3458),
.Y(n_5397)
);

CKINVDCx5p33_ASAP7_75t_R g5398 ( 
.A(n_888),
.Y(n_5398)
);

CKINVDCx5p33_ASAP7_75t_R g5399 ( 
.A(n_129),
.Y(n_5399)
);

INVx1_ASAP7_75t_L g5400 ( 
.A(n_151),
.Y(n_5400)
);

CKINVDCx5p33_ASAP7_75t_R g5401 ( 
.A(n_617),
.Y(n_5401)
);

INVx1_ASAP7_75t_L g5402 ( 
.A(n_3964),
.Y(n_5402)
);

INVx2_ASAP7_75t_L g5403 ( 
.A(n_1371),
.Y(n_5403)
);

BUFx2_ASAP7_75t_L g5404 ( 
.A(n_2179),
.Y(n_5404)
);

BUFx3_ASAP7_75t_L g5405 ( 
.A(n_829),
.Y(n_5405)
);

CKINVDCx5p33_ASAP7_75t_R g5406 ( 
.A(n_854),
.Y(n_5406)
);

CKINVDCx5p33_ASAP7_75t_R g5407 ( 
.A(n_1288),
.Y(n_5407)
);

BUFx5_ASAP7_75t_L g5408 ( 
.A(n_3870),
.Y(n_5408)
);

CKINVDCx5p33_ASAP7_75t_R g5409 ( 
.A(n_1833),
.Y(n_5409)
);

INVx2_ASAP7_75t_SL g5410 ( 
.A(n_2464),
.Y(n_5410)
);

INVx1_ASAP7_75t_L g5411 ( 
.A(n_3311),
.Y(n_5411)
);

CKINVDCx20_ASAP7_75t_R g5412 ( 
.A(n_1732),
.Y(n_5412)
);

CKINVDCx5p33_ASAP7_75t_R g5413 ( 
.A(n_436),
.Y(n_5413)
);

CKINVDCx11_ASAP7_75t_R g5414 ( 
.A(n_3062),
.Y(n_5414)
);

CKINVDCx20_ASAP7_75t_R g5415 ( 
.A(n_788),
.Y(n_5415)
);

CKINVDCx20_ASAP7_75t_R g5416 ( 
.A(n_3475),
.Y(n_5416)
);

INVx2_ASAP7_75t_SL g5417 ( 
.A(n_2553),
.Y(n_5417)
);

CKINVDCx5p33_ASAP7_75t_R g5418 ( 
.A(n_2784),
.Y(n_5418)
);

CKINVDCx5p33_ASAP7_75t_R g5419 ( 
.A(n_2836),
.Y(n_5419)
);

CKINVDCx5p33_ASAP7_75t_R g5420 ( 
.A(n_2187),
.Y(n_5420)
);

CKINVDCx5p33_ASAP7_75t_R g5421 ( 
.A(n_4066),
.Y(n_5421)
);

INVx1_ASAP7_75t_L g5422 ( 
.A(n_1086),
.Y(n_5422)
);

INVx1_ASAP7_75t_L g5423 ( 
.A(n_158),
.Y(n_5423)
);

BUFx2_ASAP7_75t_SL g5424 ( 
.A(n_69),
.Y(n_5424)
);

CKINVDCx5p33_ASAP7_75t_R g5425 ( 
.A(n_958),
.Y(n_5425)
);

CKINVDCx5p33_ASAP7_75t_R g5426 ( 
.A(n_765),
.Y(n_5426)
);

INVx1_ASAP7_75t_L g5427 ( 
.A(n_355),
.Y(n_5427)
);

CKINVDCx5p33_ASAP7_75t_R g5428 ( 
.A(n_1982),
.Y(n_5428)
);

CKINVDCx20_ASAP7_75t_R g5429 ( 
.A(n_2932),
.Y(n_5429)
);

INVx1_ASAP7_75t_L g5430 ( 
.A(n_3967),
.Y(n_5430)
);

INVx1_ASAP7_75t_L g5431 ( 
.A(n_3915),
.Y(n_5431)
);

CKINVDCx5p33_ASAP7_75t_R g5432 ( 
.A(n_1384),
.Y(n_5432)
);

INVx1_ASAP7_75t_L g5433 ( 
.A(n_3270),
.Y(n_5433)
);

CKINVDCx20_ASAP7_75t_R g5434 ( 
.A(n_2230),
.Y(n_5434)
);

CKINVDCx5p33_ASAP7_75t_R g5435 ( 
.A(n_4003),
.Y(n_5435)
);

INVx1_ASAP7_75t_L g5436 ( 
.A(n_93),
.Y(n_5436)
);

CKINVDCx5p33_ASAP7_75t_R g5437 ( 
.A(n_2660),
.Y(n_5437)
);

BUFx10_ASAP7_75t_L g5438 ( 
.A(n_3968),
.Y(n_5438)
);

CKINVDCx5p33_ASAP7_75t_R g5439 ( 
.A(n_3428),
.Y(n_5439)
);

CKINVDCx5p33_ASAP7_75t_R g5440 ( 
.A(n_1485),
.Y(n_5440)
);

BUFx2_ASAP7_75t_L g5441 ( 
.A(n_4027),
.Y(n_5441)
);

BUFx10_ASAP7_75t_L g5442 ( 
.A(n_3162),
.Y(n_5442)
);

CKINVDCx5p33_ASAP7_75t_R g5443 ( 
.A(n_988),
.Y(n_5443)
);

CKINVDCx5p33_ASAP7_75t_R g5444 ( 
.A(n_2064),
.Y(n_5444)
);

CKINVDCx5p33_ASAP7_75t_R g5445 ( 
.A(n_1983),
.Y(n_5445)
);

CKINVDCx5p33_ASAP7_75t_R g5446 ( 
.A(n_1333),
.Y(n_5446)
);

CKINVDCx5p33_ASAP7_75t_R g5447 ( 
.A(n_3892),
.Y(n_5447)
);

CKINVDCx5p33_ASAP7_75t_R g5448 ( 
.A(n_519),
.Y(n_5448)
);

INVx1_ASAP7_75t_L g5449 ( 
.A(n_2295),
.Y(n_5449)
);

BUFx10_ASAP7_75t_L g5450 ( 
.A(n_3241),
.Y(n_5450)
);

CKINVDCx5p33_ASAP7_75t_R g5451 ( 
.A(n_1356),
.Y(n_5451)
);

INVx2_ASAP7_75t_L g5452 ( 
.A(n_980),
.Y(n_5452)
);

CKINVDCx5p33_ASAP7_75t_R g5453 ( 
.A(n_304),
.Y(n_5453)
);

INVx1_ASAP7_75t_L g5454 ( 
.A(n_3707),
.Y(n_5454)
);

INVx1_ASAP7_75t_L g5455 ( 
.A(n_3928),
.Y(n_5455)
);

CKINVDCx5p33_ASAP7_75t_R g5456 ( 
.A(n_3722),
.Y(n_5456)
);

CKINVDCx16_ASAP7_75t_R g5457 ( 
.A(n_3951),
.Y(n_5457)
);

INVx2_ASAP7_75t_L g5458 ( 
.A(n_4004),
.Y(n_5458)
);

BUFx8_ASAP7_75t_SL g5459 ( 
.A(n_428),
.Y(n_5459)
);

INVx1_ASAP7_75t_L g5460 ( 
.A(n_4066),
.Y(n_5460)
);

INVx1_ASAP7_75t_L g5461 ( 
.A(n_1962),
.Y(n_5461)
);

CKINVDCx5p33_ASAP7_75t_R g5462 ( 
.A(n_3829),
.Y(n_5462)
);

CKINVDCx5p33_ASAP7_75t_R g5463 ( 
.A(n_1034),
.Y(n_5463)
);

CKINVDCx5p33_ASAP7_75t_R g5464 ( 
.A(n_1290),
.Y(n_5464)
);

CKINVDCx5p33_ASAP7_75t_R g5465 ( 
.A(n_3936),
.Y(n_5465)
);

CKINVDCx5p33_ASAP7_75t_R g5466 ( 
.A(n_100),
.Y(n_5466)
);

BUFx3_ASAP7_75t_L g5467 ( 
.A(n_1105),
.Y(n_5467)
);

CKINVDCx5p33_ASAP7_75t_R g5468 ( 
.A(n_3849),
.Y(n_5468)
);

INVx2_ASAP7_75t_L g5469 ( 
.A(n_1772),
.Y(n_5469)
);

INVx1_ASAP7_75t_L g5470 ( 
.A(n_4019),
.Y(n_5470)
);

CKINVDCx5p33_ASAP7_75t_R g5471 ( 
.A(n_507),
.Y(n_5471)
);

CKINVDCx5p33_ASAP7_75t_R g5472 ( 
.A(n_3972),
.Y(n_5472)
);

BUFx3_ASAP7_75t_L g5473 ( 
.A(n_3438),
.Y(n_5473)
);

BUFx6f_ASAP7_75t_L g5474 ( 
.A(n_2560),
.Y(n_5474)
);

CKINVDCx16_ASAP7_75t_R g5475 ( 
.A(n_3953),
.Y(n_5475)
);

CKINVDCx5p33_ASAP7_75t_R g5476 ( 
.A(n_3730),
.Y(n_5476)
);

INVx1_ASAP7_75t_L g5477 ( 
.A(n_194),
.Y(n_5477)
);

INVx1_ASAP7_75t_L g5478 ( 
.A(n_2327),
.Y(n_5478)
);

CKINVDCx5p33_ASAP7_75t_R g5479 ( 
.A(n_3335),
.Y(n_5479)
);

INVx1_ASAP7_75t_L g5480 ( 
.A(n_3920),
.Y(n_5480)
);

CKINVDCx5p33_ASAP7_75t_R g5481 ( 
.A(n_3950),
.Y(n_5481)
);

CKINVDCx5p33_ASAP7_75t_R g5482 ( 
.A(n_2261),
.Y(n_5482)
);

CKINVDCx5p33_ASAP7_75t_R g5483 ( 
.A(n_3875),
.Y(n_5483)
);

CKINVDCx20_ASAP7_75t_R g5484 ( 
.A(n_11),
.Y(n_5484)
);

INVx1_ASAP7_75t_L g5485 ( 
.A(n_558),
.Y(n_5485)
);

INVx1_ASAP7_75t_L g5486 ( 
.A(n_78),
.Y(n_5486)
);

INVx1_ASAP7_75t_L g5487 ( 
.A(n_3343),
.Y(n_5487)
);

INVx2_ASAP7_75t_SL g5488 ( 
.A(n_203),
.Y(n_5488)
);

INVx1_ASAP7_75t_L g5489 ( 
.A(n_4034),
.Y(n_5489)
);

INVx2_ASAP7_75t_L g5490 ( 
.A(n_576),
.Y(n_5490)
);

INVx1_ASAP7_75t_L g5491 ( 
.A(n_3598),
.Y(n_5491)
);

CKINVDCx5p33_ASAP7_75t_R g5492 ( 
.A(n_1805),
.Y(n_5492)
);

CKINVDCx5p33_ASAP7_75t_R g5493 ( 
.A(n_2045),
.Y(n_5493)
);

INVx1_ASAP7_75t_L g5494 ( 
.A(n_942),
.Y(n_5494)
);

CKINVDCx5p33_ASAP7_75t_R g5495 ( 
.A(n_3104),
.Y(n_5495)
);

INVx2_ASAP7_75t_L g5496 ( 
.A(n_1138),
.Y(n_5496)
);

CKINVDCx20_ASAP7_75t_R g5497 ( 
.A(n_1301),
.Y(n_5497)
);

CKINVDCx5p33_ASAP7_75t_R g5498 ( 
.A(n_3262),
.Y(n_5498)
);

CKINVDCx5p33_ASAP7_75t_R g5499 ( 
.A(n_3874),
.Y(n_5499)
);

INVx1_ASAP7_75t_L g5500 ( 
.A(n_3542),
.Y(n_5500)
);

INVx2_ASAP7_75t_L g5501 ( 
.A(n_3938),
.Y(n_5501)
);

INVx1_ASAP7_75t_SL g5502 ( 
.A(n_3568),
.Y(n_5502)
);

CKINVDCx16_ASAP7_75t_R g5503 ( 
.A(n_1942),
.Y(n_5503)
);

CKINVDCx5p33_ASAP7_75t_R g5504 ( 
.A(n_373),
.Y(n_5504)
);

INVx1_ASAP7_75t_L g5505 ( 
.A(n_4012),
.Y(n_5505)
);

CKINVDCx20_ASAP7_75t_R g5506 ( 
.A(n_3965),
.Y(n_5506)
);

CKINVDCx5p33_ASAP7_75t_R g5507 ( 
.A(n_2463),
.Y(n_5507)
);

CKINVDCx5p33_ASAP7_75t_R g5508 ( 
.A(n_2604),
.Y(n_5508)
);

BUFx10_ASAP7_75t_L g5509 ( 
.A(n_766),
.Y(n_5509)
);

INVx1_ASAP7_75t_SL g5510 ( 
.A(n_1417),
.Y(n_5510)
);

CKINVDCx5p33_ASAP7_75t_R g5511 ( 
.A(n_122),
.Y(n_5511)
);

CKINVDCx5p33_ASAP7_75t_R g5512 ( 
.A(n_362),
.Y(n_5512)
);

CKINVDCx5p33_ASAP7_75t_R g5513 ( 
.A(n_3772),
.Y(n_5513)
);

INVx1_ASAP7_75t_L g5514 ( 
.A(n_1335),
.Y(n_5514)
);

CKINVDCx5p33_ASAP7_75t_R g5515 ( 
.A(n_3865),
.Y(n_5515)
);

INVx1_ASAP7_75t_L g5516 ( 
.A(n_4013),
.Y(n_5516)
);

BUFx6f_ASAP7_75t_L g5517 ( 
.A(n_431),
.Y(n_5517)
);

INVx1_ASAP7_75t_L g5518 ( 
.A(n_768),
.Y(n_5518)
);

CKINVDCx5p33_ASAP7_75t_R g5519 ( 
.A(n_3472),
.Y(n_5519)
);

CKINVDCx16_ASAP7_75t_R g5520 ( 
.A(n_79),
.Y(n_5520)
);

INVx1_ASAP7_75t_L g5521 ( 
.A(n_2411),
.Y(n_5521)
);

CKINVDCx5p33_ASAP7_75t_R g5522 ( 
.A(n_198),
.Y(n_5522)
);

CKINVDCx5p33_ASAP7_75t_R g5523 ( 
.A(n_2040),
.Y(n_5523)
);

INVx1_ASAP7_75t_L g5524 ( 
.A(n_641),
.Y(n_5524)
);

INVx1_ASAP7_75t_L g5525 ( 
.A(n_4171),
.Y(n_5525)
);

NAND2xp5_ASAP7_75t_L g5526 ( 
.A(n_4132),
.B(n_0),
.Y(n_5526)
);

INVx1_ASAP7_75t_L g5527 ( 
.A(n_4171),
.Y(n_5527)
);

INVx1_ASAP7_75t_L g5528 ( 
.A(n_4171),
.Y(n_5528)
);

INVx1_ASAP7_75t_L g5529 ( 
.A(n_4171),
.Y(n_5529)
);

INVx1_ASAP7_75t_L g5530 ( 
.A(n_4171),
.Y(n_5530)
);

CKINVDCx5p33_ASAP7_75t_R g5531 ( 
.A(n_5414),
.Y(n_5531)
);

NOR2xp67_ASAP7_75t_L g5532 ( 
.A(n_4256),
.B(n_0),
.Y(n_5532)
);

BUFx3_ASAP7_75t_L g5533 ( 
.A(n_4397),
.Y(n_5533)
);

INVx1_ASAP7_75t_L g5534 ( 
.A(n_4221),
.Y(n_5534)
);

BUFx6f_ASAP7_75t_L g5535 ( 
.A(n_4625),
.Y(n_5535)
);

INVx1_ASAP7_75t_L g5536 ( 
.A(n_4221),
.Y(n_5536)
);

CKINVDCx5p33_ASAP7_75t_R g5537 ( 
.A(n_4126),
.Y(n_5537)
);

CKINVDCx5p33_ASAP7_75t_R g5538 ( 
.A(n_4227),
.Y(n_5538)
);

INVx1_ASAP7_75t_L g5539 ( 
.A(n_4221),
.Y(n_5539)
);

CKINVDCx5p33_ASAP7_75t_R g5540 ( 
.A(n_4522),
.Y(n_5540)
);

INVx1_ASAP7_75t_L g5541 ( 
.A(n_4221),
.Y(n_5541)
);

INVx1_ASAP7_75t_L g5542 ( 
.A(n_4221),
.Y(n_5542)
);

CKINVDCx20_ASAP7_75t_R g5543 ( 
.A(n_4478),
.Y(n_5543)
);

HB1xp67_ASAP7_75t_L g5544 ( 
.A(n_5520),
.Y(n_5544)
);

CKINVDCx5p33_ASAP7_75t_R g5545 ( 
.A(n_4571),
.Y(n_5545)
);

INVxp67_ASAP7_75t_L g5546 ( 
.A(n_4301),
.Y(n_5546)
);

INVx1_ASAP7_75t_L g5547 ( 
.A(n_4485),
.Y(n_5547)
);

INVx1_ASAP7_75t_SL g5548 ( 
.A(n_5032),
.Y(n_5548)
);

CKINVDCx16_ASAP7_75t_R g5549 ( 
.A(n_4115),
.Y(n_5549)
);

INVx1_ASAP7_75t_SL g5550 ( 
.A(n_4119),
.Y(n_5550)
);

CKINVDCx5p33_ASAP7_75t_R g5551 ( 
.A(n_5225),
.Y(n_5551)
);

CKINVDCx20_ASAP7_75t_R g5552 ( 
.A(n_4613),
.Y(n_5552)
);

INVx1_ASAP7_75t_L g5553 ( 
.A(n_4485),
.Y(n_5553)
);

CKINVDCx5p33_ASAP7_75t_R g5554 ( 
.A(n_5332),
.Y(n_5554)
);

CKINVDCx5p33_ASAP7_75t_R g5555 ( 
.A(n_5459),
.Y(n_5555)
);

CKINVDCx5p33_ASAP7_75t_R g5556 ( 
.A(n_4960),
.Y(n_5556)
);

INVx1_ASAP7_75t_L g5557 ( 
.A(n_4485),
.Y(n_5557)
);

CKINVDCx5p33_ASAP7_75t_R g5558 ( 
.A(n_5010),
.Y(n_5558)
);

CKINVDCx5p33_ASAP7_75t_R g5559 ( 
.A(n_5199),
.Y(n_5559)
);

CKINVDCx5p33_ASAP7_75t_R g5560 ( 
.A(n_5238),
.Y(n_5560)
);

INVx2_ASAP7_75t_L g5561 ( 
.A(n_4485),
.Y(n_5561)
);

CKINVDCx5p33_ASAP7_75t_R g5562 ( 
.A(n_4167),
.Y(n_5562)
);

OR2x2_ASAP7_75t_L g5563 ( 
.A(n_4710),
.B(n_0),
.Y(n_5563)
);

INVx1_ASAP7_75t_SL g5564 ( 
.A(n_4233),
.Y(n_5564)
);

BUFx2_ASAP7_75t_L g5565 ( 
.A(n_4277),
.Y(n_5565)
);

CKINVDCx5p33_ASAP7_75t_R g5566 ( 
.A(n_4206),
.Y(n_5566)
);

CKINVDCx5p33_ASAP7_75t_R g5567 ( 
.A(n_4283),
.Y(n_5567)
);

INVx1_ASAP7_75t_L g5568 ( 
.A(n_4485),
.Y(n_5568)
);

CKINVDCx5p33_ASAP7_75t_R g5569 ( 
.A(n_4483),
.Y(n_5569)
);

CKINVDCx5p33_ASAP7_75t_R g5570 ( 
.A(n_4559),
.Y(n_5570)
);

BUFx3_ASAP7_75t_L g5571 ( 
.A(n_4425),
.Y(n_5571)
);

INVx1_ASAP7_75t_L g5572 ( 
.A(n_4488),
.Y(n_5572)
);

INVx2_ASAP7_75t_SL g5573 ( 
.A(n_4318),
.Y(n_5573)
);

CKINVDCx5p33_ASAP7_75t_R g5574 ( 
.A(n_4682),
.Y(n_5574)
);

CKINVDCx5p33_ASAP7_75t_R g5575 ( 
.A(n_4690),
.Y(n_5575)
);

INVx1_ASAP7_75t_L g5576 ( 
.A(n_4488),
.Y(n_5576)
);

INVx1_ASAP7_75t_L g5577 ( 
.A(n_4488),
.Y(n_5577)
);

CKINVDCx5p33_ASAP7_75t_R g5578 ( 
.A(n_4798),
.Y(n_5578)
);

CKINVDCx5p33_ASAP7_75t_R g5579 ( 
.A(n_4833),
.Y(n_5579)
);

CKINVDCx5p33_ASAP7_75t_R g5580 ( 
.A(n_4856),
.Y(n_5580)
);

INVx1_ASAP7_75t_L g5581 ( 
.A(n_4488),
.Y(n_5581)
);

BUFx2_ASAP7_75t_L g5582 ( 
.A(n_4297),
.Y(n_5582)
);

BUFx10_ASAP7_75t_L g5583 ( 
.A(n_4235),
.Y(n_5583)
);

INVx1_ASAP7_75t_L g5584 ( 
.A(n_4488),
.Y(n_5584)
);

CKINVDCx5p33_ASAP7_75t_R g5585 ( 
.A(n_4892),
.Y(n_5585)
);

INVx2_ASAP7_75t_L g5586 ( 
.A(n_4611),
.Y(n_5586)
);

CKINVDCx5p33_ASAP7_75t_R g5587 ( 
.A(n_4932),
.Y(n_5587)
);

CKINVDCx20_ASAP7_75t_R g5588 ( 
.A(n_4976),
.Y(n_5588)
);

OR2x2_ASAP7_75t_L g5589 ( 
.A(n_4389),
.B(n_1),
.Y(n_5589)
);

CKINVDCx20_ASAP7_75t_R g5590 ( 
.A(n_5042),
.Y(n_5590)
);

INVx1_ASAP7_75t_L g5591 ( 
.A(n_4611),
.Y(n_5591)
);

INVx1_ASAP7_75t_L g5592 ( 
.A(n_4611),
.Y(n_5592)
);

INVx1_ASAP7_75t_L g5593 ( 
.A(n_4611),
.Y(n_5593)
);

INVx1_ASAP7_75t_SL g5594 ( 
.A(n_4429),
.Y(n_5594)
);

INVx1_ASAP7_75t_L g5595 ( 
.A(n_4611),
.Y(n_5595)
);

INVx1_ASAP7_75t_L g5596 ( 
.A(n_4836),
.Y(n_5596)
);

NOR2xp67_ASAP7_75t_L g5597 ( 
.A(n_4256),
.B(n_1),
.Y(n_5597)
);

INVx1_ASAP7_75t_L g5598 ( 
.A(n_4836),
.Y(n_5598)
);

INVx2_ASAP7_75t_SL g5599 ( 
.A(n_4318),
.Y(n_5599)
);

INVx1_ASAP7_75t_L g5600 ( 
.A(n_4836),
.Y(n_5600)
);

INVx1_ASAP7_75t_L g5601 ( 
.A(n_4836),
.Y(n_5601)
);

CKINVDCx5p33_ASAP7_75t_R g5602 ( 
.A(n_5067),
.Y(n_5602)
);

INVx1_ASAP7_75t_L g5603 ( 
.A(n_4836),
.Y(n_5603)
);

INVx1_ASAP7_75t_L g5604 ( 
.A(n_4891),
.Y(n_5604)
);

INVx1_ASAP7_75t_L g5605 ( 
.A(n_4891),
.Y(n_5605)
);

INVx2_ASAP7_75t_L g5606 ( 
.A(n_4891),
.Y(n_5606)
);

CKINVDCx5p33_ASAP7_75t_R g5607 ( 
.A(n_5071),
.Y(n_5607)
);

INVx2_ASAP7_75t_L g5608 ( 
.A(n_4891),
.Y(n_5608)
);

CKINVDCx16_ASAP7_75t_R g5609 ( 
.A(n_5187),
.Y(n_5609)
);

CKINVDCx5p33_ASAP7_75t_R g5610 ( 
.A(n_5352),
.Y(n_5610)
);

INVx1_ASAP7_75t_L g5611 ( 
.A(n_4891),
.Y(n_5611)
);

INVx1_ASAP7_75t_L g5612 ( 
.A(n_4922),
.Y(n_5612)
);

CKINVDCx5p33_ASAP7_75t_R g5613 ( 
.A(n_5457),
.Y(n_5613)
);

BUFx6f_ASAP7_75t_L g5614 ( 
.A(n_4625),
.Y(n_5614)
);

INVx1_ASAP7_75t_L g5615 ( 
.A(n_4922),
.Y(n_5615)
);

INVx2_ASAP7_75t_SL g5616 ( 
.A(n_4974),
.Y(n_5616)
);

CKINVDCx20_ASAP7_75t_R g5617 ( 
.A(n_5475),
.Y(n_5617)
);

INVx1_ASAP7_75t_L g5618 ( 
.A(n_4922),
.Y(n_5618)
);

CKINVDCx5p33_ASAP7_75t_R g5619 ( 
.A(n_5503),
.Y(n_5619)
);

CKINVDCx5p33_ASAP7_75t_R g5620 ( 
.A(n_4243),
.Y(n_5620)
);

CKINVDCx5p33_ASAP7_75t_R g5621 ( 
.A(n_4244),
.Y(n_5621)
);

INVx2_ASAP7_75t_L g5622 ( 
.A(n_4922),
.Y(n_5622)
);

INVx1_ASAP7_75t_L g5623 ( 
.A(n_4922),
.Y(n_5623)
);

CKINVDCx5p33_ASAP7_75t_R g5624 ( 
.A(n_4263),
.Y(n_5624)
);

CKINVDCx5p33_ASAP7_75t_R g5625 ( 
.A(n_4265),
.Y(n_5625)
);

INVx1_ASAP7_75t_SL g5626 ( 
.A(n_4466),
.Y(n_5626)
);

INVx1_ASAP7_75t_L g5627 ( 
.A(n_5408),
.Y(n_5627)
);

CKINVDCx5p33_ASAP7_75t_R g5628 ( 
.A(n_4281),
.Y(n_5628)
);

INVx1_ASAP7_75t_L g5629 ( 
.A(n_5408),
.Y(n_5629)
);

INVx1_ASAP7_75t_L g5630 ( 
.A(n_5408),
.Y(n_5630)
);

CKINVDCx5p33_ASAP7_75t_R g5631 ( 
.A(n_4345),
.Y(n_5631)
);

INVx1_ASAP7_75t_L g5632 ( 
.A(n_5408),
.Y(n_5632)
);

INVx2_ASAP7_75t_L g5633 ( 
.A(n_5408),
.Y(n_5633)
);

CKINVDCx16_ASAP7_75t_R g5634 ( 
.A(n_4588),
.Y(n_5634)
);

CKINVDCx5p33_ASAP7_75t_R g5635 ( 
.A(n_4370),
.Y(n_5635)
);

INVx2_ASAP7_75t_L g5636 ( 
.A(n_4130),
.Y(n_5636)
);

INVx1_ASAP7_75t_L g5637 ( 
.A(n_4163),
.Y(n_5637)
);

CKINVDCx5p33_ASAP7_75t_R g5638 ( 
.A(n_4410),
.Y(n_5638)
);

CKINVDCx5p33_ASAP7_75t_R g5639 ( 
.A(n_4462),
.Y(n_5639)
);

INVx1_ASAP7_75t_L g5640 ( 
.A(n_4213),
.Y(n_5640)
);

CKINVDCx5p33_ASAP7_75t_R g5641 ( 
.A(n_4502),
.Y(n_5641)
);

CKINVDCx5p33_ASAP7_75t_R g5642 ( 
.A(n_4527),
.Y(n_5642)
);

CKINVDCx5p33_ASAP7_75t_R g5643 ( 
.A(n_4543),
.Y(n_5643)
);

CKINVDCx20_ASAP7_75t_R g5644 ( 
.A(n_4100),
.Y(n_5644)
);

INVx2_ASAP7_75t_L g5645 ( 
.A(n_4266),
.Y(n_5645)
);

CKINVDCx5p33_ASAP7_75t_R g5646 ( 
.A(n_4546),
.Y(n_5646)
);

CKINVDCx16_ASAP7_75t_R g5647 ( 
.A(n_5143),
.Y(n_5647)
);

INVxp67_ASAP7_75t_L g5648 ( 
.A(n_4495),
.Y(n_5648)
);

CKINVDCx5p33_ASAP7_75t_R g5649 ( 
.A(n_4596),
.Y(n_5649)
);

INVx1_ASAP7_75t_L g5650 ( 
.A(n_4284),
.Y(n_5650)
);

CKINVDCx5p33_ASAP7_75t_R g5651 ( 
.A(n_4668),
.Y(n_5651)
);

CKINVDCx5p33_ASAP7_75t_R g5652 ( 
.A(n_4683),
.Y(n_5652)
);

CKINVDCx16_ASAP7_75t_R g5653 ( 
.A(n_4974),
.Y(n_5653)
);

INVx1_ASAP7_75t_L g5654 ( 
.A(n_4300),
.Y(n_5654)
);

HB1xp67_ASAP7_75t_L g5655 ( 
.A(n_4174),
.Y(n_5655)
);

CKINVDCx20_ASAP7_75t_R g5656 ( 
.A(n_4108),
.Y(n_5656)
);

BUFx6f_ASAP7_75t_L g5657 ( 
.A(n_4625),
.Y(n_5657)
);

INVx1_ASAP7_75t_L g5658 ( 
.A(n_4326),
.Y(n_5658)
);

BUFx5_ASAP7_75t_L g5659 ( 
.A(n_4097),
.Y(n_5659)
);

BUFx5_ASAP7_75t_L g5660 ( 
.A(n_4098),
.Y(n_5660)
);

BUFx10_ASAP7_75t_L g5661 ( 
.A(n_4997),
.Y(n_5661)
);

INVx1_ASAP7_75t_L g5662 ( 
.A(n_4413),
.Y(n_5662)
);

INVx1_ASAP7_75t_L g5663 ( 
.A(n_4551),
.Y(n_5663)
);

CKINVDCx20_ASAP7_75t_R g5664 ( 
.A(n_4120),
.Y(n_5664)
);

INVx1_ASAP7_75t_L g5665 ( 
.A(n_4557),
.Y(n_5665)
);

INVx1_ASAP7_75t_L g5666 ( 
.A(n_4643),
.Y(n_5666)
);

CKINVDCx16_ASAP7_75t_R g5667 ( 
.A(n_5098),
.Y(n_5667)
);

CKINVDCx5p33_ASAP7_75t_R g5668 ( 
.A(n_4702),
.Y(n_5668)
);

CKINVDCx5p33_ASAP7_75t_R g5669 ( 
.A(n_4726),
.Y(n_5669)
);

CKINVDCx5p33_ASAP7_75t_R g5670 ( 
.A(n_4732),
.Y(n_5670)
);

INVx1_ASAP7_75t_L g5671 ( 
.A(n_4715),
.Y(n_5671)
);

CKINVDCx5p33_ASAP7_75t_R g5672 ( 
.A(n_4783),
.Y(n_5672)
);

CKINVDCx5p33_ASAP7_75t_R g5673 ( 
.A(n_4790),
.Y(n_5673)
);

INVx1_ASAP7_75t_L g5674 ( 
.A(n_4773),
.Y(n_5674)
);

CKINVDCx5p33_ASAP7_75t_R g5675 ( 
.A(n_4847),
.Y(n_5675)
);

CKINVDCx16_ASAP7_75t_R g5676 ( 
.A(n_5098),
.Y(n_5676)
);

INVx1_ASAP7_75t_L g5677 ( 
.A(n_4849),
.Y(n_5677)
);

INVx1_ASAP7_75t_L g5678 ( 
.A(n_4879),
.Y(n_5678)
);

INVx1_ASAP7_75t_L g5679 ( 
.A(n_4910),
.Y(n_5679)
);

CKINVDCx20_ASAP7_75t_R g5680 ( 
.A(n_4150),
.Y(n_5680)
);

BUFx2_ASAP7_75t_L g5681 ( 
.A(n_4667),
.Y(n_5681)
);

INVx1_ASAP7_75t_L g5682 ( 
.A(n_4943),
.Y(n_5682)
);

INVx1_ASAP7_75t_L g5683 ( 
.A(n_4950),
.Y(n_5683)
);

CKINVDCx5p33_ASAP7_75t_R g5684 ( 
.A(n_4877),
.Y(n_5684)
);

INVx1_ASAP7_75t_L g5685 ( 
.A(n_4989),
.Y(n_5685)
);

INVx1_ASAP7_75t_L g5686 ( 
.A(n_5045),
.Y(n_5686)
);

CKINVDCx5p33_ASAP7_75t_R g5687 ( 
.A(n_4883),
.Y(n_5687)
);

CKINVDCx5p33_ASAP7_75t_R g5688 ( 
.A(n_4911),
.Y(n_5688)
);

INVx2_ASAP7_75t_L g5689 ( 
.A(n_5088),
.Y(n_5689)
);

INVx2_ASAP7_75t_L g5690 ( 
.A(n_5131),
.Y(n_5690)
);

INVx1_ASAP7_75t_L g5691 ( 
.A(n_5163),
.Y(n_5691)
);

CKINVDCx16_ASAP7_75t_R g5692 ( 
.A(n_4254),
.Y(n_5692)
);

OR2x2_ASAP7_75t_L g5693 ( 
.A(n_4692),
.B(n_2),
.Y(n_5693)
);

CKINVDCx5p33_ASAP7_75t_R g5694 ( 
.A(n_4955),
.Y(n_5694)
);

CKINVDCx5p33_ASAP7_75t_R g5695 ( 
.A(n_4995),
.Y(n_5695)
);

CKINVDCx5p33_ASAP7_75t_R g5696 ( 
.A(n_5030),
.Y(n_5696)
);

INVx1_ASAP7_75t_L g5697 ( 
.A(n_5205),
.Y(n_5697)
);

CKINVDCx20_ASAP7_75t_R g5698 ( 
.A(n_4151),
.Y(n_5698)
);

NOR2xp67_ASAP7_75t_L g5699 ( 
.A(n_4431),
.B(n_2),
.Y(n_5699)
);

CKINVDCx5p33_ASAP7_75t_R g5700 ( 
.A(n_5126),
.Y(n_5700)
);

INVx1_ASAP7_75t_L g5701 ( 
.A(n_5333),
.Y(n_5701)
);

INVxp33_ASAP7_75t_R g5702 ( 
.A(n_4254),
.Y(n_5702)
);

INVx1_ASAP7_75t_L g5703 ( 
.A(n_5339),
.Y(n_5703)
);

BUFx5_ASAP7_75t_L g5704 ( 
.A(n_4103),
.Y(n_5704)
);

CKINVDCx5p33_ASAP7_75t_R g5705 ( 
.A(n_5141),
.Y(n_5705)
);

INVx1_ASAP7_75t_L g5706 ( 
.A(n_5400),
.Y(n_5706)
);

INVx1_ASAP7_75t_L g5707 ( 
.A(n_5423),
.Y(n_5707)
);

CKINVDCx20_ASAP7_75t_R g5708 ( 
.A(n_4177),
.Y(n_5708)
);

INVx1_ASAP7_75t_L g5709 ( 
.A(n_5436),
.Y(n_5709)
);

INVx1_ASAP7_75t_L g5710 ( 
.A(n_5477),
.Y(n_5710)
);

INVx1_ASAP7_75t_L g5711 ( 
.A(n_5486),
.Y(n_5711)
);

INVx1_ASAP7_75t_L g5712 ( 
.A(n_4468),
.Y(n_5712)
);

CKINVDCx5p33_ASAP7_75t_R g5713 ( 
.A(n_5148),
.Y(n_5713)
);

CKINVDCx5p33_ASAP7_75t_R g5714 ( 
.A(n_5228),
.Y(n_5714)
);

CKINVDCx5p33_ASAP7_75t_R g5715 ( 
.A(n_5235),
.Y(n_5715)
);

CKINVDCx5p33_ASAP7_75t_R g5716 ( 
.A(n_5271),
.Y(n_5716)
);

CKINVDCx5p33_ASAP7_75t_R g5717 ( 
.A(n_5305),
.Y(n_5717)
);

INVx1_ASAP7_75t_L g5718 ( 
.A(n_4561),
.Y(n_5718)
);

INVx1_ASAP7_75t_L g5719 ( 
.A(n_4754),
.Y(n_5719)
);

CKINVDCx5p33_ASAP7_75t_R g5720 ( 
.A(n_5315),
.Y(n_5720)
);

INVx1_ASAP7_75t_L g5721 ( 
.A(n_4993),
.Y(n_5721)
);

CKINVDCx5p33_ASAP7_75t_R g5722 ( 
.A(n_5320),
.Y(n_5722)
);

NOR2xp67_ASAP7_75t_L g5723 ( 
.A(n_4431),
.B(n_2),
.Y(n_5723)
);

CKINVDCx5p33_ASAP7_75t_R g5724 ( 
.A(n_5338),
.Y(n_5724)
);

NOR2xp67_ASAP7_75t_L g5725 ( 
.A(n_4270),
.B(n_3),
.Y(n_5725)
);

CKINVDCx5p33_ASAP7_75t_R g5726 ( 
.A(n_5364),
.Y(n_5726)
);

INVx2_ASAP7_75t_SL g5727 ( 
.A(n_4287),
.Y(n_5727)
);

INVx1_ASAP7_75t_L g5728 ( 
.A(n_4942),
.Y(n_5728)
);

CKINVDCx5p33_ASAP7_75t_R g5729 ( 
.A(n_5399),
.Y(n_5729)
);

INVx1_ASAP7_75t_L g5730 ( 
.A(n_4942),
.Y(n_5730)
);

INVx1_ASAP7_75t_SL g5731 ( 
.A(n_4748),
.Y(n_5731)
);

INVx1_ASAP7_75t_L g5732 ( 
.A(n_4942),
.Y(n_5732)
);

NOR2xp33_ASAP7_75t_L g5733 ( 
.A(n_4699),
.B(n_5019),
.Y(n_5733)
);

INVx2_ASAP7_75t_L g5734 ( 
.A(n_4107),
.Y(n_5734)
);

INVx1_ASAP7_75t_L g5735 ( 
.A(n_4865),
.Y(n_5735)
);

CKINVDCx5p33_ASAP7_75t_R g5736 ( 
.A(n_5466),
.Y(n_5736)
);

CKINVDCx5p33_ASAP7_75t_R g5737 ( 
.A(n_5511),
.Y(n_5737)
);

CKINVDCx5p33_ASAP7_75t_R g5738 ( 
.A(n_5522),
.Y(n_5738)
);

CKINVDCx5p33_ASAP7_75t_R g5739 ( 
.A(n_5512),
.Y(n_5739)
);

INVx2_ASAP7_75t_L g5740 ( 
.A(n_5015),
.Y(n_5740)
);

BUFx3_ASAP7_75t_L g5741 ( 
.A(n_4116),
.Y(n_5741)
);

BUFx2_ASAP7_75t_SL g5742 ( 
.A(n_4191),
.Y(n_5742)
);

INVx1_ASAP7_75t_L g5743 ( 
.A(n_4101),
.Y(n_5743)
);

INVx1_ASAP7_75t_L g5744 ( 
.A(n_4101),
.Y(n_5744)
);

NOR2xp67_ASAP7_75t_L g5745 ( 
.A(n_4338),
.B(n_3),
.Y(n_5745)
);

CKINVDCx5p33_ASAP7_75t_R g5746 ( 
.A(n_5519),
.Y(n_5746)
);

CKINVDCx5p33_ASAP7_75t_R g5747 ( 
.A(n_5523),
.Y(n_5747)
);

CKINVDCx5p33_ASAP7_75t_R g5748 ( 
.A(n_4099),
.Y(n_5748)
);

CKINVDCx20_ASAP7_75t_R g5749 ( 
.A(n_4209),
.Y(n_5749)
);

INVx1_ASAP7_75t_SL g5750 ( 
.A(n_5101),
.Y(n_5750)
);

CKINVDCx5p33_ASAP7_75t_R g5751 ( 
.A(n_4102),
.Y(n_5751)
);

CKINVDCx5p33_ASAP7_75t_R g5752 ( 
.A(n_4104),
.Y(n_5752)
);

CKINVDCx5p33_ASAP7_75t_R g5753 ( 
.A(n_4105),
.Y(n_5753)
);

CKINVDCx5p33_ASAP7_75t_R g5754 ( 
.A(n_5504),
.Y(n_5754)
);

INVx1_ASAP7_75t_L g5755 ( 
.A(n_4101),
.Y(n_5755)
);

INVx2_ASAP7_75t_L g5756 ( 
.A(n_5517),
.Y(n_5756)
);

INVx1_ASAP7_75t_L g5757 ( 
.A(n_4109),
.Y(n_5757)
);

INVx1_ASAP7_75t_L g5758 ( 
.A(n_4109),
.Y(n_5758)
);

CKINVDCx5p33_ASAP7_75t_R g5759 ( 
.A(n_5507),
.Y(n_5759)
);

INVx1_ASAP7_75t_L g5760 ( 
.A(n_4109),
.Y(n_5760)
);

CKINVDCx5p33_ASAP7_75t_R g5761 ( 
.A(n_5508),
.Y(n_5761)
);

CKINVDCx16_ASAP7_75t_R g5762 ( 
.A(n_5509),
.Y(n_5762)
);

CKINVDCx5p33_ASAP7_75t_R g5763 ( 
.A(n_5513),
.Y(n_5763)
);

CKINVDCx5p33_ASAP7_75t_R g5764 ( 
.A(n_5515),
.Y(n_5764)
);

CKINVDCx5p33_ASAP7_75t_R g5765 ( 
.A(n_4106),
.Y(n_5765)
);

CKINVDCx20_ASAP7_75t_R g5766 ( 
.A(n_4249),
.Y(n_5766)
);

INVx2_ASAP7_75t_L g5767 ( 
.A(n_5517),
.Y(n_5767)
);

INVx1_ASAP7_75t_L g5768 ( 
.A(n_4181),
.Y(n_5768)
);

INVxp67_ASAP7_75t_SL g5769 ( 
.A(n_4188),
.Y(n_5769)
);

CKINVDCx5p33_ASAP7_75t_R g5770 ( 
.A(n_4110),
.Y(n_5770)
);

NOR2xp33_ASAP7_75t_L g5771 ( 
.A(n_5214),
.B(n_3),
.Y(n_5771)
);

CKINVDCx5p33_ASAP7_75t_R g5772 ( 
.A(n_4111),
.Y(n_5772)
);

INVx1_ASAP7_75t_L g5773 ( 
.A(n_4181),
.Y(n_5773)
);

BUFx5_ASAP7_75t_L g5774 ( 
.A(n_4114),
.Y(n_5774)
);

INVx1_ASAP7_75t_L g5775 ( 
.A(n_4181),
.Y(n_5775)
);

CKINVDCx5p33_ASAP7_75t_R g5776 ( 
.A(n_4112),
.Y(n_5776)
);

INVx1_ASAP7_75t_L g5777 ( 
.A(n_4198),
.Y(n_5777)
);

INVx1_ASAP7_75t_SL g5778 ( 
.A(n_5221),
.Y(n_5778)
);

INVx1_ASAP7_75t_L g5779 ( 
.A(n_4198),
.Y(n_5779)
);

CKINVDCx5p33_ASAP7_75t_R g5780 ( 
.A(n_5499),
.Y(n_5780)
);

INVx1_ASAP7_75t_L g5781 ( 
.A(n_4198),
.Y(n_5781)
);

CKINVDCx20_ASAP7_75t_R g5782 ( 
.A(n_4257),
.Y(n_5782)
);

BUFx3_ASAP7_75t_L g5783 ( 
.A(n_4133),
.Y(n_5783)
);

INVx1_ASAP7_75t_L g5784 ( 
.A(n_4199),
.Y(n_5784)
);

INVx1_ASAP7_75t_L g5785 ( 
.A(n_4199),
.Y(n_5785)
);

CKINVDCx5p33_ASAP7_75t_R g5786 ( 
.A(n_4113),
.Y(n_5786)
);

INVx1_ASAP7_75t_L g5787 ( 
.A(n_4199),
.Y(n_5787)
);

BUFx5_ASAP7_75t_L g5788 ( 
.A(n_4117),
.Y(n_5788)
);

NOR2xp67_ASAP7_75t_L g5789 ( 
.A(n_4500),
.B(n_4),
.Y(n_5789)
);

CKINVDCx20_ASAP7_75t_R g5790 ( 
.A(n_4280),
.Y(n_5790)
);

CKINVDCx5p33_ASAP7_75t_R g5791 ( 
.A(n_4118),
.Y(n_5791)
);

CKINVDCx5p33_ASAP7_75t_R g5792 ( 
.A(n_4124),
.Y(n_5792)
);

NOR2xp67_ASAP7_75t_L g5793 ( 
.A(n_4553),
.B(n_4),
.Y(n_5793)
);

INVx1_ASAP7_75t_L g5794 ( 
.A(n_4237),
.Y(n_5794)
);

INVx2_ASAP7_75t_L g5795 ( 
.A(n_4237),
.Y(n_5795)
);

INVx2_ASAP7_75t_L g5796 ( 
.A(n_4237),
.Y(n_5796)
);

CKINVDCx14_ASAP7_75t_R g5797 ( 
.A(n_5297),
.Y(n_5797)
);

HB1xp67_ASAP7_75t_L g5798 ( 
.A(n_4269),
.Y(n_5798)
);

INVx1_ASAP7_75t_L g5799 ( 
.A(n_4250),
.Y(n_5799)
);

BUFx2_ASAP7_75t_L g5800 ( 
.A(n_5301),
.Y(n_5800)
);

INVx1_ASAP7_75t_L g5801 ( 
.A(n_4250),
.Y(n_5801)
);

XOR2xp5_ASAP7_75t_L g5802 ( 
.A(n_4313),
.B(n_4),
.Y(n_5802)
);

CKINVDCx5p33_ASAP7_75t_R g5803 ( 
.A(n_4125),
.Y(n_5803)
);

INVx1_ASAP7_75t_L g5804 ( 
.A(n_4250),
.Y(n_5804)
);

CKINVDCx20_ASAP7_75t_R g5805 ( 
.A(n_4320),
.Y(n_5805)
);

BUFx3_ASAP7_75t_L g5806 ( 
.A(n_4158),
.Y(n_5806)
);

BUFx3_ASAP7_75t_L g5807 ( 
.A(n_4241),
.Y(n_5807)
);

INVx1_ASAP7_75t_L g5808 ( 
.A(n_4251),
.Y(n_5808)
);

CKINVDCx5p33_ASAP7_75t_R g5809 ( 
.A(n_4131),
.Y(n_5809)
);

INVx2_ASAP7_75t_L g5810 ( 
.A(n_5517),
.Y(n_5810)
);

CKINVDCx5p33_ASAP7_75t_R g5811 ( 
.A(n_4137),
.Y(n_5811)
);

CKINVDCx20_ASAP7_75t_R g5812 ( 
.A(n_4348),
.Y(n_5812)
);

INVx1_ASAP7_75t_L g5813 ( 
.A(n_4251),
.Y(n_5813)
);

CKINVDCx5p33_ASAP7_75t_R g5814 ( 
.A(n_4139),
.Y(n_5814)
);

INVx1_ASAP7_75t_L g5815 ( 
.A(n_4251),
.Y(n_5815)
);

INVx1_ASAP7_75t_L g5816 ( 
.A(n_4299),
.Y(n_5816)
);

INVx1_ASAP7_75t_L g5817 ( 
.A(n_4299),
.Y(n_5817)
);

INVx1_ASAP7_75t_L g5818 ( 
.A(n_4299),
.Y(n_5818)
);

CKINVDCx5p33_ASAP7_75t_R g5819 ( 
.A(n_4141),
.Y(n_5819)
);

INVx1_ASAP7_75t_L g5820 ( 
.A(n_4347),
.Y(n_5820)
);

INVx1_ASAP7_75t_L g5821 ( 
.A(n_4347),
.Y(n_5821)
);

INVx2_ASAP7_75t_L g5822 ( 
.A(n_4347),
.Y(n_5822)
);

INVx2_ASAP7_75t_L g5823 ( 
.A(n_4366),
.Y(n_5823)
);

CKINVDCx5p33_ASAP7_75t_R g5824 ( 
.A(n_5498),
.Y(n_5824)
);

INVx1_ASAP7_75t_L g5825 ( 
.A(n_4366),
.Y(n_5825)
);

CKINVDCx5p33_ASAP7_75t_R g5826 ( 
.A(n_4142),
.Y(n_5826)
);

BUFx5_ASAP7_75t_L g5827 ( 
.A(n_4121),
.Y(n_5827)
);

CKINVDCx5p33_ASAP7_75t_R g5828 ( 
.A(n_4143),
.Y(n_5828)
);

HB1xp67_ASAP7_75t_L g5829 ( 
.A(n_4469),
.Y(n_5829)
);

INVx1_ASAP7_75t_L g5830 ( 
.A(n_4366),
.Y(n_5830)
);

BUFx2_ASAP7_75t_SL g5831 ( 
.A(n_4212),
.Y(n_5831)
);

INVx2_ASAP7_75t_SL g5832 ( 
.A(n_4287),
.Y(n_5832)
);

CKINVDCx20_ASAP7_75t_R g5833 ( 
.A(n_4371),
.Y(n_5833)
);

INVx1_ASAP7_75t_L g5834 ( 
.A(n_4394),
.Y(n_5834)
);

INVx1_ASAP7_75t_L g5835 ( 
.A(n_4394),
.Y(n_5835)
);

CKINVDCx5p33_ASAP7_75t_R g5836 ( 
.A(n_4144),
.Y(n_5836)
);

CKINVDCx20_ASAP7_75t_R g5837 ( 
.A(n_4380),
.Y(n_5837)
);

CKINVDCx5p33_ASAP7_75t_R g5838 ( 
.A(n_4145),
.Y(n_5838)
);

CKINVDCx5p33_ASAP7_75t_R g5839 ( 
.A(n_4148),
.Y(n_5839)
);

BUFx6f_ASAP7_75t_L g5840 ( 
.A(n_4394),
.Y(n_5840)
);

CKINVDCx16_ASAP7_75t_R g5841 ( 
.A(n_4560),
.Y(n_5841)
);

CKINVDCx5p33_ASAP7_75t_R g5842 ( 
.A(n_4149),
.Y(n_5842)
);

INVx1_ASAP7_75t_SL g5843 ( 
.A(n_5303),
.Y(n_5843)
);

INVx1_ASAP7_75t_L g5844 ( 
.A(n_4453),
.Y(n_5844)
);

INVx1_ASAP7_75t_L g5845 ( 
.A(n_4453),
.Y(n_5845)
);

INVx1_ASAP7_75t_L g5846 ( 
.A(n_4453),
.Y(n_5846)
);

CKINVDCx5p33_ASAP7_75t_R g5847 ( 
.A(n_4153),
.Y(n_5847)
);

INVx1_ASAP7_75t_L g5848 ( 
.A(n_4490),
.Y(n_5848)
);

INVx1_ASAP7_75t_L g5849 ( 
.A(n_4490),
.Y(n_5849)
);

CKINVDCx5p33_ASAP7_75t_R g5850 ( 
.A(n_4154),
.Y(n_5850)
);

INVx1_ASAP7_75t_L g5851 ( 
.A(n_4490),
.Y(n_5851)
);

INVx1_ASAP7_75t_L g5852 ( 
.A(n_4552),
.Y(n_5852)
);

INVx1_ASAP7_75t_L g5853 ( 
.A(n_4552),
.Y(n_5853)
);

CKINVDCx5p33_ASAP7_75t_R g5854 ( 
.A(n_4155),
.Y(n_5854)
);

INVx1_ASAP7_75t_L g5855 ( 
.A(n_4552),
.Y(n_5855)
);

INVx1_ASAP7_75t_L g5856 ( 
.A(n_4666),
.Y(n_5856)
);

INVx1_ASAP7_75t_L g5857 ( 
.A(n_4666),
.Y(n_5857)
);

BUFx2_ASAP7_75t_L g5858 ( 
.A(n_5404),
.Y(n_5858)
);

CKINVDCx5p33_ASAP7_75t_R g5859 ( 
.A(n_4156),
.Y(n_5859)
);

INVx2_ASAP7_75t_SL g5860 ( 
.A(n_4560),
.Y(n_5860)
);

INVx1_ASAP7_75t_SL g5861 ( 
.A(n_5441),
.Y(n_5861)
);

CKINVDCx5p33_ASAP7_75t_R g5862 ( 
.A(n_4157),
.Y(n_5862)
);

INVx1_ASAP7_75t_L g5863 ( 
.A(n_4666),
.Y(n_5863)
);

CKINVDCx5p33_ASAP7_75t_R g5864 ( 
.A(n_4160),
.Y(n_5864)
);

BUFx10_ASAP7_75t_L g5865 ( 
.A(n_4578),
.Y(n_5865)
);

CKINVDCx5p33_ASAP7_75t_R g5866 ( 
.A(n_4162),
.Y(n_5866)
);

BUFx6f_ASAP7_75t_L g5867 ( 
.A(n_4671),
.Y(n_5867)
);

INVx1_ASAP7_75t_SL g5868 ( 
.A(n_4814),
.Y(n_5868)
);

CKINVDCx5p33_ASAP7_75t_R g5869 ( 
.A(n_5495),
.Y(n_5869)
);

INVx1_ASAP7_75t_L g5870 ( 
.A(n_4671),
.Y(n_5870)
);

BUFx3_ASAP7_75t_L g5871 ( 
.A(n_4258),
.Y(n_5871)
);

CKINVDCx5p33_ASAP7_75t_R g5872 ( 
.A(n_4168),
.Y(n_5872)
);

OR2x2_ASAP7_75t_L g5873 ( 
.A(n_4443),
.B(n_5488),
.Y(n_5873)
);

INVx1_ASAP7_75t_L g5874 ( 
.A(n_4671),
.Y(n_5874)
);

CKINVDCx5p33_ASAP7_75t_R g5875 ( 
.A(n_4169),
.Y(n_5875)
);

INVx1_ASAP7_75t_L g5876 ( 
.A(n_4746),
.Y(n_5876)
);

INVx2_ASAP7_75t_L g5877 ( 
.A(n_4746),
.Y(n_5877)
);

CKINVDCx20_ASAP7_75t_R g5878 ( 
.A(n_4403),
.Y(n_5878)
);

INVx1_ASAP7_75t_L g5879 ( 
.A(n_4746),
.Y(n_5879)
);

CKINVDCx5p33_ASAP7_75t_R g5880 ( 
.A(n_4170),
.Y(n_5880)
);

CKINVDCx5p33_ASAP7_75t_R g5881 ( 
.A(n_4176),
.Y(n_5881)
);

INVx1_ASAP7_75t_SL g5882 ( 
.A(n_4917),
.Y(n_5882)
);

INVx1_ASAP7_75t_L g5883 ( 
.A(n_4792),
.Y(n_5883)
);

CKINVDCx5p33_ASAP7_75t_R g5884 ( 
.A(n_4178),
.Y(n_5884)
);

INVx1_ASAP7_75t_L g5885 ( 
.A(n_4792),
.Y(n_5885)
);

BUFx3_ASAP7_75t_L g5886 ( 
.A(n_4292),
.Y(n_5886)
);

INVx1_ASAP7_75t_L g5887 ( 
.A(n_4792),
.Y(n_5887)
);

INVx1_ASAP7_75t_L g5888 ( 
.A(n_4799),
.Y(n_5888)
);

CKINVDCx5p33_ASAP7_75t_R g5889 ( 
.A(n_4180),
.Y(n_5889)
);

CKINVDCx5p33_ASAP7_75t_R g5890 ( 
.A(n_4183),
.Y(n_5890)
);

CKINVDCx5p33_ASAP7_75t_R g5891 ( 
.A(n_4187),
.Y(n_5891)
);

INVx2_ASAP7_75t_L g5892 ( 
.A(n_4799),
.Y(n_5892)
);

CKINVDCx5p33_ASAP7_75t_R g5893 ( 
.A(n_4190),
.Y(n_5893)
);

CKINVDCx5p33_ASAP7_75t_R g5894 ( 
.A(n_4192),
.Y(n_5894)
);

INVx1_ASAP7_75t_L g5895 ( 
.A(n_4799),
.Y(n_5895)
);

CKINVDCx5p33_ASAP7_75t_R g5896 ( 
.A(n_4193),
.Y(n_5896)
);

BUFx5_ASAP7_75t_L g5897 ( 
.A(n_4122),
.Y(n_5897)
);

CKINVDCx5p33_ASAP7_75t_R g5898 ( 
.A(n_4194),
.Y(n_5898)
);

INVx2_ASAP7_75t_L g5899 ( 
.A(n_4806),
.Y(n_5899)
);

CKINVDCx5p33_ASAP7_75t_R g5900 ( 
.A(n_4197),
.Y(n_5900)
);

CKINVDCx20_ASAP7_75t_R g5901 ( 
.A(n_4406),
.Y(n_5901)
);

CKINVDCx5p33_ASAP7_75t_R g5902 ( 
.A(n_4203),
.Y(n_5902)
);

CKINVDCx5p33_ASAP7_75t_R g5903 ( 
.A(n_4204),
.Y(n_5903)
);

INVx1_ASAP7_75t_L g5904 ( 
.A(n_4806),
.Y(n_5904)
);

INVx1_ASAP7_75t_L g5905 ( 
.A(n_4806),
.Y(n_5905)
);

CKINVDCx20_ASAP7_75t_R g5906 ( 
.A(n_4445),
.Y(n_5906)
);

CKINVDCx5p33_ASAP7_75t_R g5907 ( 
.A(n_4207),
.Y(n_5907)
);

INVx1_ASAP7_75t_L g5908 ( 
.A(n_4854),
.Y(n_5908)
);

INVx2_ASAP7_75t_L g5909 ( 
.A(n_4854),
.Y(n_5909)
);

CKINVDCx5p33_ASAP7_75t_R g5910 ( 
.A(n_4208),
.Y(n_5910)
);

CKINVDCx5p33_ASAP7_75t_R g5911 ( 
.A(n_4211),
.Y(n_5911)
);

CKINVDCx5p33_ASAP7_75t_R g5912 ( 
.A(n_4215),
.Y(n_5912)
);

INVx1_ASAP7_75t_L g5913 ( 
.A(n_4854),
.Y(n_5913)
);

CKINVDCx20_ASAP7_75t_R g5914 ( 
.A(n_4496),
.Y(n_5914)
);

BUFx3_ASAP7_75t_L g5915 ( 
.A(n_4304),
.Y(n_5915)
);

INVx1_ASAP7_75t_L g5916 ( 
.A(n_4878),
.Y(n_5916)
);

INVx1_ASAP7_75t_L g5917 ( 
.A(n_4878),
.Y(n_5917)
);

CKINVDCx5p33_ASAP7_75t_R g5918 ( 
.A(n_4216),
.Y(n_5918)
);

INVx1_ASAP7_75t_L g5919 ( 
.A(n_4878),
.Y(n_5919)
);

CKINVDCx5p33_ASAP7_75t_R g5920 ( 
.A(n_4218),
.Y(n_5920)
);

CKINVDCx5p33_ASAP7_75t_R g5921 ( 
.A(n_4219),
.Y(n_5921)
);

INVx1_ASAP7_75t_L g5922 ( 
.A(n_4894),
.Y(n_5922)
);

INVx1_ASAP7_75t_L g5923 ( 
.A(n_4894),
.Y(n_5923)
);

CKINVDCx5p33_ASAP7_75t_R g5924 ( 
.A(n_4220),
.Y(n_5924)
);

INVx1_ASAP7_75t_L g5925 ( 
.A(n_4894),
.Y(n_5925)
);

CKINVDCx20_ASAP7_75t_R g5926 ( 
.A(n_4498),
.Y(n_5926)
);

INVx1_ASAP7_75t_L g5927 ( 
.A(n_5014),
.Y(n_5927)
);

CKINVDCx5p33_ASAP7_75t_R g5928 ( 
.A(n_4222),
.Y(n_5928)
);

INVx1_ASAP7_75t_SL g5929 ( 
.A(n_5201),
.Y(n_5929)
);

CKINVDCx5p33_ASAP7_75t_R g5930 ( 
.A(n_4223),
.Y(n_5930)
);

CKINVDCx5p33_ASAP7_75t_R g5931 ( 
.A(n_4224),
.Y(n_5931)
);

INVx1_ASAP7_75t_L g5932 ( 
.A(n_5014),
.Y(n_5932)
);

CKINVDCx20_ASAP7_75t_R g5933 ( 
.A(n_4503),
.Y(n_5933)
);

INVxp33_ASAP7_75t_SL g5934 ( 
.A(n_4743),
.Y(n_5934)
);

CKINVDCx5p33_ASAP7_75t_R g5935 ( 
.A(n_4225),
.Y(n_5935)
);

INVx2_ASAP7_75t_L g5936 ( 
.A(n_5014),
.Y(n_5936)
);

CKINVDCx16_ASAP7_75t_R g5937 ( 
.A(n_5509),
.Y(n_5937)
);

BUFx3_ASAP7_75t_L g5938 ( 
.A(n_4337),
.Y(n_5938)
);

INVx1_ASAP7_75t_L g5939 ( 
.A(n_5031),
.Y(n_5939)
);

INVx1_ASAP7_75t_L g5940 ( 
.A(n_5031),
.Y(n_5940)
);

INVx1_ASAP7_75t_L g5941 ( 
.A(n_5031),
.Y(n_5941)
);

CKINVDCx5p33_ASAP7_75t_R g5942 ( 
.A(n_4228),
.Y(n_5942)
);

CKINVDCx5p33_ASAP7_75t_R g5943 ( 
.A(n_4230),
.Y(n_5943)
);

INVx1_ASAP7_75t_L g5944 ( 
.A(n_5053),
.Y(n_5944)
);

HB1xp67_ASAP7_75t_L g5945 ( 
.A(n_4908),
.Y(n_5945)
);

INVx1_ASAP7_75t_L g5946 ( 
.A(n_5053),
.Y(n_5946)
);

CKINVDCx5p33_ASAP7_75t_R g5947 ( 
.A(n_4231),
.Y(n_5947)
);

CKINVDCx5p33_ASAP7_75t_R g5948 ( 
.A(n_4232),
.Y(n_5948)
);

BUFx6f_ASAP7_75t_L g5949 ( 
.A(n_5053),
.Y(n_5949)
);

INVx1_ASAP7_75t_L g5950 ( 
.A(n_5087),
.Y(n_5950)
);

INVx1_ASAP7_75t_L g5951 ( 
.A(n_5087),
.Y(n_5951)
);

CKINVDCx5p33_ASAP7_75t_R g5952 ( 
.A(n_4236),
.Y(n_5952)
);

INVx1_ASAP7_75t_L g5953 ( 
.A(n_5087),
.Y(n_5953)
);

INVx1_ASAP7_75t_L g5954 ( 
.A(n_5094),
.Y(n_5954)
);

BUFx6f_ASAP7_75t_L g5955 ( 
.A(n_5094),
.Y(n_5955)
);

CKINVDCx5p33_ASAP7_75t_R g5956 ( 
.A(n_4238),
.Y(n_5956)
);

INVx2_ASAP7_75t_L g5957 ( 
.A(n_5094),
.Y(n_5957)
);

INVx1_ASAP7_75t_L g5958 ( 
.A(n_5120),
.Y(n_5958)
);

BUFx6f_ASAP7_75t_L g5959 ( 
.A(n_5120),
.Y(n_5959)
);

INVx1_ASAP7_75t_L g5960 ( 
.A(n_5120),
.Y(n_5960)
);

CKINVDCx5p33_ASAP7_75t_R g5961 ( 
.A(n_4239),
.Y(n_5961)
);

INVx2_ASAP7_75t_SL g5962 ( 
.A(n_4584),
.Y(n_5962)
);

CKINVDCx5p33_ASAP7_75t_R g5963 ( 
.A(n_4240),
.Y(n_5963)
);

BUFx6f_ASAP7_75t_L g5964 ( 
.A(n_5121),
.Y(n_5964)
);

CKINVDCx5p33_ASAP7_75t_R g5965 ( 
.A(n_4242),
.Y(n_5965)
);

INVx2_ASAP7_75t_L g5966 ( 
.A(n_5121),
.Y(n_5966)
);

BUFx2_ASAP7_75t_L g5967 ( 
.A(n_4382),
.Y(n_5967)
);

NOR2xp67_ASAP7_75t_L g5968 ( 
.A(n_4771),
.B(n_5),
.Y(n_5968)
);

CKINVDCx5p33_ASAP7_75t_R g5969 ( 
.A(n_4246),
.Y(n_5969)
);

CKINVDCx20_ASAP7_75t_R g5970 ( 
.A(n_5644),
.Y(n_5970)
);

INVx1_ASAP7_75t_L g5971 ( 
.A(n_5535),
.Y(n_5971)
);

INVx1_ASAP7_75t_L g5972 ( 
.A(n_5535),
.Y(n_5972)
);

INVx1_ASAP7_75t_L g5973 ( 
.A(n_5614),
.Y(n_5973)
);

CKINVDCx5p33_ASAP7_75t_R g5974 ( 
.A(n_5739),
.Y(n_5974)
);

CKINVDCx5p33_ASAP7_75t_R g5975 ( 
.A(n_5746),
.Y(n_5975)
);

INVx1_ASAP7_75t_L g5976 ( 
.A(n_5614),
.Y(n_5976)
);

INVx1_ASAP7_75t_L g5977 ( 
.A(n_5657),
.Y(n_5977)
);

INVx1_ASAP7_75t_L g5978 ( 
.A(n_5657),
.Y(n_5978)
);

INVxp67_ASAP7_75t_SL g5979 ( 
.A(n_5741),
.Y(n_5979)
);

INVx1_ASAP7_75t_L g5980 ( 
.A(n_5840),
.Y(n_5980)
);

CKINVDCx5p33_ASAP7_75t_R g5981 ( 
.A(n_5747),
.Y(n_5981)
);

INVx1_ASAP7_75t_L g5982 ( 
.A(n_5840),
.Y(n_5982)
);

INVx1_ASAP7_75t_L g5983 ( 
.A(n_5867),
.Y(n_5983)
);

CKINVDCx5p33_ASAP7_75t_R g5984 ( 
.A(n_5748),
.Y(n_5984)
);

INVx1_ASAP7_75t_L g5985 ( 
.A(n_5867),
.Y(n_5985)
);

CKINVDCx20_ASAP7_75t_R g5986 ( 
.A(n_5656),
.Y(n_5986)
);

INVx1_ASAP7_75t_L g5987 ( 
.A(n_5949),
.Y(n_5987)
);

INVx1_ASAP7_75t_L g5988 ( 
.A(n_5949),
.Y(n_5988)
);

CKINVDCx5p33_ASAP7_75t_R g5989 ( 
.A(n_5751),
.Y(n_5989)
);

HB1xp67_ASAP7_75t_L g5990 ( 
.A(n_5562),
.Y(n_5990)
);

CKINVDCx5p33_ASAP7_75t_R g5991 ( 
.A(n_5752),
.Y(n_5991)
);

INVx1_ASAP7_75t_L g5992 ( 
.A(n_5955),
.Y(n_5992)
);

INVx1_ASAP7_75t_L g5993 ( 
.A(n_5955),
.Y(n_5993)
);

CKINVDCx5p33_ASAP7_75t_R g5994 ( 
.A(n_5753),
.Y(n_5994)
);

INVx2_ASAP7_75t_SL g5995 ( 
.A(n_5583),
.Y(n_5995)
);

CKINVDCx5p33_ASAP7_75t_R g5996 ( 
.A(n_5754),
.Y(n_5996)
);

INVx1_ASAP7_75t_L g5997 ( 
.A(n_5959),
.Y(n_5997)
);

CKINVDCx20_ASAP7_75t_R g5998 ( 
.A(n_5664),
.Y(n_5998)
);

INVx1_ASAP7_75t_L g5999 ( 
.A(n_5959),
.Y(n_5999)
);

CKINVDCx5p33_ASAP7_75t_R g6000 ( 
.A(n_5759),
.Y(n_6000)
);

HB1xp67_ASAP7_75t_L g6001 ( 
.A(n_5566),
.Y(n_6001)
);

INVx2_ASAP7_75t_L g6002 ( 
.A(n_5756),
.Y(n_6002)
);

INVx1_ASAP7_75t_L g6003 ( 
.A(n_5964),
.Y(n_6003)
);

INVx1_ASAP7_75t_L g6004 ( 
.A(n_5964),
.Y(n_6004)
);

BUFx5_ASAP7_75t_L g6005 ( 
.A(n_5525),
.Y(n_6005)
);

INVx1_ASAP7_75t_L g6006 ( 
.A(n_5728),
.Y(n_6006)
);

INVx1_ASAP7_75t_L g6007 ( 
.A(n_5730),
.Y(n_6007)
);

INVx1_ASAP7_75t_L g6008 ( 
.A(n_5732),
.Y(n_6008)
);

INVx1_ASAP7_75t_L g6009 ( 
.A(n_5767),
.Y(n_6009)
);

CKINVDCx5p33_ASAP7_75t_R g6010 ( 
.A(n_5761),
.Y(n_6010)
);

INVx1_ASAP7_75t_L g6011 ( 
.A(n_5795),
.Y(n_6011)
);

INVx1_ASAP7_75t_L g6012 ( 
.A(n_5796),
.Y(n_6012)
);

CKINVDCx20_ASAP7_75t_R g6013 ( 
.A(n_5680),
.Y(n_6013)
);

CKINVDCx5p33_ASAP7_75t_R g6014 ( 
.A(n_5763),
.Y(n_6014)
);

INVx1_ASAP7_75t_L g6015 ( 
.A(n_5810),
.Y(n_6015)
);

INVx1_ASAP7_75t_L g6016 ( 
.A(n_5822),
.Y(n_6016)
);

INVx1_ASAP7_75t_L g6017 ( 
.A(n_5823),
.Y(n_6017)
);

CKINVDCx5p33_ASAP7_75t_R g6018 ( 
.A(n_5764),
.Y(n_6018)
);

INVx1_ASAP7_75t_L g6019 ( 
.A(n_5877),
.Y(n_6019)
);

CKINVDCx20_ASAP7_75t_R g6020 ( 
.A(n_5698),
.Y(n_6020)
);

INVx1_ASAP7_75t_L g6021 ( 
.A(n_5892),
.Y(n_6021)
);

INVxp67_ASAP7_75t_SL g6022 ( 
.A(n_5783),
.Y(n_6022)
);

INVx1_ASAP7_75t_L g6023 ( 
.A(n_5899),
.Y(n_6023)
);

INVx1_ASAP7_75t_L g6024 ( 
.A(n_5909),
.Y(n_6024)
);

INVx1_ASAP7_75t_L g6025 ( 
.A(n_5936),
.Y(n_6025)
);

INVx1_ASAP7_75t_L g6026 ( 
.A(n_5957),
.Y(n_6026)
);

CKINVDCx5p33_ASAP7_75t_R g6027 ( 
.A(n_5765),
.Y(n_6027)
);

INVx1_ASAP7_75t_L g6028 ( 
.A(n_5966),
.Y(n_6028)
);

CKINVDCx5p33_ASAP7_75t_R g6029 ( 
.A(n_5770),
.Y(n_6029)
);

BUFx2_ASAP7_75t_L g6030 ( 
.A(n_5588),
.Y(n_6030)
);

INVx1_ASAP7_75t_L g6031 ( 
.A(n_5743),
.Y(n_6031)
);

INVxp33_ASAP7_75t_SL g6032 ( 
.A(n_5537),
.Y(n_6032)
);

CKINVDCx20_ASAP7_75t_R g6033 ( 
.A(n_5708),
.Y(n_6033)
);

INVx1_ASAP7_75t_L g6034 ( 
.A(n_5744),
.Y(n_6034)
);

INVx1_ASAP7_75t_L g6035 ( 
.A(n_5755),
.Y(n_6035)
);

CKINVDCx5p33_ASAP7_75t_R g6036 ( 
.A(n_5772),
.Y(n_6036)
);

INVx2_ASAP7_75t_L g6037 ( 
.A(n_5757),
.Y(n_6037)
);

CKINVDCx5p33_ASAP7_75t_R g6038 ( 
.A(n_5776),
.Y(n_6038)
);

INVx1_ASAP7_75t_L g6039 ( 
.A(n_5758),
.Y(n_6039)
);

INVxp67_ASAP7_75t_L g6040 ( 
.A(n_5544),
.Y(n_6040)
);

INVxp67_ASAP7_75t_L g6041 ( 
.A(n_5967),
.Y(n_6041)
);

INVx1_ASAP7_75t_L g6042 ( 
.A(n_5760),
.Y(n_6042)
);

CKINVDCx20_ASAP7_75t_R g6043 ( 
.A(n_5749),
.Y(n_6043)
);

INVx1_ASAP7_75t_L g6044 ( 
.A(n_5768),
.Y(n_6044)
);

CKINVDCx5p33_ASAP7_75t_R g6045 ( 
.A(n_5780),
.Y(n_6045)
);

INVx1_ASAP7_75t_L g6046 ( 
.A(n_5773),
.Y(n_6046)
);

INVx1_ASAP7_75t_L g6047 ( 
.A(n_5775),
.Y(n_6047)
);

HB1xp67_ASAP7_75t_L g6048 ( 
.A(n_5567),
.Y(n_6048)
);

CKINVDCx5p33_ASAP7_75t_R g6049 ( 
.A(n_5786),
.Y(n_6049)
);

INVx1_ASAP7_75t_L g6050 ( 
.A(n_5777),
.Y(n_6050)
);

CKINVDCx5p33_ASAP7_75t_R g6051 ( 
.A(n_5791),
.Y(n_6051)
);

INVx1_ASAP7_75t_L g6052 ( 
.A(n_5779),
.Y(n_6052)
);

CKINVDCx20_ASAP7_75t_R g6053 ( 
.A(n_5766),
.Y(n_6053)
);

INVx1_ASAP7_75t_L g6054 ( 
.A(n_5781),
.Y(n_6054)
);

INVx1_ASAP7_75t_L g6055 ( 
.A(n_5784),
.Y(n_6055)
);

INVx1_ASAP7_75t_L g6056 ( 
.A(n_5785),
.Y(n_6056)
);

INVx1_ASAP7_75t_L g6057 ( 
.A(n_5787),
.Y(n_6057)
);

INVx1_ASAP7_75t_SL g6058 ( 
.A(n_5868),
.Y(n_6058)
);

INVx1_ASAP7_75t_L g6059 ( 
.A(n_5794),
.Y(n_6059)
);

CKINVDCx5p33_ASAP7_75t_R g6060 ( 
.A(n_5792),
.Y(n_6060)
);

CKINVDCx20_ASAP7_75t_R g6061 ( 
.A(n_5782),
.Y(n_6061)
);

INVx1_ASAP7_75t_L g6062 ( 
.A(n_5799),
.Y(n_6062)
);

INVx1_ASAP7_75t_L g6063 ( 
.A(n_5801),
.Y(n_6063)
);

INVxp33_ASAP7_75t_L g6064 ( 
.A(n_5733),
.Y(n_6064)
);

INVx1_ASAP7_75t_L g6065 ( 
.A(n_5804),
.Y(n_6065)
);

CKINVDCx20_ASAP7_75t_R g6066 ( 
.A(n_5790),
.Y(n_6066)
);

INVx1_ASAP7_75t_L g6067 ( 
.A(n_5808),
.Y(n_6067)
);

CKINVDCx5p33_ASAP7_75t_R g6068 ( 
.A(n_5803),
.Y(n_6068)
);

INVx1_ASAP7_75t_L g6069 ( 
.A(n_5813),
.Y(n_6069)
);

INVx2_ASAP7_75t_L g6070 ( 
.A(n_5815),
.Y(n_6070)
);

CKINVDCx5p33_ASAP7_75t_R g6071 ( 
.A(n_5809),
.Y(n_6071)
);

INVx1_ASAP7_75t_L g6072 ( 
.A(n_5816),
.Y(n_6072)
);

INVx1_ASAP7_75t_L g6073 ( 
.A(n_5817),
.Y(n_6073)
);

INVxp67_ASAP7_75t_SL g6074 ( 
.A(n_5806),
.Y(n_6074)
);

INVxp67_ASAP7_75t_SL g6075 ( 
.A(n_5807),
.Y(n_6075)
);

HB1xp67_ASAP7_75t_L g6076 ( 
.A(n_5569),
.Y(n_6076)
);

CKINVDCx5p33_ASAP7_75t_R g6077 ( 
.A(n_5811),
.Y(n_6077)
);

CKINVDCx16_ASAP7_75t_R g6078 ( 
.A(n_5634),
.Y(n_6078)
);

INVx2_ASAP7_75t_L g6079 ( 
.A(n_5818),
.Y(n_6079)
);

INVx1_ASAP7_75t_SL g6080 ( 
.A(n_5882),
.Y(n_6080)
);

INVx1_ASAP7_75t_L g6081 ( 
.A(n_5820),
.Y(n_6081)
);

CKINVDCx5p33_ASAP7_75t_R g6082 ( 
.A(n_5814),
.Y(n_6082)
);

INVx1_ASAP7_75t_L g6083 ( 
.A(n_5821),
.Y(n_6083)
);

INVx1_ASAP7_75t_L g6084 ( 
.A(n_5825),
.Y(n_6084)
);

INVxp67_ASAP7_75t_L g6085 ( 
.A(n_5727),
.Y(n_6085)
);

CKINVDCx20_ASAP7_75t_R g6086 ( 
.A(n_5805),
.Y(n_6086)
);

CKINVDCx5p33_ASAP7_75t_R g6087 ( 
.A(n_5819),
.Y(n_6087)
);

INVx1_ASAP7_75t_L g6088 ( 
.A(n_5830),
.Y(n_6088)
);

INVx1_ASAP7_75t_L g6089 ( 
.A(n_5834),
.Y(n_6089)
);

INVx1_ASAP7_75t_L g6090 ( 
.A(n_5835),
.Y(n_6090)
);

INVx1_ASAP7_75t_L g6091 ( 
.A(n_5844),
.Y(n_6091)
);

CKINVDCx5p33_ASAP7_75t_R g6092 ( 
.A(n_5824),
.Y(n_6092)
);

INVx1_ASAP7_75t_L g6093 ( 
.A(n_5845),
.Y(n_6093)
);

INVx1_ASAP7_75t_L g6094 ( 
.A(n_5846),
.Y(n_6094)
);

HB1xp67_ASAP7_75t_L g6095 ( 
.A(n_5570),
.Y(n_6095)
);

HB1xp67_ASAP7_75t_L g6096 ( 
.A(n_5574),
.Y(n_6096)
);

INVx2_ASAP7_75t_L g6097 ( 
.A(n_5848),
.Y(n_6097)
);

INVx1_ASAP7_75t_L g6098 ( 
.A(n_5849),
.Y(n_6098)
);

INVx1_ASAP7_75t_L g6099 ( 
.A(n_5851),
.Y(n_6099)
);

CKINVDCx5p33_ASAP7_75t_R g6100 ( 
.A(n_5826),
.Y(n_6100)
);

CKINVDCx5p33_ASAP7_75t_R g6101 ( 
.A(n_5828),
.Y(n_6101)
);

INVxp33_ASAP7_75t_SL g6102 ( 
.A(n_5538),
.Y(n_6102)
);

CKINVDCx5p33_ASAP7_75t_R g6103 ( 
.A(n_5836),
.Y(n_6103)
);

INVx1_ASAP7_75t_L g6104 ( 
.A(n_5852),
.Y(n_6104)
);

CKINVDCx5p33_ASAP7_75t_R g6105 ( 
.A(n_5838),
.Y(n_6105)
);

INVx1_ASAP7_75t_L g6106 ( 
.A(n_5853),
.Y(n_6106)
);

INVx1_ASAP7_75t_L g6107 ( 
.A(n_5855),
.Y(n_6107)
);

INVx1_ASAP7_75t_SL g6108 ( 
.A(n_5929),
.Y(n_6108)
);

INVx1_ASAP7_75t_L g6109 ( 
.A(n_5856),
.Y(n_6109)
);

CKINVDCx5p33_ASAP7_75t_R g6110 ( 
.A(n_5839),
.Y(n_6110)
);

INVx1_ASAP7_75t_L g6111 ( 
.A(n_5857),
.Y(n_6111)
);

INVx1_ASAP7_75t_L g6112 ( 
.A(n_5863),
.Y(n_6112)
);

INVxp67_ASAP7_75t_SL g6113 ( 
.A(n_5871),
.Y(n_6113)
);

CKINVDCx20_ASAP7_75t_R g6114 ( 
.A(n_5812),
.Y(n_6114)
);

INVx1_ASAP7_75t_L g6115 ( 
.A(n_5870),
.Y(n_6115)
);

INVxp67_ASAP7_75t_L g6116 ( 
.A(n_5832),
.Y(n_6116)
);

INVx1_ASAP7_75t_L g6117 ( 
.A(n_5874),
.Y(n_6117)
);

INVx1_ASAP7_75t_SL g6118 ( 
.A(n_5647),
.Y(n_6118)
);

INVx1_ASAP7_75t_L g6119 ( 
.A(n_5876),
.Y(n_6119)
);

INVx2_ASAP7_75t_L g6120 ( 
.A(n_5879),
.Y(n_6120)
);

INVx1_ASAP7_75t_L g6121 ( 
.A(n_5883),
.Y(n_6121)
);

CKINVDCx16_ASAP7_75t_R g6122 ( 
.A(n_5543),
.Y(n_6122)
);

INVx1_ASAP7_75t_L g6123 ( 
.A(n_5885),
.Y(n_6123)
);

INVx1_ASAP7_75t_L g6124 ( 
.A(n_5887),
.Y(n_6124)
);

CKINVDCx5p33_ASAP7_75t_R g6125 ( 
.A(n_5842),
.Y(n_6125)
);

CKINVDCx14_ASAP7_75t_R g6126 ( 
.A(n_5797),
.Y(n_6126)
);

INVx2_ASAP7_75t_L g6127 ( 
.A(n_5888),
.Y(n_6127)
);

INVx1_ASAP7_75t_L g6128 ( 
.A(n_5895),
.Y(n_6128)
);

INVx1_ASAP7_75t_L g6129 ( 
.A(n_5904),
.Y(n_6129)
);

INVx1_ASAP7_75t_L g6130 ( 
.A(n_5905),
.Y(n_6130)
);

CKINVDCx16_ASAP7_75t_R g6131 ( 
.A(n_5552),
.Y(n_6131)
);

INVx1_ASAP7_75t_L g6132 ( 
.A(n_5908),
.Y(n_6132)
);

INVxp67_ASAP7_75t_L g6133 ( 
.A(n_5860),
.Y(n_6133)
);

CKINVDCx20_ASAP7_75t_R g6134 ( 
.A(n_5833),
.Y(n_6134)
);

CKINVDCx5p33_ASAP7_75t_R g6135 ( 
.A(n_5847),
.Y(n_6135)
);

CKINVDCx20_ASAP7_75t_R g6136 ( 
.A(n_5837),
.Y(n_6136)
);

INVxp67_ASAP7_75t_L g6137 ( 
.A(n_5962),
.Y(n_6137)
);

CKINVDCx20_ASAP7_75t_R g6138 ( 
.A(n_5878),
.Y(n_6138)
);

INVx1_ASAP7_75t_L g6139 ( 
.A(n_5913),
.Y(n_6139)
);

INVx1_ASAP7_75t_L g6140 ( 
.A(n_5916),
.Y(n_6140)
);

BUFx3_ASAP7_75t_L g6141 ( 
.A(n_5533),
.Y(n_6141)
);

INVx1_ASAP7_75t_L g6142 ( 
.A(n_5917),
.Y(n_6142)
);

INVxp33_ASAP7_75t_SL g6143 ( 
.A(n_5540),
.Y(n_6143)
);

CKINVDCx5p33_ASAP7_75t_R g6144 ( 
.A(n_5850),
.Y(n_6144)
);

INVx1_ASAP7_75t_L g6145 ( 
.A(n_5919),
.Y(n_6145)
);

INVx1_ASAP7_75t_L g6146 ( 
.A(n_5922),
.Y(n_6146)
);

INVx1_ASAP7_75t_L g6147 ( 
.A(n_5923),
.Y(n_6147)
);

INVx1_ASAP7_75t_L g6148 ( 
.A(n_5925),
.Y(n_6148)
);

CKINVDCx20_ASAP7_75t_R g6149 ( 
.A(n_5901),
.Y(n_6149)
);

INVx1_ASAP7_75t_L g6150 ( 
.A(n_5927),
.Y(n_6150)
);

INVx1_ASAP7_75t_L g6151 ( 
.A(n_5932),
.Y(n_6151)
);

BUFx2_ASAP7_75t_L g6152 ( 
.A(n_5590),
.Y(n_6152)
);

INVx1_ASAP7_75t_L g6153 ( 
.A(n_5939),
.Y(n_6153)
);

INVx1_ASAP7_75t_L g6154 ( 
.A(n_5940),
.Y(n_6154)
);

INVx1_ASAP7_75t_L g6155 ( 
.A(n_5941),
.Y(n_6155)
);

INVx1_ASAP7_75t_L g6156 ( 
.A(n_5944),
.Y(n_6156)
);

CKINVDCx5p33_ASAP7_75t_R g6157 ( 
.A(n_5854),
.Y(n_6157)
);

INVx1_ASAP7_75t_L g6158 ( 
.A(n_5946),
.Y(n_6158)
);

CKINVDCx5p33_ASAP7_75t_R g6159 ( 
.A(n_5859),
.Y(n_6159)
);

INVx1_ASAP7_75t_L g6160 ( 
.A(n_5950),
.Y(n_6160)
);

CKINVDCx20_ASAP7_75t_R g6161 ( 
.A(n_5906),
.Y(n_6161)
);

INVx1_ASAP7_75t_L g6162 ( 
.A(n_5951),
.Y(n_6162)
);

INVx1_ASAP7_75t_L g6163 ( 
.A(n_5953),
.Y(n_6163)
);

CKINVDCx16_ASAP7_75t_R g6164 ( 
.A(n_5549),
.Y(n_6164)
);

INVxp33_ASAP7_75t_L g6165 ( 
.A(n_5655),
.Y(n_6165)
);

INVx1_ASAP7_75t_L g6166 ( 
.A(n_5954),
.Y(n_6166)
);

CKINVDCx20_ASAP7_75t_R g6167 ( 
.A(n_5914),
.Y(n_6167)
);

CKINVDCx20_ASAP7_75t_R g6168 ( 
.A(n_5926),
.Y(n_6168)
);

CKINVDCx5p33_ASAP7_75t_R g6169 ( 
.A(n_5862),
.Y(n_6169)
);

INVxp33_ASAP7_75t_SL g6170 ( 
.A(n_5545),
.Y(n_6170)
);

INVx1_ASAP7_75t_L g6171 ( 
.A(n_5958),
.Y(n_6171)
);

INVx1_ASAP7_75t_L g6172 ( 
.A(n_5960),
.Y(n_6172)
);

BUFx3_ASAP7_75t_L g6173 ( 
.A(n_5571),
.Y(n_6173)
);

INVx1_ASAP7_75t_L g6174 ( 
.A(n_5527),
.Y(n_6174)
);

INVx1_ASAP7_75t_L g6175 ( 
.A(n_5528),
.Y(n_6175)
);

INVx1_ASAP7_75t_L g6176 ( 
.A(n_5529),
.Y(n_6176)
);

CKINVDCx20_ASAP7_75t_R g6177 ( 
.A(n_5933),
.Y(n_6177)
);

CKINVDCx16_ASAP7_75t_R g6178 ( 
.A(n_5609),
.Y(n_6178)
);

BUFx3_ASAP7_75t_L g6179 ( 
.A(n_5886),
.Y(n_6179)
);

CKINVDCx5p33_ASAP7_75t_R g6180 ( 
.A(n_5864),
.Y(n_6180)
);

CKINVDCx5p33_ASAP7_75t_R g6181 ( 
.A(n_5866),
.Y(n_6181)
);

INVx1_ASAP7_75t_L g6182 ( 
.A(n_5530),
.Y(n_6182)
);

INVx1_ASAP7_75t_L g6183 ( 
.A(n_5534),
.Y(n_6183)
);

INVx1_ASAP7_75t_L g6184 ( 
.A(n_5536),
.Y(n_6184)
);

INVx1_ASAP7_75t_L g6185 ( 
.A(n_5539),
.Y(n_6185)
);

INVx1_ASAP7_75t_L g6186 ( 
.A(n_5541),
.Y(n_6186)
);

INVx1_ASAP7_75t_L g6187 ( 
.A(n_5542),
.Y(n_6187)
);

INVx2_ASAP7_75t_L g6188 ( 
.A(n_5561),
.Y(n_6188)
);

INVx1_ASAP7_75t_L g6189 ( 
.A(n_5547),
.Y(n_6189)
);

INVx1_ASAP7_75t_L g6190 ( 
.A(n_5553),
.Y(n_6190)
);

INVxp67_ASAP7_75t_SL g6191 ( 
.A(n_5915),
.Y(n_6191)
);

CKINVDCx5p33_ASAP7_75t_R g6192 ( 
.A(n_5869),
.Y(n_6192)
);

BUFx3_ASAP7_75t_L g6193 ( 
.A(n_5938),
.Y(n_6193)
);

HB1xp67_ASAP7_75t_L g6194 ( 
.A(n_5575),
.Y(n_6194)
);

INVx1_ASAP7_75t_L g6195 ( 
.A(n_5557),
.Y(n_6195)
);

INVxp67_ASAP7_75t_SL g6196 ( 
.A(n_5526),
.Y(n_6196)
);

INVx1_ASAP7_75t_L g6197 ( 
.A(n_5568),
.Y(n_6197)
);

INVxp67_ASAP7_75t_SL g6198 ( 
.A(n_5771),
.Y(n_6198)
);

INVx2_ASAP7_75t_L g6199 ( 
.A(n_5586),
.Y(n_6199)
);

INVxp67_ASAP7_75t_L g6200 ( 
.A(n_5565),
.Y(n_6200)
);

CKINVDCx5p33_ASAP7_75t_R g6201 ( 
.A(n_5872),
.Y(n_6201)
);

INVx1_ASAP7_75t_L g6202 ( 
.A(n_5572),
.Y(n_6202)
);

INVxp33_ASAP7_75t_SL g6203 ( 
.A(n_5551),
.Y(n_6203)
);

CKINVDCx5p33_ASAP7_75t_R g6204 ( 
.A(n_5875),
.Y(n_6204)
);

INVx1_ASAP7_75t_L g6205 ( 
.A(n_5576),
.Y(n_6205)
);

INVx1_ASAP7_75t_L g6206 ( 
.A(n_5577),
.Y(n_6206)
);

INVxp67_ASAP7_75t_L g6207 ( 
.A(n_5582),
.Y(n_6207)
);

INVx1_ASAP7_75t_L g6208 ( 
.A(n_5581),
.Y(n_6208)
);

INVx1_ASAP7_75t_L g6209 ( 
.A(n_5584),
.Y(n_6209)
);

INVx1_ASAP7_75t_L g6210 ( 
.A(n_5591),
.Y(n_6210)
);

INVxp67_ASAP7_75t_L g6211 ( 
.A(n_5681),
.Y(n_6211)
);

INVx1_ASAP7_75t_L g6212 ( 
.A(n_5592),
.Y(n_6212)
);

INVx1_ASAP7_75t_L g6213 ( 
.A(n_5593),
.Y(n_6213)
);

INVx1_ASAP7_75t_L g6214 ( 
.A(n_5595),
.Y(n_6214)
);

INVx2_ASAP7_75t_L g6215 ( 
.A(n_5606),
.Y(n_6215)
);

CKINVDCx5p33_ASAP7_75t_R g6216 ( 
.A(n_5880),
.Y(n_6216)
);

CKINVDCx20_ASAP7_75t_R g6217 ( 
.A(n_5617),
.Y(n_6217)
);

INVxp67_ASAP7_75t_SL g6218 ( 
.A(n_5532),
.Y(n_6218)
);

INVx1_ASAP7_75t_L g6219 ( 
.A(n_5596),
.Y(n_6219)
);

INVx2_ASAP7_75t_SL g6220 ( 
.A(n_5661),
.Y(n_6220)
);

INVxp33_ASAP7_75t_SL g6221 ( 
.A(n_5554),
.Y(n_6221)
);

INVxp67_ASAP7_75t_SL g6222 ( 
.A(n_5597),
.Y(n_6222)
);

INVxp67_ASAP7_75t_L g6223 ( 
.A(n_5800),
.Y(n_6223)
);

INVx1_ASAP7_75t_L g6224 ( 
.A(n_5598),
.Y(n_6224)
);

CKINVDCx20_ASAP7_75t_R g6225 ( 
.A(n_5578),
.Y(n_6225)
);

INVxp67_ASAP7_75t_SL g6226 ( 
.A(n_5699),
.Y(n_6226)
);

CKINVDCx5p33_ASAP7_75t_R g6227 ( 
.A(n_5881),
.Y(n_6227)
);

INVxp67_ASAP7_75t_L g6228 ( 
.A(n_5858),
.Y(n_6228)
);

INVxp67_ASAP7_75t_SL g6229 ( 
.A(n_5723),
.Y(n_6229)
);

INVx1_ASAP7_75t_L g6230 ( 
.A(n_5600),
.Y(n_6230)
);

INVxp67_ASAP7_75t_L g6231 ( 
.A(n_5742),
.Y(n_6231)
);

INVx1_ASAP7_75t_L g6232 ( 
.A(n_5601),
.Y(n_6232)
);

CKINVDCx16_ASAP7_75t_R g6233 ( 
.A(n_5653),
.Y(n_6233)
);

INVx1_ASAP7_75t_L g6234 ( 
.A(n_5603),
.Y(n_6234)
);

CKINVDCx5p33_ASAP7_75t_R g6235 ( 
.A(n_5884),
.Y(n_6235)
);

HB1xp67_ASAP7_75t_L g6236 ( 
.A(n_5579),
.Y(n_6236)
);

INVxp67_ASAP7_75t_L g6237 ( 
.A(n_5831),
.Y(n_6237)
);

BUFx10_ASAP7_75t_L g6238 ( 
.A(n_5555),
.Y(n_6238)
);

CKINVDCx5p33_ASAP7_75t_R g6239 ( 
.A(n_5889),
.Y(n_6239)
);

CKINVDCx5p33_ASAP7_75t_R g6240 ( 
.A(n_5890),
.Y(n_6240)
);

INVx1_ASAP7_75t_L g6241 ( 
.A(n_5604),
.Y(n_6241)
);

INVx1_ASAP7_75t_L g6242 ( 
.A(n_5605),
.Y(n_6242)
);

INVx1_ASAP7_75t_L g6243 ( 
.A(n_5611),
.Y(n_6243)
);

HB1xp67_ASAP7_75t_L g6244 ( 
.A(n_5580),
.Y(n_6244)
);

INVx2_ASAP7_75t_L g6245 ( 
.A(n_5608),
.Y(n_6245)
);

INVx1_ASAP7_75t_L g6246 ( 
.A(n_5612),
.Y(n_6246)
);

INVxp67_ASAP7_75t_L g6247 ( 
.A(n_5573),
.Y(n_6247)
);

INVx1_ASAP7_75t_L g6248 ( 
.A(n_5615),
.Y(n_6248)
);

INVxp33_ASAP7_75t_SL g6249 ( 
.A(n_5531),
.Y(n_6249)
);

INVx1_ASAP7_75t_L g6250 ( 
.A(n_5618),
.Y(n_6250)
);

INVx2_ASAP7_75t_L g6251 ( 
.A(n_5622),
.Y(n_6251)
);

HB1xp67_ASAP7_75t_L g6252 ( 
.A(n_5585),
.Y(n_6252)
);

INVx1_ASAP7_75t_L g6253 ( 
.A(n_5623),
.Y(n_6253)
);

CKINVDCx20_ASAP7_75t_R g6254 ( 
.A(n_5587),
.Y(n_6254)
);

INVx1_ASAP7_75t_L g6255 ( 
.A(n_5627),
.Y(n_6255)
);

INVx1_ASAP7_75t_L g6256 ( 
.A(n_5629),
.Y(n_6256)
);

CKINVDCx5p33_ASAP7_75t_R g6257 ( 
.A(n_5891),
.Y(n_6257)
);

INVx1_ASAP7_75t_L g6258 ( 
.A(n_5630),
.Y(n_6258)
);

INVx1_ASAP7_75t_L g6259 ( 
.A(n_5632),
.Y(n_6259)
);

CKINVDCx16_ASAP7_75t_R g6260 ( 
.A(n_5667),
.Y(n_6260)
);

INVxp67_ASAP7_75t_SL g6261 ( 
.A(n_5712),
.Y(n_6261)
);

CKINVDCx5p33_ASAP7_75t_R g6262 ( 
.A(n_5893),
.Y(n_6262)
);

INVx1_ASAP7_75t_L g6263 ( 
.A(n_5637),
.Y(n_6263)
);

INVxp67_ASAP7_75t_L g6264 ( 
.A(n_5599),
.Y(n_6264)
);

INVx1_ASAP7_75t_L g6265 ( 
.A(n_5640),
.Y(n_6265)
);

CKINVDCx20_ASAP7_75t_R g6266 ( 
.A(n_5602),
.Y(n_6266)
);

CKINVDCx20_ASAP7_75t_R g6267 ( 
.A(n_5607),
.Y(n_6267)
);

INVx1_ASAP7_75t_L g6268 ( 
.A(n_5650),
.Y(n_6268)
);

INVx1_ASAP7_75t_L g6269 ( 
.A(n_5654),
.Y(n_6269)
);

INVx1_ASAP7_75t_L g6270 ( 
.A(n_5658),
.Y(n_6270)
);

CKINVDCx20_ASAP7_75t_R g6271 ( 
.A(n_5610),
.Y(n_6271)
);

INVx1_ASAP7_75t_L g6272 ( 
.A(n_5662),
.Y(n_6272)
);

INVxp67_ASAP7_75t_SL g6273 ( 
.A(n_5718),
.Y(n_6273)
);

CKINVDCx5p33_ASAP7_75t_R g6274 ( 
.A(n_5894),
.Y(n_6274)
);

INVx3_ASAP7_75t_L g6275 ( 
.A(n_5734),
.Y(n_6275)
);

INVx1_ASAP7_75t_L g6276 ( 
.A(n_5663),
.Y(n_6276)
);

CKINVDCx5p33_ASAP7_75t_R g6277 ( 
.A(n_5896),
.Y(n_6277)
);

CKINVDCx5p33_ASAP7_75t_R g6278 ( 
.A(n_5898),
.Y(n_6278)
);

CKINVDCx5p33_ASAP7_75t_R g6279 ( 
.A(n_5900),
.Y(n_6279)
);

CKINVDCx5p33_ASAP7_75t_R g6280 ( 
.A(n_5902),
.Y(n_6280)
);

INVxp67_ASAP7_75t_SL g6281 ( 
.A(n_5719),
.Y(n_6281)
);

INVxp33_ASAP7_75t_L g6282 ( 
.A(n_5798),
.Y(n_6282)
);

CKINVDCx20_ASAP7_75t_R g6283 ( 
.A(n_5613),
.Y(n_6283)
);

CKINVDCx20_ASAP7_75t_R g6284 ( 
.A(n_5619),
.Y(n_6284)
);

INVxp33_ASAP7_75t_SL g6285 ( 
.A(n_5556),
.Y(n_6285)
);

CKINVDCx16_ASAP7_75t_R g6286 ( 
.A(n_5676),
.Y(n_6286)
);

INVx1_ASAP7_75t_L g6287 ( 
.A(n_5665),
.Y(n_6287)
);

INVxp67_ASAP7_75t_SL g6288 ( 
.A(n_5721),
.Y(n_6288)
);

CKINVDCx5p33_ASAP7_75t_R g6289 ( 
.A(n_5903),
.Y(n_6289)
);

CKINVDCx5p33_ASAP7_75t_R g6290 ( 
.A(n_5907),
.Y(n_6290)
);

CKINVDCx5p33_ASAP7_75t_R g6291 ( 
.A(n_5910),
.Y(n_6291)
);

CKINVDCx5p33_ASAP7_75t_R g6292 ( 
.A(n_5911),
.Y(n_6292)
);

INVx1_ASAP7_75t_L g6293 ( 
.A(n_5666),
.Y(n_6293)
);

CKINVDCx5p33_ASAP7_75t_R g6294 ( 
.A(n_5912),
.Y(n_6294)
);

HB1xp67_ASAP7_75t_L g6295 ( 
.A(n_5918),
.Y(n_6295)
);

CKINVDCx20_ASAP7_75t_R g6296 ( 
.A(n_5920),
.Y(n_6296)
);

CKINVDCx5p33_ASAP7_75t_R g6297 ( 
.A(n_5921),
.Y(n_6297)
);

INVx1_ASAP7_75t_L g6298 ( 
.A(n_5671),
.Y(n_6298)
);

INVxp67_ASAP7_75t_SL g6299 ( 
.A(n_5873),
.Y(n_6299)
);

INVx1_ASAP7_75t_L g6300 ( 
.A(n_5674),
.Y(n_6300)
);

INVx1_ASAP7_75t_L g6301 ( 
.A(n_5677),
.Y(n_6301)
);

BUFx6f_ASAP7_75t_SL g6302 ( 
.A(n_5865),
.Y(n_6302)
);

INVx2_ASAP7_75t_L g6303 ( 
.A(n_5633),
.Y(n_6303)
);

INVxp67_ASAP7_75t_L g6304 ( 
.A(n_5616),
.Y(n_6304)
);

INVx1_ASAP7_75t_L g6305 ( 
.A(n_5678),
.Y(n_6305)
);

BUFx2_ASAP7_75t_L g6306 ( 
.A(n_5924),
.Y(n_6306)
);

CKINVDCx5p33_ASAP7_75t_R g6307 ( 
.A(n_5928),
.Y(n_6307)
);

HB1xp67_ASAP7_75t_L g6308 ( 
.A(n_5930),
.Y(n_6308)
);

HB1xp67_ASAP7_75t_L g6309 ( 
.A(n_5931),
.Y(n_6309)
);

INVx1_ASAP7_75t_L g6310 ( 
.A(n_5679),
.Y(n_6310)
);

INVx1_ASAP7_75t_L g6311 ( 
.A(n_5682),
.Y(n_6311)
);

CKINVDCx20_ASAP7_75t_R g6312 ( 
.A(n_5935),
.Y(n_6312)
);

INVx1_ASAP7_75t_L g6313 ( 
.A(n_5683),
.Y(n_6313)
);

INVx1_ASAP7_75t_L g6314 ( 
.A(n_5685),
.Y(n_6314)
);

CKINVDCx20_ASAP7_75t_R g6315 ( 
.A(n_5942),
.Y(n_6315)
);

INVx1_ASAP7_75t_L g6316 ( 
.A(n_5686),
.Y(n_6316)
);

CKINVDCx5p33_ASAP7_75t_R g6317 ( 
.A(n_5943),
.Y(n_6317)
);

CKINVDCx5p33_ASAP7_75t_R g6318 ( 
.A(n_5947),
.Y(n_6318)
);

INVx1_ASAP7_75t_L g6319 ( 
.A(n_5691),
.Y(n_6319)
);

CKINVDCx5p33_ASAP7_75t_R g6320 ( 
.A(n_5948),
.Y(n_6320)
);

INVx1_ASAP7_75t_L g6321 ( 
.A(n_5697),
.Y(n_6321)
);

HB1xp67_ASAP7_75t_L g6322 ( 
.A(n_5952),
.Y(n_6322)
);

INVx1_ASAP7_75t_L g6323 ( 
.A(n_5701),
.Y(n_6323)
);

INVxp33_ASAP7_75t_L g6324 ( 
.A(n_5829),
.Y(n_6324)
);

CKINVDCx20_ASAP7_75t_R g6325 ( 
.A(n_5956),
.Y(n_6325)
);

INVxp67_ASAP7_75t_SL g6326 ( 
.A(n_5945),
.Y(n_6326)
);

INVx1_ASAP7_75t_L g6327 ( 
.A(n_5703),
.Y(n_6327)
);

INVx1_ASAP7_75t_L g6328 ( 
.A(n_5706),
.Y(n_6328)
);

INVx1_ASAP7_75t_L g6329 ( 
.A(n_5707),
.Y(n_6329)
);

CKINVDCx5p33_ASAP7_75t_R g6330 ( 
.A(n_5961),
.Y(n_6330)
);

INVxp33_ASAP7_75t_SL g6331 ( 
.A(n_5558),
.Y(n_6331)
);

INVx1_ASAP7_75t_L g6332 ( 
.A(n_5709),
.Y(n_6332)
);

CKINVDCx16_ASAP7_75t_R g6333 ( 
.A(n_5692),
.Y(n_6333)
);

CKINVDCx20_ASAP7_75t_R g6334 ( 
.A(n_5963),
.Y(n_6334)
);

CKINVDCx5p33_ASAP7_75t_R g6335 ( 
.A(n_5965),
.Y(n_6335)
);

INVx1_ASAP7_75t_L g6336 ( 
.A(n_5710),
.Y(n_6336)
);

CKINVDCx5p33_ASAP7_75t_R g6337 ( 
.A(n_5969),
.Y(n_6337)
);

INVx2_ASAP7_75t_L g6338 ( 
.A(n_5636),
.Y(n_6338)
);

CKINVDCx20_ASAP7_75t_R g6339 ( 
.A(n_5559),
.Y(n_6339)
);

CKINVDCx5p33_ASAP7_75t_R g6340 ( 
.A(n_5620),
.Y(n_6340)
);

CKINVDCx5p33_ASAP7_75t_R g6341 ( 
.A(n_5621),
.Y(n_6341)
);

INVx1_ASAP7_75t_L g6342 ( 
.A(n_5711),
.Y(n_6342)
);

INVx1_ASAP7_75t_L g6343 ( 
.A(n_5645),
.Y(n_6343)
);

INVx1_ASAP7_75t_L g6344 ( 
.A(n_5689),
.Y(n_6344)
);

CKINVDCx5p33_ASAP7_75t_R g6345 ( 
.A(n_5624),
.Y(n_6345)
);

INVx1_ASAP7_75t_L g6346 ( 
.A(n_5690),
.Y(n_6346)
);

INVxp67_ASAP7_75t_SL g6347 ( 
.A(n_5546),
.Y(n_6347)
);

INVx1_ASAP7_75t_L g6348 ( 
.A(n_5740),
.Y(n_6348)
);

HB1xp67_ASAP7_75t_L g6349 ( 
.A(n_5625),
.Y(n_6349)
);

CKINVDCx5p33_ASAP7_75t_R g6350 ( 
.A(n_5628),
.Y(n_6350)
);

INVx1_ASAP7_75t_L g6351 ( 
.A(n_5659),
.Y(n_6351)
);

CKINVDCx5p33_ASAP7_75t_R g6352 ( 
.A(n_5631),
.Y(n_6352)
);

INVxp33_ASAP7_75t_SL g6353 ( 
.A(n_5560),
.Y(n_6353)
);

INVx1_ASAP7_75t_L g6354 ( 
.A(n_5659),
.Y(n_6354)
);

INVx1_ASAP7_75t_L g6355 ( 
.A(n_5659),
.Y(n_6355)
);

CKINVDCx20_ASAP7_75t_R g6356 ( 
.A(n_5635),
.Y(n_6356)
);

BUFx2_ASAP7_75t_L g6357 ( 
.A(n_5638),
.Y(n_6357)
);

INVx1_ASAP7_75t_L g6358 ( 
.A(n_5659),
.Y(n_6358)
);

CKINVDCx20_ASAP7_75t_R g6359 ( 
.A(n_5639),
.Y(n_6359)
);

CKINVDCx16_ASAP7_75t_R g6360 ( 
.A(n_5762),
.Y(n_6360)
);

CKINVDCx5p33_ASAP7_75t_R g6361 ( 
.A(n_5641),
.Y(n_6361)
);

CKINVDCx5p33_ASAP7_75t_R g6362 ( 
.A(n_5642),
.Y(n_6362)
);

INVx1_ASAP7_75t_L g6363 ( 
.A(n_5660),
.Y(n_6363)
);

INVx1_ASAP7_75t_L g6364 ( 
.A(n_5660),
.Y(n_6364)
);

INVxp67_ASAP7_75t_L g6365 ( 
.A(n_5548),
.Y(n_6365)
);

HB1xp67_ASAP7_75t_L g6366 ( 
.A(n_5643),
.Y(n_6366)
);

CKINVDCx5p33_ASAP7_75t_R g6367 ( 
.A(n_5646),
.Y(n_6367)
);

INVx1_ASAP7_75t_L g6368 ( 
.A(n_5660),
.Y(n_6368)
);

CKINVDCx5p33_ASAP7_75t_R g6369 ( 
.A(n_5649),
.Y(n_6369)
);

INVx1_ASAP7_75t_L g6370 ( 
.A(n_5660),
.Y(n_6370)
);

INVx1_ASAP7_75t_L g6371 ( 
.A(n_5704),
.Y(n_6371)
);

CKINVDCx5p33_ASAP7_75t_R g6372 ( 
.A(n_5651),
.Y(n_6372)
);

CKINVDCx5p33_ASAP7_75t_R g6373 ( 
.A(n_5652),
.Y(n_6373)
);

INVx1_ASAP7_75t_L g6374 ( 
.A(n_5704),
.Y(n_6374)
);

INVx1_ASAP7_75t_L g6375 ( 
.A(n_5704),
.Y(n_6375)
);

INVx1_ASAP7_75t_L g6376 ( 
.A(n_5704),
.Y(n_6376)
);

BUFx3_ASAP7_75t_L g6377 ( 
.A(n_5774),
.Y(n_6377)
);

INVx1_ASAP7_75t_L g6378 ( 
.A(n_5774),
.Y(n_6378)
);

INVx1_ASAP7_75t_L g6379 ( 
.A(n_5774),
.Y(n_6379)
);

CKINVDCx5p33_ASAP7_75t_R g6380 ( 
.A(n_5668),
.Y(n_6380)
);

INVx1_ASAP7_75t_L g6381 ( 
.A(n_5774),
.Y(n_6381)
);

CKINVDCx5p33_ASAP7_75t_R g6382 ( 
.A(n_5669),
.Y(n_6382)
);

INVx1_ASAP7_75t_L g6383 ( 
.A(n_5788),
.Y(n_6383)
);

CKINVDCx14_ASAP7_75t_R g6384 ( 
.A(n_5670),
.Y(n_6384)
);

INVx1_ASAP7_75t_L g6385 ( 
.A(n_5788),
.Y(n_6385)
);

INVx1_ASAP7_75t_L g6386 ( 
.A(n_5788),
.Y(n_6386)
);

INVx1_ASAP7_75t_L g6387 ( 
.A(n_5788),
.Y(n_6387)
);

INVx1_ASAP7_75t_L g6388 ( 
.A(n_5827),
.Y(n_6388)
);

INVx1_ASAP7_75t_L g6389 ( 
.A(n_5827),
.Y(n_6389)
);

CKINVDCx5p33_ASAP7_75t_R g6390 ( 
.A(n_5672),
.Y(n_6390)
);

INVxp67_ASAP7_75t_L g6391 ( 
.A(n_5550),
.Y(n_6391)
);

CKINVDCx20_ASAP7_75t_R g6392 ( 
.A(n_5673),
.Y(n_6392)
);

CKINVDCx20_ASAP7_75t_R g6393 ( 
.A(n_5675),
.Y(n_6393)
);

INVx2_ASAP7_75t_L g6394 ( 
.A(n_5827),
.Y(n_6394)
);

INVx1_ASAP7_75t_L g6395 ( 
.A(n_5827),
.Y(n_6395)
);

INVxp67_ASAP7_75t_L g6396 ( 
.A(n_5564),
.Y(n_6396)
);

INVx1_ASAP7_75t_L g6397 ( 
.A(n_5897),
.Y(n_6397)
);

INVxp67_ASAP7_75t_SL g6398 ( 
.A(n_5769),
.Y(n_6398)
);

CKINVDCx20_ASAP7_75t_R g6399 ( 
.A(n_5684),
.Y(n_6399)
);

INVx1_ASAP7_75t_L g6400 ( 
.A(n_5897),
.Y(n_6400)
);

INVx1_ASAP7_75t_L g6401 ( 
.A(n_5897),
.Y(n_6401)
);

CKINVDCx20_ASAP7_75t_R g6402 ( 
.A(n_5687),
.Y(n_6402)
);

INVx1_ASAP7_75t_L g6403 ( 
.A(n_5897),
.Y(n_6403)
);

INVxp67_ASAP7_75t_SL g6404 ( 
.A(n_5589),
.Y(n_6404)
);

CKINVDCx20_ASAP7_75t_R g6405 ( 
.A(n_5688),
.Y(n_6405)
);

BUFx2_ASAP7_75t_SL g6406 ( 
.A(n_5594),
.Y(n_6406)
);

CKINVDCx20_ASAP7_75t_R g6407 ( 
.A(n_5694),
.Y(n_6407)
);

INVx1_ASAP7_75t_L g6408 ( 
.A(n_5735),
.Y(n_6408)
);

INVx1_ASAP7_75t_L g6409 ( 
.A(n_5725),
.Y(n_6409)
);

INVx1_ASAP7_75t_L g6410 ( 
.A(n_5745),
.Y(n_6410)
);

CKINVDCx20_ASAP7_75t_R g6411 ( 
.A(n_5695),
.Y(n_6411)
);

INVx1_ASAP7_75t_L g6412 ( 
.A(n_5789),
.Y(n_6412)
);

CKINVDCx16_ASAP7_75t_R g6413 ( 
.A(n_5841),
.Y(n_6413)
);

INVx1_ASAP7_75t_L g6414 ( 
.A(n_5793),
.Y(n_6414)
);

INVx1_ASAP7_75t_L g6415 ( 
.A(n_5968),
.Y(n_6415)
);

INVx1_ASAP7_75t_L g6416 ( 
.A(n_5696),
.Y(n_6416)
);

INVx1_ASAP7_75t_L g6417 ( 
.A(n_5700),
.Y(n_6417)
);

INVx1_ASAP7_75t_L g6418 ( 
.A(n_5705),
.Y(n_6418)
);

INVx2_ASAP7_75t_L g6419 ( 
.A(n_5563),
.Y(n_6419)
);

INVx2_ASAP7_75t_L g6420 ( 
.A(n_5693),
.Y(n_6420)
);

INVxp33_ASAP7_75t_SL g6421 ( 
.A(n_5713),
.Y(n_6421)
);

INVx1_ASAP7_75t_L g6422 ( 
.A(n_5714),
.Y(n_6422)
);

INVx2_ASAP7_75t_L g6423 ( 
.A(n_5715),
.Y(n_6423)
);

INVx1_ASAP7_75t_L g6424 ( 
.A(n_5716),
.Y(n_6424)
);

INVx1_ASAP7_75t_L g6425 ( 
.A(n_5717),
.Y(n_6425)
);

INVx1_ASAP7_75t_L g6426 ( 
.A(n_5720),
.Y(n_6426)
);

HB1xp67_ASAP7_75t_L g6427 ( 
.A(n_5722),
.Y(n_6427)
);

CKINVDCx5p33_ASAP7_75t_R g6428 ( 
.A(n_5724),
.Y(n_6428)
);

INVxp67_ASAP7_75t_L g6429 ( 
.A(n_5626),
.Y(n_6429)
);

CKINVDCx5p33_ASAP7_75t_R g6430 ( 
.A(n_5726),
.Y(n_6430)
);

CKINVDCx5p33_ASAP7_75t_R g6431 ( 
.A(n_5729),
.Y(n_6431)
);

CKINVDCx20_ASAP7_75t_R g6432 ( 
.A(n_5736),
.Y(n_6432)
);

BUFx3_ASAP7_75t_L g6433 ( 
.A(n_5737),
.Y(n_6433)
);

CKINVDCx20_ASAP7_75t_R g6434 ( 
.A(n_5738),
.Y(n_6434)
);

INVx1_ASAP7_75t_L g6435 ( 
.A(n_5648),
.Y(n_6435)
);

CKINVDCx20_ASAP7_75t_R g6436 ( 
.A(n_5937),
.Y(n_6436)
);

CKINVDCx20_ASAP7_75t_R g6437 ( 
.A(n_5731),
.Y(n_6437)
);

INVx1_ASAP7_75t_L g6438 ( 
.A(n_5934),
.Y(n_6438)
);

CKINVDCx5p33_ASAP7_75t_R g6439 ( 
.A(n_5750),
.Y(n_6439)
);

INVx1_ASAP7_75t_L g6440 ( 
.A(n_5778),
.Y(n_6440)
);

INVx1_ASAP7_75t_L g6441 ( 
.A(n_5843),
.Y(n_6441)
);

INVx1_ASAP7_75t_L g6442 ( 
.A(n_5861),
.Y(n_6442)
);

INVx1_ASAP7_75t_L g6443 ( 
.A(n_5802),
.Y(n_6443)
);

INVx1_ASAP7_75t_L g6444 ( 
.A(n_5702),
.Y(n_6444)
);

INVx1_ASAP7_75t_L g6445 ( 
.A(n_5535),
.Y(n_6445)
);

INVxp33_ASAP7_75t_SL g6446 ( 
.A(n_5537),
.Y(n_6446)
);

CKINVDCx20_ASAP7_75t_R g6447 ( 
.A(n_5644),
.Y(n_6447)
);

INVx1_ASAP7_75t_L g6448 ( 
.A(n_5535),
.Y(n_6448)
);

INVx1_ASAP7_75t_L g6449 ( 
.A(n_5535),
.Y(n_6449)
);

CKINVDCx16_ASAP7_75t_R g6450 ( 
.A(n_5634),
.Y(n_6450)
);

CKINVDCx20_ASAP7_75t_R g6451 ( 
.A(n_5644),
.Y(n_6451)
);

CKINVDCx20_ASAP7_75t_R g6452 ( 
.A(n_5644),
.Y(n_6452)
);

INVx1_ASAP7_75t_L g6453 ( 
.A(n_5535),
.Y(n_6453)
);

INVx1_ASAP7_75t_L g6454 ( 
.A(n_5535),
.Y(n_6454)
);

INVx1_ASAP7_75t_L g6455 ( 
.A(n_5535),
.Y(n_6455)
);

INVx2_ASAP7_75t_L g6456 ( 
.A(n_5756),
.Y(n_6456)
);

INVxp67_ASAP7_75t_SL g6457 ( 
.A(n_5741),
.Y(n_6457)
);

INVx1_ASAP7_75t_L g6458 ( 
.A(n_5535),
.Y(n_6458)
);

HB1xp67_ASAP7_75t_L g6459 ( 
.A(n_5562),
.Y(n_6459)
);

CKINVDCx20_ASAP7_75t_R g6460 ( 
.A(n_5644),
.Y(n_6460)
);

CKINVDCx5p33_ASAP7_75t_R g6461 ( 
.A(n_5739),
.Y(n_6461)
);

INVxp67_ASAP7_75t_SL g6462 ( 
.A(n_5741),
.Y(n_6462)
);

INVx1_ASAP7_75t_L g6463 ( 
.A(n_5535),
.Y(n_6463)
);

CKINVDCx16_ASAP7_75t_R g6464 ( 
.A(n_5634),
.Y(n_6464)
);

INVxp67_ASAP7_75t_SL g6465 ( 
.A(n_5741),
.Y(n_6465)
);

CKINVDCx16_ASAP7_75t_R g6466 ( 
.A(n_5634),
.Y(n_6466)
);

CKINVDCx5p33_ASAP7_75t_R g6467 ( 
.A(n_5739),
.Y(n_6467)
);

CKINVDCx20_ASAP7_75t_R g6468 ( 
.A(n_5644),
.Y(n_6468)
);

HB1xp67_ASAP7_75t_L g6469 ( 
.A(n_5562),
.Y(n_6469)
);

CKINVDCx20_ASAP7_75t_R g6470 ( 
.A(n_5644),
.Y(n_6470)
);

HB1xp67_ASAP7_75t_L g6471 ( 
.A(n_5562),
.Y(n_6471)
);

HB1xp67_ASAP7_75t_L g6472 ( 
.A(n_5562),
.Y(n_6472)
);

INVx1_ASAP7_75t_L g6473 ( 
.A(n_5535),
.Y(n_6473)
);

CKINVDCx5p33_ASAP7_75t_R g6474 ( 
.A(n_5739),
.Y(n_6474)
);

CKINVDCx20_ASAP7_75t_R g6475 ( 
.A(n_5644),
.Y(n_6475)
);

INVx1_ASAP7_75t_L g6476 ( 
.A(n_5535),
.Y(n_6476)
);

CKINVDCx16_ASAP7_75t_R g6477 ( 
.A(n_5634),
.Y(n_6477)
);

CKINVDCx20_ASAP7_75t_R g6478 ( 
.A(n_5644),
.Y(n_6478)
);

INVx1_ASAP7_75t_L g6479 ( 
.A(n_5535),
.Y(n_6479)
);

INVx1_ASAP7_75t_L g6480 ( 
.A(n_5535),
.Y(n_6480)
);

CKINVDCx5p33_ASAP7_75t_R g6481 ( 
.A(n_5739),
.Y(n_6481)
);

INVx1_ASAP7_75t_L g6482 ( 
.A(n_5535),
.Y(n_6482)
);

INVxp67_ASAP7_75t_L g6483 ( 
.A(n_5544),
.Y(n_6483)
);

INVxp67_ASAP7_75t_L g6484 ( 
.A(n_5544),
.Y(n_6484)
);

CKINVDCx5p33_ASAP7_75t_R g6485 ( 
.A(n_5739),
.Y(n_6485)
);

BUFx6f_ASAP7_75t_L g6486 ( 
.A(n_6141),
.Y(n_6486)
);

INVx1_ASAP7_75t_L g6487 ( 
.A(n_6263),
.Y(n_6487)
);

INVx2_ASAP7_75t_L g6488 ( 
.A(n_6002),
.Y(n_6488)
);

BUFx6f_ASAP7_75t_L g6489 ( 
.A(n_6173),
.Y(n_6489)
);

BUFx8_ASAP7_75t_SL g6490 ( 
.A(n_6436),
.Y(n_6490)
);

INVx2_ASAP7_75t_L g6491 ( 
.A(n_6456),
.Y(n_6491)
);

AND2x4_ASAP7_75t_L g6492 ( 
.A(n_6179),
.B(n_4451),
.Y(n_6492)
);

BUFx6f_ASAP7_75t_L g6493 ( 
.A(n_6193),
.Y(n_6493)
);

INVx2_ASAP7_75t_L g6494 ( 
.A(n_6188),
.Y(n_6494)
);

AND2x2_ASAP7_75t_L g6495 ( 
.A(n_6406),
.B(n_5115),
.Y(n_6495)
);

INVx2_ASAP7_75t_SL g6496 ( 
.A(n_6439),
.Y(n_6496)
);

INVx2_ASAP7_75t_L g6497 ( 
.A(n_6199),
.Y(n_6497)
);

BUFx6f_ASAP7_75t_L g6498 ( 
.A(n_6338),
.Y(n_6498)
);

BUFx3_ASAP7_75t_L g6499 ( 
.A(n_6433),
.Y(n_6499)
);

BUFx8_ASAP7_75t_SL g6500 ( 
.A(n_6437),
.Y(n_6500)
);

CKINVDCx8_ASAP7_75t_R g6501 ( 
.A(n_6078),
.Y(n_6501)
);

CKINVDCx6p67_ASAP7_75t_R g6502 ( 
.A(n_6302),
.Y(n_6502)
);

NAND2xp5_ASAP7_75t_L g6503 ( 
.A(n_6196),
.B(n_5121),
.Y(n_6503)
);

INVx3_ASAP7_75t_L g6504 ( 
.A(n_6275),
.Y(n_6504)
);

AND2x4_ASAP7_75t_L g6505 ( 
.A(n_6218),
.B(n_4480),
.Y(n_6505)
);

AND2x2_ASAP7_75t_SL g6506 ( 
.A(n_6450),
.B(n_5152),
.Y(n_6506)
);

BUFx3_ASAP7_75t_L g6507 ( 
.A(n_6296),
.Y(n_6507)
);

INVx3_ASAP7_75t_L g6508 ( 
.A(n_6275),
.Y(n_6508)
);

INVx1_ASAP7_75t_L g6509 ( 
.A(n_6265),
.Y(n_6509)
);

AND2x4_ASAP7_75t_L g6510 ( 
.A(n_6222),
.B(n_4518),
.Y(n_6510)
);

INVx1_ASAP7_75t_L g6511 ( 
.A(n_6268),
.Y(n_6511)
);

INVx2_ASAP7_75t_L g6512 ( 
.A(n_6215),
.Y(n_6512)
);

OA21x2_ASAP7_75t_L g6513 ( 
.A1(n_6394),
.A2(n_4317),
.B(n_4184),
.Y(n_6513)
);

BUFx12f_ASAP7_75t_L g6514 ( 
.A(n_6238),
.Y(n_6514)
);

CKINVDCx5p33_ASAP7_75t_R g6515 ( 
.A(n_5974),
.Y(n_6515)
);

INVx2_ASAP7_75t_L g6516 ( 
.A(n_6245),
.Y(n_6516)
);

BUFx6f_ASAP7_75t_L g6517 ( 
.A(n_5980),
.Y(n_6517)
);

BUFx6f_ASAP7_75t_L g6518 ( 
.A(n_5982),
.Y(n_6518)
);

BUFx6f_ASAP7_75t_L g6519 ( 
.A(n_5983),
.Y(n_6519)
);

BUFx12f_ASAP7_75t_L g6520 ( 
.A(n_6238),
.Y(n_6520)
);

AND2x4_ASAP7_75t_L g6521 ( 
.A(n_6226),
.B(n_4532),
.Y(n_6521)
);

AND2x4_ASAP7_75t_L g6522 ( 
.A(n_6229),
.B(n_4632),
.Y(n_6522)
);

OA21x2_ASAP7_75t_L g6523 ( 
.A1(n_6351),
.A2(n_5159),
.B(n_4362),
.Y(n_6523)
);

NAND2xp5_ASAP7_75t_L g6524 ( 
.A(n_6377),
.B(n_5169),
.Y(n_6524)
);

OAI22x1_ASAP7_75t_SL g6525 ( 
.A1(n_6443),
.A2(n_5484),
.B1(n_4540),
.B2(n_4554),
.Y(n_6525)
);

BUFx3_ASAP7_75t_L g6526 ( 
.A(n_6312),
.Y(n_6526)
);

AOI22xp5_ASAP7_75t_L g6527 ( 
.A1(n_6198),
.A2(n_4179),
.B1(n_4319),
.B2(n_4147),
.Y(n_6527)
);

INVx1_ASAP7_75t_L g6528 ( 
.A(n_6269),
.Y(n_6528)
);

INVx2_ASAP7_75t_L g6529 ( 
.A(n_6251),
.Y(n_6529)
);

INVx1_ASAP7_75t_L g6530 ( 
.A(n_6270),
.Y(n_6530)
);

AND2x4_ASAP7_75t_L g6531 ( 
.A(n_5979),
.B(n_4677),
.Y(n_6531)
);

INVx1_ASAP7_75t_L g6532 ( 
.A(n_6272),
.Y(n_6532)
);

INVx1_ASAP7_75t_L g6533 ( 
.A(n_6276),
.Y(n_6533)
);

CKINVDCx5p33_ASAP7_75t_R g6534 ( 
.A(n_5975),
.Y(n_6534)
);

AND2x2_ASAP7_75t_L g6535 ( 
.A(n_6391),
.B(n_5307),
.Y(n_6535)
);

OAI22x1_ASAP7_75t_R g6536 ( 
.A1(n_6217),
.A2(n_4567),
.B1(n_4579),
.B2(n_4511),
.Y(n_6536)
);

NAND2xp5_ASAP7_75t_L g6537 ( 
.A(n_6005),
.B(n_5169),
.Y(n_6537)
);

BUFx6f_ASAP7_75t_L g6538 ( 
.A(n_5985),
.Y(n_6538)
);

BUFx6f_ASAP7_75t_L g6539 ( 
.A(n_5987),
.Y(n_6539)
);

AND2x2_ASAP7_75t_L g6540 ( 
.A(n_6396),
.B(n_5345),
.Y(n_6540)
);

AND2x4_ASAP7_75t_L g6541 ( 
.A(n_6022),
.B(n_4696),
.Y(n_6541)
);

INVx2_ASAP7_75t_L g6542 ( 
.A(n_6303),
.Y(n_6542)
);

NOR2x1_ASAP7_75t_L g6543 ( 
.A(n_6416),
.B(n_4723),
.Y(n_6543)
);

BUFx8_ASAP7_75t_L g6544 ( 
.A(n_6302),
.Y(n_6544)
);

INVx2_ASAP7_75t_L g6545 ( 
.A(n_6037),
.Y(n_6545)
);

NOR2xp33_ASAP7_75t_L g6546 ( 
.A(n_6064),
.B(n_5371),
.Y(n_6546)
);

INVx2_ASAP7_75t_L g6547 ( 
.A(n_6070),
.Y(n_6547)
);

INVx1_ASAP7_75t_L g6548 ( 
.A(n_6287),
.Y(n_6548)
);

AND2x2_ASAP7_75t_L g6549 ( 
.A(n_6429),
.B(n_4584),
.Y(n_6549)
);

AND2x2_ASAP7_75t_L g6550 ( 
.A(n_6365),
.B(n_4593),
.Y(n_6550)
);

INVx2_ASAP7_75t_L g6551 ( 
.A(n_6079),
.Y(n_6551)
);

BUFx6f_ASAP7_75t_L g6552 ( 
.A(n_5988),
.Y(n_6552)
);

OAI21x1_ASAP7_75t_L g6553 ( 
.A1(n_6354),
.A2(n_4173),
.B(n_4161),
.Y(n_6553)
);

INVx1_ASAP7_75t_L g6554 ( 
.A(n_6293),
.Y(n_6554)
);

AND2x2_ASAP7_75t_L g6555 ( 
.A(n_6440),
.B(n_4593),
.Y(n_6555)
);

INVx1_ASAP7_75t_L g6556 ( 
.A(n_6298),
.Y(n_6556)
);

AND2x2_ASAP7_75t_L g6557 ( 
.A(n_6441),
.B(n_4605),
.Y(n_6557)
);

AND2x2_ASAP7_75t_L g6558 ( 
.A(n_6442),
.B(n_4605),
.Y(n_6558)
);

HB1xp67_ASAP7_75t_L g6559 ( 
.A(n_6058),
.Y(n_6559)
);

INVx1_ASAP7_75t_L g6560 ( 
.A(n_6300),
.Y(n_6560)
);

BUFx6f_ASAP7_75t_L g6561 ( 
.A(n_5992),
.Y(n_6561)
);

INVx1_ASAP7_75t_L g6562 ( 
.A(n_6301),
.Y(n_6562)
);

INVx6_ASAP7_75t_L g6563 ( 
.A(n_6164),
.Y(n_6563)
);

INVxp33_ASAP7_75t_SL g6564 ( 
.A(n_6080),
.Y(n_6564)
);

BUFx6f_ASAP7_75t_L g6565 ( 
.A(n_5993),
.Y(n_6565)
);

BUFx6f_ASAP7_75t_L g6566 ( 
.A(n_5997),
.Y(n_6566)
);

INVx5_ASAP7_75t_L g6567 ( 
.A(n_6178),
.Y(n_6567)
);

CKINVDCx5p33_ASAP7_75t_R g6568 ( 
.A(n_5981),
.Y(n_6568)
);

BUFx6f_ASAP7_75t_L g6569 ( 
.A(n_5999),
.Y(n_6569)
);

AND2x4_ASAP7_75t_L g6570 ( 
.A(n_6074),
.B(n_4752),
.Y(n_6570)
);

BUFx3_ASAP7_75t_L g6571 ( 
.A(n_6315),
.Y(n_6571)
);

AND2x2_ASAP7_75t_L g6572 ( 
.A(n_6347),
.B(n_4650),
.Y(n_6572)
);

BUFx6f_ASAP7_75t_L g6573 ( 
.A(n_6003),
.Y(n_6573)
);

INVx3_ASAP7_75t_L g6574 ( 
.A(n_6004),
.Y(n_6574)
);

INVx2_ASAP7_75t_L g6575 ( 
.A(n_6097),
.Y(n_6575)
);

BUFx6f_ASAP7_75t_L g6576 ( 
.A(n_5971),
.Y(n_6576)
);

INVx4_ASAP7_75t_L g6577 ( 
.A(n_5984),
.Y(n_6577)
);

INVxp33_ASAP7_75t_SL g6578 ( 
.A(n_6108),
.Y(n_6578)
);

NAND2xp5_ASAP7_75t_L g6579 ( 
.A(n_6005),
.B(n_5169),
.Y(n_6579)
);

NOR2x1_ASAP7_75t_L g6580 ( 
.A(n_6417),
.B(n_6418),
.Y(n_6580)
);

BUFx3_ASAP7_75t_L g6581 ( 
.A(n_6325),
.Y(n_6581)
);

CKINVDCx6p67_ASAP7_75t_R g6582 ( 
.A(n_6233),
.Y(n_6582)
);

CKINVDCx5p33_ASAP7_75t_R g6583 ( 
.A(n_5989),
.Y(n_6583)
);

INVx1_ASAP7_75t_L g6584 ( 
.A(n_6305),
.Y(n_6584)
);

AND2x2_ASAP7_75t_L g6585 ( 
.A(n_6231),
.B(n_4650),
.Y(n_6585)
);

INVx2_ASAP7_75t_L g6586 ( 
.A(n_6120),
.Y(n_6586)
);

INVx1_ASAP7_75t_L g6587 ( 
.A(n_6310),
.Y(n_6587)
);

AND2x2_ASAP7_75t_L g6588 ( 
.A(n_6237),
.B(n_6404),
.Y(n_6588)
);

INVx1_ASAP7_75t_L g6589 ( 
.A(n_6311),
.Y(n_6589)
);

CKINVDCx6p67_ASAP7_75t_R g6590 ( 
.A(n_6260),
.Y(n_6590)
);

BUFx6f_ASAP7_75t_L g6591 ( 
.A(n_5972),
.Y(n_6591)
);

INVx2_ASAP7_75t_L g6592 ( 
.A(n_6127),
.Y(n_6592)
);

OA21x2_ASAP7_75t_L g6593 ( 
.A1(n_6355),
.A2(n_4822),
.B(n_4778),
.Y(n_6593)
);

INVx1_ASAP7_75t_L g6594 ( 
.A(n_6313),
.Y(n_6594)
);

HB1xp67_ASAP7_75t_L g6595 ( 
.A(n_6041),
.Y(n_6595)
);

OAI22xp5_ASAP7_75t_SL g6596 ( 
.A1(n_6225),
.A2(n_4590),
.B1(n_4601),
.B2(n_4581),
.Y(n_6596)
);

INVx1_ASAP7_75t_L g6597 ( 
.A(n_6314),
.Y(n_6597)
);

BUFx6f_ASAP7_75t_L g6598 ( 
.A(n_5973),
.Y(n_6598)
);

INVx3_ASAP7_75t_L g6599 ( 
.A(n_5976),
.Y(n_6599)
);

BUFx12f_ASAP7_75t_L g6600 ( 
.A(n_6340),
.Y(n_6600)
);

INVx2_ASAP7_75t_SL g6601 ( 
.A(n_6420),
.Y(n_6601)
);

BUFx2_ASAP7_75t_L g6602 ( 
.A(n_6254),
.Y(n_6602)
);

INVx2_ASAP7_75t_L g6603 ( 
.A(n_6006),
.Y(n_6603)
);

CKINVDCx5p33_ASAP7_75t_R g6604 ( 
.A(n_5991),
.Y(n_6604)
);

AOI22xp5_ASAP7_75t_L g6605 ( 
.A1(n_6398),
.A2(n_4336),
.B1(n_4357),
.B2(n_4330),
.Y(n_6605)
);

AND2x4_ASAP7_75t_L g6606 ( 
.A(n_6075),
.B(n_4791),
.Y(n_6606)
);

INVx3_ASAP7_75t_L g6607 ( 
.A(n_5977),
.Y(n_6607)
);

CKINVDCx5p33_ASAP7_75t_R g6608 ( 
.A(n_5994),
.Y(n_6608)
);

CKINVDCx5p33_ASAP7_75t_R g6609 ( 
.A(n_5996),
.Y(n_6609)
);

OAI22x1_ASAP7_75t_SL g6610 ( 
.A1(n_6444),
.A2(n_4615),
.B1(n_4617),
.B2(n_4614),
.Y(n_6610)
);

BUFx6f_ASAP7_75t_L g6611 ( 
.A(n_5978),
.Y(n_6611)
);

OA21x2_ASAP7_75t_L g6612 ( 
.A1(n_6358),
.A2(n_4959),
.B(n_4931),
.Y(n_6612)
);

INVx1_ASAP7_75t_L g6613 ( 
.A(n_6316),
.Y(n_6613)
);

INVx1_ASAP7_75t_L g6614 ( 
.A(n_6319),
.Y(n_6614)
);

INVx1_ASAP7_75t_L g6615 ( 
.A(n_6321),
.Y(n_6615)
);

INVx1_ASAP7_75t_L g6616 ( 
.A(n_6323),
.Y(n_6616)
);

INVx1_ASAP7_75t_L g6617 ( 
.A(n_6327),
.Y(n_6617)
);

INVx5_ASAP7_75t_L g6618 ( 
.A(n_5995),
.Y(n_6618)
);

INVx1_ASAP7_75t_L g6619 ( 
.A(n_6328),
.Y(n_6619)
);

AOI22xp5_ASAP7_75t_L g6620 ( 
.A1(n_6422),
.A2(n_4409),
.B1(n_4501),
.B2(n_4359),
.Y(n_6620)
);

BUFx12f_ASAP7_75t_L g6621 ( 
.A(n_6341),
.Y(n_6621)
);

AND2x2_ASAP7_75t_L g6622 ( 
.A(n_6126),
.B(n_6299),
.Y(n_6622)
);

NAND2xp5_ASAP7_75t_L g6623 ( 
.A(n_6005),
.B(n_5190),
.Y(n_6623)
);

INVx2_ASAP7_75t_L g6624 ( 
.A(n_6007),
.Y(n_6624)
);

HB1xp67_ASAP7_75t_L g6625 ( 
.A(n_6200),
.Y(n_6625)
);

OAI21x1_ASAP7_75t_L g6626 ( 
.A1(n_6363),
.A2(n_4189),
.B(n_4175),
.Y(n_6626)
);

AOI22xp5_ASAP7_75t_L g6627 ( 
.A1(n_6424),
.A2(n_4609),
.B1(n_4674),
.B2(n_4570),
.Y(n_6627)
);

NAND2xp5_ASAP7_75t_L g6628 ( 
.A(n_6005),
.B(n_5190),
.Y(n_6628)
);

AND2x2_ASAP7_75t_L g6629 ( 
.A(n_6384),
.B(n_4714),
.Y(n_6629)
);

INVx1_ASAP7_75t_L g6630 ( 
.A(n_6329),
.Y(n_6630)
);

NOR2xp33_ASAP7_75t_SL g6631 ( 
.A(n_6421),
.B(n_4623),
.Y(n_6631)
);

AND2x4_ASAP7_75t_L g6632 ( 
.A(n_6113),
.B(n_4815),
.Y(n_6632)
);

INVx1_ASAP7_75t_L g6633 ( 
.A(n_6332),
.Y(n_6633)
);

OAI21x1_ASAP7_75t_L g6634 ( 
.A1(n_6364),
.A2(n_4278),
.B(n_4196),
.Y(n_6634)
);

INVx1_ASAP7_75t_L g6635 ( 
.A(n_6336),
.Y(n_6635)
);

BUFx6f_ASAP7_75t_L g6636 ( 
.A(n_6445),
.Y(n_6636)
);

BUFx6f_ASAP7_75t_L g6637 ( 
.A(n_6448),
.Y(n_6637)
);

BUFx12f_ASAP7_75t_L g6638 ( 
.A(n_6345),
.Y(n_6638)
);

INVx2_ASAP7_75t_L g6639 ( 
.A(n_6008),
.Y(n_6639)
);

NAND2xp5_ASAP7_75t_L g6640 ( 
.A(n_6005),
.B(n_5190),
.Y(n_6640)
);

INVx2_ASAP7_75t_L g6641 ( 
.A(n_6348),
.Y(n_6641)
);

INVx5_ASAP7_75t_L g6642 ( 
.A(n_6220),
.Y(n_6642)
);

HB1xp67_ASAP7_75t_L g6643 ( 
.A(n_6207),
.Y(n_6643)
);

BUFx2_ASAP7_75t_L g6644 ( 
.A(n_6266),
.Y(n_6644)
);

AOI22xp5_ASAP7_75t_L g6645 ( 
.A1(n_6425),
.A2(n_4705),
.B1(n_4736),
.B2(n_4687),
.Y(n_6645)
);

BUFx8_ASAP7_75t_SL g6646 ( 
.A(n_5970),
.Y(n_6646)
);

INVx2_ASAP7_75t_L g6647 ( 
.A(n_6031),
.Y(n_6647)
);

BUFx6f_ASAP7_75t_L g6648 ( 
.A(n_6449),
.Y(n_6648)
);

INVx1_ASAP7_75t_L g6649 ( 
.A(n_6342),
.Y(n_6649)
);

INVx2_ASAP7_75t_L g6650 ( 
.A(n_6034),
.Y(n_6650)
);

INVx5_ASAP7_75t_L g6651 ( 
.A(n_6286),
.Y(n_6651)
);

INVx1_ASAP7_75t_L g6652 ( 
.A(n_6174),
.Y(n_6652)
);

BUFx6f_ASAP7_75t_L g6653 ( 
.A(n_6453),
.Y(n_6653)
);

HB1xp67_ASAP7_75t_L g6654 ( 
.A(n_6211),
.Y(n_6654)
);

AND2x4_ASAP7_75t_L g6655 ( 
.A(n_6191),
.B(n_4818),
.Y(n_6655)
);

BUFx12f_ASAP7_75t_L g6656 ( 
.A(n_6350),
.Y(n_6656)
);

AND2x4_ASAP7_75t_L g6657 ( 
.A(n_6457),
.B(n_4829),
.Y(n_6657)
);

INVx2_ASAP7_75t_L g6658 ( 
.A(n_6035),
.Y(n_6658)
);

HB1xp67_ASAP7_75t_L g6659 ( 
.A(n_6223),
.Y(n_6659)
);

BUFx3_ASAP7_75t_L g6660 ( 
.A(n_6334),
.Y(n_6660)
);

INVx1_ASAP7_75t_L g6661 ( 
.A(n_6175),
.Y(n_6661)
);

AND2x2_ASAP7_75t_L g6662 ( 
.A(n_6165),
.B(n_6282),
.Y(n_6662)
);

INVx1_ASAP7_75t_L g6663 ( 
.A(n_6176),
.Y(n_6663)
);

CKINVDCx8_ASAP7_75t_R g6664 ( 
.A(n_6464),
.Y(n_6664)
);

INVx2_ASAP7_75t_L g6665 ( 
.A(n_6039),
.Y(n_6665)
);

INVx2_ASAP7_75t_L g6666 ( 
.A(n_6042),
.Y(n_6666)
);

INVx3_ASAP7_75t_L g6667 ( 
.A(n_6454),
.Y(n_6667)
);

INVx2_ASAP7_75t_L g6668 ( 
.A(n_6044),
.Y(n_6668)
);

CKINVDCx20_ASAP7_75t_R g6669 ( 
.A(n_5986),
.Y(n_6669)
);

BUFx6f_ASAP7_75t_L g6670 ( 
.A(n_6455),
.Y(n_6670)
);

INVx1_ASAP7_75t_L g6671 ( 
.A(n_6182),
.Y(n_6671)
);

AOI22x1_ASAP7_75t_SL g6672 ( 
.A1(n_5998),
.A2(n_4712),
.B1(n_4729),
.B2(n_4641),
.Y(n_6672)
);

BUFx6f_ASAP7_75t_L g6673 ( 
.A(n_6458),
.Y(n_6673)
);

INVx2_ASAP7_75t_L g6674 ( 
.A(n_6046),
.Y(n_6674)
);

INVx1_ASAP7_75t_L g6675 ( 
.A(n_6183),
.Y(n_6675)
);

AND2x4_ASAP7_75t_L g6676 ( 
.A(n_6462),
.B(n_4862),
.Y(n_6676)
);

INVx1_ASAP7_75t_L g6677 ( 
.A(n_6184),
.Y(n_6677)
);

INVx2_ASAP7_75t_SL g6678 ( 
.A(n_6419),
.Y(n_6678)
);

OAI22x1_ASAP7_75t_R g6679 ( 
.A1(n_6013),
.A2(n_4735),
.B1(n_4789),
.B2(n_4734),
.Y(n_6679)
);

INVx1_ASAP7_75t_L g6680 ( 
.A(n_6185),
.Y(n_6680)
);

BUFx6f_ASAP7_75t_L g6681 ( 
.A(n_6463),
.Y(n_6681)
);

OAI22xp5_ASAP7_75t_L g6682 ( 
.A1(n_6426),
.A2(n_5341),
.B1(n_4247),
.B2(n_4255),
.Y(n_6682)
);

INVx2_ASAP7_75t_L g6683 ( 
.A(n_6047),
.Y(n_6683)
);

INVx2_ASAP7_75t_L g6684 ( 
.A(n_6050),
.Y(n_6684)
);

INVx2_ASAP7_75t_L g6685 ( 
.A(n_6052),
.Y(n_6685)
);

INVx5_ASAP7_75t_L g6686 ( 
.A(n_6333),
.Y(n_6686)
);

NAND2xp5_ASAP7_75t_L g6687 ( 
.A(n_6186),
.B(n_5229),
.Y(n_6687)
);

OAI21x1_ASAP7_75t_L g6688 ( 
.A1(n_6368),
.A2(n_6371),
.B(n_6370),
.Y(n_6688)
);

NAND2xp5_ASAP7_75t_L g6689 ( 
.A(n_6187),
.B(n_6189),
.Y(n_6689)
);

CKINVDCx16_ASAP7_75t_R g6690 ( 
.A(n_6466),
.Y(n_6690)
);

AND2x2_ASAP7_75t_L g6691 ( 
.A(n_6324),
.B(n_4714),
.Y(n_6691)
);

BUFx6f_ASAP7_75t_L g6692 ( 
.A(n_6473),
.Y(n_6692)
);

NAND2xp5_ASAP7_75t_L g6693 ( 
.A(n_6190),
.B(n_5229),
.Y(n_6693)
);

CKINVDCx5p33_ASAP7_75t_R g6694 ( 
.A(n_6000),
.Y(n_6694)
);

INVxp67_ASAP7_75t_L g6695 ( 
.A(n_6438),
.Y(n_6695)
);

INVx1_ASAP7_75t_L g6696 ( 
.A(n_6195),
.Y(n_6696)
);

NOR2x1_ASAP7_75t_L g6697 ( 
.A(n_6423),
.B(n_4866),
.Y(n_6697)
);

AOI22xp5_ASAP7_75t_L g6698 ( 
.A1(n_6326),
.A2(n_4781),
.B1(n_4843),
.B2(n_4751),
.Y(n_6698)
);

INVx2_ASAP7_75t_SL g6699 ( 
.A(n_6435),
.Y(n_6699)
);

INVx2_ASAP7_75t_L g6700 ( 
.A(n_6054),
.Y(n_6700)
);

INVx2_ASAP7_75t_L g6701 ( 
.A(n_6055),
.Y(n_6701)
);

AND2x4_ASAP7_75t_L g6702 ( 
.A(n_6465),
.B(n_4871),
.Y(n_6702)
);

BUFx6f_ASAP7_75t_L g6703 ( 
.A(n_6476),
.Y(n_6703)
);

AND2x2_ASAP7_75t_L g6704 ( 
.A(n_6357),
.B(n_4780),
.Y(n_6704)
);

NAND2xp5_ASAP7_75t_L g6705 ( 
.A(n_6197),
.B(n_5229),
.Y(n_6705)
);

AND2x2_ASAP7_75t_L g6706 ( 
.A(n_6306),
.B(n_4780),
.Y(n_6706)
);

INVx1_ASAP7_75t_L g6707 ( 
.A(n_6202),
.Y(n_6707)
);

INVx2_ASAP7_75t_L g6708 ( 
.A(n_6056),
.Y(n_6708)
);

INVx2_ASAP7_75t_L g6709 ( 
.A(n_6057),
.Y(n_6709)
);

OAI22xp5_ASAP7_75t_L g6710 ( 
.A1(n_6040),
.A2(n_4248),
.B1(n_4261),
.B2(n_4259),
.Y(n_6710)
);

BUFx6f_ASAP7_75t_L g6711 ( 
.A(n_6479),
.Y(n_6711)
);

INVx3_ASAP7_75t_L g6712 ( 
.A(n_6480),
.Y(n_6712)
);

INVx2_ASAP7_75t_L g6713 ( 
.A(n_6059),
.Y(n_6713)
);

CKINVDCx5p33_ASAP7_75t_R g6714 ( 
.A(n_6010),
.Y(n_6714)
);

AND2x2_ASAP7_75t_L g6715 ( 
.A(n_6409),
.B(n_4941),
.Y(n_6715)
);

NAND2xp5_ASAP7_75t_L g6716 ( 
.A(n_6205),
.B(n_5244),
.Y(n_6716)
);

AND2x2_ASAP7_75t_L g6717 ( 
.A(n_6410),
.B(n_4941),
.Y(n_6717)
);

INVx5_ASAP7_75t_L g6718 ( 
.A(n_6360),
.Y(n_6718)
);

OA21x2_ASAP7_75t_L g6719 ( 
.A1(n_6374),
.A2(n_4127),
.B(n_4123),
.Y(n_6719)
);

INVx1_ASAP7_75t_L g6720 ( 
.A(n_6206),
.Y(n_6720)
);

BUFx6f_ASAP7_75t_L g6721 ( 
.A(n_6482),
.Y(n_6721)
);

NAND2xp5_ASAP7_75t_L g6722 ( 
.A(n_6208),
.B(n_5244),
.Y(n_6722)
);

INVxp33_ASAP7_75t_SL g6723 ( 
.A(n_6014),
.Y(n_6723)
);

INVx1_ASAP7_75t_L g6724 ( 
.A(n_6209),
.Y(n_6724)
);

BUFx6f_ASAP7_75t_L g6725 ( 
.A(n_6408),
.Y(n_6725)
);

CKINVDCx5p33_ASAP7_75t_R g6726 ( 
.A(n_6018),
.Y(n_6726)
);

INVx2_ASAP7_75t_L g6727 ( 
.A(n_6062),
.Y(n_6727)
);

BUFx6f_ASAP7_75t_L g6728 ( 
.A(n_6063),
.Y(n_6728)
);

INVx2_ASAP7_75t_L g6729 ( 
.A(n_6065),
.Y(n_6729)
);

NAND2xp5_ASAP7_75t_L g6730 ( 
.A(n_6210),
.B(n_5244),
.Y(n_6730)
);

INVx2_ASAP7_75t_L g6731 ( 
.A(n_6067),
.Y(n_6731)
);

AND2x6_ASAP7_75t_L g6732 ( 
.A(n_6412),
.B(n_4888),
.Y(n_6732)
);

INVx2_ASAP7_75t_L g6733 ( 
.A(n_6069),
.Y(n_6733)
);

BUFx6f_ASAP7_75t_L g6734 ( 
.A(n_6072),
.Y(n_6734)
);

BUFx3_ASAP7_75t_L g6735 ( 
.A(n_6356),
.Y(n_6735)
);

INVx1_ASAP7_75t_L g6736 ( 
.A(n_6212),
.Y(n_6736)
);

INVx5_ASAP7_75t_L g6737 ( 
.A(n_6413),
.Y(n_6737)
);

NAND2xp5_ASAP7_75t_SL g6738 ( 
.A(n_6027),
.B(n_5295),
.Y(n_6738)
);

INVx3_ASAP7_75t_L g6739 ( 
.A(n_6213),
.Y(n_6739)
);

INVx1_ASAP7_75t_L g6740 ( 
.A(n_6214),
.Y(n_6740)
);

BUFx8_ASAP7_75t_SL g6741 ( 
.A(n_6020),
.Y(n_6741)
);

AND2x6_ASAP7_75t_L g6742 ( 
.A(n_6414),
.B(n_4895),
.Y(n_6742)
);

INVx4_ASAP7_75t_L g6743 ( 
.A(n_6029),
.Y(n_6743)
);

HB1xp67_ASAP7_75t_L g6744 ( 
.A(n_6228),
.Y(n_6744)
);

BUFx6f_ASAP7_75t_L g6745 ( 
.A(n_6073),
.Y(n_6745)
);

INVx1_ASAP7_75t_L g6746 ( 
.A(n_6219),
.Y(n_6746)
);

INVx2_ASAP7_75t_L g6747 ( 
.A(n_6081),
.Y(n_6747)
);

CKINVDCx5p33_ASAP7_75t_R g6748 ( 
.A(n_6036),
.Y(n_6748)
);

AND2x2_ASAP7_75t_L g6749 ( 
.A(n_6415),
.B(n_4994),
.Y(n_6749)
);

INVx2_ASAP7_75t_L g6750 ( 
.A(n_6083),
.Y(n_6750)
);

INVx1_ASAP7_75t_L g6751 ( 
.A(n_6224),
.Y(n_6751)
);

OAI21x1_ASAP7_75t_L g6752 ( 
.A1(n_6375),
.A2(n_4308),
.B(n_4282),
.Y(n_6752)
);

AND2x2_ASAP7_75t_L g6753 ( 
.A(n_6247),
.B(n_4994),
.Y(n_6753)
);

INVx2_ASAP7_75t_L g6754 ( 
.A(n_6084),
.Y(n_6754)
);

NOR2xp33_ASAP7_75t_L g6755 ( 
.A(n_6038),
.B(n_4229),
.Y(n_6755)
);

AND2x4_ASAP7_75t_L g6756 ( 
.A(n_6261),
.B(n_4904),
.Y(n_6756)
);

BUFx6f_ASAP7_75t_L g6757 ( 
.A(n_6088),
.Y(n_6757)
);

CKINVDCx5p33_ASAP7_75t_R g6758 ( 
.A(n_6045),
.Y(n_6758)
);

INVx6_ASAP7_75t_L g6759 ( 
.A(n_6477),
.Y(n_6759)
);

INVx1_ASAP7_75t_L g6760 ( 
.A(n_6230),
.Y(n_6760)
);

NAND2xp5_ASAP7_75t_L g6761 ( 
.A(n_6232),
.B(n_5295),
.Y(n_6761)
);

INVx2_ASAP7_75t_L g6762 ( 
.A(n_6089),
.Y(n_6762)
);

NAND2xp5_ASAP7_75t_L g6763 ( 
.A(n_6234),
.B(n_5295),
.Y(n_6763)
);

OAI22xp5_ASAP7_75t_L g6764 ( 
.A1(n_6483),
.A2(n_4264),
.B1(n_4268),
.B2(n_4262),
.Y(n_6764)
);

INVx2_ASAP7_75t_L g6765 ( 
.A(n_6090),
.Y(n_6765)
);

BUFx6f_ASAP7_75t_L g6766 ( 
.A(n_6091),
.Y(n_6766)
);

OAI21x1_ASAP7_75t_L g6767 ( 
.A1(n_6376),
.A2(n_4396),
.B(n_4346),
.Y(n_6767)
);

NAND2xp5_ASAP7_75t_L g6768 ( 
.A(n_6241),
.B(n_5306),
.Y(n_6768)
);

BUFx6f_ASAP7_75t_L g6769 ( 
.A(n_6093),
.Y(n_6769)
);

BUFx6f_ASAP7_75t_L g6770 ( 
.A(n_6094),
.Y(n_6770)
);

AND2x4_ASAP7_75t_L g6771 ( 
.A(n_6273),
.B(n_5132),
.Y(n_6771)
);

HB1xp67_ASAP7_75t_L g6772 ( 
.A(n_6484),
.Y(n_6772)
);

AOI22x1_ASAP7_75t_SL g6773 ( 
.A1(n_6033),
.A2(n_4809),
.B1(n_4812),
.B2(n_4793),
.Y(n_6773)
);

INVx2_ASAP7_75t_L g6774 ( 
.A(n_6098),
.Y(n_6774)
);

HB1xp67_ASAP7_75t_L g6775 ( 
.A(n_6118),
.Y(n_6775)
);

INVx1_ASAP7_75t_L g6776 ( 
.A(n_6242),
.Y(n_6776)
);

INVx1_ASAP7_75t_L g6777 ( 
.A(n_6243),
.Y(n_6777)
);

INVx3_ASAP7_75t_L g6778 ( 
.A(n_6246),
.Y(n_6778)
);

AND2x4_ASAP7_75t_L g6779 ( 
.A(n_6281),
.B(n_5243),
.Y(n_6779)
);

NOR2xp33_ASAP7_75t_L g6780 ( 
.A(n_6049),
.B(n_6051),
.Y(n_6780)
);

OAI21x1_ASAP7_75t_L g6781 ( 
.A1(n_6378),
.A2(n_4417),
.B(n_4404),
.Y(n_6781)
);

OA21x2_ASAP7_75t_L g6782 ( 
.A1(n_6379),
.A2(n_4129),
.B(n_4128),
.Y(n_6782)
);

BUFx6f_ASAP7_75t_L g6783 ( 
.A(n_6099),
.Y(n_6783)
);

BUFx6f_ASAP7_75t_L g6784 ( 
.A(n_6104),
.Y(n_6784)
);

INVx1_ASAP7_75t_L g6785 ( 
.A(n_6248),
.Y(n_6785)
);

INVx1_ASAP7_75t_L g6786 ( 
.A(n_6250),
.Y(n_6786)
);

INVx1_ASAP7_75t_L g6787 ( 
.A(n_6253),
.Y(n_6787)
);

INVx2_ASAP7_75t_L g6788 ( 
.A(n_6106),
.Y(n_6788)
);

INVx3_ASAP7_75t_L g6789 ( 
.A(n_6255),
.Y(n_6789)
);

INVx3_ASAP7_75t_L g6790 ( 
.A(n_6256),
.Y(n_6790)
);

OAI22xp5_ASAP7_75t_SL g6791 ( 
.A1(n_6267),
.A2(n_4828),
.B1(n_4848),
.B2(n_4819),
.Y(n_6791)
);

INVx2_ASAP7_75t_L g6792 ( 
.A(n_6107),
.Y(n_6792)
);

AOI22xp5_ASAP7_75t_L g6793 ( 
.A1(n_6295),
.A2(n_4967),
.B1(n_4972),
.B2(n_4846),
.Y(n_6793)
);

OAI21x1_ASAP7_75t_L g6794 ( 
.A1(n_6381),
.A2(n_4439),
.B(n_4432),
.Y(n_6794)
);

AND2x2_ASAP7_75t_L g6795 ( 
.A(n_6264),
.B(n_4999),
.Y(n_6795)
);

NAND2xp5_ASAP7_75t_L g6796 ( 
.A(n_6258),
.B(n_5306),
.Y(n_6796)
);

INVx2_ASAP7_75t_L g6797 ( 
.A(n_6109),
.Y(n_6797)
);

OAI21x1_ASAP7_75t_L g6798 ( 
.A1(n_6383),
.A2(n_4489),
.B(n_4463),
.Y(n_6798)
);

CKINVDCx20_ASAP7_75t_R g6799 ( 
.A(n_6043),
.Y(n_6799)
);

INVx2_ASAP7_75t_L g6800 ( 
.A(n_6111),
.Y(n_6800)
);

BUFx3_ASAP7_75t_L g6801 ( 
.A(n_6359),
.Y(n_6801)
);

CKINVDCx11_ASAP7_75t_R g6802 ( 
.A(n_6053),
.Y(n_6802)
);

INVx1_ASAP7_75t_L g6803 ( 
.A(n_6259),
.Y(n_6803)
);

INVx2_ASAP7_75t_L g6804 ( 
.A(n_6112),
.Y(n_6804)
);

BUFx6f_ASAP7_75t_L g6805 ( 
.A(n_6115),
.Y(n_6805)
);

BUFx3_ASAP7_75t_L g6806 ( 
.A(n_6392),
.Y(n_6806)
);

INVx1_ASAP7_75t_L g6807 ( 
.A(n_6385),
.Y(n_6807)
);

NAND2xp5_ASAP7_75t_L g6808 ( 
.A(n_6386),
.B(n_5306),
.Y(n_6808)
);

INVx1_ASAP7_75t_L g6809 ( 
.A(n_6387),
.Y(n_6809)
);

BUFx12f_ASAP7_75t_L g6810 ( 
.A(n_6352),
.Y(n_6810)
);

CKINVDCx5p33_ASAP7_75t_R g6811 ( 
.A(n_6060),
.Y(n_6811)
);

INVx2_ASAP7_75t_L g6812 ( 
.A(n_6117),
.Y(n_6812)
);

CKINVDCx16_ASAP7_75t_R g6813 ( 
.A(n_6122),
.Y(n_6813)
);

AND2x2_ASAP7_75t_L g6814 ( 
.A(n_6304),
.B(n_4999),
.Y(n_6814)
);

BUFx3_ASAP7_75t_L g6815 ( 
.A(n_6393),
.Y(n_6815)
);

INVx3_ASAP7_75t_L g6816 ( 
.A(n_6119),
.Y(n_6816)
);

AND2x2_ASAP7_75t_L g6817 ( 
.A(n_6288),
.B(n_5012),
.Y(n_6817)
);

INVx2_ASAP7_75t_L g6818 ( 
.A(n_6121),
.Y(n_6818)
);

NAND2xp5_ASAP7_75t_L g6819 ( 
.A(n_6388),
.B(n_5368),
.Y(n_6819)
);

INVx2_ASAP7_75t_L g6820 ( 
.A(n_6123),
.Y(n_6820)
);

BUFx6f_ASAP7_75t_L g6821 ( 
.A(n_6124),
.Y(n_6821)
);

HB1xp67_ASAP7_75t_L g6822 ( 
.A(n_6085),
.Y(n_6822)
);

INVx5_ASAP7_75t_L g6823 ( 
.A(n_6030),
.Y(n_6823)
);

AND2x2_ASAP7_75t_L g6824 ( 
.A(n_6116),
.B(n_5012),
.Y(n_6824)
);

BUFx2_ASAP7_75t_L g6825 ( 
.A(n_6271),
.Y(n_6825)
);

OAI22xp5_ASAP7_75t_L g6826 ( 
.A1(n_6308),
.A2(n_6322),
.B1(n_6309),
.B2(n_6349),
.Y(n_6826)
);

BUFx6f_ASAP7_75t_L g6827 ( 
.A(n_6128),
.Y(n_6827)
);

NAND2xp5_ASAP7_75t_L g6828 ( 
.A(n_6389),
.B(n_6395),
.Y(n_6828)
);

OAI22x1_ASAP7_75t_SL g6829 ( 
.A1(n_6061),
.A2(n_4873),
.B1(n_4906),
.B2(n_4850),
.Y(n_6829)
);

INVx6_ASAP7_75t_L g6830 ( 
.A(n_6131),
.Y(n_6830)
);

OA21x2_ASAP7_75t_L g6831 ( 
.A1(n_6397),
.A2(n_4135),
.B(n_4134),
.Y(n_6831)
);

BUFx6f_ASAP7_75t_L g6832 ( 
.A(n_6129),
.Y(n_6832)
);

AND2x4_ASAP7_75t_L g6833 ( 
.A(n_6133),
.B(n_5281),
.Y(n_6833)
);

NAND2xp5_ASAP7_75t_L g6834 ( 
.A(n_6400),
.B(n_5368),
.Y(n_6834)
);

BUFx6f_ASAP7_75t_L g6835 ( 
.A(n_6130),
.Y(n_6835)
);

AND2x2_ASAP7_75t_L g6836 ( 
.A(n_6137),
.B(n_5023),
.Y(n_6836)
);

BUFx2_ASAP7_75t_L g6837 ( 
.A(n_6283),
.Y(n_6837)
);

OAI22xp5_ASAP7_75t_L g6838 ( 
.A1(n_6366),
.A2(n_4279),
.B1(n_4285),
.B2(n_4271),
.Y(n_6838)
);

AND2x4_ASAP7_75t_L g6839 ( 
.A(n_6427),
.B(n_5405),
.Y(n_6839)
);

INVx2_ASAP7_75t_L g6840 ( 
.A(n_6132),
.Y(n_6840)
);

NOR2xp33_ASAP7_75t_SL g6841 ( 
.A(n_6361),
.B(n_4934),
.Y(n_6841)
);

CKINVDCx5p33_ASAP7_75t_R g6842 ( 
.A(n_6068),
.Y(n_6842)
);

INVx2_ASAP7_75t_L g6843 ( 
.A(n_6139),
.Y(n_6843)
);

INVx1_ASAP7_75t_L g6844 ( 
.A(n_6401),
.Y(n_6844)
);

INVx3_ASAP7_75t_L g6845 ( 
.A(n_6140),
.Y(n_6845)
);

INVx2_ASAP7_75t_L g6846 ( 
.A(n_6142),
.Y(n_6846)
);

INVx1_ASAP7_75t_L g6847 ( 
.A(n_6403),
.Y(n_6847)
);

BUFx12f_ASAP7_75t_L g6848 ( 
.A(n_6362),
.Y(n_6848)
);

BUFx6f_ASAP7_75t_L g6849 ( 
.A(n_6145),
.Y(n_6849)
);

INVx2_ASAP7_75t_L g6850 ( 
.A(n_6146),
.Y(n_6850)
);

INVx1_ASAP7_75t_L g6851 ( 
.A(n_6147),
.Y(n_6851)
);

INVx2_ASAP7_75t_L g6852 ( 
.A(n_6148),
.Y(n_6852)
);

INVx5_ASAP7_75t_L g6853 ( 
.A(n_6152),
.Y(n_6853)
);

NAND2xp5_ASAP7_75t_L g6854 ( 
.A(n_6150),
.B(n_5368),
.Y(n_6854)
);

AND2x4_ASAP7_75t_L g6855 ( 
.A(n_6151),
.B(n_5467),
.Y(n_6855)
);

INVx1_ASAP7_75t_L g6856 ( 
.A(n_6153),
.Y(n_6856)
);

AOI22xp5_ASAP7_75t_L g6857 ( 
.A1(n_6071),
.A2(n_5005),
.B1(n_5013),
.B2(n_5001),
.Y(n_6857)
);

INVx2_ASAP7_75t_L g6858 ( 
.A(n_6154),
.Y(n_6858)
);

INVx1_ASAP7_75t_L g6859 ( 
.A(n_6155),
.Y(n_6859)
);

BUFx6f_ASAP7_75t_L g6860 ( 
.A(n_6156),
.Y(n_6860)
);

BUFx6f_ASAP7_75t_L g6861 ( 
.A(n_6158),
.Y(n_6861)
);

OA21x2_ASAP7_75t_L g6862 ( 
.A1(n_6160),
.A2(n_4138),
.B(n_4136),
.Y(n_6862)
);

INVx3_ASAP7_75t_L g6863 ( 
.A(n_6162),
.Y(n_6863)
);

INVx2_ASAP7_75t_L g6864 ( 
.A(n_6163),
.Y(n_6864)
);

INVx1_ASAP7_75t_L g6865 ( 
.A(n_6166),
.Y(n_6865)
);

BUFx3_ASAP7_75t_L g6866 ( 
.A(n_6399),
.Y(n_6866)
);

INVx3_ASAP7_75t_L g6867 ( 
.A(n_6171),
.Y(n_6867)
);

AOI22xp5_ASAP7_75t_L g6868 ( 
.A1(n_6077),
.A2(n_5108),
.B1(n_5176),
.B2(n_5074),
.Y(n_6868)
);

BUFx6f_ASAP7_75t_L g6869 ( 
.A(n_6172),
.Y(n_6869)
);

NAND2xp5_ASAP7_75t_L g6870 ( 
.A(n_6009),
.B(n_5392),
.Y(n_6870)
);

BUFx3_ASAP7_75t_L g6871 ( 
.A(n_6402),
.Y(n_6871)
);

BUFx6f_ASAP7_75t_L g6872 ( 
.A(n_6343),
.Y(n_6872)
);

INVx3_ASAP7_75t_L g6873 ( 
.A(n_6344),
.Y(n_6873)
);

INVx1_ASAP7_75t_L g6874 ( 
.A(n_6346),
.Y(n_6874)
);

INVx3_ASAP7_75t_L g6875 ( 
.A(n_6011),
.Y(n_6875)
);

AND2x4_ASAP7_75t_L g6876 ( 
.A(n_5990),
.B(n_5473),
.Y(n_6876)
);

BUFx12f_ASAP7_75t_L g6877 ( 
.A(n_6367),
.Y(n_6877)
);

INVx1_ASAP7_75t_L g6878 ( 
.A(n_6012),
.Y(n_6878)
);

OA21x2_ASAP7_75t_L g6879 ( 
.A1(n_6015),
.A2(n_4146),
.B(n_4140),
.Y(n_6879)
);

INVx2_ASAP7_75t_L g6880 ( 
.A(n_6016),
.Y(n_6880)
);

INVx4_ASAP7_75t_L g6881 ( 
.A(n_6082),
.Y(n_6881)
);

AOI22xp5_ASAP7_75t_L g6882 ( 
.A1(n_6087),
.A2(n_5224),
.B1(n_5231),
.B2(n_5184),
.Y(n_6882)
);

BUFx6f_ASAP7_75t_L g6883 ( 
.A(n_6017),
.Y(n_6883)
);

INVx3_ASAP7_75t_L g6884 ( 
.A(n_6019),
.Y(n_6884)
);

INVx1_ASAP7_75t_L g6885 ( 
.A(n_6021),
.Y(n_6885)
);

AND2x4_ASAP7_75t_L g6886 ( 
.A(n_6001),
.B(n_4291),
.Y(n_6886)
);

INVx2_ASAP7_75t_L g6887 ( 
.A(n_6023),
.Y(n_6887)
);

INVx2_ASAP7_75t_L g6888 ( 
.A(n_6024),
.Y(n_6888)
);

NAND2xp5_ASAP7_75t_L g6889 ( 
.A(n_6025),
.B(n_5392),
.Y(n_6889)
);

INVx1_ASAP7_75t_L g6890 ( 
.A(n_6026),
.Y(n_6890)
);

INVx1_ASAP7_75t_L g6891 ( 
.A(n_6028),
.Y(n_6891)
);

INVx2_ASAP7_75t_L g6892 ( 
.A(n_6092),
.Y(n_6892)
);

BUFx6f_ASAP7_75t_L g6893 ( 
.A(n_6369),
.Y(n_6893)
);

INVx3_ASAP7_75t_L g6894 ( 
.A(n_6100),
.Y(n_6894)
);

INVx1_ASAP7_75t_L g6895 ( 
.A(n_6048),
.Y(n_6895)
);

BUFx6f_ASAP7_75t_L g6896 ( 
.A(n_6372),
.Y(n_6896)
);

INVx3_ASAP7_75t_L g6897 ( 
.A(n_6101),
.Y(n_6897)
);

AND2x4_ASAP7_75t_L g6898 ( 
.A(n_6076),
.B(n_4312),
.Y(n_6898)
);

INVx2_ASAP7_75t_L g6899 ( 
.A(n_6103),
.Y(n_6899)
);

INVx2_ASAP7_75t_L g6900 ( 
.A(n_6105),
.Y(n_6900)
);

BUFx6f_ASAP7_75t_L g6901 ( 
.A(n_6373),
.Y(n_6901)
);

BUFx6f_ASAP7_75t_L g6902 ( 
.A(n_6380),
.Y(n_6902)
);

INVx1_ASAP7_75t_L g6903 ( 
.A(n_6095),
.Y(n_6903)
);

INVx5_ASAP7_75t_L g6904 ( 
.A(n_6032),
.Y(n_6904)
);

BUFx8_ASAP7_75t_L g6905 ( 
.A(n_6249),
.Y(n_6905)
);

INVx6_ASAP7_75t_L g6906 ( 
.A(n_6066),
.Y(n_6906)
);

BUFx6f_ASAP7_75t_L g6907 ( 
.A(n_6382),
.Y(n_6907)
);

OA21x2_ASAP7_75t_L g6908 ( 
.A1(n_6485),
.A2(n_4159),
.B(n_4152),
.Y(n_6908)
);

BUFx8_ASAP7_75t_L g6909 ( 
.A(n_6086),
.Y(n_6909)
);

BUFx6f_ASAP7_75t_L g6910 ( 
.A(n_6390),
.Y(n_6910)
);

CKINVDCx6p67_ASAP7_75t_R g6911 ( 
.A(n_6284),
.Y(n_6911)
);

INVx1_ASAP7_75t_L g6912 ( 
.A(n_6096),
.Y(n_6912)
);

INVx1_ASAP7_75t_L g6913 ( 
.A(n_6194),
.Y(n_6913)
);

OAI22xp5_ASAP7_75t_SL g6914 ( 
.A1(n_6405),
.A2(n_4969),
.B1(n_4975),
.B2(n_4957),
.Y(n_6914)
);

CKINVDCx20_ASAP7_75t_R g6915 ( 
.A(n_6114),
.Y(n_6915)
);

INVx1_ASAP7_75t_L g6916 ( 
.A(n_6236),
.Y(n_6916)
);

AND2x2_ASAP7_75t_L g6917 ( 
.A(n_6428),
.B(n_6430),
.Y(n_6917)
);

OA21x2_ASAP7_75t_L g6918 ( 
.A1(n_6110),
.A2(n_4166),
.B(n_4164),
.Y(n_6918)
);

AND2x2_ASAP7_75t_L g6919 ( 
.A(n_6431),
.B(n_5023),
.Y(n_6919)
);

NOR2xp33_ASAP7_75t_L g6920 ( 
.A(n_6125),
.B(n_4424),
.Y(n_6920)
);

INVx2_ASAP7_75t_L g6921 ( 
.A(n_6135),
.Y(n_6921)
);

INVx1_ASAP7_75t_L g6922 ( 
.A(n_6244),
.Y(n_6922)
);

BUFx8_ASAP7_75t_L g6923 ( 
.A(n_6134),
.Y(n_6923)
);

BUFx8_ASAP7_75t_SL g6924 ( 
.A(n_6136),
.Y(n_6924)
);

HB1xp67_ASAP7_75t_L g6925 ( 
.A(n_6252),
.Y(n_6925)
);

BUFx6f_ASAP7_75t_L g6926 ( 
.A(n_6144),
.Y(n_6926)
);

AND2x2_ASAP7_75t_L g6927 ( 
.A(n_6157),
.B(n_5070),
.Y(n_6927)
);

BUFx3_ASAP7_75t_L g6928 ( 
.A(n_6407),
.Y(n_6928)
);

CKINVDCx16_ASAP7_75t_R g6929 ( 
.A(n_6138),
.Y(n_6929)
);

INVx3_ASAP7_75t_L g6930 ( 
.A(n_6159),
.Y(n_6930)
);

INVx2_ASAP7_75t_L g6931 ( 
.A(n_6169),
.Y(n_6931)
);

INVx2_ASAP7_75t_L g6932 ( 
.A(n_6180),
.Y(n_6932)
);

BUFx3_ASAP7_75t_L g6933 ( 
.A(n_6411),
.Y(n_6933)
);

INVx1_ASAP7_75t_L g6934 ( 
.A(n_6459),
.Y(n_6934)
);

AND2x4_ASAP7_75t_L g6935 ( 
.A(n_6469),
.B(n_4494),
.Y(n_6935)
);

OA21x2_ASAP7_75t_L g6936 ( 
.A1(n_6181),
.A2(n_4182),
.B(n_4172),
.Y(n_6936)
);

INVx2_ASAP7_75t_L g6937 ( 
.A(n_6192),
.Y(n_6937)
);

BUFx6f_ASAP7_75t_L g6938 ( 
.A(n_6201),
.Y(n_6938)
);

INVx3_ASAP7_75t_L g6939 ( 
.A(n_6204),
.Y(n_6939)
);

AND2x2_ASAP7_75t_L g6940 ( 
.A(n_6216),
.B(n_5070),
.Y(n_6940)
);

INVx2_ASAP7_75t_L g6941 ( 
.A(n_6227),
.Y(n_6941)
);

BUFx6f_ASAP7_75t_L g6942 ( 
.A(n_6235),
.Y(n_6942)
);

BUFx2_ASAP7_75t_L g6943 ( 
.A(n_6432),
.Y(n_6943)
);

NOR2xp33_ASAP7_75t_SL g6944 ( 
.A(n_6239),
.B(n_4981),
.Y(n_6944)
);

INVx1_ASAP7_75t_L g6945 ( 
.A(n_6471),
.Y(n_6945)
);

OAI22xp5_ASAP7_75t_L g6946 ( 
.A1(n_6240),
.A2(n_6262),
.B1(n_6274),
.B2(n_6257),
.Y(n_6946)
);

INVx2_ASAP7_75t_L g6947 ( 
.A(n_6277),
.Y(n_6947)
);

INVx1_ASAP7_75t_L g6948 ( 
.A(n_6472),
.Y(n_6948)
);

NAND2xp5_ASAP7_75t_L g6949 ( 
.A(n_6278),
.B(n_5392),
.Y(n_6949)
);

BUFx6f_ASAP7_75t_L g6950 ( 
.A(n_6279),
.Y(n_6950)
);

NAND2xp5_ASAP7_75t_L g6951 ( 
.A(n_6280),
.B(n_5474),
.Y(n_6951)
);

HB1xp67_ASAP7_75t_L g6952 ( 
.A(n_6289),
.Y(n_6952)
);

INVx1_ASAP7_75t_L g6953 ( 
.A(n_6290),
.Y(n_6953)
);

CKINVDCx16_ASAP7_75t_R g6954 ( 
.A(n_6149),
.Y(n_6954)
);

BUFx8_ASAP7_75t_L g6955 ( 
.A(n_6161),
.Y(n_6955)
);

INVx5_ASAP7_75t_L g6956 ( 
.A(n_6102),
.Y(n_6956)
);

INVx1_ASAP7_75t_L g6957 ( 
.A(n_6291),
.Y(n_6957)
);

OA21x2_ASAP7_75t_L g6958 ( 
.A1(n_6481),
.A2(n_4186),
.B(n_4185),
.Y(n_6958)
);

INVx1_ASAP7_75t_L g6959 ( 
.A(n_6292),
.Y(n_6959)
);

BUFx3_ASAP7_75t_L g6960 ( 
.A(n_6434),
.Y(n_6960)
);

BUFx6f_ASAP7_75t_L g6961 ( 
.A(n_6294),
.Y(n_6961)
);

BUFx6f_ASAP7_75t_L g6962 ( 
.A(n_6297),
.Y(n_6962)
);

BUFx6f_ASAP7_75t_L g6963 ( 
.A(n_6307),
.Y(n_6963)
);

INVx2_ASAP7_75t_L g6964 ( 
.A(n_6317),
.Y(n_6964)
);

INVx1_ASAP7_75t_L g6965 ( 
.A(n_6318),
.Y(n_6965)
);

INVx3_ASAP7_75t_L g6966 ( 
.A(n_6320),
.Y(n_6966)
);

BUFx6f_ASAP7_75t_L g6967 ( 
.A(n_6330),
.Y(n_6967)
);

BUFx6f_ASAP7_75t_L g6968 ( 
.A(n_6335),
.Y(n_6968)
);

INVxp33_ASAP7_75t_SL g6969 ( 
.A(n_6337),
.Y(n_6969)
);

AND2x2_ASAP7_75t_L g6970 ( 
.A(n_6461),
.B(n_5116),
.Y(n_6970)
);

BUFx6f_ASAP7_75t_L g6971 ( 
.A(n_6467),
.Y(n_6971)
);

INVx1_ASAP7_75t_L g6972 ( 
.A(n_6474),
.Y(n_6972)
);

AND2x2_ASAP7_75t_L g6973 ( 
.A(n_6339),
.B(n_5116),
.Y(n_6973)
);

INVx2_ASAP7_75t_L g6974 ( 
.A(n_6167),
.Y(n_6974)
);

NAND2xp5_ASAP7_75t_L g6975 ( 
.A(n_6285),
.B(n_5474),
.Y(n_6975)
);

INVx1_ASAP7_75t_L g6976 ( 
.A(n_6331),
.Y(n_6976)
);

INVx1_ASAP7_75t_L g6977 ( 
.A(n_6353),
.Y(n_6977)
);

BUFx6f_ASAP7_75t_L g6978 ( 
.A(n_6168),
.Y(n_6978)
);

BUFx6f_ASAP7_75t_L g6979 ( 
.A(n_6177),
.Y(n_6979)
);

INVx2_ASAP7_75t_L g6980 ( 
.A(n_6447),
.Y(n_6980)
);

AOI22x1_ASAP7_75t_SL g6981 ( 
.A1(n_6451),
.A2(n_5022),
.B1(n_5033),
.B2(n_5017),
.Y(n_6981)
);

INVx1_ASAP7_75t_L g6982 ( 
.A(n_6143),
.Y(n_6982)
);

INVx5_ASAP7_75t_L g6983 ( 
.A(n_6170),
.Y(n_6983)
);

INVx2_ASAP7_75t_L g6984 ( 
.A(n_6452),
.Y(n_6984)
);

BUFx3_ASAP7_75t_L g6985 ( 
.A(n_6460),
.Y(n_6985)
);

INVx2_ASAP7_75t_L g6986 ( 
.A(n_6468),
.Y(n_6986)
);

AND2x6_ASAP7_75t_L g6987 ( 
.A(n_6203),
.B(n_5254),
.Y(n_6987)
);

BUFx6f_ASAP7_75t_L g6988 ( 
.A(n_6470),
.Y(n_6988)
);

INVx1_ASAP7_75t_L g6989 ( 
.A(n_6221),
.Y(n_6989)
);

NOR2x1_ASAP7_75t_L g6990 ( 
.A(n_6478),
.B(n_4165),
.Y(n_6990)
);

OAI21x1_ASAP7_75t_L g6991 ( 
.A1(n_6446),
.A2(n_4541),
.B(n_4534),
.Y(n_6991)
);

NAND2xp5_ASAP7_75t_L g6992 ( 
.A(n_6475),
.B(n_5474),
.Y(n_6992)
);

AOI22xp5_ASAP7_75t_L g6993 ( 
.A1(n_6196),
.A2(n_5369),
.B1(n_5374),
.B2(n_5296),
.Y(n_6993)
);

OA21x2_ASAP7_75t_L g6994 ( 
.A1(n_6394),
.A2(n_4200),
.B(n_4195),
.Y(n_6994)
);

INVx6_ASAP7_75t_L g6995 ( 
.A(n_6238),
.Y(n_6995)
);

INVx1_ASAP7_75t_L g6996 ( 
.A(n_6263),
.Y(n_6996)
);

INVx2_ASAP7_75t_L g6997 ( 
.A(n_6002),
.Y(n_6997)
);

BUFx6f_ASAP7_75t_L g6998 ( 
.A(n_6141),
.Y(n_6998)
);

INVx1_ASAP7_75t_L g6999 ( 
.A(n_6263),
.Y(n_6999)
);

INVx2_ASAP7_75t_L g7000 ( 
.A(n_6002),
.Y(n_7000)
);

INVx2_ASAP7_75t_L g7001 ( 
.A(n_6002),
.Y(n_7001)
);

BUFx6f_ASAP7_75t_L g7002 ( 
.A(n_6141),
.Y(n_7002)
);

BUFx6f_ASAP7_75t_L g7003 ( 
.A(n_6141),
.Y(n_7003)
);

INVx6_ASAP7_75t_L g7004 ( 
.A(n_6238),
.Y(n_7004)
);

BUFx2_ASAP7_75t_L g7005 ( 
.A(n_6437),
.Y(n_7005)
);

BUFx12f_ASAP7_75t_L g7006 ( 
.A(n_6439),
.Y(n_7006)
);

BUFx6f_ASAP7_75t_L g7007 ( 
.A(n_6141),
.Y(n_7007)
);

INVx1_ASAP7_75t_L g7008 ( 
.A(n_6263),
.Y(n_7008)
);

AND2x4_ASAP7_75t_L g7009 ( 
.A(n_6141),
.B(n_4700),
.Y(n_7009)
);

INVx2_ASAP7_75t_L g7010 ( 
.A(n_6002),
.Y(n_7010)
);

INVx3_ASAP7_75t_L g7011 ( 
.A(n_6141),
.Y(n_7011)
);

INVx1_ASAP7_75t_L g7012 ( 
.A(n_6263),
.Y(n_7012)
);

HB1xp67_ASAP7_75t_L g7013 ( 
.A(n_6365),
.Y(n_7013)
);

BUFx6f_ASAP7_75t_L g7014 ( 
.A(n_6141),
.Y(n_7014)
);

BUFx6f_ASAP7_75t_L g7015 ( 
.A(n_6141),
.Y(n_7015)
);

BUFx6f_ASAP7_75t_L g7016 ( 
.A(n_6141),
.Y(n_7016)
);

BUFx6f_ASAP7_75t_L g7017 ( 
.A(n_6141),
.Y(n_7017)
);

AOI22xp5_ASAP7_75t_L g7018 ( 
.A1(n_6196),
.A2(n_5510),
.B1(n_5502),
.B2(n_4293),
.Y(n_7018)
);

AOI22xp5_ASAP7_75t_L g7019 ( 
.A1(n_6196),
.A2(n_4294),
.B1(n_4295),
.B2(n_4290),
.Y(n_7019)
);

BUFx6f_ASAP7_75t_L g7020 ( 
.A(n_6141),
.Y(n_7020)
);

BUFx6f_ASAP7_75t_L g7021 ( 
.A(n_6141),
.Y(n_7021)
);

INVx3_ASAP7_75t_L g7022 ( 
.A(n_6141),
.Y(n_7022)
);

INVx1_ASAP7_75t_L g7023 ( 
.A(n_6263),
.Y(n_7023)
);

AND2x6_ASAP7_75t_L g7024 ( 
.A(n_6416),
.B(n_4201),
.Y(n_7024)
);

INVx2_ASAP7_75t_L g7025 ( 
.A(n_6002),
.Y(n_7025)
);

INVx6_ASAP7_75t_L g7026 ( 
.A(n_6238),
.Y(n_7026)
);

AND2x2_ASAP7_75t_L g7027 ( 
.A(n_6406),
.B(n_5123),
.Y(n_7027)
);

CKINVDCx14_ASAP7_75t_R g7028 ( 
.A(n_6126),
.Y(n_7028)
);

AND2x4_ASAP7_75t_L g7029 ( 
.A(n_6141),
.B(n_4744),
.Y(n_7029)
);

BUFx2_ASAP7_75t_L g7030 ( 
.A(n_6437),
.Y(n_7030)
);

BUFx6f_ASAP7_75t_L g7031 ( 
.A(n_6141),
.Y(n_7031)
);

INVx3_ASAP7_75t_L g7032 ( 
.A(n_6141),
.Y(n_7032)
);

INVx2_ASAP7_75t_L g7033 ( 
.A(n_6002),
.Y(n_7033)
);

NAND2xp5_ASAP7_75t_L g7034 ( 
.A(n_6196),
.B(n_4757),
.Y(n_7034)
);

OAI21x1_ASAP7_75t_L g7035 ( 
.A1(n_6394),
.A2(n_4548),
.B(n_4544),
.Y(n_7035)
);

INVx2_ASAP7_75t_L g7036 ( 
.A(n_6002),
.Y(n_7036)
);

BUFx3_ASAP7_75t_L g7037 ( 
.A(n_6141),
.Y(n_7037)
);

OAI21x1_ASAP7_75t_L g7038 ( 
.A1(n_6394),
.A2(n_4580),
.B(n_4550),
.Y(n_7038)
);

AND2x4_ASAP7_75t_L g7039 ( 
.A(n_6141),
.B(n_4788),
.Y(n_7039)
);

NAND2xp5_ASAP7_75t_SL g7040 ( 
.A(n_6439),
.B(n_4298),
.Y(n_7040)
);

INVx2_ASAP7_75t_L g7041 ( 
.A(n_6002),
.Y(n_7041)
);

AND2x2_ASAP7_75t_L g7042 ( 
.A(n_6406),
.B(n_5123),
.Y(n_7042)
);

OA21x2_ASAP7_75t_L g7043 ( 
.A1(n_6394),
.A2(n_4205),
.B(n_4202),
.Y(n_7043)
);

INVx1_ASAP7_75t_L g7044 ( 
.A(n_6263),
.Y(n_7044)
);

INVxp67_ASAP7_75t_L g7045 ( 
.A(n_6406),
.Y(n_7045)
);

CKINVDCx5p33_ASAP7_75t_R g7046 ( 
.A(n_5974),
.Y(n_7046)
);

INVxp33_ASAP7_75t_SL g7047 ( 
.A(n_6406),
.Y(n_7047)
);

INVx2_ASAP7_75t_L g7048 ( 
.A(n_6002),
.Y(n_7048)
);

CKINVDCx14_ASAP7_75t_R g7049 ( 
.A(n_6126),
.Y(n_7049)
);

INVx2_ASAP7_75t_L g7050 ( 
.A(n_6002),
.Y(n_7050)
);

NAND2xp5_ASAP7_75t_L g7051 ( 
.A(n_6196),
.B(n_4795),
.Y(n_7051)
);

OA21x2_ASAP7_75t_L g7052 ( 
.A1(n_6394),
.A2(n_4214),
.B(n_4210),
.Y(n_7052)
);

INVx2_ASAP7_75t_L g7053 ( 
.A(n_6002),
.Y(n_7053)
);

INVx6_ASAP7_75t_L g7054 ( 
.A(n_6238),
.Y(n_7054)
);

AOI22xp5_ASAP7_75t_L g7055 ( 
.A1(n_6196),
.A2(n_4303),
.B1(n_4305),
.B2(n_4302),
.Y(n_7055)
);

INVx1_ASAP7_75t_L g7056 ( 
.A(n_6263),
.Y(n_7056)
);

INVx2_ASAP7_75t_L g7057 ( 
.A(n_6002),
.Y(n_7057)
);

BUFx6f_ASAP7_75t_L g7058 ( 
.A(n_6141),
.Y(n_7058)
);

INVx2_ASAP7_75t_L g7059 ( 
.A(n_6002),
.Y(n_7059)
);

AND2x2_ASAP7_75t_L g7060 ( 
.A(n_6406),
.B(n_5164),
.Y(n_7060)
);

AND2x4_ASAP7_75t_L g7061 ( 
.A(n_6141),
.B(n_4839),
.Y(n_7061)
);

INVx1_ASAP7_75t_L g7062 ( 
.A(n_6263),
.Y(n_7062)
);

BUFx6f_ASAP7_75t_L g7063 ( 
.A(n_6141),
.Y(n_7063)
);

BUFx2_ASAP7_75t_L g7064 ( 
.A(n_6437),
.Y(n_7064)
);

INVx1_ASAP7_75t_L g7065 ( 
.A(n_6263),
.Y(n_7065)
);

INVx2_ASAP7_75t_L g7066 ( 
.A(n_6494),
.Y(n_7066)
);

CKINVDCx5p33_ASAP7_75t_R g7067 ( 
.A(n_6646),
.Y(n_7067)
);

CKINVDCx5p33_ASAP7_75t_R g7068 ( 
.A(n_6741),
.Y(n_7068)
);

INVx2_ASAP7_75t_L g7069 ( 
.A(n_6497),
.Y(n_7069)
);

INVx1_ASAP7_75t_L g7070 ( 
.A(n_6487),
.Y(n_7070)
);

CKINVDCx5p33_ASAP7_75t_R g7071 ( 
.A(n_6924),
.Y(n_7071)
);

INVx2_ASAP7_75t_L g7072 ( 
.A(n_6512),
.Y(n_7072)
);

INVx1_ASAP7_75t_L g7073 ( 
.A(n_7056),
.Y(n_7073)
);

INVx1_ASAP7_75t_L g7074 ( 
.A(n_7062),
.Y(n_7074)
);

OAI21x1_ASAP7_75t_L g7075 ( 
.A1(n_6688),
.A2(n_4654),
.B(n_4603),
.Y(n_7075)
);

CKINVDCx5p33_ASAP7_75t_R g7076 ( 
.A(n_6515),
.Y(n_7076)
);

INVx1_ASAP7_75t_L g7077 ( 
.A(n_7065),
.Y(n_7077)
);

INVx1_ASAP7_75t_L g7078 ( 
.A(n_6509),
.Y(n_7078)
);

INVx1_ASAP7_75t_L g7079 ( 
.A(n_6511),
.Y(n_7079)
);

HB1xp67_ASAP7_75t_L g7080 ( 
.A(n_6559),
.Y(n_7080)
);

BUFx6f_ASAP7_75t_L g7081 ( 
.A(n_6486),
.Y(n_7081)
);

BUFx10_ASAP7_75t_L g7082 ( 
.A(n_6995),
.Y(n_7082)
);

BUFx12f_ASAP7_75t_L g7083 ( 
.A(n_6802),
.Y(n_7083)
);

INVx3_ASAP7_75t_L g7084 ( 
.A(n_6498),
.Y(n_7084)
);

CKINVDCx5p33_ASAP7_75t_R g7085 ( 
.A(n_6534),
.Y(n_7085)
);

INVx6_ASAP7_75t_L g7086 ( 
.A(n_6909),
.Y(n_7086)
);

INVx3_ASAP7_75t_L g7087 ( 
.A(n_6504),
.Y(n_7087)
);

INVx1_ASAP7_75t_L g7088 ( 
.A(n_6528),
.Y(n_7088)
);

INVx1_ASAP7_75t_L g7089 ( 
.A(n_6530),
.Y(n_7089)
);

INVx1_ASAP7_75t_L g7090 ( 
.A(n_6532),
.Y(n_7090)
);

AND2x4_ASAP7_75t_L g7091 ( 
.A(n_7037),
.B(n_4217),
.Y(n_7091)
);

NAND2xp5_ASAP7_75t_L g7092 ( 
.A(n_6807),
.B(n_4853),
.Y(n_7092)
);

INVx1_ASAP7_75t_L g7093 ( 
.A(n_6533),
.Y(n_7093)
);

OA21x2_ASAP7_75t_L g7094 ( 
.A1(n_6553),
.A2(n_4234),
.B(n_4226),
.Y(n_7094)
);

HB1xp67_ASAP7_75t_L g7095 ( 
.A(n_6662),
.Y(n_7095)
);

NAND2xp5_ASAP7_75t_L g7096 ( 
.A(n_6809),
.B(n_6844),
.Y(n_7096)
);

NAND2xp5_ASAP7_75t_L g7097 ( 
.A(n_6847),
.B(n_4925),
.Y(n_7097)
);

CKINVDCx5p33_ASAP7_75t_R g7098 ( 
.A(n_6568),
.Y(n_7098)
);

INVx1_ASAP7_75t_L g7099 ( 
.A(n_6548),
.Y(n_7099)
);

CKINVDCx16_ASAP7_75t_R g7100 ( 
.A(n_6690),
.Y(n_7100)
);

BUFx6f_ASAP7_75t_L g7101 ( 
.A(n_6489),
.Y(n_7101)
);

INVx2_ASAP7_75t_L g7102 ( 
.A(n_6516),
.Y(n_7102)
);

BUFx3_ASAP7_75t_L g7103 ( 
.A(n_6493),
.Y(n_7103)
);

INVx3_ASAP7_75t_L g7104 ( 
.A(n_6508),
.Y(n_7104)
);

INVx6_ASAP7_75t_L g7105 ( 
.A(n_6923),
.Y(n_7105)
);

INVx1_ASAP7_75t_L g7106 ( 
.A(n_6554),
.Y(n_7106)
);

INVx2_ASAP7_75t_L g7107 ( 
.A(n_6529),
.Y(n_7107)
);

CKINVDCx20_ASAP7_75t_R g7108 ( 
.A(n_6669),
.Y(n_7108)
);

OA21x2_ASAP7_75t_L g7109 ( 
.A1(n_6626),
.A2(n_4252),
.B(n_4245),
.Y(n_7109)
);

NAND2xp5_ASAP7_75t_L g7110 ( 
.A(n_6503),
.B(n_4929),
.Y(n_7110)
);

INVx1_ASAP7_75t_L g7111 ( 
.A(n_6556),
.Y(n_7111)
);

CKINVDCx5p33_ASAP7_75t_R g7112 ( 
.A(n_6583),
.Y(n_7112)
);

INVx1_ASAP7_75t_L g7113 ( 
.A(n_6560),
.Y(n_7113)
);

NAND2xp5_ASAP7_75t_L g7114 ( 
.A(n_6588),
.B(n_5024),
.Y(n_7114)
);

INVx3_ASAP7_75t_L g7115 ( 
.A(n_6998),
.Y(n_7115)
);

NAND2xp5_ASAP7_75t_L g7116 ( 
.A(n_6652),
.B(n_5083),
.Y(n_7116)
);

INVx1_ASAP7_75t_L g7117 ( 
.A(n_6562),
.Y(n_7117)
);

CKINVDCx5p33_ASAP7_75t_R g7118 ( 
.A(n_6604),
.Y(n_7118)
);

CKINVDCx5p33_ASAP7_75t_R g7119 ( 
.A(n_6608),
.Y(n_7119)
);

CKINVDCx5p33_ASAP7_75t_R g7120 ( 
.A(n_6609),
.Y(n_7120)
);

BUFx8_ASAP7_75t_L g7121 ( 
.A(n_7005),
.Y(n_7121)
);

INVx2_ASAP7_75t_L g7122 ( 
.A(n_6542),
.Y(n_7122)
);

INVx2_ASAP7_75t_L g7123 ( 
.A(n_6488),
.Y(n_7123)
);

NOR2xp33_ASAP7_75t_R g7124 ( 
.A(n_7028),
.B(n_5050),
.Y(n_7124)
);

INVx1_ASAP7_75t_L g7125 ( 
.A(n_6584),
.Y(n_7125)
);

HB1xp67_ASAP7_75t_L g7126 ( 
.A(n_7013),
.Y(n_7126)
);

INVx3_ASAP7_75t_L g7127 ( 
.A(n_7002),
.Y(n_7127)
);

AND2x2_ASAP7_75t_L g7128 ( 
.A(n_7027),
.B(n_5164),
.Y(n_7128)
);

NAND2xp5_ASAP7_75t_SL g7129 ( 
.A(n_7047),
.B(n_4306),
.Y(n_7129)
);

INVx1_ASAP7_75t_L g7130 ( 
.A(n_6587),
.Y(n_7130)
);

INVx2_ASAP7_75t_L g7131 ( 
.A(n_6491),
.Y(n_7131)
);

CKINVDCx5p33_ASAP7_75t_R g7132 ( 
.A(n_6694),
.Y(n_7132)
);

BUFx2_ASAP7_75t_L g7133 ( 
.A(n_7030),
.Y(n_7133)
);

INVx1_ASAP7_75t_L g7134 ( 
.A(n_6589),
.Y(n_7134)
);

INVx2_ASAP7_75t_L g7135 ( 
.A(n_6997),
.Y(n_7135)
);

INVx2_ASAP7_75t_L g7136 ( 
.A(n_7000),
.Y(n_7136)
);

CKINVDCx20_ASAP7_75t_R g7137 ( 
.A(n_6799),
.Y(n_7137)
);

AND2x4_ASAP7_75t_L g7138 ( 
.A(n_7011),
.B(n_7022),
.Y(n_7138)
);

BUFx3_ASAP7_75t_L g7139 ( 
.A(n_7003),
.Y(n_7139)
);

INVx1_ASAP7_75t_L g7140 ( 
.A(n_6594),
.Y(n_7140)
);

CKINVDCx5p33_ASAP7_75t_R g7141 ( 
.A(n_6714),
.Y(n_7141)
);

CKINVDCx5p33_ASAP7_75t_R g7142 ( 
.A(n_6726),
.Y(n_7142)
);

INVx3_ASAP7_75t_L g7143 ( 
.A(n_7007),
.Y(n_7143)
);

INVx2_ASAP7_75t_L g7144 ( 
.A(n_7001),
.Y(n_7144)
);

CKINVDCx5p33_ASAP7_75t_R g7145 ( 
.A(n_6748),
.Y(n_7145)
);

CKINVDCx5p33_ASAP7_75t_R g7146 ( 
.A(n_6758),
.Y(n_7146)
);

CKINVDCx20_ASAP7_75t_R g7147 ( 
.A(n_6915),
.Y(n_7147)
);

OAI21x1_ASAP7_75t_L g7148 ( 
.A1(n_6634),
.A2(n_4738),
.B(n_4724),
.Y(n_7148)
);

NOR2xp33_ASAP7_75t_R g7149 ( 
.A(n_7049),
.B(n_5089),
.Y(n_7149)
);

CKINVDCx20_ASAP7_75t_R g7150 ( 
.A(n_6955),
.Y(n_7150)
);

INVx2_ASAP7_75t_L g7151 ( 
.A(n_7010),
.Y(n_7151)
);

INVx1_ASAP7_75t_L g7152 ( 
.A(n_6597),
.Y(n_7152)
);

INVx1_ASAP7_75t_L g7153 ( 
.A(n_6613),
.Y(n_7153)
);

INVx2_ASAP7_75t_L g7154 ( 
.A(n_7025),
.Y(n_7154)
);

CKINVDCx5p33_ASAP7_75t_R g7155 ( 
.A(n_6811),
.Y(n_7155)
);

INVx1_ASAP7_75t_L g7156 ( 
.A(n_6614),
.Y(n_7156)
);

CKINVDCx5p33_ASAP7_75t_R g7157 ( 
.A(n_6842),
.Y(n_7157)
);

CKINVDCx5p33_ASAP7_75t_R g7158 ( 
.A(n_7046),
.Y(n_7158)
);

NAND2xp5_ASAP7_75t_L g7159 ( 
.A(n_6661),
.B(n_5237),
.Y(n_7159)
);

INVx1_ASAP7_75t_L g7160 ( 
.A(n_6615),
.Y(n_7160)
);

CKINVDCx5p33_ASAP7_75t_R g7161 ( 
.A(n_6500),
.Y(n_7161)
);

AND2x2_ASAP7_75t_L g7162 ( 
.A(n_7042),
.B(n_5196),
.Y(n_7162)
);

INVx3_ASAP7_75t_L g7163 ( 
.A(n_7014),
.Y(n_7163)
);

BUFx3_ASAP7_75t_L g7164 ( 
.A(n_7015),
.Y(n_7164)
);

INVx1_ASAP7_75t_L g7165 ( 
.A(n_6616),
.Y(n_7165)
);

CKINVDCx5p33_ASAP7_75t_R g7166 ( 
.A(n_6723),
.Y(n_7166)
);

NAND2xp5_ASAP7_75t_SL g7167 ( 
.A(n_7060),
.B(n_4307),
.Y(n_7167)
);

BUFx6f_ASAP7_75t_L g7168 ( 
.A(n_7016),
.Y(n_7168)
);

INVx1_ASAP7_75t_L g7169 ( 
.A(n_6617),
.Y(n_7169)
);

HB1xp67_ASAP7_75t_L g7170 ( 
.A(n_6564),
.Y(n_7170)
);

HB1xp67_ASAP7_75t_L g7171 ( 
.A(n_6578),
.Y(n_7171)
);

INVx1_ASAP7_75t_L g7172 ( 
.A(n_6619),
.Y(n_7172)
);

CKINVDCx5p33_ASAP7_75t_R g7173 ( 
.A(n_6969),
.Y(n_7173)
);

INVx1_ASAP7_75t_L g7174 ( 
.A(n_6630),
.Y(n_7174)
);

INVx1_ASAP7_75t_L g7175 ( 
.A(n_6633),
.Y(n_7175)
);

HB1xp67_ASAP7_75t_L g7176 ( 
.A(n_6992),
.Y(n_7176)
);

INVx2_ASAP7_75t_L g7177 ( 
.A(n_7033),
.Y(n_7177)
);

CKINVDCx5p33_ASAP7_75t_R g7178 ( 
.A(n_6490),
.Y(n_7178)
);

CKINVDCx5p33_ASAP7_75t_R g7179 ( 
.A(n_6600),
.Y(n_7179)
);

INVx1_ASAP7_75t_L g7180 ( 
.A(n_6635),
.Y(n_7180)
);

INVx1_ASAP7_75t_L g7181 ( 
.A(n_6649),
.Y(n_7181)
);

CKINVDCx5p33_ASAP7_75t_R g7182 ( 
.A(n_6621),
.Y(n_7182)
);

INVx2_ASAP7_75t_L g7183 ( 
.A(n_7036),
.Y(n_7183)
);

INVx1_ASAP7_75t_L g7184 ( 
.A(n_6996),
.Y(n_7184)
);

NOR2xp33_ASAP7_75t_L g7185 ( 
.A(n_7045),
.B(n_4309),
.Y(n_7185)
);

INVx2_ASAP7_75t_SL g7186 ( 
.A(n_6492),
.Y(n_7186)
);

INVxp33_ASAP7_75t_L g7187 ( 
.A(n_6549),
.Y(n_7187)
);

INVx1_ASAP7_75t_L g7188 ( 
.A(n_6999),
.Y(n_7188)
);

CKINVDCx5p33_ASAP7_75t_R g7189 ( 
.A(n_6638),
.Y(n_7189)
);

INVx1_ASAP7_75t_L g7190 ( 
.A(n_7008),
.Y(n_7190)
);

INVx1_ASAP7_75t_L g7191 ( 
.A(n_7012),
.Y(n_7191)
);

INVx1_ASAP7_75t_L g7192 ( 
.A(n_7023),
.Y(n_7192)
);

CKINVDCx5p33_ASAP7_75t_R g7193 ( 
.A(n_6656),
.Y(n_7193)
);

NOR2xp33_ASAP7_75t_L g7194 ( 
.A(n_6695),
.B(n_6755),
.Y(n_7194)
);

INVx1_ASAP7_75t_L g7195 ( 
.A(n_7044),
.Y(n_7195)
);

INVx2_ASAP7_75t_L g7196 ( 
.A(n_7041),
.Y(n_7196)
);

CKINVDCx5p33_ASAP7_75t_R g7197 ( 
.A(n_6810),
.Y(n_7197)
);

INVx1_ASAP7_75t_L g7198 ( 
.A(n_6851),
.Y(n_7198)
);

INVx2_ASAP7_75t_L g7199 ( 
.A(n_7048),
.Y(n_7199)
);

CKINVDCx20_ASAP7_75t_R g7200 ( 
.A(n_6929),
.Y(n_7200)
);

CKINVDCx5p33_ASAP7_75t_R g7201 ( 
.A(n_6848),
.Y(n_7201)
);

CKINVDCx5p33_ASAP7_75t_R g7202 ( 
.A(n_6877),
.Y(n_7202)
);

NAND2xp5_ASAP7_75t_L g7203 ( 
.A(n_6663),
.B(n_5396),
.Y(n_7203)
);

INVx2_ASAP7_75t_L g7204 ( 
.A(n_7050),
.Y(n_7204)
);

INVxp67_ASAP7_75t_L g7205 ( 
.A(n_6550),
.Y(n_7205)
);

INVx2_ASAP7_75t_L g7206 ( 
.A(n_7053),
.Y(n_7206)
);

INVx1_ASAP7_75t_L g7207 ( 
.A(n_6856),
.Y(n_7207)
);

BUFx6f_ASAP7_75t_L g7208 ( 
.A(n_7017),
.Y(n_7208)
);

NOR2xp33_ASAP7_75t_R g7209 ( 
.A(n_6813),
.B(n_5103),
.Y(n_7209)
);

BUFx6f_ASAP7_75t_L g7210 ( 
.A(n_7020),
.Y(n_7210)
);

NAND2xp5_ASAP7_75t_L g7211 ( 
.A(n_6671),
.B(n_5410),
.Y(n_7211)
);

CKINVDCx5p33_ASAP7_75t_R g7212 ( 
.A(n_7006),
.Y(n_7212)
);

INVx1_ASAP7_75t_L g7213 ( 
.A(n_6859),
.Y(n_7213)
);

CKINVDCx5p33_ASAP7_75t_R g7214 ( 
.A(n_6954),
.Y(n_7214)
);

HB1xp67_ASAP7_75t_L g7215 ( 
.A(n_7064),
.Y(n_7215)
);

INVx1_ASAP7_75t_L g7216 ( 
.A(n_6865),
.Y(n_7216)
);

NAND2xp5_ASAP7_75t_L g7217 ( 
.A(n_6675),
.B(n_5417),
.Y(n_7217)
);

CKINVDCx20_ASAP7_75t_R g7218 ( 
.A(n_6911),
.Y(n_7218)
);

NAND2xp5_ASAP7_75t_SL g7219 ( 
.A(n_6496),
.B(n_4310),
.Y(n_7219)
);

INVxp67_ASAP7_75t_L g7220 ( 
.A(n_6495),
.Y(n_7220)
);

NOR2xp33_ASAP7_75t_R g7221 ( 
.A(n_6501),
.B(n_6664),
.Y(n_7221)
);

BUFx6f_ASAP7_75t_L g7222 ( 
.A(n_7021),
.Y(n_7222)
);

BUFx6f_ASAP7_75t_L g7223 ( 
.A(n_7031),
.Y(n_7223)
);

INVx1_ASAP7_75t_SL g7224 ( 
.A(n_6775),
.Y(n_7224)
);

INVx2_ASAP7_75t_L g7225 ( 
.A(n_7057),
.Y(n_7225)
);

NOR2xp67_ASAP7_75t_L g7226 ( 
.A(n_6618),
.B(n_4316),
.Y(n_7226)
);

CKINVDCx5p33_ASAP7_75t_R g7227 ( 
.A(n_6893),
.Y(n_7227)
);

BUFx6f_ASAP7_75t_L g7228 ( 
.A(n_7058),
.Y(n_7228)
);

AND2x2_ASAP7_75t_L g7229 ( 
.A(n_6601),
.B(n_5196),
.Y(n_7229)
);

INVx2_ASAP7_75t_L g7230 ( 
.A(n_7059),
.Y(n_7230)
);

INVx1_ASAP7_75t_L g7231 ( 
.A(n_6874),
.Y(n_7231)
);

CKINVDCx5p33_ASAP7_75t_R g7232 ( 
.A(n_6896),
.Y(n_7232)
);

INVx1_ASAP7_75t_L g7233 ( 
.A(n_6641),
.Y(n_7233)
);

CKINVDCx5p33_ASAP7_75t_R g7234 ( 
.A(n_6901),
.Y(n_7234)
);

BUFx2_ASAP7_75t_L g7235 ( 
.A(n_6625),
.Y(n_7235)
);

INVx1_ASAP7_75t_L g7236 ( 
.A(n_6677),
.Y(n_7236)
);

BUFx2_ASAP7_75t_L g7237 ( 
.A(n_6643),
.Y(n_7237)
);

INVx1_ASAP7_75t_L g7238 ( 
.A(n_6680),
.Y(n_7238)
);

NOR2xp33_ASAP7_75t_L g7239 ( 
.A(n_6920),
.B(n_4321),
.Y(n_7239)
);

CKINVDCx5p33_ASAP7_75t_R g7240 ( 
.A(n_6902),
.Y(n_7240)
);

BUFx6f_ASAP7_75t_L g7241 ( 
.A(n_7063),
.Y(n_7241)
);

INVx2_ASAP7_75t_L g7242 ( 
.A(n_6545),
.Y(n_7242)
);

BUFx6f_ASAP7_75t_L g7243 ( 
.A(n_6978),
.Y(n_7243)
);

INVx4_ASAP7_75t_L g7244 ( 
.A(n_7004),
.Y(n_7244)
);

NOR2xp33_ASAP7_75t_R g7245 ( 
.A(n_6563),
.B(n_5144),
.Y(n_7245)
);

INVx1_ASAP7_75t_L g7246 ( 
.A(n_6696),
.Y(n_7246)
);

INVx2_ASAP7_75t_L g7247 ( 
.A(n_6547),
.Y(n_7247)
);

AND2x2_ASAP7_75t_L g7248 ( 
.A(n_6678),
.B(n_5286),
.Y(n_7248)
);

AND2x2_ASAP7_75t_L g7249 ( 
.A(n_6535),
.B(n_5286),
.Y(n_7249)
);

CKINVDCx5p33_ASAP7_75t_R g7250 ( 
.A(n_6907),
.Y(n_7250)
);

CKINVDCx20_ASAP7_75t_R g7251 ( 
.A(n_6582),
.Y(n_7251)
);

INVx2_ASAP7_75t_L g7252 ( 
.A(n_6551),
.Y(n_7252)
);

INVx1_ASAP7_75t_L g7253 ( 
.A(n_6707),
.Y(n_7253)
);

INVx2_ASAP7_75t_L g7254 ( 
.A(n_6575),
.Y(n_7254)
);

BUFx6f_ASAP7_75t_L g7255 ( 
.A(n_6979),
.Y(n_7255)
);

INVx2_ASAP7_75t_L g7256 ( 
.A(n_6586),
.Y(n_7256)
);

CKINVDCx5p33_ASAP7_75t_R g7257 ( 
.A(n_6910),
.Y(n_7257)
);

CKINVDCx20_ASAP7_75t_R g7258 ( 
.A(n_6590),
.Y(n_7258)
);

OAI21x1_ASAP7_75t_L g7259 ( 
.A1(n_6752),
.A2(n_4750),
.B(n_4742),
.Y(n_7259)
);

NAND2xp5_ASAP7_75t_SL g7260 ( 
.A(n_7034),
.B(n_4322),
.Y(n_7260)
);

INVx1_ASAP7_75t_SL g7261 ( 
.A(n_6691),
.Y(n_7261)
);

NOR2xp33_ASAP7_75t_L g7262 ( 
.A(n_6949),
.B(n_4323),
.Y(n_7262)
);

CKINVDCx20_ASAP7_75t_R g7263 ( 
.A(n_6985),
.Y(n_7263)
);

AND2x2_ASAP7_75t_L g7264 ( 
.A(n_6540),
.B(n_5290),
.Y(n_7264)
);

INVx1_ASAP7_75t_L g7265 ( 
.A(n_6720),
.Y(n_7265)
);

INVx1_ASAP7_75t_L g7266 ( 
.A(n_6724),
.Y(n_7266)
);

HB1xp67_ASAP7_75t_L g7267 ( 
.A(n_6876),
.Y(n_7267)
);

INVx1_ASAP7_75t_L g7268 ( 
.A(n_6736),
.Y(n_7268)
);

INVx1_ASAP7_75t_L g7269 ( 
.A(n_6740),
.Y(n_7269)
);

INVx2_ASAP7_75t_L g7270 ( 
.A(n_6592),
.Y(n_7270)
);

INVx2_ASAP7_75t_L g7271 ( 
.A(n_6880),
.Y(n_7271)
);

INVx2_ASAP7_75t_L g7272 ( 
.A(n_6887),
.Y(n_7272)
);

CKINVDCx5p33_ASAP7_75t_R g7273 ( 
.A(n_6926),
.Y(n_7273)
);

BUFx6f_ASAP7_75t_L g7274 ( 
.A(n_6988),
.Y(n_7274)
);

INVx2_ASAP7_75t_L g7275 ( 
.A(n_6888),
.Y(n_7275)
);

CKINVDCx5p33_ASAP7_75t_R g7276 ( 
.A(n_6938),
.Y(n_7276)
);

INVx3_ASAP7_75t_L g7277 ( 
.A(n_6872),
.Y(n_7277)
);

BUFx6f_ASAP7_75t_L g7278 ( 
.A(n_6994),
.Y(n_7278)
);

CKINVDCx20_ASAP7_75t_R g7279 ( 
.A(n_6507),
.Y(n_7279)
);

INVx1_ASAP7_75t_L g7280 ( 
.A(n_6746),
.Y(n_7280)
);

INVx1_ASAP7_75t_L g7281 ( 
.A(n_6751),
.Y(n_7281)
);

INVx1_ASAP7_75t_L g7282 ( 
.A(n_6760),
.Y(n_7282)
);

CKINVDCx20_ASAP7_75t_R g7283 ( 
.A(n_6526),
.Y(n_7283)
);

CKINVDCx5p33_ASAP7_75t_R g7284 ( 
.A(n_6942),
.Y(n_7284)
);

CKINVDCx5p33_ASAP7_75t_R g7285 ( 
.A(n_6950),
.Y(n_7285)
);

CKINVDCx5p33_ASAP7_75t_R g7286 ( 
.A(n_6961),
.Y(n_7286)
);

INVx1_ASAP7_75t_L g7287 ( 
.A(n_6776),
.Y(n_7287)
);

BUFx6f_ASAP7_75t_L g7288 ( 
.A(n_7043),
.Y(n_7288)
);

NOR2xp33_ASAP7_75t_L g7289 ( 
.A(n_6951),
.B(n_4324),
.Y(n_7289)
);

CKINVDCx5p33_ASAP7_75t_R g7290 ( 
.A(n_6962),
.Y(n_7290)
);

INVx2_ASAP7_75t_L g7291 ( 
.A(n_6603),
.Y(n_7291)
);

OA21x2_ASAP7_75t_L g7292 ( 
.A1(n_6767),
.A2(n_4260),
.B(n_4253),
.Y(n_7292)
);

INVx3_ASAP7_75t_L g7293 ( 
.A(n_6517),
.Y(n_7293)
);

INVx2_ASAP7_75t_L g7294 ( 
.A(n_6624),
.Y(n_7294)
);

CKINVDCx20_ASAP7_75t_R g7295 ( 
.A(n_6571),
.Y(n_7295)
);

AND2x2_ASAP7_75t_L g7296 ( 
.A(n_6555),
.B(n_5290),
.Y(n_7296)
);

INVx1_ASAP7_75t_L g7297 ( 
.A(n_6777),
.Y(n_7297)
);

CKINVDCx5p33_ASAP7_75t_R g7298 ( 
.A(n_6963),
.Y(n_7298)
);

INVx1_ASAP7_75t_L g7299 ( 
.A(n_6785),
.Y(n_7299)
);

NOR2xp33_ASAP7_75t_L g7300 ( 
.A(n_6546),
.B(n_4327),
.Y(n_7300)
);

BUFx3_ASAP7_75t_L g7301 ( 
.A(n_6906),
.Y(n_7301)
);

HB1xp67_ASAP7_75t_L g7302 ( 
.A(n_6654),
.Y(n_7302)
);

CKINVDCx20_ASAP7_75t_R g7303 ( 
.A(n_6581),
.Y(n_7303)
);

CKINVDCx5p33_ASAP7_75t_R g7304 ( 
.A(n_6967),
.Y(n_7304)
);

CKINVDCx5p33_ASAP7_75t_R g7305 ( 
.A(n_6968),
.Y(n_7305)
);

INVx3_ASAP7_75t_L g7306 ( 
.A(n_6518),
.Y(n_7306)
);

CKINVDCx5p33_ASAP7_75t_R g7307 ( 
.A(n_6971),
.Y(n_7307)
);

CKINVDCx5p33_ASAP7_75t_R g7308 ( 
.A(n_6780),
.Y(n_7308)
);

CKINVDCx20_ASAP7_75t_R g7309 ( 
.A(n_6660),
.Y(n_7309)
);

CKINVDCx5p33_ASAP7_75t_R g7310 ( 
.A(n_6946),
.Y(n_7310)
);

CKINVDCx5p33_ASAP7_75t_R g7311 ( 
.A(n_6735),
.Y(n_7311)
);

AND2x2_ASAP7_75t_L g7312 ( 
.A(n_6557),
.B(n_5325),
.Y(n_7312)
);

INVx1_ASAP7_75t_L g7313 ( 
.A(n_6786),
.Y(n_7313)
);

AND2x4_ASAP7_75t_L g7314 ( 
.A(n_7032),
.B(n_4267),
.Y(n_7314)
);

CKINVDCx16_ASAP7_75t_R g7315 ( 
.A(n_6841),
.Y(n_7315)
);

INVx1_ASAP7_75t_L g7316 ( 
.A(n_6787),
.Y(n_7316)
);

INVx5_ASAP7_75t_L g7317 ( 
.A(n_6759),
.Y(n_7317)
);

INVx2_ASAP7_75t_L g7318 ( 
.A(n_6639),
.Y(n_7318)
);

NAND2xp5_ASAP7_75t_L g7319 ( 
.A(n_6803),
.B(n_6828),
.Y(n_7319)
);

CKINVDCx5p33_ASAP7_75t_R g7320 ( 
.A(n_6801),
.Y(n_7320)
);

AND2x4_ASAP7_75t_L g7321 ( 
.A(n_6855),
.B(n_4272),
.Y(n_7321)
);

CKINVDCx20_ASAP7_75t_R g7322 ( 
.A(n_6806),
.Y(n_7322)
);

INVx1_ASAP7_75t_L g7323 ( 
.A(n_6878),
.Y(n_7323)
);

BUFx6f_ASAP7_75t_L g7324 ( 
.A(n_7052),
.Y(n_7324)
);

INVx1_ASAP7_75t_L g7325 ( 
.A(n_6885),
.Y(n_7325)
);

OAI22xp5_ASAP7_75t_SL g7326 ( 
.A1(n_6914),
.A2(n_5150),
.B1(n_5171),
.B2(n_5149),
.Y(n_7326)
);

CKINVDCx5p33_ASAP7_75t_R g7327 ( 
.A(n_6815),
.Y(n_7327)
);

NAND2xp5_ASAP7_75t_L g7328 ( 
.A(n_7051),
.B(n_5424),
.Y(n_7328)
);

CKINVDCx5p33_ASAP7_75t_R g7329 ( 
.A(n_6866),
.Y(n_7329)
);

INVx1_ASAP7_75t_L g7330 ( 
.A(n_6890),
.Y(n_7330)
);

HB1xp67_ASAP7_75t_L g7331 ( 
.A(n_6659),
.Y(n_7331)
);

INVx4_ASAP7_75t_L g7332 ( 
.A(n_7026),
.Y(n_7332)
);

INVx1_ASAP7_75t_L g7333 ( 
.A(n_6891),
.Y(n_7333)
);

INVx2_ASAP7_75t_L g7334 ( 
.A(n_6647),
.Y(n_7334)
);

AND2x4_ASAP7_75t_L g7335 ( 
.A(n_6567),
.B(n_4273),
.Y(n_7335)
);

NAND2xp5_ASAP7_75t_L g7336 ( 
.A(n_6739),
.B(n_6778),
.Y(n_7336)
);

NAND2xp5_ASAP7_75t_L g7337 ( 
.A(n_6789),
.B(n_6790),
.Y(n_7337)
);

INVx1_ASAP7_75t_L g7338 ( 
.A(n_6873),
.Y(n_7338)
);

INVx2_ASAP7_75t_L g7339 ( 
.A(n_6650),
.Y(n_7339)
);

INVx1_ASAP7_75t_L g7340 ( 
.A(n_6513),
.Y(n_7340)
);

INVx2_ASAP7_75t_L g7341 ( 
.A(n_6658),
.Y(n_7341)
);

INVx1_ASAP7_75t_L g7342 ( 
.A(n_6665),
.Y(n_7342)
);

INVx1_ASAP7_75t_L g7343 ( 
.A(n_6666),
.Y(n_7343)
);

INVx1_ASAP7_75t_L g7344 ( 
.A(n_6668),
.Y(n_7344)
);

INVx1_ASAP7_75t_L g7345 ( 
.A(n_6674),
.Y(n_7345)
);

INVx2_ASAP7_75t_L g7346 ( 
.A(n_6683),
.Y(n_7346)
);

NAND2xp33_ASAP7_75t_SL g7347 ( 
.A(n_6919),
.B(n_5188),
.Y(n_7347)
);

CKINVDCx5p33_ASAP7_75t_R g7348 ( 
.A(n_6871),
.Y(n_7348)
);

INVx2_ASAP7_75t_L g7349 ( 
.A(n_6684),
.Y(n_7349)
);

INVx1_ASAP7_75t_L g7350 ( 
.A(n_6685),
.Y(n_7350)
);

INVx1_ASAP7_75t_L g7351 ( 
.A(n_6700),
.Y(n_7351)
);

INVx1_ASAP7_75t_L g7352 ( 
.A(n_6701),
.Y(n_7352)
);

CKINVDCx20_ASAP7_75t_R g7353 ( 
.A(n_6928),
.Y(n_7353)
);

INVx2_ASAP7_75t_L g7354 ( 
.A(n_6708),
.Y(n_7354)
);

INVx2_ASAP7_75t_L g7355 ( 
.A(n_6709),
.Y(n_7355)
);

INVx3_ASAP7_75t_L g7356 ( 
.A(n_6519),
.Y(n_7356)
);

INVx1_ASAP7_75t_L g7357 ( 
.A(n_6713),
.Y(n_7357)
);

AND2x4_ASAP7_75t_L g7358 ( 
.A(n_6499),
.B(n_4274),
.Y(n_7358)
);

CKINVDCx5p33_ASAP7_75t_R g7359 ( 
.A(n_6933),
.Y(n_7359)
);

AND2x2_ASAP7_75t_L g7360 ( 
.A(n_6558),
.B(n_6572),
.Y(n_7360)
);

INVx2_ASAP7_75t_L g7361 ( 
.A(n_6727),
.Y(n_7361)
);

HB1xp67_ASAP7_75t_L g7362 ( 
.A(n_6744),
.Y(n_7362)
);

CKINVDCx5p33_ASAP7_75t_R g7363 ( 
.A(n_6960),
.Y(n_7363)
);

AND2x4_ASAP7_75t_L g7364 ( 
.A(n_6505),
.B(n_4275),
.Y(n_7364)
);

NAND2xp5_ASAP7_75t_L g7365 ( 
.A(n_6689),
.B(n_4332),
.Y(n_7365)
);

CKINVDCx16_ASAP7_75t_R g7366 ( 
.A(n_6944),
.Y(n_7366)
);

CKINVDCx5p33_ASAP7_75t_R g7367 ( 
.A(n_6514),
.Y(n_7367)
);

INVx1_ASAP7_75t_L g7368 ( 
.A(n_6729),
.Y(n_7368)
);

INVx1_ASAP7_75t_L g7369 ( 
.A(n_6731),
.Y(n_7369)
);

OA21x2_ASAP7_75t_L g7370 ( 
.A1(n_6781),
.A2(n_4286),
.B(n_4276),
.Y(n_7370)
);

OAI21x1_ASAP7_75t_L g7371 ( 
.A1(n_6794),
.A2(n_4796),
.B(n_4753),
.Y(n_7371)
);

AND2x4_ASAP7_75t_L g7372 ( 
.A(n_6510),
.B(n_4288),
.Y(n_7372)
);

INVx2_ASAP7_75t_L g7373 ( 
.A(n_6733),
.Y(n_7373)
);

CKINVDCx5p33_ASAP7_75t_R g7374 ( 
.A(n_6520),
.Y(n_7374)
);

INVx1_ASAP7_75t_L g7375 ( 
.A(n_6747),
.Y(n_7375)
);

INVx1_ASAP7_75t_L g7376 ( 
.A(n_6750),
.Y(n_7376)
);

INVx1_ASAP7_75t_L g7377 ( 
.A(n_6754),
.Y(n_7377)
);

INVx1_ASAP7_75t_L g7378 ( 
.A(n_6762),
.Y(n_7378)
);

BUFx2_ASAP7_75t_L g7379 ( 
.A(n_6772),
.Y(n_7379)
);

INVx1_ASAP7_75t_L g7380 ( 
.A(n_6765),
.Y(n_7380)
);

CKINVDCx5p33_ASAP7_75t_R g7381 ( 
.A(n_6577),
.Y(n_7381)
);

CKINVDCx5p33_ASAP7_75t_R g7382 ( 
.A(n_6743),
.Y(n_7382)
);

INVx1_ASAP7_75t_L g7383 ( 
.A(n_6774),
.Y(n_7383)
);

CKINVDCx5p33_ASAP7_75t_R g7384 ( 
.A(n_6881),
.Y(n_7384)
);

CKINVDCx20_ASAP7_75t_R g7385 ( 
.A(n_6943),
.Y(n_7385)
);

INVx1_ASAP7_75t_L g7386 ( 
.A(n_6788),
.Y(n_7386)
);

INVx2_ASAP7_75t_L g7387 ( 
.A(n_6792),
.Y(n_7387)
);

NAND2xp5_ASAP7_75t_L g7388 ( 
.A(n_6524),
.B(n_4333),
.Y(n_7388)
);

BUFx6f_ASAP7_75t_L g7389 ( 
.A(n_6538),
.Y(n_7389)
);

CKINVDCx20_ASAP7_75t_R g7390 ( 
.A(n_6830),
.Y(n_7390)
);

CKINVDCx5p33_ASAP7_75t_R g7391 ( 
.A(n_6905),
.Y(n_7391)
);

CKINVDCx20_ASAP7_75t_R g7392 ( 
.A(n_6602),
.Y(n_7392)
);

HB1xp67_ASAP7_75t_L g7393 ( 
.A(n_6839),
.Y(n_7393)
);

BUFx6f_ASAP7_75t_L g7394 ( 
.A(n_6539),
.Y(n_7394)
);

INVx2_ASAP7_75t_L g7395 ( 
.A(n_6797),
.Y(n_7395)
);

CKINVDCx20_ASAP7_75t_R g7396 ( 
.A(n_6644),
.Y(n_7396)
);

INVx2_ASAP7_75t_L g7397 ( 
.A(n_6800),
.Y(n_7397)
);

INVx2_ASAP7_75t_L g7398 ( 
.A(n_6804),
.Y(n_7398)
);

INVx2_ASAP7_75t_L g7399 ( 
.A(n_6812),
.Y(n_7399)
);

AND2x6_ASAP7_75t_L g7400 ( 
.A(n_6580),
.B(n_4289),
.Y(n_7400)
);

INVxp67_ASAP7_75t_L g7401 ( 
.A(n_6753),
.Y(n_7401)
);

OA21x2_ASAP7_75t_L g7402 ( 
.A1(n_6798),
.A2(n_4311),
.B(n_4296),
.Y(n_7402)
);

BUFx2_ASAP7_75t_L g7403 ( 
.A(n_6595),
.Y(n_7403)
);

INVx1_ASAP7_75t_L g7404 ( 
.A(n_6818),
.Y(n_7404)
);

INVx2_ASAP7_75t_L g7405 ( 
.A(n_6820),
.Y(n_7405)
);

INVx1_ASAP7_75t_L g7406 ( 
.A(n_6840),
.Y(n_7406)
);

INVx1_ASAP7_75t_L g7407 ( 
.A(n_6843),
.Y(n_7407)
);

INVx2_ASAP7_75t_L g7408 ( 
.A(n_6846),
.Y(n_7408)
);

INVx2_ASAP7_75t_L g7409 ( 
.A(n_6850),
.Y(n_7409)
);

INVx1_ASAP7_75t_L g7410 ( 
.A(n_6852),
.Y(n_7410)
);

INVx3_ASAP7_75t_L g7411 ( 
.A(n_6552),
.Y(n_7411)
);

BUFx6f_ASAP7_75t_L g7412 ( 
.A(n_6561),
.Y(n_7412)
);

CKINVDCx20_ASAP7_75t_R g7413 ( 
.A(n_6825),
.Y(n_7413)
);

INVx2_ASAP7_75t_L g7414 ( 
.A(n_6858),
.Y(n_7414)
);

NAND2xp5_ASAP7_75t_L g7415 ( 
.A(n_6593),
.B(n_4335),
.Y(n_7415)
);

NAND2xp5_ASAP7_75t_L g7416 ( 
.A(n_6612),
.B(n_6523),
.Y(n_7416)
);

CKINVDCx20_ASAP7_75t_R g7417 ( 
.A(n_6837),
.Y(n_7417)
);

AND2x2_ASAP7_75t_L g7418 ( 
.A(n_6715),
.B(n_5325),
.Y(n_7418)
);

CKINVDCx5p33_ASAP7_75t_R g7419 ( 
.A(n_7054),
.Y(n_7419)
);

INVx1_ASAP7_75t_L g7420 ( 
.A(n_6864),
.Y(n_7420)
);

AND2x2_ASAP7_75t_L g7421 ( 
.A(n_6717),
.B(n_5337),
.Y(n_7421)
);

INVx1_ASAP7_75t_L g7422 ( 
.A(n_6875),
.Y(n_7422)
);

INVx1_ASAP7_75t_L g7423 ( 
.A(n_6884),
.Y(n_7423)
);

AND2x4_ASAP7_75t_L g7424 ( 
.A(n_6521),
.B(n_4314),
.Y(n_7424)
);

HB1xp67_ASAP7_75t_L g7425 ( 
.A(n_6908),
.Y(n_7425)
);

INVx1_ASAP7_75t_L g7426 ( 
.A(n_6816),
.Y(n_7426)
);

NOR2xp67_ASAP7_75t_L g7427 ( 
.A(n_6642),
.B(n_4340),
.Y(n_7427)
);

CKINVDCx5p33_ASAP7_75t_R g7428 ( 
.A(n_6894),
.Y(n_7428)
);

NAND2xp5_ASAP7_75t_SL g7429 ( 
.A(n_6699),
.B(n_4343),
.Y(n_7429)
);

CKINVDCx5p33_ASAP7_75t_R g7430 ( 
.A(n_6897),
.Y(n_7430)
);

CKINVDCx5p33_ASAP7_75t_R g7431 ( 
.A(n_6930),
.Y(n_7431)
);

INVx3_ASAP7_75t_L g7432 ( 
.A(n_6565),
.Y(n_7432)
);

INVx1_ASAP7_75t_L g7433 ( 
.A(n_6845),
.Y(n_7433)
);

INVx2_ASAP7_75t_L g7434 ( 
.A(n_7035),
.Y(n_7434)
);

INVx1_ASAP7_75t_SL g7435 ( 
.A(n_6704),
.Y(n_7435)
);

NOR2xp33_ASAP7_75t_L g7436 ( 
.A(n_7040),
.B(n_4349),
.Y(n_7436)
);

BUFx6f_ASAP7_75t_L g7437 ( 
.A(n_6566),
.Y(n_7437)
);

INVx2_ASAP7_75t_L g7438 ( 
.A(n_7038),
.Y(n_7438)
);

CKINVDCx20_ASAP7_75t_R g7439 ( 
.A(n_6651),
.Y(n_7439)
);

NAND2xp5_ASAP7_75t_L g7440 ( 
.A(n_6817),
.B(n_4351),
.Y(n_7440)
);

CKINVDCx5p33_ASAP7_75t_R g7441 ( 
.A(n_6939),
.Y(n_7441)
);

INVx1_ASAP7_75t_L g7442 ( 
.A(n_6863),
.Y(n_7442)
);

INVx1_ASAP7_75t_L g7443 ( 
.A(n_6867),
.Y(n_7443)
);

INVx1_ASAP7_75t_L g7444 ( 
.A(n_6862),
.Y(n_7444)
);

CKINVDCx20_ASAP7_75t_R g7445 ( 
.A(n_6686),
.Y(n_7445)
);

CKINVDCx11_ASAP7_75t_R g7446 ( 
.A(n_6502),
.Y(n_7446)
);

INVx2_ASAP7_75t_L g7447 ( 
.A(n_6883),
.Y(n_7447)
);

INVx1_ASAP7_75t_L g7448 ( 
.A(n_6879),
.Y(n_7448)
);

INVx1_ASAP7_75t_L g7449 ( 
.A(n_6574),
.Y(n_7449)
);

NOR2xp33_ASAP7_75t_L g7450 ( 
.A(n_6975),
.B(n_4352),
.Y(n_7450)
);

CKINVDCx5p33_ASAP7_75t_R g7451 ( 
.A(n_6966),
.Y(n_7451)
);

INVx2_ASAP7_75t_L g7452 ( 
.A(n_6599),
.Y(n_7452)
);

NOR2xp33_ASAP7_75t_R g7453 ( 
.A(n_6718),
.B(n_5192),
.Y(n_7453)
);

INVx4_ASAP7_75t_L g7454 ( 
.A(n_6737),
.Y(n_7454)
);

NAND2xp5_ASAP7_75t_SL g7455 ( 
.A(n_6706),
.B(n_4353),
.Y(n_7455)
);

OAI21x1_ASAP7_75t_L g7456 ( 
.A1(n_6991),
.A2(n_4813),
.B(n_4802),
.Y(n_7456)
);

AND2x2_ASAP7_75t_L g7457 ( 
.A(n_6749),
.B(n_5337),
.Y(n_7457)
);

INVx3_ASAP7_75t_L g7458 ( 
.A(n_6569),
.Y(n_7458)
);

INVx2_ASAP7_75t_L g7459 ( 
.A(n_6607),
.Y(n_7459)
);

CKINVDCx20_ASAP7_75t_R g7460 ( 
.A(n_6952),
.Y(n_7460)
);

INVx1_ASAP7_75t_L g7461 ( 
.A(n_6667),
.Y(n_7461)
);

INVx1_ASAP7_75t_L g7462 ( 
.A(n_6712),
.Y(n_7462)
);

CKINVDCx20_ASAP7_75t_R g7463 ( 
.A(n_6904),
.Y(n_7463)
);

INVx1_ASAP7_75t_L g7464 ( 
.A(n_6870),
.Y(n_7464)
);

NAND2xp5_ASAP7_75t_L g7465 ( 
.A(n_6756),
.B(n_4354),
.Y(n_7465)
);

INVx1_ASAP7_75t_L g7466 ( 
.A(n_6889),
.Y(n_7466)
);

INVx1_ASAP7_75t_L g7467 ( 
.A(n_6854),
.Y(n_7467)
);

NOR2xp67_ASAP7_75t_L g7468 ( 
.A(n_6956),
.B(n_6983),
.Y(n_7468)
);

BUFx6f_ASAP7_75t_L g7469 ( 
.A(n_6573),
.Y(n_7469)
);

INVx1_ASAP7_75t_L g7470 ( 
.A(n_6522),
.Y(n_7470)
);

INVx1_ASAP7_75t_L g7471 ( 
.A(n_6719),
.Y(n_7471)
);

INVx3_ASAP7_75t_L g7472 ( 
.A(n_6576),
.Y(n_7472)
);

CKINVDCx5p33_ASAP7_75t_R g7473 ( 
.A(n_6917),
.Y(n_7473)
);

INVx1_ASAP7_75t_L g7474 ( 
.A(n_6782),
.Y(n_7474)
);

AND2x2_ASAP7_75t_L g7475 ( 
.A(n_6585),
.B(n_5438),
.Y(n_7475)
);

BUFx10_ASAP7_75t_L g7476 ( 
.A(n_6833),
.Y(n_7476)
);

INVx1_ASAP7_75t_L g7477 ( 
.A(n_6831),
.Y(n_7477)
);

INVx1_ASAP7_75t_L g7478 ( 
.A(n_6687),
.Y(n_7478)
);

INVx2_ASAP7_75t_L g7479 ( 
.A(n_6725),
.Y(n_7479)
);

CKINVDCx5p33_ASAP7_75t_R g7480 ( 
.A(n_6892),
.Y(n_7480)
);

CKINVDCx5p33_ASAP7_75t_R g7481 ( 
.A(n_6899),
.Y(n_7481)
);

CKINVDCx5p33_ASAP7_75t_R g7482 ( 
.A(n_6900),
.Y(n_7482)
);

CKINVDCx5p33_ASAP7_75t_R g7483 ( 
.A(n_6921),
.Y(n_7483)
);

AND2x4_ASAP7_75t_L g7484 ( 
.A(n_7009),
.B(n_4315),
.Y(n_7484)
);

AND2x4_ASAP7_75t_L g7485 ( 
.A(n_7029),
.B(n_4325),
.Y(n_7485)
);

HB1xp67_ASAP7_75t_L g7486 ( 
.A(n_6918),
.Y(n_7486)
);

INVx1_ASAP7_75t_L g7487 ( 
.A(n_6693),
.Y(n_7487)
);

CKINVDCx5p33_ASAP7_75t_R g7488 ( 
.A(n_6931),
.Y(n_7488)
);

INVx1_ASAP7_75t_L g7489 ( 
.A(n_6705),
.Y(n_7489)
);

INVx2_ASAP7_75t_L g7490 ( 
.A(n_6728),
.Y(n_7490)
);

INVx1_ASAP7_75t_L g7491 ( 
.A(n_6716),
.Y(n_7491)
);

AND2x4_ASAP7_75t_L g7492 ( 
.A(n_7039),
.B(n_4328),
.Y(n_7492)
);

CKINVDCx5p33_ASAP7_75t_R g7493 ( 
.A(n_6932),
.Y(n_7493)
);

INVx1_ASAP7_75t_L g7494 ( 
.A(n_6722),
.Y(n_7494)
);

INVx1_ASAP7_75t_L g7495 ( 
.A(n_6730),
.Y(n_7495)
);

CKINVDCx20_ASAP7_75t_R g7496 ( 
.A(n_6823),
.Y(n_7496)
);

NOR2xp33_ASAP7_75t_R g7497 ( 
.A(n_6976),
.B(n_5216),
.Y(n_7497)
);

CKINVDCx5p33_ASAP7_75t_R g7498 ( 
.A(n_6937),
.Y(n_7498)
);

INVx2_ASAP7_75t_L g7499 ( 
.A(n_6734),
.Y(n_7499)
);

INVx1_ASAP7_75t_L g7500 ( 
.A(n_6761),
.Y(n_7500)
);

HB1xp67_ASAP7_75t_L g7501 ( 
.A(n_6936),
.Y(n_7501)
);

INVx1_ASAP7_75t_L g7502 ( 
.A(n_6763),
.Y(n_7502)
);

CKINVDCx5p33_ASAP7_75t_R g7503 ( 
.A(n_6941),
.Y(n_7503)
);

INVx1_ASAP7_75t_L g7504 ( 
.A(n_6768),
.Y(n_7504)
);

BUFx6f_ASAP7_75t_L g7505 ( 
.A(n_6591),
.Y(n_7505)
);

INVx1_ASAP7_75t_L g7506 ( 
.A(n_6796),
.Y(n_7506)
);

INVx1_ASAP7_75t_L g7507 ( 
.A(n_6771),
.Y(n_7507)
);

INVx1_ASAP7_75t_L g7508 ( 
.A(n_6779),
.Y(n_7508)
);

NAND2xp5_ASAP7_75t_SL g7509 ( 
.A(n_6629),
.B(n_4355),
.Y(n_7509)
);

INVx2_ASAP7_75t_L g7510 ( 
.A(n_6745),
.Y(n_7510)
);

CKINVDCx16_ASAP7_75t_R g7511 ( 
.A(n_6631),
.Y(n_7511)
);

NOR2xp33_ASAP7_75t_R g7512 ( 
.A(n_6977),
.B(n_5233),
.Y(n_7512)
);

INVx1_ASAP7_75t_SL g7513 ( 
.A(n_6795),
.Y(n_7513)
);

NAND3xp33_ASAP7_75t_L g7514 ( 
.A(n_7019),
.B(n_4358),
.C(n_4356),
.Y(n_7514)
);

INVx1_ASAP7_75t_SL g7515 ( 
.A(n_6814),
.Y(n_7515)
);

INVx1_ASAP7_75t_L g7516 ( 
.A(n_6808),
.Y(n_7516)
);

INVx4_ASAP7_75t_L g7517 ( 
.A(n_6853),
.Y(n_7517)
);

BUFx6f_ASAP7_75t_L g7518 ( 
.A(n_6598),
.Y(n_7518)
);

CKINVDCx5p33_ASAP7_75t_R g7519 ( 
.A(n_6947),
.Y(n_7519)
);

CKINVDCx5p33_ASAP7_75t_R g7520 ( 
.A(n_6964),
.Y(n_7520)
);

OAI21x1_ASAP7_75t_L g7521 ( 
.A1(n_6537),
.A2(n_4840),
.B(n_4831),
.Y(n_7521)
);

CKINVDCx5p33_ASAP7_75t_R g7522 ( 
.A(n_6953),
.Y(n_7522)
);

CKINVDCx5p33_ASAP7_75t_R g7523 ( 
.A(n_6957),
.Y(n_7523)
);

INVx1_ASAP7_75t_L g7524 ( 
.A(n_6819),
.Y(n_7524)
);

INVxp67_ASAP7_75t_L g7525 ( 
.A(n_6824),
.Y(n_7525)
);

INVx2_ASAP7_75t_L g7526 ( 
.A(n_6757),
.Y(n_7526)
);

INVx4_ASAP7_75t_L g7527 ( 
.A(n_6766),
.Y(n_7527)
);

CKINVDCx16_ASAP7_75t_R g7528 ( 
.A(n_6536),
.Y(n_7528)
);

CKINVDCx5p33_ASAP7_75t_R g7529 ( 
.A(n_6959),
.Y(n_7529)
);

AND2x2_ASAP7_75t_L g7530 ( 
.A(n_6836),
.B(n_5438),
.Y(n_7530)
);

CKINVDCx5p33_ASAP7_75t_R g7531 ( 
.A(n_6965),
.Y(n_7531)
);

NAND2x1_ASAP7_75t_L g7532 ( 
.A(n_6579),
.B(n_4428),
.Y(n_7532)
);

OAI21x1_ASAP7_75t_L g7533 ( 
.A1(n_6623),
.A2(n_4924),
.B(n_4881),
.Y(n_7533)
);

OA21x2_ASAP7_75t_L g7534 ( 
.A1(n_6628),
.A2(n_4331),
.B(n_4329),
.Y(n_7534)
);

HB1xp67_ASAP7_75t_L g7535 ( 
.A(n_6958),
.Y(n_7535)
);

HB1xp67_ASAP7_75t_L g7536 ( 
.A(n_6886),
.Y(n_7536)
);

NOR2xp33_ASAP7_75t_L g7537 ( 
.A(n_6822),
.B(n_4360),
.Y(n_7537)
);

BUFx6f_ASAP7_75t_L g7538 ( 
.A(n_6611),
.Y(n_7538)
);

CKINVDCx5p33_ASAP7_75t_R g7539 ( 
.A(n_6972),
.Y(n_7539)
);

INVx1_ASAP7_75t_L g7540 ( 
.A(n_6834),
.Y(n_7540)
);

AND3x2_ASAP7_75t_L g7541 ( 
.A(n_6927),
.B(n_4949),
.C(n_4933),
.Y(n_7541)
);

CKINVDCx20_ASAP7_75t_R g7542 ( 
.A(n_6925),
.Y(n_7542)
);

INVx3_ASAP7_75t_L g7543 ( 
.A(n_6636),
.Y(n_7543)
);

CKINVDCx20_ASAP7_75t_R g7544 ( 
.A(n_6596),
.Y(n_7544)
);

NAND2xp5_ASAP7_75t_L g7545 ( 
.A(n_6531),
.B(n_4361),
.Y(n_7545)
);

INVx2_ASAP7_75t_L g7546 ( 
.A(n_6769),
.Y(n_7546)
);

INVx1_ASAP7_75t_L g7547 ( 
.A(n_6770),
.Y(n_7547)
);

INVx2_ASAP7_75t_L g7548 ( 
.A(n_6783),
.Y(n_7548)
);

NAND2xp5_ASAP7_75t_L g7549 ( 
.A(n_6541),
.B(n_4364),
.Y(n_7549)
);

HB1xp67_ASAP7_75t_L g7550 ( 
.A(n_6898),
.Y(n_7550)
);

INVx2_ASAP7_75t_L g7551 ( 
.A(n_6784),
.Y(n_7551)
);

INVx1_ASAP7_75t_L g7552 ( 
.A(n_6805),
.Y(n_7552)
);

NAND2xp5_ASAP7_75t_L g7553 ( 
.A(n_6570),
.B(n_4365),
.Y(n_7553)
);

BUFx6f_ASAP7_75t_L g7554 ( 
.A(n_6637),
.Y(n_7554)
);

NAND2xp5_ASAP7_75t_SL g7555 ( 
.A(n_6622),
.B(n_4368),
.Y(n_7555)
);

INVx2_ASAP7_75t_L g7556 ( 
.A(n_6821),
.Y(n_7556)
);

NOR2xp33_ASAP7_75t_L g7557 ( 
.A(n_6940),
.B(n_4369),
.Y(n_7557)
);

AND2x2_ASAP7_75t_L g7558 ( 
.A(n_6970),
.B(n_5442),
.Y(n_7558)
);

CKINVDCx5p33_ASAP7_75t_R g7559 ( 
.A(n_6544),
.Y(n_7559)
);

INVx2_ASAP7_75t_L g7560 ( 
.A(n_6827),
.Y(n_7560)
);

INVx1_ASAP7_75t_L g7561 ( 
.A(n_6832),
.Y(n_7561)
);

INVx1_ASAP7_75t_L g7562 ( 
.A(n_6835),
.Y(n_7562)
);

BUFx2_ASAP7_75t_SL g7563 ( 
.A(n_6974),
.Y(n_7563)
);

HB1xp67_ASAP7_75t_L g7564 ( 
.A(n_6935),
.Y(n_7564)
);

INVx3_ASAP7_75t_L g7565 ( 
.A(n_6648),
.Y(n_7565)
);

NOR2xp33_ASAP7_75t_L g7566 ( 
.A(n_6838),
.B(n_7055),
.Y(n_7566)
);

INVxp33_ASAP7_75t_SL g7567 ( 
.A(n_6791),
.Y(n_7567)
);

INVx1_ASAP7_75t_L g7568 ( 
.A(n_6849),
.Y(n_7568)
);

BUFx2_ASAP7_75t_L g7569 ( 
.A(n_6987),
.Y(n_7569)
);

INVx3_ASAP7_75t_L g7570 ( 
.A(n_6653),
.Y(n_7570)
);

INVx2_ASAP7_75t_L g7571 ( 
.A(n_6860),
.Y(n_7571)
);

HB1xp67_ASAP7_75t_L g7572 ( 
.A(n_6606),
.Y(n_7572)
);

INVx1_ASAP7_75t_L g7573 ( 
.A(n_6861),
.Y(n_7573)
);

CKINVDCx5p33_ASAP7_75t_R g7574 ( 
.A(n_6980),
.Y(n_7574)
);

INVx1_ASAP7_75t_L g7575 ( 
.A(n_6869),
.Y(n_7575)
);

BUFx2_ASAP7_75t_L g7576 ( 
.A(n_6987),
.Y(n_7576)
);

CKINVDCx5p33_ASAP7_75t_R g7577 ( 
.A(n_6984),
.Y(n_7577)
);

BUFx2_ASAP7_75t_L g7578 ( 
.A(n_6973),
.Y(n_7578)
);

INVx2_ASAP7_75t_L g7579 ( 
.A(n_6670),
.Y(n_7579)
);

BUFx6f_ASAP7_75t_L g7580 ( 
.A(n_6673),
.Y(n_7580)
);

BUFx3_ASAP7_75t_L g7581 ( 
.A(n_6632),
.Y(n_7581)
);

NAND2xp5_ASAP7_75t_L g7582 ( 
.A(n_6655),
.B(n_4372),
.Y(n_7582)
);

INVx1_ASAP7_75t_L g7583 ( 
.A(n_6657),
.Y(n_7583)
);

INVx1_ASAP7_75t_L g7584 ( 
.A(n_6676),
.Y(n_7584)
);

CKINVDCx5p33_ASAP7_75t_R g7585 ( 
.A(n_6986),
.Y(n_7585)
);

CKINVDCx5p33_ASAP7_75t_R g7586 ( 
.A(n_6826),
.Y(n_7586)
);

INVx1_ASAP7_75t_L g7587 ( 
.A(n_6702),
.Y(n_7587)
);

CKINVDCx20_ASAP7_75t_R g7588 ( 
.A(n_6982),
.Y(n_7588)
);

CKINVDCx5p33_ASAP7_75t_R g7589 ( 
.A(n_6989),
.Y(n_7589)
);

NAND2xp5_ASAP7_75t_L g7590 ( 
.A(n_7024),
.B(n_4373),
.Y(n_7590)
);

BUFx6f_ASAP7_75t_L g7591 ( 
.A(n_6681),
.Y(n_7591)
);

INVx1_ASAP7_75t_L g7592 ( 
.A(n_6692),
.Y(n_7592)
);

INVx1_ASAP7_75t_L g7593 ( 
.A(n_6703),
.Y(n_7593)
);

INVx1_ASAP7_75t_L g7594 ( 
.A(n_6711),
.Y(n_7594)
);

OAI21x1_ASAP7_75t_L g7595 ( 
.A1(n_6640),
.A2(n_5063),
.B(n_5029),
.Y(n_7595)
);

NAND2xp5_ASAP7_75t_L g7596 ( 
.A(n_7024),
.B(n_4374),
.Y(n_7596)
);

NAND2xp5_ASAP7_75t_SL g7597 ( 
.A(n_7018),
.B(n_4377),
.Y(n_7597)
);

HB1xp67_ASAP7_75t_L g7598 ( 
.A(n_7061),
.Y(n_7598)
);

INVx1_ASAP7_75t_L g7599 ( 
.A(n_6721),
.Y(n_7599)
);

INVx2_ASAP7_75t_L g7600 ( 
.A(n_6697),
.Y(n_7600)
);

CKINVDCx16_ASAP7_75t_R g7601 ( 
.A(n_6679),
.Y(n_7601)
);

NAND2xp5_ASAP7_75t_SL g7602 ( 
.A(n_6543),
.B(n_4379),
.Y(n_7602)
);

INVx1_ASAP7_75t_L g7603 ( 
.A(n_6895),
.Y(n_7603)
);

INVx1_ASAP7_75t_L g7604 ( 
.A(n_6903),
.Y(n_7604)
);

INVx2_ASAP7_75t_L g7605 ( 
.A(n_6990),
.Y(n_7605)
);

INVx1_ASAP7_75t_L g7606 ( 
.A(n_6912),
.Y(n_7606)
);

CKINVDCx5p33_ASAP7_75t_R g7607 ( 
.A(n_6506),
.Y(n_7607)
);

INVx2_ASAP7_75t_L g7608 ( 
.A(n_6738),
.Y(n_7608)
);

AND2x2_ASAP7_75t_L g7609 ( 
.A(n_6993),
.B(n_5442),
.Y(n_7609)
);

CKINVDCx5p33_ASAP7_75t_R g7610 ( 
.A(n_6829),
.Y(n_7610)
);

INVx2_ASAP7_75t_L g7611 ( 
.A(n_6913),
.Y(n_7611)
);

BUFx6f_ASAP7_75t_L g7612 ( 
.A(n_6732),
.Y(n_7612)
);

CKINVDCx20_ASAP7_75t_R g7613 ( 
.A(n_6916),
.Y(n_7613)
);

INVx1_ASAP7_75t_L g7614 ( 
.A(n_6922),
.Y(n_7614)
);

NAND2xp5_ASAP7_75t_L g7615 ( 
.A(n_6732),
.B(n_4381),
.Y(n_7615)
);

INVx1_ASAP7_75t_L g7616 ( 
.A(n_6934),
.Y(n_7616)
);

INVx1_ASAP7_75t_L g7617 ( 
.A(n_6945),
.Y(n_7617)
);

BUFx6f_ASAP7_75t_L g7618 ( 
.A(n_6742),
.Y(n_7618)
);

INVx3_ASAP7_75t_L g7619 ( 
.A(n_6948),
.Y(n_7619)
);

INVx2_ASAP7_75t_L g7620 ( 
.A(n_6742),
.Y(n_7620)
);

NAND2xp5_ASAP7_75t_L g7621 ( 
.A(n_6682),
.B(n_4383),
.Y(n_7621)
);

INVx1_ASAP7_75t_L g7622 ( 
.A(n_6605),
.Y(n_7622)
);

OAI22xp5_ASAP7_75t_SL g7623 ( 
.A1(n_6857),
.A2(n_5236),
.B1(n_5239),
.B2(n_5234),
.Y(n_7623)
);

INVx2_ASAP7_75t_L g7624 ( 
.A(n_6620),
.Y(n_7624)
);

CKINVDCx16_ASAP7_75t_R g7625 ( 
.A(n_6672),
.Y(n_7625)
);

CKINVDCx20_ASAP7_75t_R g7626 ( 
.A(n_6773),
.Y(n_7626)
);

NAND2xp5_ASAP7_75t_L g7627 ( 
.A(n_6527),
.B(n_4384),
.Y(n_7627)
);

INVx2_ASAP7_75t_L g7628 ( 
.A(n_7066),
.Y(n_7628)
);

INVx1_ASAP7_75t_L g7629 ( 
.A(n_7070),
.Y(n_7629)
);

BUFx6f_ASAP7_75t_L g7630 ( 
.A(n_7243),
.Y(n_7630)
);

INVx1_ASAP7_75t_L g7631 ( 
.A(n_7073),
.Y(n_7631)
);

CKINVDCx6p67_ASAP7_75t_R g7632 ( 
.A(n_7317),
.Y(n_7632)
);

INVx2_ASAP7_75t_SL g7633 ( 
.A(n_7080),
.Y(n_7633)
);

AOI22xp33_ASAP7_75t_L g7634 ( 
.A1(n_7566),
.A2(n_6645),
.B1(n_6627),
.B2(n_6868),
.Y(n_7634)
);

OR2x2_ASAP7_75t_L g7635 ( 
.A(n_7224),
.B(n_6882),
.Y(n_7635)
);

INVx1_ASAP7_75t_L g7636 ( 
.A(n_7074),
.Y(n_7636)
);

INVx1_ASAP7_75t_L g7637 ( 
.A(n_7077),
.Y(n_7637)
);

INVx2_ASAP7_75t_L g7638 ( 
.A(n_7069),
.Y(n_7638)
);

INVx1_ASAP7_75t_L g7639 ( 
.A(n_7078),
.Y(n_7639)
);

INVx1_ASAP7_75t_L g7640 ( 
.A(n_7079),
.Y(n_7640)
);

INVx2_ASAP7_75t_L g7641 ( 
.A(n_7072),
.Y(n_7641)
);

NAND2xp33_ASAP7_75t_L g7642 ( 
.A(n_7381),
.B(n_6793),
.Y(n_7642)
);

NAND2xp5_ASAP7_75t_SL g7643 ( 
.A(n_7360),
.B(n_6698),
.Y(n_7643)
);

INVx2_ASAP7_75t_L g7644 ( 
.A(n_7102),
.Y(n_7644)
);

AOI22xp5_ASAP7_75t_L g7645 ( 
.A1(n_7300),
.A2(n_6764),
.B1(n_6710),
.B2(n_5268),
.Y(n_7645)
);

NAND2xp5_ASAP7_75t_SL g7646 ( 
.A(n_7220),
.B(n_5248),
.Y(n_7646)
);

INVx2_ASAP7_75t_L g7647 ( 
.A(n_7107),
.Y(n_7647)
);

INVx1_ASAP7_75t_L g7648 ( 
.A(n_7088),
.Y(n_7648)
);

NOR2xp33_ASAP7_75t_L g7649 ( 
.A(n_7194),
.B(n_6525),
.Y(n_7649)
);

INVx2_ASAP7_75t_L g7650 ( 
.A(n_7122),
.Y(n_7650)
);

INVx2_ASAP7_75t_L g7651 ( 
.A(n_7123),
.Y(n_7651)
);

INVxp33_ASAP7_75t_SL g7652 ( 
.A(n_7419),
.Y(n_7652)
);

INVx1_ASAP7_75t_L g7653 ( 
.A(n_7089),
.Y(n_7653)
);

NAND2xp5_ASAP7_75t_SL g7654 ( 
.A(n_7480),
.B(n_5367),
.Y(n_7654)
);

NAND2xp5_ASAP7_75t_SL g7655 ( 
.A(n_7481),
.B(n_5372),
.Y(n_7655)
);

NAND2xp5_ASAP7_75t_SL g7656 ( 
.A(n_7482),
.B(n_5395),
.Y(n_7656)
);

INVx1_ASAP7_75t_L g7657 ( 
.A(n_7090),
.Y(n_7657)
);

INVxp33_ASAP7_75t_L g7658 ( 
.A(n_7170),
.Y(n_7658)
);

NAND2xp5_ASAP7_75t_L g7659 ( 
.A(n_7319),
.B(n_4386),
.Y(n_7659)
);

INVx2_ASAP7_75t_L g7660 ( 
.A(n_7131),
.Y(n_7660)
);

INVx3_ASAP7_75t_L g7661 ( 
.A(n_7389),
.Y(n_7661)
);

NAND2xp5_ASAP7_75t_SL g7662 ( 
.A(n_7483),
.B(n_5412),
.Y(n_7662)
);

AND2x2_ASAP7_75t_L g7663 ( 
.A(n_7128),
.B(n_5450),
.Y(n_7663)
);

INVx1_ASAP7_75t_L g7664 ( 
.A(n_7093),
.Y(n_7664)
);

INVx2_ASAP7_75t_SL g7665 ( 
.A(n_7379),
.Y(n_7665)
);

INVx1_ASAP7_75t_L g7666 ( 
.A(n_7099),
.Y(n_7666)
);

AO21x2_ASAP7_75t_L g7667 ( 
.A1(n_7416),
.A2(n_4339),
.B(n_4334),
.Y(n_7667)
);

INVx5_ASAP7_75t_L g7668 ( 
.A(n_7082),
.Y(n_7668)
);

BUFx3_ASAP7_75t_L g7669 ( 
.A(n_7243),
.Y(n_7669)
);

INVx2_ASAP7_75t_L g7670 ( 
.A(n_7135),
.Y(n_7670)
);

INVx1_ASAP7_75t_L g7671 ( 
.A(n_7106),
.Y(n_7671)
);

INVx1_ASAP7_75t_L g7672 ( 
.A(n_7111),
.Y(n_7672)
);

BUFx2_ASAP7_75t_L g7673 ( 
.A(n_7235),
.Y(n_7673)
);

NAND2xp5_ASAP7_75t_L g7674 ( 
.A(n_7239),
.B(n_4499),
.Y(n_7674)
);

INVx2_ASAP7_75t_L g7675 ( 
.A(n_7136),
.Y(n_7675)
);

NAND2xp33_ASAP7_75t_L g7676 ( 
.A(n_7382),
.B(n_4385),
.Y(n_7676)
);

INVx1_ASAP7_75t_L g7677 ( 
.A(n_7113),
.Y(n_7677)
);

INVx2_ASAP7_75t_SL g7678 ( 
.A(n_7126),
.Y(n_7678)
);

AND2x2_ASAP7_75t_L g7679 ( 
.A(n_7162),
.B(n_5450),
.Y(n_7679)
);

INVx1_ASAP7_75t_L g7680 ( 
.A(n_7117),
.Y(n_7680)
);

NAND3xp33_ASAP7_75t_L g7681 ( 
.A(n_7537),
.B(n_6981),
.C(n_4388),
.Y(n_7681)
);

NAND2xp33_ASAP7_75t_SL g7682 ( 
.A(n_7612),
.B(n_5415),
.Y(n_7682)
);

NAND2xp5_ASAP7_75t_L g7683 ( 
.A(n_7262),
.B(n_4387),
.Y(n_7683)
);

INVx2_ASAP7_75t_L g7684 ( 
.A(n_7144),
.Y(n_7684)
);

INVx1_ASAP7_75t_L g7685 ( 
.A(n_7125),
.Y(n_7685)
);

BUFx8_ASAP7_75t_SL g7686 ( 
.A(n_7083),
.Y(n_7686)
);

NAND2xp5_ASAP7_75t_L g7687 ( 
.A(n_7289),
.B(n_4390),
.Y(n_7687)
);

NAND3xp33_ASAP7_75t_L g7688 ( 
.A(n_7557),
.B(n_7436),
.C(n_7205),
.Y(n_7688)
);

NAND3xp33_ASAP7_75t_L g7689 ( 
.A(n_7440),
.B(n_4392),
.C(n_4391),
.Y(n_7689)
);

INVx1_ASAP7_75t_L g7690 ( 
.A(n_7130),
.Y(n_7690)
);

AND2x2_ASAP7_75t_L g7691 ( 
.A(n_7261),
.B(n_4399),
.Y(n_7691)
);

INVx2_ASAP7_75t_L g7692 ( 
.A(n_7151),
.Y(n_7692)
);

NAND2xp5_ASAP7_75t_SL g7693 ( 
.A(n_7488),
.B(n_7493),
.Y(n_7693)
);

NAND3xp33_ASAP7_75t_L g7694 ( 
.A(n_7603),
.B(n_7606),
.C(n_7604),
.Y(n_7694)
);

NAND2xp5_ASAP7_75t_L g7695 ( 
.A(n_7467),
.B(n_4401),
.Y(n_7695)
);

AND2x2_ASAP7_75t_L g7696 ( 
.A(n_7249),
.B(n_4405),
.Y(n_7696)
);

INVx1_ASAP7_75t_L g7697 ( 
.A(n_7134),
.Y(n_7697)
);

INVx2_ASAP7_75t_L g7698 ( 
.A(n_7154),
.Y(n_7698)
);

NAND3xp33_ASAP7_75t_SL g7699 ( 
.A(n_7586),
.B(n_5429),
.C(n_5416),
.Y(n_7699)
);

BUFx3_ASAP7_75t_L g7700 ( 
.A(n_7255),
.Y(n_7700)
);

INVx2_ASAP7_75t_L g7701 ( 
.A(n_7177),
.Y(n_7701)
);

INVx2_ASAP7_75t_L g7702 ( 
.A(n_7183),
.Y(n_7702)
);

INVx2_ASAP7_75t_L g7703 ( 
.A(n_7196),
.Y(n_7703)
);

INVx2_ASAP7_75t_L g7704 ( 
.A(n_7199),
.Y(n_7704)
);

INVx4_ASAP7_75t_L g7705 ( 
.A(n_7317),
.Y(n_7705)
);

NOR2xp33_ASAP7_75t_L g7706 ( 
.A(n_7308),
.B(n_6610),
.Y(n_7706)
);

INVx3_ASAP7_75t_L g7707 ( 
.A(n_7389),
.Y(n_7707)
);

NAND2xp5_ASAP7_75t_L g7708 ( 
.A(n_7478),
.B(n_4407),
.Y(n_7708)
);

BUFx2_ASAP7_75t_L g7709 ( 
.A(n_7237),
.Y(n_7709)
);

INVx2_ASAP7_75t_L g7710 ( 
.A(n_7204),
.Y(n_7710)
);

BUFx10_ASAP7_75t_L g7711 ( 
.A(n_7086),
.Y(n_7711)
);

NAND2xp5_ASAP7_75t_SL g7712 ( 
.A(n_7498),
.B(n_5434),
.Y(n_7712)
);

INVx1_ASAP7_75t_L g7713 ( 
.A(n_7140),
.Y(n_7713)
);

INVx2_ASAP7_75t_L g7714 ( 
.A(n_7206),
.Y(n_7714)
);

INVx2_ASAP7_75t_L g7715 ( 
.A(n_7225),
.Y(n_7715)
);

BUFx6f_ASAP7_75t_L g7716 ( 
.A(n_7255),
.Y(n_7716)
);

INVx2_ASAP7_75t_L g7717 ( 
.A(n_7230),
.Y(n_7717)
);

NAND2xp5_ASAP7_75t_L g7718 ( 
.A(n_7487),
.B(n_4408),
.Y(n_7718)
);

INVx2_ASAP7_75t_L g7719 ( 
.A(n_7242),
.Y(n_7719)
);

INVx2_ASAP7_75t_L g7720 ( 
.A(n_7247),
.Y(n_7720)
);

BUFx10_ASAP7_75t_L g7721 ( 
.A(n_7105),
.Y(n_7721)
);

INVx5_ASAP7_75t_L g7722 ( 
.A(n_7244),
.Y(n_7722)
);

NAND2xp5_ASAP7_75t_L g7723 ( 
.A(n_7489),
.B(n_4411),
.Y(n_7723)
);

NOR2xp33_ASAP7_75t_L g7724 ( 
.A(n_7187),
.B(n_5497),
.Y(n_7724)
);

INVxp67_ASAP7_75t_L g7725 ( 
.A(n_7171),
.Y(n_7725)
);

INVx1_ASAP7_75t_L g7726 ( 
.A(n_7152),
.Y(n_7726)
);

INVx2_ASAP7_75t_SL g7727 ( 
.A(n_7302),
.Y(n_7727)
);

NAND2xp5_ASAP7_75t_SL g7728 ( 
.A(n_7503),
.B(n_5506),
.Y(n_7728)
);

INVxp33_ASAP7_75t_SL g7729 ( 
.A(n_7221),
.Y(n_7729)
);

NAND2xp5_ASAP7_75t_L g7730 ( 
.A(n_7491),
.B(n_4414),
.Y(n_7730)
);

INVx1_ASAP7_75t_SL g7731 ( 
.A(n_7403),
.Y(n_7731)
);

INVx1_ASAP7_75t_L g7732 ( 
.A(n_7153),
.Y(n_7732)
);

INVx2_ASAP7_75t_L g7733 ( 
.A(n_7252),
.Y(n_7733)
);

BUFx6f_ASAP7_75t_L g7734 ( 
.A(n_7274),
.Y(n_7734)
);

INVx2_ASAP7_75t_L g7735 ( 
.A(n_7254),
.Y(n_7735)
);

NOR2xp33_ASAP7_75t_L g7736 ( 
.A(n_7435),
.B(n_4415),
.Y(n_7736)
);

AOI22xp33_ASAP7_75t_L g7737 ( 
.A1(n_7444),
.A2(n_5165),
.B1(n_5212),
.B2(n_5066),
.Y(n_7737)
);

NAND2xp5_ASAP7_75t_L g7738 ( 
.A(n_7494),
.B(n_4419),
.Y(n_7738)
);

INVx2_ASAP7_75t_L g7739 ( 
.A(n_7256),
.Y(n_7739)
);

INVx3_ASAP7_75t_L g7740 ( 
.A(n_7394),
.Y(n_7740)
);

NAND2xp5_ASAP7_75t_SL g7741 ( 
.A(n_7519),
.B(n_4422),
.Y(n_7741)
);

INVx3_ASAP7_75t_L g7742 ( 
.A(n_7394),
.Y(n_7742)
);

NAND2xp5_ASAP7_75t_L g7743 ( 
.A(n_7495),
.B(n_4426),
.Y(n_7743)
);

INVx1_ASAP7_75t_SL g7744 ( 
.A(n_7331),
.Y(n_7744)
);

NAND2xp5_ASAP7_75t_L g7745 ( 
.A(n_7500),
.B(n_4427),
.Y(n_7745)
);

INVx2_ASAP7_75t_L g7746 ( 
.A(n_7270),
.Y(n_7746)
);

INVx2_ASAP7_75t_SL g7747 ( 
.A(n_7362),
.Y(n_7747)
);

NAND2xp33_ASAP7_75t_SL g7748 ( 
.A(n_7612),
.B(n_4430),
.Y(n_7748)
);

INVx2_ASAP7_75t_L g7749 ( 
.A(n_7156),
.Y(n_7749)
);

INVx1_ASAP7_75t_L g7750 ( 
.A(n_7160),
.Y(n_7750)
);

INVxp67_ASAP7_75t_L g7751 ( 
.A(n_7229),
.Y(n_7751)
);

INVx2_ASAP7_75t_L g7752 ( 
.A(n_7165),
.Y(n_7752)
);

INVx2_ASAP7_75t_L g7753 ( 
.A(n_7169),
.Y(n_7753)
);

NAND2xp5_ASAP7_75t_SL g7754 ( 
.A(n_7520),
.B(n_4433),
.Y(n_7754)
);

INVx2_ASAP7_75t_L g7755 ( 
.A(n_7172),
.Y(n_7755)
);

INVx2_ASAP7_75t_L g7756 ( 
.A(n_7174),
.Y(n_7756)
);

INVx2_ASAP7_75t_SL g7757 ( 
.A(n_7248),
.Y(n_7757)
);

INVx2_ASAP7_75t_L g7758 ( 
.A(n_7175),
.Y(n_7758)
);

NAND2xp5_ASAP7_75t_L g7759 ( 
.A(n_7502),
.B(n_4437),
.Y(n_7759)
);

NOR2xp33_ASAP7_75t_L g7760 ( 
.A(n_7513),
.B(n_4440),
.Y(n_7760)
);

NOR2xp33_ASAP7_75t_L g7761 ( 
.A(n_7515),
.B(n_4441),
.Y(n_7761)
);

INVx2_ASAP7_75t_L g7762 ( 
.A(n_7180),
.Y(n_7762)
);

INVx3_ASAP7_75t_L g7763 ( 
.A(n_7412),
.Y(n_7763)
);

BUFx6f_ASAP7_75t_L g7764 ( 
.A(n_7274),
.Y(n_7764)
);

INVx2_ASAP7_75t_L g7765 ( 
.A(n_7181),
.Y(n_7765)
);

BUFx6f_ASAP7_75t_L g7766 ( 
.A(n_7081),
.Y(n_7766)
);

NAND2xp5_ASAP7_75t_SL g7767 ( 
.A(n_7315),
.B(n_4442),
.Y(n_7767)
);

NAND2xp5_ASAP7_75t_L g7768 ( 
.A(n_7504),
.B(n_4446),
.Y(n_7768)
);

INVx2_ASAP7_75t_L g7769 ( 
.A(n_7184),
.Y(n_7769)
);

INVx2_ASAP7_75t_L g7770 ( 
.A(n_7188),
.Y(n_7770)
);

INVx2_ASAP7_75t_L g7771 ( 
.A(n_7190),
.Y(n_7771)
);

INVx1_ASAP7_75t_L g7772 ( 
.A(n_7191),
.Y(n_7772)
);

AOI22xp5_ASAP7_75t_L g7773 ( 
.A1(n_7401),
.A2(n_4448),
.B1(n_4449),
.B2(n_4447),
.Y(n_7773)
);

INVx2_ASAP7_75t_L g7774 ( 
.A(n_7192),
.Y(n_7774)
);

INVx2_ASAP7_75t_SL g7775 ( 
.A(n_7095),
.Y(n_7775)
);

INVx3_ASAP7_75t_L g7776 ( 
.A(n_7412),
.Y(n_7776)
);

INVx1_ASAP7_75t_L g7777 ( 
.A(n_7195),
.Y(n_7777)
);

CKINVDCx5p33_ASAP7_75t_R g7778 ( 
.A(n_7076),
.Y(n_7778)
);

INVx1_ASAP7_75t_L g7779 ( 
.A(n_7198),
.Y(n_7779)
);

BUFx6f_ASAP7_75t_L g7780 ( 
.A(n_7081),
.Y(n_7780)
);

INVx1_ASAP7_75t_L g7781 ( 
.A(n_7207),
.Y(n_7781)
);

INVx2_ASAP7_75t_L g7782 ( 
.A(n_7213),
.Y(n_7782)
);

INVx2_ASAP7_75t_L g7783 ( 
.A(n_7216),
.Y(n_7783)
);

INVx1_ASAP7_75t_L g7784 ( 
.A(n_7236),
.Y(n_7784)
);

INVx1_ASAP7_75t_L g7785 ( 
.A(n_7238),
.Y(n_7785)
);

NOR2xp33_ASAP7_75t_L g7786 ( 
.A(n_7176),
.B(n_4454),
.Y(n_7786)
);

INVx2_ASAP7_75t_L g7787 ( 
.A(n_7246),
.Y(n_7787)
);

OAI22xp33_ASAP7_75t_L g7788 ( 
.A1(n_7622),
.A2(n_4456),
.B1(n_4461),
.B2(n_4455),
.Y(n_7788)
);

INVx3_ASAP7_75t_L g7789 ( 
.A(n_7437),
.Y(n_7789)
);

INVx1_ASAP7_75t_L g7790 ( 
.A(n_7253),
.Y(n_7790)
);

INVx2_ASAP7_75t_L g7791 ( 
.A(n_7265),
.Y(n_7791)
);

INVx2_ASAP7_75t_L g7792 ( 
.A(n_7266),
.Y(n_7792)
);

INVx3_ASAP7_75t_L g7793 ( 
.A(n_7437),
.Y(n_7793)
);

NAND2xp5_ASAP7_75t_L g7794 ( 
.A(n_7506),
.B(n_4465),
.Y(n_7794)
);

INVx3_ASAP7_75t_L g7795 ( 
.A(n_7469),
.Y(n_7795)
);

CKINVDCx5p33_ASAP7_75t_R g7796 ( 
.A(n_7085),
.Y(n_7796)
);

NOR2xp33_ASAP7_75t_L g7797 ( 
.A(n_7525),
.B(n_4467),
.Y(n_7797)
);

NAND2xp5_ASAP7_75t_L g7798 ( 
.A(n_7450),
.B(n_4471),
.Y(n_7798)
);

INVx2_ASAP7_75t_L g7799 ( 
.A(n_7268),
.Y(n_7799)
);

INVx8_ASAP7_75t_L g7800 ( 
.A(n_7390),
.Y(n_7800)
);

INVx3_ASAP7_75t_L g7801 ( 
.A(n_7469),
.Y(n_7801)
);

OR2x2_ASAP7_75t_L g7802 ( 
.A(n_7133),
.B(n_4473),
.Y(n_7802)
);

INVx1_ASAP7_75t_L g7803 ( 
.A(n_7269),
.Y(n_7803)
);

NAND2xp5_ASAP7_75t_L g7804 ( 
.A(n_7464),
.B(n_4475),
.Y(n_7804)
);

BUFx3_ASAP7_75t_L g7805 ( 
.A(n_7101),
.Y(n_7805)
);

INVx1_ASAP7_75t_L g7806 ( 
.A(n_7280),
.Y(n_7806)
);

INVx2_ASAP7_75t_L g7807 ( 
.A(n_7281),
.Y(n_7807)
);

INVx2_ASAP7_75t_L g7808 ( 
.A(n_7282),
.Y(n_7808)
);

NOR2xp33_ASAP7_75t_L g7809 ( 
.A(n_7619),
.B(n_4479),
.Y(n_7809)
);

XNOR2xp5_ASAP7_75t_L g7810 ( 
.A(n_7108),
.B(n_4481),
.Y(n_7810)
);

INVx2_ASAP7_75t_L g7811 ( 
.A(n_7287),
.Y(n_7811)
);

INVx1_ASAP7_75t_SL g7812 ( 
.A(n_7542),
.Y(n_7812)
);

INVx2_ASAP7_75t_SL g7813 ( 
.A(n_7091),
.Y(n_7813)
);

INVx2_ASAP7_75t_L g7814 ( 
.A(n_7297),
.Y(n_7814)
);

INVx1_ASAP7_75t_L g7815 ( 
.A(n_7299),
.Y(n_7815)
);

OR2x2_ASAP7_75t_L g7816 ( 
.A(n_7215),
.B(n_4482),
.Y(n_7816)
);

INVx1_ASAP7_75t_L g7817 ( 
.A(n_7313),
.Y(n_7817)
);

NAND2xp33_ASAP7_75t_SL g7818 ( 
.A(n_7618),
.B(n_4484),
.Y(n_7818)
);

INVx1_ASAP7_75t_L g7819 ( 
.A(n_7316),
.Y(n_7819)
);

INVx1_ASAP7_75t_L g7820 ( 
.A(n_7231),
.Y(n_7820)
);

BUFx4f_ASAP7_75t_L g7821 ( 
.A(n_7618),
.Y(n_7821)
);

CKINVDCx5p33_ASAP7_75t_R g7822 ( 
.A(n_7098),
.Y(n_7822)
);

INVx2_ASAP7_75t_L g7823 ( 
.A(n_7323),
.Y(n_7823)
);

NOR2xp33_ASAP7_75t_L g7824 ( 
.A(n_7589),
.B(n_4486),
.Y(n_7824)
);

INVx2_ASAP7_75t_L g7825 ( 
.A(n_7325),
.Y(n_7825)
);

INVx2_ASAP7_75t_L g7826 ( 
.A(n_7330),
.Y(n_7826)
);

INVxp33_ASAP7_75t_L g7827 ( 
.A(n_7245),
.Y(n_7827)
);

INVx1_ASAP7_75t_L g7828 ( 
.A(n_7333),
.Y(n_7828)
);

NAND2xp5_ASAP7_75t_L g7829 ( 
.A(n_7466),
.B(n_4493),
.Y(n_7829)
);

NAND2xp5_ASAP7_75t_SL g7830 ( 
.A(n_7366),
.B(n_4497),
.Y(n_7830)
);

INVx2_ASAP7_75t_L g7831 ( 
.A(n_7291),
.Y(n_7831)
);

INVx2_ASAP7_75t_L g7832 ( 
.A(n_7294),
.Y(n_7832)
);

INVx2_ASAP7_75t_L g7833 ( 
.A(n_7318),
.Y(n_7833)
);

INVx8_ASAP7_75t_L g7834 ( 
.A(n_7227),
.Y(n_7834)
);

INVx2_ASAP7_75t_L g7835 ( 
.A(n_7334),
.Y(n_7835)
);

INVx3_ASAP7_75t_L g7836 ( 
.A(n_7505),
.Y(n_7836)
);

NOR2xp33_ASAP7_75t_L g7837 ( 
.A(n_7522),
.B(n_7523),
.Y(n_7837)
);

INVx1_ASAP7_75t_L g7838 ( 
.A(n_7342),
.Y(n_7838)
);

INVx2_ASAP7_75t_L g7839 ( 
.A(n_7339),
.Y(n_7839)
);

INVx1_ASAP7_75t_L g7840 ( 
.A(n_7343),
.Y(n_7840)
);

INVx2_ASAP7_75t_L g7841 ( 
.A(n_7341),
.Y(n_7841)
);

INVx1_ASAP7_75t_L g7842 ( 
.A(n_7344),
.Y(n_7842)
);

INVx1_ASAP7_75t_L g7843 ( 
.A(n_7345),
.Y(n_7843)
);

BUFx6f_ASAP7_75t_L g7844 ( 
.A(n_7101),
.Y(n_7844)
);

INVx1_ASAP7_75t_L g7845 ( 
.A(n_7350),
.Y(n_7845)
);

INVx2_ASAP7_75t_SL g7846 ( 
.A(n_7358),
.Y(n_7846)
);

INVx1_ASAP7_75t_L g7847 ( 
.A(n_7351),
.Y(n_7847)
);

INVx1_ASAP7_75t_L g7848 ( 
.A(n_7352),
.Y(n_7848)
);

INVx1_ASAP7_75t_L g7849 ( 
.A(n_7357),
.Y(n_7849)
);

INVx2_ASAP7_75t_L g7850 ( 
.A(n_7346),
.Y(n_7850)
);

BUFx6f_ASAP7_75t_L g7851 ( 
.A(n_7168),
.Y(n_7851)
);

NAND3xp33_ASAP7_75t_L g7852 ( 
.A(n_7614),
.B(n_4505),
.C(n_4504),
.Y(n_7852)
);

BUFx10_ASAP7_75t_L g7853 ( 
.A(n_7112),
.Y(n_7853)
);

NAND2xp5_ASAP7_75t_SL g7854 ( 
.A(n_7511),
.B(n_4507),
.Y(n_7854)
);

INVx2_ASAP7_75t_L g7855 ( 
.A(n_7349),
.Y(n_7855)
);

INVx1_ASAP7_75t_L g7856 ( 
.A(n_7368),
.Y(n_7856)
);

NAND2xp5_ASAP7_75t_L g7857 ( 
.A(n_7328),
.B(n_4508),
.Y(n_7857)
);

INVx2_ASAP7_75t_L g7858 ( 
.A(n_7354),
.Y(n_7858)
);

NOR2xp33_ASAP7_75t_L g7859 ( 
.A(n_7529),
.B(n_4512),
.Y(n_7859)
);

INVx1_ASAP7_75t_L g7860 ( 
.A(n_7369),
.Y(n_7860)
);

INVx1_ASAP7_75t_L g7861 ( 
.A(n_7375),
.Y(n_7861)
);

INVx2_ASAP7_75t_L g7862 ( 
.A(n_7355),
.Y(n_7862)
);

INVx1_ASAP7_75t_L g7863 ( 
.A(n_7376),
.Y(n_7863)
);

INVx1_ASAP7_75t_L g7864 ( 
.A(n_7377),
.Y(n_7864)
);

NAND3xp33_ASAP7_75t_L g7865 ( 
.A(n_7616),
.B(n_4515),
.C(n_4514),
.Y(n_7865)
);

INVx2_ASAP7_75t_L g7866 ( 
.A(n_7361),
.Y(n_7866)
);

INVx1_ASAP7_75t_L g7867 ( 
.A(n_7378),
.Y(n_7867)
);

INVx1_ASAP7_75t_L g7868 ( 
.A(n_7380),
.Y(n_7868)
);

NOR2xp33_ASAP7_75t_L g7869 ( 
.A(n_7531),
.B(n_4516),
.Y(n_7869)
);

NAND2xp5_ASAP7_75t_SL g7870 ( 
.A(n_7539),
.B(n_4517),
.Y(n_7870)
);

INVx2_ASAP7_75t_L g7871 ( 
.A(n_7373),
.Y(n_7871)
);

BUFx6f_ASAP7_75t_L g7872 ( 
.A(n_7168),
.Y(n_7872)
);

INVx2_ASAP7_75t_L g7873 ( 
.A(n_7387),
.Y(n_7873)
);

INVx3_ASAP7_75t_L g7874 ( 
.A(n_7505),
.Y(n_7874)
);

INVx2_ASAP7_75t_L g7875 ( 
.A(n_7395),
.Y(n_7875)
);

INVx4_ASAP7_75t_L g7876 ( 
.A(n_7232),
.Y(n_7876)
);

INVx2_ASAP7_75t_L g7877 ( 
.A(n_7397),
.Y(n_7877)
);

INVx2_ASAP7_75t_L g7878 ( 
.A(n_7398),
.Y(n_7878)
);

INVx2_ASAP7_75t_SL g7879 ( 
.A(n_7314),
.Y(n_7879)
);

INVx1_ASAP7_75t_L g7880 ( 
.A(n_7383),
.Y(n_7880)
);

INVx2_ASAP7_75t_L g7881 ( 
.A(n_7399),
.Y(n_7881)
);

INVx2_ASAP7_75t_L g7882 ( 
.A(n_7405),
.Y(n_7882)
);

AOI22xp33_ASAP7_75t_L g7883 ( 
.A1(n_7340),
.A2(n_5257),
.B1(n_5324),
.B2(n_5226),
.Y(n_7883)
);

INVx2_ASAP7_75t_L g7884 ( 
.A(n_7408),
.Y(n_7884)
);

NAND2xp33_ASAP7_75t_L g7885 ( 
.A(n_7384),
.B(n_4519),
.Y(n_7885)
);

BUFx2_ASAP7_75t_L g7886 ( 
.A(n_7613),
.Y(n_7886)
);

INVx2_ASAP7_75t_L g7887 ( 
.A(n_7409),
.Y(n_7887)
);

INVx2_ASAP7_75t_SL g7888 ( 
.A(n_7335),
.Y(n_7888)
);

INVx2_ASAP7_75t_L g7889 ( 
.A(n_7414),
.Y(n_7889)
);

INVx3_ASAP7_75t_L g7890 ( 
.A(n_7518),
.Y(n_7890)
);

NAND2xp5_ASAP7_75t_SL g7891 ( 
.A(n_7336),
.B(n_4520),
.Y(n_7891)
);

INVx2_ASAP7_75t_L g7892 ( 
.A(n_7271),
.Y(n_7892)
);

INVx2_ASAP7_75t_SL g7893 ( 
.A(n_7611),
.Y(n_7893)
);

INVx2_ASAP7_75t_L g7894 ( 
.A(n_7272),
.Y(n_7894)
);

NAND2xp5_ASAP7_75t_L g7895 ( 
.A(n_7516),
.B(n_4523),
.Y(n_7895)
);

AND3x2_ASAP7_75t_L g7896 ( 
.A(n_7578),
.B(n_4342),
.C(n_4341),
.Y(n_7896)
);

INVx2_ASAP7_75t_SL g7897 ( 
.A(n_7364),
.Y(n_7897)
);

NAND2xp5_ASAP7_75t_SL g7898 ( 
.A(n_7337),
.B(n_4525),
.Y(n_7898)
);

NAND2xp5_ASAP7_75t_L g7899 ( 
.A(n_7524),
.B(n_4526),
.Y(n_7899)
);

INVx2_ASAP7_75t_L g7900 ( 
.A(n_7275),
.Y(n_7900)
);

INVx1_ASAP7_75t_L g7901 ( 
.A(n_7386),
.Y(n_7901)
);

INVx2_ASAP7_75t_L g7902 ( 
.A(n_7404),
.Y(n_7902)
);

NOR2xp33_ASAP7_75t_L g7903 ( 
.A(n_7574),
.B(n_4530),
.Y(n_7903)
);

AOI21x1_ASAP7_75t_L g7904 ( 
.A1(n_7471),
.A2(n_4350),
.B(n_4344),
.Y(n_7904)
);

INVx2_ASAP7_75t_L g7905 ( 
.A(n_7406),
.Y(n_7905)
);

INVx1_ASAP7_75t_L g7906 ( 
.A(n_7407),
.Y(n_7906)
);

INVx1_ASAP7_75t_L g7907 ( 
.A(n_7410),
.Y(n_7907)
);

INVx1_ASAP7_75t_L g7908 ( 
.A(n_7420),
.Y(n_7908)
);

BUFx6f_ASAP7_75t_SL g7909 ( 
.A(n_7332),
.Y(n_7909)
);

INVx1_ASAP7_75t_L g7910 ( 
.A(n_7096),
.Y(n_7910)
);

AOI22xp5_ASAP7_75t_L g7911 ( 
.A1(n_7425),
.A2(n_4533),
.B1(n_4535),
.B2(n_4531),
.Y(n_7911)
);

INVx2_ASAP7_75t_L g7912 ( 
.A(n_7233),
.Y(n_7912)
);

NAND2xp5_ASAP7_75t_L g7913 ( 
.A(n_7540),
.B(n_4536),
.Y(n_7913)
);

INVx1_ASAP7_75t_L g7914 ( 
.A(n_7338),
.Y(n_7914)
);

INVx2_ASAP7_75t_L g7915 ( 
.A(n_7278),
.Y(n_7915)
);

INVx2_ASAP7_75t_L g7916 ( 
.A(n_7278),
.Y(n_7916)
);

INVx8_ASAP7_75t_L g7917 ( 
.A(n_7234),
.Y(n_7917)
);

INVx1_ASAP7_75t_L g7918 ( 
.A(n_7422),
.Y(n_7918)
);

INVx2_ASAP7_75t_L g7919 ( 
.A(n_7288),
.Y(n_7919)
);

INVx5_ASAP7_75t_L g7920 ( 
.A(n_7454),
.Y(n_7920)
);

INVx2_ASAP7_75t_L g7921 ( 
.A(n_7288),
.Y(n_7921)
);

INVx2_ASAP7_75t_L g7922 ( 
.A(n_7324),
.Y(n_7922)
);

INVx2_ASAP7_75t_L g7923 ( 
.A(n_7324),
.Y(n_7923)
);

INVx3_ASAP7_75t_L g7924 ( 
.A(n_7518),
.Y(n_7924)
);

AO21x2_ASAP7_75t_L g7925 ( 
.A1(n_7474),
.A2(n_4367),
.B(n_4363),
.Y(n_7925)
);

BUFx6f_ASAP7_75t_L g7926 ( 
.A(n_7208),
.Y(n_7926)
);

NOR3xp33_ASAP7_75t_L g7927 ( 
.A(n_7623),
.B(n_4538),
.C(n_4537),
.Y(n_7927)
);

INVx1_ASAP7_75t_L g7928 ( 
.A(n_7423),
.Y(n_7928)
);

NAND2xp5_ASAP7_75t_L g7929 ( 
.A(n_7114),
.B(n_4545),
.Y(n_7929)
);

NAND2xp5_ASAP7_75t_SL g7930 ( 
.A(n_7428),
.B(n_4547),
.Y(n_7930)
);

AND2x6_ASAP7_75t_L g7931 ( 
.A(n_7620),
.B(n_7448),
.Y(n_7931)
);

NOR2xp33_ASAP7_75t_L g7932 ( 
.A(n_7577),
.B(n_4549),
.Y(n_7932)
);

AOI21x1_ASAP7_75t_L g7933 ( 
.A1(n_7477),
.A2(n_4376),
.B(n_4375),
.Y(n_7933)
);

INVx1_ASAP7_75t_L g7934 ( 
.A(n_7449),
.Y(n_7934)
);

INVx2_ASAP7_75t_L g7935 ( 
.A(n_7452),
.Y(n_7935)
);

BUFx2_ASAP7_75t_L g7936 ( 
.A(n_7385),
.Y(n_7936)
);

INVx1_ASAP7_75t_SL g7937 ( 
.A(n_7392),
.Y(n_7937)
);

INVx2_ASAP7_75t_L g7938 ( 
.A(n_7459),
.Y(n_7938)
);

INVx3_ASAP7_75t_L g7939 ( 
.A(n_7538),
.Y(n_7939)
);

NOR2xp33_ASAP7_75t_L g7940 ( 
.A(n_7585),
.B(n_4555),
.Y(n_7940)
);

INVx2_ASAP7_75t_L g7941 ( 
.A(n_7087),
.Y(n_7941)
);

BUFx3_ASAP7_75t_L g7942 ( 
.A(n_7208),
.Y(n_7942)
);

INVx1_ASAP7_75t_L g7943 ( 
.A(n_7461),
.Y(n_7943)
);

AOI21x1_ASAP7_75t_L g7944 ( 
.A1(n_7434),
.A2(n_7438),
.B(n_7110),
.Y(n_7944)
);

AO21x2_ASAP7_75t_L g7945 ( 
.A1(n_7456),
.A2(n_4393),
.B(n_4378),
.Y(n_7945)
);

NOR2xp33_ASAP7_75t_L g7946 ( 
.A(n_7185),
.B(n_4558),
.Y(n_7946)
);

INVx3_ASAP7_75t_L g7947 ( 
.A(n_7538),
.Y(n_7947)
);

INVx1_ASAP7_75t_L g7948 ( 
.A(n_7462),
.Y(n_7948)
);

INVx2_ASAP7_75t_L g7949 ( 
.A(n_7104),
.Y(n_7949)
);

NAND2xp5_ASAP7_75t_SL g7950 ( 
.A(n_7430),
.B(n_4562),
.Y(n_7950)
);

INVx1_ASAP7_75t_L g7951 ( 
.A(n_7426),
.Y(n_7951)
);

NAND2xp5_ASAP7_75t_L g7952 ( 
.A(n_7365),
.B(n_7264),
.Y(n_7952)
);

INVx3_ASAP7_75t_L g7953 ( 
.A(n_7554),
.Y(n_7953)
);

INVx2_ASAP7_75t_L g7954 ( 
.A(n_7433),
.Y(n_7954)
);

INVx2_ASAP7_75t_SL g7955 ( 
.A(n_7372),
.Y(n_7955)
);

NAND2xp5_ASAP7_75t_SL g7956 ( 
.A(n_7431),
.B(n_4563),
.Y(n_7956)
);

INVx1_ASAP7_75t_L g7957 ( 
.A(n_7442),
.Y(n_7957)
);

INVx2_ASAP7_75t_SL g7958 ( 
.A(n_7424),
.Y(n_7958)
);

NAND3xp33_ASAP7_75t_L g7959 ( 
.A(n_7617),
.B(n_4568),
.C(n_4565),
.Y(n_7959)
);

NAND2xp33_ASAP7_75t_L g7960 ( 
.A(n_7400),
.B(n_4569),
.Y(n_7960)
);

INVx2_ASAP7_75t_L g7961 ( 
.A(n_7443),
.Y(n_7961)
);

INVx2_ASAP7_75t_L g7962 ( 
.A(n_7534),
.Y(n_7962)
);

NOR2x1p5_ASAP7_75t_L g7963 ( 
.A(n_7240),
.B(n_4572),
.Y(n_7963)
);

INVx2_ASAP7_75t_L g7964 ( 
.A(n_7075),
.Y(n_7964)
);

INVxp33_ASAP7_75t_L g7965 ( 
.A(n_7209),
.Y(n_7965)
);

NAND2xp5_ASAP7_75t_SL g7966 ( 
.A(n_7441),
.B(n_4576),
.Y(n_7966)
);

INVx1_ASAP7_75t_L g7967 ( 
.A(n_7092),
.Y(n_7967)
);

NAND2xp5_ASAP7_75t_SL g7968 ( 
.A(n_7451),
.B(n_4577),
.Y(n_7968)
);

BUFx4f_ASAP7_75t_L g7969 ( 
.A(n_7210),
.Y(n_7969)
);

INVx2_ASAP7_75t_L g7970 ( 
.A(n_7447),
.Y(n_7970)
);

INVx5_ASAP7_75t_L g7971 ( 
.A(n_7100),
.Y(n_7971)
);

NOR2xp33_ASAP7_75t_L g7972 ( 
.A(n_7624),
.B(n_4585),
.Y(n_7972)
);

INVx1_ASAP7_75t_L g7973 ( 
.A(n_7097),
.Y(n_7973)
);

INVx1_ASAP7_75t_L g7974 ( 
.A(n_7116),
.Y(n_7974)
);

BUFx4f_ASAP7_75t_L g7975 ( 
.A(n_7210),
.Y(n_7975)
);

INVxp67_ASAP7_75t_L g7976 ( 
.A(n_7296),
.Y(n_7976)
);

INVx2_ASAP7_75t_L g7977 ( 
.A(n_7094),
.Y(n_7977)
);

NAND2xp5_ASAP7_75t_SL g7978 ( 
.A(n_7605),
.B(n_4587),
.Y(n_7978)
);

AND3x2_ASAP7_75t_L g7979 ( 
.A(n_7569),
.B(n_4398),
.C(n_4395),
.Y(n_7979)
);

INVx2_ASAP7_75t_L g7980 ( 
.A(n_7109),
.Y(n_7980)
);

NAND2xp5_ASAP7_75t_SL g7981 ( 
.A(n_7558),
.B(n_4589),
.Y(n_7981)
);

INVx1_ASAP7_75t_L g7982 ( 
.A(n_7159),
.Y(n_7982)
);

INVx2_ASAP7_75t_L g7983 ( 
.A(n_7292),
.Y(n_7983)
);

INVx2_ASAP7_75t_L g7984 ( 
.A(n_7370),
.Y(n_7984)
);

INVx2_ASAP7_75t_L g7985 ( 
.A(n_7402),
.Y(n_7985)
);

NAND2xp5_ASAP7_75t_L g7986 ( 
.A(n_7388),
.B(n_7475),
.Y(n_7986)
);

OR2x2_ASAP7_75t_L g7987 ( 
.A(n_7627),
.B(n_4591),
.Y(n_7987)
);

INVx1_ASAP7_75t_L g7988 ( 
.A(n_7203),
.Y(n_7988)
);

INVx1_ASAP7_75t_L g7989 ( 
.A(n_7211),
.Y(n_7989)
);

INVx1_ASAP7_75t_L g7990 ( 
.A(n_7217),
.Y(n_7990)
);

INVx2_ASAP7_75t_L g7991 ( 
.A(n_7479),
.Y(n_7991)
);

INVx2_ASAP7_75t_L g7992 ( 
.A(n_7490),
.Y(n_7992)
);

INVx2_ASAP7_75t_L g7993 ( 
.A(n_7499),
.Y(n_7993)
);

INVx2_ASAP7_75t_L g7994 ( 
.A(n_7510),
.Y(n_7994)
);

INVx2_ASAP7_75t_L g7995 ( 
.A(n_7526),
.Y(n_7995)
);

INVx2_ASAP7_75t_L g7996 ( 
.A(n_7546),
.Y(n_7996)
);

INVx2_ASAP7_75t_SL g7997 ( 
.A(n_7554),
.Y(n_7997)
);

NAND2xp5_ASAP7_75t_L g7998 ( 
.A(n_7400),
.B(n_4592),
.Y(n_7998)
);

NAND3xp33_ASAP7_75t_L g7999 ( 
.A(n_7514),
.B(n_4595),
.C(n_4594),
.Y(n_7999)
);

NAND2xp5_ASAP7_75t_L g8000 ( 
.A(n_7400),
.B(n_4600),
.Y(n_8000)
);

INVx1_ASAP7_75t_L g8001 ( 
.A(n_7507),
.Y(n_8001)
);

INVx1_ASAP7_75t_L g8002 ( 
.A(n_7508),
.Y(n_8002)
);

INVx2_ASAP7_75t_SL g8003 ( 
.A(n_7580),
.Y(n_8003)
);

INVx1_ASAP7_75t_L g8004 ( 
.A(n_7583),
.Y(n_8004)
);

NAND2xp5_ASAP7_75t_L g8005 ( 
.A(n_7312),
.B(n_7415),
.Y(n_8005)
);

INVx1_ASAP7_75t_L g8006 ( 
.A(n_7584),
.Y(n_8006)
);

INVx1_ASAP7_75t_L g8007 ( 
.A(n_7587),
.Y(n_8007)
);

INVx2_ASAP7_75t_L g8008 ( 
.A(n_7548),
.Y(n_8008)
);

NOR2xp33_ASAP7_75t_L g8009 ( 
.A(n_7167),
.B(n_4602),
.Y(n_8009)
);

INVx1_ASAP7_75t_L g8010 ( 
.A(n_7470),
.Y(n_8010)
);

INVx2_ASAP7_75t_L g8011 ( 
.A(n_7551),
.Y(n_8011)
);

INVx1_ASAP7_75t_L g8012 ( 
.A(n_7486),
.Y(n_8012)
);

INVx8_ASAP7_75t_L g8013 ( 
.A(n_7250),
.Y(n_8013)
);

INVx2_ASAP7_75t_L g8014 ( 
.A(n_7556),
.Y(n_8014)
);

INVx2_ASAP7_75t_L g8015 ( 
.A(n_7560),
.Y(n_8015)
);

INVx2_ASAP7_75t_L g8016 ( 
.A(n_7571),
.Y(n_8016)
);

AND2x6_ASAP7_75t_L g8017 ( 
.A(n_7608),
.B(n_4400),
.Y(n_8017)
);

INVx3_ASAP7_75t_L g8018 ( 
.A(n_7580),
.Y(n_8018)
);

CKINVDCx6p67_ASAP7_75t_R g8019 ( 
.A(n_7446),
.Y(n_8019)
);

INVx2_ASAP7_75t_L g8020 ( 
.A(n_7521),
.Y(n_8020)
);

NOR2xp33_ASAP7_75t_L g8021 ( 
.A(n_7129),
.B(n_4604),
.Y(n_8021)
);

BUFx4f_ASAP7_75t_L g8022 ( 
.A(n_7222),
.Y(n_8022)
);

AOI22xp5_ASAP7_75t_L g8023 ( 
.A1(n_7501),
.A2(n_4608),
.B1(n_4610),
.B2(n_4607),
.Y(n_8023)
);

INVx2_ASAP7_75t_L g8024 ( 
.A(n_7533),
.Y(n_8024)
);

BUFx6f_ASAP7_75t_SL g8025 ( 
.A(n_7301),
.Y(n_8025)
);

INVx1_ASAP7_75t_L g8026 ( 
.A(n_7535),
.Y(n_8026)
);

INVx1_ASAP7_75t_L g8027 ( 
.A(n_7547),
.Y(n_8027)
);

INVx1_ASAP7_75t_L g8028 ( 
.A(n_7552),
.Y(n_8028)
);

NAND2xp5_ASAP7_75t_SL g8029 ( 
.A(n_7310),
.B(n_4612),
.Y(n_8029)
);

INVx3_ASAP7_75t_L g8030 ( 
.A(n_7591),
.Y(n_8030)
);

INVx1_ASAP7_75t_L g8031 ( 
.A(n_7561),
.Y(n_8031)
);

INVx1_ASAP7_75t_L g8032 ( 
.A(n_7562),
.Y(n_8032)
);

INVx2_ASAP7_75t_L g8033 ( 
.A(n_7595),
.Y(n_8033)
);

INVx2_ASAP7_75t_L g8034 ( 
.A(n_7138),
.Y(n_8034)
);

INVx1_ASAP7_75t_L g8035 ( 
.A(n_7568),
.Y(n_8035)
);

OR2x6_ASAP7_75t_L g8036 ( 
.A(n_7468),
.B(n_4402),
.Y(n_8036)
);

INVx1_ASAP7_75t_L g8037 ( 
.A(n_7573),
.Y(n_8037)
);

NAND2xp5_ASAP7_75t_L g8038 ( 
.A(n_7530),
.B(n_4616),
.Y(n_8038)
);

BUFx3_ASAP7_75t_L g8039 ( 
.A(n_7222),
.Y(n_8039)
);

BUFx6f_ASAP7_75t_L g8040 ( 
.A(n_7223),
.Y(n_8040)
);

CKINVDCx5p33_ASAP7_75t_R g8041 ( 
.A(n_7118),
.Y(n_8041)
);

AO21x2_ASAP7_75t_L g8042 ( 
.A1(n_7148),
.A2(n_4416),
.B(n_4412),
.Y(n_8042)
);

INVx2_ASAP7_75t_SL g8043 ( 
.A(n_7591),
.Y(n_8043)
);

AND2x2_ASAP7_75t_L g8044 ( 
.A(n_7418),
.B(n_4618),
.Y(n_8044)
);

INVx2_ASAP7_75t_L g8045 ( 
.A(n_7575),
.Y(n_8045)
);

BUFx2_ASAP7_75t_L g8046 ( 
.A(n_7396),
.Y(n_8046)
);

AO21x2_ASAP7_75t_L g8047 ( 
.A1(n_7259),
.A2(n_4420),
.B(n_4418),
.Y(n_8047)
);

INVx1_ASAP7_75t_L g8048 ( 
.A(n_7572),
.Y(n_8048)
);

BUFx6f_ASAP7_75t_SL g8049 ( 
.A(n_7517),
.Y(n_8049)
);

NAND2xp5_ASAP7_75t_SL g8050 ( 
.A(n_7421),
.B(n_7457),
.Y(n_8050)
);

AND2x6_ASAP7_75t_L g8051 ( 
.A(n_7600),
.B(n_4421),
.Y(n_8051)
);

AOI21x1_ASAP7_75t_L g8052 ( 
.A1(n_7532),
.A2(n_4434),
.B(n_4423),
.Y(n_8052)
);

NAND2xp5_ASAP7_75t_SL g8053 ( 
.A(n_7473),
.B(n_4622),
.Y(n_8053)
);

AND2x4_ASAP7_75t_L g8054 ( 
.A(n_7103),
.B(n_4435),
.Y(n_8054)
);

INVx2_ASAP7_75t_L g8055 ( 
.A(n_7371),
.Y(n_8055)
);

OAI22xp33_ASAP7_75t_L g8056 ( 
.A1(n_7621),
.A2(n_4627),
.B1(n_4628),
.B2(n_4624),
.Y(n_8056)
);

NAND2xp33_ASAP7_75t_SL g8057 ( 
.A(n_7257),
.B(n_4630),
.Y(n_8057)
);

NAND2xp5_ASAP7_75t_SL g8058 ( 
.A(n_7273),
.B(n_4634),
.Y(n_8058)
);

INVx3_ASAP7_75t_L g8059 ( 
.A(n_7223),
.Y(n_8059)
);

INVx2_ASAP7_75t_L g8060 ( 
.A(n_7579),
.Y(n_8060)
);

INVx2_ASAP7_75t_L g8061 ( 
.A(n_7321),
.Y(n_8061)
);

INVx3_ASAP7_75t_L g8062 ( 
.A(n_7228),
.Y(n_8062)
);

NAND2xp5_ASAP7_75t_L g8063 ( 
.A(n_7260),
.B(n_4635),
.Y(n_8063)
);

NAND2xp5_ASAP7_75t_SL g8064 ( 
.A(n_7276),
.B(n_4637),
.Y(n_8064)
);

NAND2xp5_ASAP7_75t_SL g8065 ( 
.A(n_7284),
.B(n_4639),
.Y(n_8065)
);

AND2x2_ASAP7_75t_L g8066 ( 
.A(n_7563),
.B(n_4642),
.Y(n_8066)
);

INVxp33_ASAP7_75t_L g8067 ( 
.A(n_7453),
.Y(n_8067)
);

NAND2xp5_ASAP7_75t_L g8068 ( 
.A(n_7465),
.B(n_4644),
.Y(n_8068)
);

NAND2xp5_ASAP7_75t_SL g8069 ( 
.A(n_7285),
.B(n_4645),
.Y(n_8069)
);

NAND2xp5_ASAP7_75t_SL g8070 ( 
.A(n_7286),
.B(n_4646),
.Y(n_8070)
);

BUFx3_ASAP7_75t_L g8071 ( 
.A(n_7228),
.Y(n_8071)
);

NAND2xp5_ASAP7_75t_L g8072 ( 
.A(n_7545),
.B(n_4647),
.Y(n_8072)
);

INVx2_ASAP7_75t_L g8073 ( 
.A(n_7084),
.Y(n_8073)
);

INVx8_ASAP7_75t_L g8074 ( 
.A(n_7290),
.Y(n_8074)
);

INVxp33_ASAP7_75t_L g8075 ( 
.A(n_7497),
.Y(n_8075)
);

NAND2xp5_ASAP7_75t_SL g8076 ( 
.A(n_7298),
.B(n_4648),
.Y(n_8076)
);

NAND2xp33_ASAP7_75t_L g8077 ( 
.A(n_7304),
.B(n_4649),
.Y(n_8077)
);

INVx2_ASAP7_75t_L g8078 ( 
.A(n_7277),
.Y(n_8078)
);

INVx1_ASAP7_75t_L g8079 ( 
.A(n_7592),
.Y(n_8079)
);

NAND2xp33_ASAP7_75t_L g8080 ( 
.A(n_7305),
.B(n_7307),
.Y(n_8080)
);

INVx2_ASAP7_75t_L g8081 ( 
.A(n_7593),
.Y(n_8081)
);

NAND2xp5_ASAP7_75t_L g8082 ( 
.A(n_7549),
.B(n_4653),
.Y(n_8082)
);

INVx2_ASAP7_75t_L g8083 ( 
.A(n_7594),
.Y(n_8083)
);

BUFx4f_ASAP7_75t_L g8084 ( 
.A(n_7241),
.Y(n_8084)
);

NAND3xp33_ASAP7_75t_L g8085 ( 
.A(n_7555),
.B(n_4656),
.C(n_4655),
.Y(n_8085)
);

INVx2_ASAP7_75t_L g8086 ( 
.A(n_7599),
.Y(n_8086)
);

NOR2xp33_ASAP7_75t_L g8087 ( 
.A(n_7597),
.B(n_4658),
.Y(n_8087)
);

INVx1_ASAP7_75t_L g8088 ( 
.A(n_7484),
.Y(n_8088)
);

INVx1_ASAP7_75t_L g8089 ( 
.A(n_7485),
.Y(n_8089)
);

OR2x2_ASAP7_75t_L g8090 ( 
.A(n_7347),
.B(n_4659),
.Y(n_8090)
);

INVxp67_ASAP7_75t_SL g8091 ( 
.A(n_7241),
.Y(n_8091)
);

BUFx6f_ASAP7_75t_L g8092 ( 
.A(n_7139),
.Y(n_8092)
);

INVx2_ASAP7_75t_L g8093 ( 
.A(n_7581),
.Y(n_8093)
);

INVx3_ASAP7_75t_L g8094 ( 
.A(n_7527),
.Y(n_8094)
);

NAND2xp5_ASAP7_75t_L g8095 ( 
.A(n_7553),
.B(n_4660),
.Y(n_8095)
);

INVx2_ASAP7_75t_L g8096 ( 
.A(n_7492),
.Y(n_8096)
);

BUFx6f_ASAP7_75t_SL g8097 ( 
.A(n_7164),
.Y(n_8097)
);

INVx1_ASAP7_75t_L g8098 ( 
.A(n_7582),
.Y(n_8098)
);

INVx1_ASAP7_75t_L g8099 ( 
.A(n_7293),
.Y(n_8099)
);

INVx1_ASAP7_75t_L g8100 ( 
.A(n_7306),
.Y(n_8100)
);

INVx4_ASAP7_75t_L g8101 ( 
.A(n_7119),
.Y(n_8101)
);

INVx2_ASAP7_75t_L g8102 ( 
.A(n_7356),
.Y(n_8102)
);

BUFx2_ASAP7_75t_L g8103 ( 
.A(n_7413),
.Y(n_8103)
);

NAND2xp5_ASAP7_75t_L g8104 ( 
.A(n_7609),
.B(n_4661),
.Y(n_8104)
);

NOR2xp33_ASAP7_75t_L g8105 ( 
.A(n_7219),
.B(n_4662),
.Y(n_8105)
);

INVx1_ASAP7_75t_L g8106 ( 
.A(n_7411),
.Y(n_8106)
);

INVx2_ASAP7_75t_L g8107 ( 
.A(n_7432),
.Y(n_8107)
);

AOI22xp33_ASAP7_75t_L g8108 ( 
.A1(n_7567),
.A2(n_5348),
.B1(n_5376),
.B2(n_5329),
.Y(n_8108)
);

INVx2_ASAP7_75t_L g8109 ( 
.A(n_7458),
.Y(n_8109)
);

INVx2_ASAP7_75t_L g8110 ( 
.A(n_7472),
.Y(n_8110)
);

INVx1_ASAP7_75t_L g8111 ( 
.A(n_7543),
.Y(n_8111)
);

NAND2xp5_ASAP7_75t_SL g8112 ( 
.A(n_7166),
.B(n_4673),
.Y(n_8112)
);

NOR2xp33_ASAP7_75t_L g8113 ( 
.A(n_7607),
.B(n_7173),
.Y(n_8113)
);

INVx1_ASAP7_75t_L g8114 ( 
.A(n_7565),
.Y(n_8114)
);

NOR2x1_ASAP7_75t_L g8115 ( 
.A(n_7576),
.B(n_7615),
.Y(n_8115)
);

INVx2_ASAP7_75t_L g8116 ( 
.A(n_7570),
.Y(n_8116)
);

INVx2_ASAP7_75t_L g8117 ( 
.A(n_7186),
.Y(n_8117)
);

AND3x2_ASAP7_75t_L g8118 ( 
.A(n_7536),
.B(n_4438),
.C(n_4436),
.Y(n_8118)
);

INVx2_ASAP7_75t_SL g8119 ( 
.A(n_7476),
.Y(n_8119)
);

NAND2xp5_ASAP7_75t_L g8120 ( 
.A(n_7590),
.B(n_4679),
.Y(n_8120)
);

INVx1_ASAP7_75t_L g8121 ( 
.A(n_7267),
.Y(n_8121)
);

INVx3_ASAP7_75t_L g8122 ( 
.A(n_7115),
.Y(n_8122)
);

INVx4_ASAP7_75t_L g8123 ( 
.A(n_7120),
.Y(n_8123)
);

INVx2_ASAP7_75t_L g8124 ( 
.A(n_7127),
.Y(n_8124)
);

INVx2_ASAP7_75t_L g8125 ( 
.A(n_7143),
.Y(n_8125)
);

INVx1_ASAP7_75t_L g8126 ( 
.A(n_7393),
.Y(n_8126)
);

CKINVDCx5p33_ASAP7_75t_R g8127 ( 
.A(n_7132),
.Y(n_8127)
);

INVx1_ASAP7_75t_L g8128 ( 
.A(n_7598),
.Y(n_8128)
);

AND3x2_ASAP7_75t_L g8129 ( 
.A(n_7550),
.B(n_7564),
.C(n_4450),
.Y(n_8129)
);

INVx2_ASAP7_75t_L g8130 ( 
.A(n_7163),
.Y(n_8130)
);

INVx2_ASAP7_75t_L g8131 ( 
.A(n_7541),
.Y(n_8131)
);

INVx2_ASAP7_75t_L g8132 ( 
.A(n_7596),
.Y(n_8132)
);

INVx3_ASAP7_75t_L g8133 ( 
.A(n_7311),
.Y(n_8133)
);

INVx3_ASAP7_75t_L g8134 ( 
.A(n_7320),
.Y(n_8134)
);

CKINVDCx5p33_ASAP7_75t_R g8135 ( 
.A(n_7141),
.Y(n_8135)
);

INVx1_ASAP7_75t_L g8136 ( 
.A(n_7429),
.Y(n_8136)
);

INVx1_ASAP7_75t_L g8137 ( 
.A(n_7602),
.Y(n_8137)
);

INVx1_ASAP7_75t_L g8138 ( 
.A(n_7455),
.Y(n_8138)
);

OAI22xp5_ASAP7_75t_L g8139 ( 
.A1(n_7509),
.A2(n_4681),
.B1(n_4686),
.B2(n_4680),
.Y(n_8139)
);

NAND2xp5_ASAP7_75t_L g8140 ( 
.A(n_7226),
.B(n_4691),
.Y(n_8140)
);

OAI22xp33_ASAP7_75t_L g8141 ( 
.A1(n_7142),
.A2(n_4694),
.B1(n_4695),
.B2(n_4693),
.Y(n_8141)
);

INVx2_ASAP7_75t_L g8142 ( 
.A(n_7327),
.Y(n_8142)
);

INVx2_ASAP7_75t_L g8143 ( 
.A(n_7329),
.Y(n_8143)
);

AOI21x1_ASAP7_75t_L g8144 ( 
.A1(n_7427),
.A2(n_4452),
.B(n_4444),
.Y(n_8144)
);

NAND2xp5_ASAP7_75t_L g8145 ( 
.A(n_7145),
.B(n_4701),
.Y(n_8145)
);

BUFx3_ASAP7_75t_L g8146 ( 
.A(n_7263),
.Y(n_8146)
);

AOI22xp33_ASAP7_75t_L g8147 ( 
.A1(n_7326),
.A2(n_5403),
.B1(n_5452),
.B2(n_5394),
.Y(n_8147)
);

CKINVDCx5p33_ASAP7_75t_R g8148 ( 
.A(n_7146),
.Y(n_8148)
);

INVx1_ASAP7_75t_L g8149 ( 
.A(n_7348),
.Y(n_8149)
);

BUFx6f_ASAP7_75t_L g8150 ( 
.A(n_7155),
.Y(n_8150)
);

NAND2xp5_ASAP7_75t_SL g8151 ( 
.A(n_7157),
.B(n_4707),
.Y(n_8151)
);

INVx3_ASAP7_75t_L g8152 ( 
.A(n_7359),
.Y(n_8152)
);

INVx2_ASAP7_75t_L g8153 ( 
.A(n_7363),
.Y(n_8153)
);

INVx2_ASAP7_75t_L g8154 ( 
.A(n_7588),
.Y(n_8154)
);

OAI22xp5_ASAP7_75t_L g8155 ( 
.A1(n_7158),
.A2(n_4711),
.B1(n_4713),
.B2(n_4709),
.Y(n_8155)
);

NAND2xp33_ASAP7_75t_L g8156 ( 
.A(n_7512),
.B(n_4716),
.Y(n_8156)
);

INVx2_ASAP7_75t_L g8157 ( 
.A(n_7279),
.Y(n_8157)
);

INVx1_ASAP7_75t_L g8158 ( 
.A(n_7460),
.Y(n_8158)
);

NAND2xp5_ASAP7_75t_SL g8159 ( 
.A(n_7124),
.B(n_4718),
.Y(n_8159)
);

BUFx3_ASAP7_75t_L g8160 ( 
.A(n_7283),
.Y(n_8160)
);

INVx2_ASAP7_75t_SL g8161 ( 
.A(n_7121),
.Y(n_8161)
);

NAND2xp5_ASAP7_75t_SL g8162 ( 
.A(n_7149),
.B(n_4719),
.Y(n_8162)
);

BUFx6f_ASAP7_75t_L g8163 ( 
.A(n_7391),
.Y(n_8163)
);

NAND2xp5_ASAP7_75t_SL g8164 ( 
.A(n_7528),
.B(n_4720),
.Y(n_8164)
);

INVx2_ASAP7_75t_L g8165 ( 
.A(n_7295),
.Y(n_8165)
);

NAND3xp33_ASAP7_75t_L g8166 ( 
.A(n_7214),
.B(n_4722),
.C(n_4721),
.Y(n_8166)
);

INVx8_ASAP7_75t_L g8167 ( 
.A(n_7439),
.Y(n_8167)
);

BUFx3_ASAP7_75t_L g8168 ( 
.A(n_7303),
.Y(n_8168)
);

INVx2_ASAP7_75t_L g8169 ( 
.A(n_7309),
.Y(n_8169)
);

INVx2_ASAP7_75t_L g8170 ( 
.A(n_7322),
.Y(n_8170)
);

INVx2_ASAP7_75t_L g8171 ( 
.A(n_7353),
.Y(n_8171)
);

NAND2xp5_ASAP7_75t_SL g8172 ( 
.A(n_7601),
.B(n_4725),
.Y(n_8172)
);

INVx1_ASAP7_75t_L g8173 ( 
.A(n_7417),
.Y(n_8173)
);

NOR2xp33_ASAP7_75t_L g8174 ( 
.A(n_7200),
.B(n_4727),
.Y(n_8174)
);

BUFx10_ASAP7_75t_L g8175 ( 
.A(n_7178),
.Y(n_8175)
);

NAND2xp5_ASAP7_75t_SL g8176 ( 
.A(n_7179),
.B(n_4728),
.Y(n_8176)
);

INVx2_ASAP7_75t_L g8177 ( 
.A(n_7496),
.Y(n_8177)
);

INVx2_ASAP7_75t_L g8178 ( 
.A(n_7445),
.Y(n_8178)
);

NAND2xp5_ASAP7_75t_SL g8179 ( 
.A(n_7182),
.B(n_4731),
.Y(n_8179)
);

INVx2_ASAP7_75t_L g8180 ( 
.A(n_7463),
.Y(n_8180)
);

INVx1_ASAP7_75t_L g8181 ( 
.A(n_7544),
.Y(n_8181)
);

INVx2_ASAP7_75t_L g8182 ( 
.A(n_7749),
.Y(n_8182)
);

INVx1_ASAP7_75t_L g8183 ( 
.A(n_7629),
.Y(n_8183)
);

AND2x2_ASAP7_75t_SL g8184 ( 
.A(n_8080),
.B(n_7625),
.Y(n_8184)
);

CKINVDCx5p33_ASAP7_75t_R g8185 ( 
.A(n_7778),
.Y(n_8185)
);

AND2x2_ASAP7_75t_L g8186 ( 
.A(n_7696),
.B(n_7212),
.Y(n_8186)
);

NAND2xp5_ASAP7_75t_L g8187 ( 
.A(n_7910),
.B(n_4733),
.Y(n_8187)
);

CKINVDCx16_ASAP7_75t_R g8188 ( 
.A(n_8025),
.Y(n_8188)
);

INVx3_ASAP7_75t_L g8189 ( 
.A(n_7630),
.Y(n_8189)
);

AOI22xp5_ASAP7_75t_L g8190 ( 
.A1(n_7946),
.A2(n_7147),
.B1(n_7137),
.B2(n_7218),
.Y(n_8190)
);

INVx1_ASAP7_75t_L g8191 ( 
.A(n_7631),
.Y(n_8191)
);

INVx2_ASAP7_75t_L g8192 ( 
.A(n_7752),
.Y(n_8192)
);

INVx2_ASAP7_75t_L g8193 ( 
.A(n_7753),
.Y(n_8193)
);

BUFx3_ASAP7_75t_L g8194 ( 
.A(n_7630),
.Y(n_8194)
);

BUFx6f_ASAP7_75t_L g8195 ( 
.A(n_7716),
.Y(n_8195)
);

INVx1_ASAP7_75t_L g8196 ( 
.A(n_7636),
.Y(n_8196)
);

INVx2_ASAP7_75t_SL g8197 ( 
.A(n_7716),
.Y(n_8197)
);

BUFx4f_ASAP7_75t_L g8198 ( 
.A(n_7632),
.Y(n_8198)
);

INVx2_ASAP7_75t_L g8199 ( 
.A(n_7755),
.Y(n_8199)
);

INVx2_ASAP7_75t_L g8200 ( 
.A(n_7756),
.Y(n_8200)
);

NOR2xp33_ASAP7_75t_L g8201 ( 
.A(n_7952),
.B(n_7067),
.Y(n_8201)
);

CKINVDCx20_ASAP7_75t_R g8202 ( 
.A(n_7686),
.Y(n_8202)
);

INVx3_ASAP7_75t_L g8203 ( 
.A(n_7734),
.Y(n_8203)
);

NOR2xp33_ASAP7_75t_L g8204 ( 
.A(n_7837),
.B(n_7688),
.Y(n_8204)
);

INVx2_ASAP7_75t_SL g8205 ( 
.A(n_7734),
.Y(n_8205)
);

BUFx6f_ASAP7_75t_L g8206 ( 
.A(n_7764),
.Y(n_8206)
);

INVx2_ASAP7_75t_SL g8207 ( 
.A(n_7764),
.Y(n_8207)
);

INVx5_ASAP7_75t_L g8208 ( 
.A(n_7834),
.Y(n_8208)
);

NAND2xp5_ASAP7_75t_SL g8209 ( 
.A(n_7986),
.B(n_7189),
.Y(n_8209)
);

INVx4_ASAP7_75t_SL g8210 ( 
.A(n_7909),
.Y(n_8210)
);

NAND2xp5_ASAP7_75t_L g8211 ( 
.A(n_7659),
.B(n_4739),
.Y(n_8211)
);

INVx1_ASAP7_75t_L g8212 ( 
.A(n_7637),
.Y(n_8212)
);

NAND2xp5_ASAP7_75t_SL g8213 ( 
.A(n_8098),
.B(n_7193),
.Y(n_8213)
);

AND2x6_ASAP7_75t_L g8214 ( 
.A(n_8150),
.B(n_4457),
.Y(n_8214)
);

INVx2_ASAP7_75t_L g8215 ( 
.A(n_7758),
.Y(n_8215)
);

OAI22xp5_ASAP7_75t_L g8216 ( 
.A1(n_7634),
.A2(n_7258),
.B1(n_7251),
.B2(n_7201),
.Y(n_8216)
);

INVx2_ASAP7_75t_L g8217 ( 
.A(n_7762),
.Y(n_8217)
);

BUFx3_ASAP7_75t_L g8218 ( 
.A(n_7834),
.Y(n_8218)
);

BUFx6f_ASAP7_75t_L g8219 ( 
.A(n_7766),
.Y(n_8219)
);

OAI22xp33_ASAP7_75t_L g8220 ( 
.A1(n_7645),
.A2(n_7674),
.B1(n_7635),
.B2(n_7798),
.Y(n_8220)
);

NOR2xp33_ASAP7_75t_L g8221 ( 
.A(n_7658),
.B(n_7068),
.Y(n_8221)
);

INVx1_ASAP7_75t_L g8222 ( 
.A(n_7639),
.Y(n_8222)
);

NAND2xp5_ASAP7_75t_SL g8223 ( 
.A(n_7757),
.B(n_7197),
.Y(n_8223)
);

OR2x6_ASAP7_75t_L g8224 ( 
.A(n_7917),
.B(n_7202),
.Y(n_8224)
);

NAND2xp5_ASAP7_75t_SL g8225 ( 
.A(n_8005),
.B(n_7071),
.Y(n_8225)
);

BUFx2_ASAP7_75t_L g8226 ( 
.A(n_7673),
.Y(n_8226)
);

INVx1_ASAP7_75t_L g8227 ( 
.A(n_7640),
.Y(n_8227)
);

INVx1_ASAP7_75t_L g8228 ( 
.A(n_7648),
.Y(n_8228)
);

AND2x2_ASAP7_75t_L g8229 ( 
.A(n_7663),
.B(n_7679),
.Y(n_8229)
);

INVx1_ASAP7_75t_L g8230 ( 
.A(n_7653),
.Y(n_8230)
);

NAND2xp5_ASAP7_75t_L g8231 ( 
.A(n_7967),
.B(n_4755),
.Y(n_8231)
);

NAND3x1_ASAP7_75t_L g8232 ( 
.A(n_7706),
.B(n_7649),
.C(n_8113),
.Y(n_8232)
);

BUFx3_ASAP7_75t_L g8233 ( 
.A(n_7917),
.Y(n_8233)
);

INVx1_ASAP7_75t_L g8234 ( 
.A(n_7657),
.Y(n_8234)
);

AND2x4_ASAP7_75t_L g8235 ( 
.A(n_7668),
.B(n_7150),
.Y(n_8235)
);

NOR2xp33_ASAP7_75t_L g8236 ( 
.A(n_7731),
.B(n_7161),
.Y(n_8236)
);

AND2x2_ASAP7_75t_L g8237 ( 
.A(n_8044),
.B(n_7367),
.Y(n_8237)
);

CKINVDCx20_ASAP7_75t_R g8238 ( 
.A(n_7796),
.Y(n_8238)
);

AND2x4_ASAP7_75t_L g8239 ( 
.A(n_7668),
.B(n_7374),
.Y(n_8239)
);

INVx1_ASAP7_75t_L g8240 ( 
.A(n_7664),
.Y(n_8240)
);

OAI22xp5_ASAP7_75t_L g8241 ( 
.A1(n_8132),
.A2(n_7915),
.B1(n_7919),
.B2(n_7916),
.Y(n_8241)
);

INVx4_ASAP7_75t_SL g8242 ( 
.A(n_8049),
.Y(n_8242)
);

NAND2xp5_ASAP7_75t_L g8243 ( 
.A(n_7973),
.B(n_4756),
.Y(n_8243)
);

NOR2xp33_ASAP7_75t_L g8244 ( 
.A(n_7693),
.B(n_7610),
.Y(n_8244)
);

INVx1_ASAP7_75t_L g8245 ( 
.A(n_7666),
.Y(n_8245)
);

INVx3_ASAP7_75t_L g8246 ( 
.A(n_8013),
.Y(n_8246)
);

INVxp33_ASAP7_75t_L g8247 ( 
.A(n_7709),
.Y(n_8247)
);

INVx2_ASAP7_75t_L g8248 ( 
.A(n_7765),
.Y(n_8248)
);

BUFx4_ASAP7_75t_L g8249 ( 
.A(n_8173),
.Y(n_8249)
);

AND2x4_ASAP7_75t_L g8250 ( 
.A(n_7669),
.B(n_7559),
.Y(n_8250)
);

INVx1_ASAP7_75t_SL g8251 ( 
.A(n_7744),
.Y(n_8251)
);

BUFx10_ASAP7_75t_L g8252 ( 
.A(n_8097),
.Y(n_8252)
);

CKINVDCx20_ASAP7_75t_R g8253 ( 
.A(n_7822),
.Y(n_8253)
);

NAND2xp5_ASAP7_75t_L g8254 ( 
.A(n_7974),
.B(n_4758),
.Y(n_8254)
);

BUFx6f_ASAP7_75t_L g8255 ( 
.A(n_7766),
.Y(n_8255)
);

AND2x6_ASAP7_75t_L g8256 ( 
.A(n_8150),
.B(n_4458),
.Y(n_8256)
);

BUFx3_ASAP7_75t_L g8257 ( 
.A(n_8013),
.Y(n_8257)
);

INVx1_ASAP7_75t_L g8258 ( 
.A(n_7671),
.Y(n_8258)
);

INVx1_ASAP7_75t_L g8259 ( 
.A(n_7672),
.Y(n_8259)
);

BUFx6f_ASAP7_75t_L g8260 ( 
.A(n_7780),
.Y(n_8260)
);

INVx1_ASAP7_75t_SL g8261 ( 
.A(n_7665),
.Y(n_8261)
);

AND2x2_ASAP7_75t_SL g8262 ( 
.A(n_7876),
.B(n_8101),
.Y(n_8262)
);

INVx1_ASAP7_75t_L g8263 ( 
.A(n_7677),
.Y(n_8263)
);

INVx1_ASAP7_75t_L g8264 ( 
.A(n_7680),
.Y(n_8264)
);

NAND2xp5_ASAP7_75t_SL g8265 ( 
.A(n_7633),
.B(n_7626),
.Y(n_8265)
);

CKINVDCx5p33_ASAP7_75t_R g8266 ( 
.A(n_8041),
.Y(n_8266)
);

INVx2_ASAP7_75t_L g8267 ( 
.A(n_7769),
.Y(n_8267)
);

AOI22xp5_ASAP7_75t_L g8268 ( 
.A1(n_8087),
.A2(n_4760),
.B1(n_4761),
.B2(n_4759),
.Y(n_8268)
);

INVx3_ASAP7_75t_L g8269 ( 
.A(n_8074),
.Y(n_8269)
);

CKINVDCx5p33_ASAP7_75t_R g8270 ( 
.A(n_8127),
.Y(n_8270)
);

NAND2xp5_ASAP7_75t_L g8271 ( 
.A(n_7982),
.B(n_4764),
.Y(n_8271)
);

AND2x4_ASAP7_75t_L g8272 ( 
.A(n_7700),
.B(n_4459),
.Y(n_8272)
);

INVx1_ASAP7_75t_L g8273 ( 
.A(n_7685),
.Y(n_8273)
);

NAND2xp5_ASAP7_75t_SL g8274 ( 
.A(n_7678),
.B(n_4768),
.Y(n_8274)
);

AND2x4_ASAP7_75t_L g8275 ( 
.A(n_7722),
.B(n_4460),
.Y(n_8275)
);

OR2x2_ASAP7_75t_L g8276 ( 
.A(n_7937),
.B(n_4769),
.Y(n_8276)
);

NAND2xp5_ASAP7_75t_SL g8277 ( 
.A(n_7727),
.B(n_4770),
.Y(n_8277)
);

INVx1_ASAP7_75t_L g8278 ( 
.A(n_7690),
.Y(n_8278)
);

INVx8_ASAP7_75t_L g8279 ( 
.A(n_8074),
.Y(n_8279)
);

INVx2_ASAP7_75t_L g8280 ( 
.A(n_7770),
.Y(n_8280)
);

INVx2_ASAP7_75t_L g8281 ( 
.A(n_7771),
.Y(n_8281)
);

INVx2_ASAP7_75t_SL g8282 ( 
.A(n_7969),
.Y(n_8282)
);

AND2x2_ASAP7_75t_SL g8283 ( 
.A(n_8123),
.B(n_7927),
.Y(n_8283)
);

AOI22xp33_ASAP7_75t_L g8284 ( 
.A1(n_8056),
.A2(n_5469),
.B1(n_5490),
.B2(n_5458),
.Y(n_8284)
);

INVx2_ASAP7_75t_L g8285 ( 
.A(n_7774),
.Y(n_8285)
);

INVx1_ASAP7_75t_L g8286 ( 
.A(n_7697),
.Y(n_8286)
);

NAND2xp5_ASAP7_75t_L g8287 ( 
.A(n_7988),
.B(n_4772),
.Y(n_8287)
);

NAND2xp5_ASAP7_75t_L g8288 ( 
.A(n_7989),
.B(n_4774),
.Y(n_8288)
);

INVx4_ASAP7_75t_L g8289 ( 
.A(n_7722),
.Y(n_8289)
);

CKINVDCx5p33_ASAP7_75t_R g8290 ( 
.A(n_8135),
.Y(n_8290)
);

INVx1_ASAP7_75t_L g8291 ( 
.A(n_7713),
.Y(n_8291)
);

INVx2_ASAP7_75t_L g8292 ( 
.A(n_7782),
.Y(n_8292)
);

NAND2xp5_ASAP7_75t_SL g8293 ( 
.A(n_7747),
.B(n_4779),
.Y(n_8293)
);

INVx4_ASAP7_75t_L g8294 ( 
.A(n_7780),
.Y(n_8294)
);

BUFx6f_ASAP7_75t_L g8295 ( 
.A(n_7844),
.Y(n_8295)
);

NAND2xp5_ASAP7_75t_SL g8296 ( 
.A(n_7751),
.B(n_4784),
.Y(n_8296)
);

INVx1_ASAP7_75t_L g8297 ( 
.A(n_7726),
.Y(n_8297)
);

BUFx2_ASAP7_75t_L g8298 ( 
.A(n_7886),
.Y(n_8298)
);

NOR2xp33_ASAP7_75t_L g8299 ( 
.A(n_7725),
.B(n_4794),
.Y(n_8299)
);

AND2x2_ASAP7_75t_L g8300 ( 
.A(n_8066),
.B(n_4800),
.Y(n_8300)
);

AND2x2_ASAP7_75t_L g8301 ( 
.A(n_7691),
.B(n_4801),
.Y(n_8301)
);

INVx8_ASAP7_75t_L g8302 ( 
.A(n_7800),
.Y(n_8302)
);

INVxp67_ASAP7_75t_L g8303 ( 
.A(n_7775),
.Y(n_8303)
);

NOR2xp33_ASAP7_75t_L g8304 ( 
.A(n_7654),
.B(n_4803),
.Y(n_8304)
);

OR2x6_ASAP7_75t_L g8305 ( 
.A(n_7800),
.B(n_4464),
.Y(n_8305)
);

INVx2_ASAP7_75t_L g8306 ( 
.A(n_7783),
.Y(n_8306)
);

INVx1_ASAP7_75t_L g8307 ( 
.A(n_7732),
.Y(n_8307)
);

OR2x6_ASAP7_75t_L g8308 ( 
.A(n_7705),
.B(n_4470),
.Y(n_8308)
);

INVx1_ASAP7_75t_L g8309 ( 
.A(n_7750),
.Y(n_8309)
);

INVx4_ASAP7_75t_L g8310 ( 
.A(n_7844),
.Y(n_8310)
);

OR2x2_ASAP7_75t_L g8311 ( 
.A(n_8157),
.B(n_4804),
.Y(n_8311)
);

AND2x6_ASAP7_75t_L g8312 ( 
.A(n_8115),
.B(n_4472),
.Y(n_8312)
);

NAND2xp5_ASAP7_75t_SL g8313 ( 
.A(n_7893),
.B(n_4807),
.Y(n_8313)
);

INVx3_ASAP7_75t_L g8314 ( 
.A(n_7851),
.Y(n_8314)
);

NOR2xp33_ASAP7_75t_L g8315 ( 
.A(n_7655),
.B(n_4810),
.Y(n_8315)
);

BUFx6f_ASAP7_75t_L g8316 ( 
.A(n_7851),
.Y(n_8316)
);

NOR2x1p5_ASAP7_75t_L g8317 ( 
.A(n_8019),
.B(n_4811),
.Y(n_8317)
);

INVx1_ASAP7_75t_L g8318 ( 
.A(n_7772),
.Y(n_8318)
);

NAND2xp5_ASAP7_75t_L g8319 ( 
.A(n_7990),
.B(n_4816),
.Y(n_8319)
);

CKINVDCx5p33_ASAP7_75t_R g8320 ( 
.A(n_8148),
.Y(n_8320)
);

NOR2xp33_ASAP7_75t_L g8321 ( 
.A(n_7656),
.B(n_4817),
.Y(n_8321)
);

INVx2_ASAP7_75t_L g8322 ( 
.A(n_7787),
.Y(n_8322)
);

NAND2xp5_ASAP7_75t_L g8323 ( 
.A(n_7683),
.B(n_4820),
.Y(n_8323)
);

NAND2xp5_ASAP7_75t_L g8324 ( 
.A(n_7687),
.B(n_4823),
.Y(n_8324)
);

NAND2xp5_ASAP7_75t_SL g8325 ( 
.A(n_7976),
.B(n_4824),
.Y(n_8325)
);

OR2x2_ASAP7_75t_L g8326 ( 
.A(n_8165),
.B(n_4825),
.Y(n_8326)
);

INVx4_ASAP7_75t_L g8327 ( 
.A(n_7872),
.Y(n_8327)
);

AND2x2_ASAP7_75t_L g8328 ( 
.A(n_7859),
.B(n_4826),
.Y(n_8328)
);

INVx2_ASAP7_75t_L g8329 ( 
.A(n_7791),
.Y(n_8329)
);

OAI22xp33_ASAP7_75t_L g8330 ( 
.A1(n_8104),
.A2(n_4830),
.B1(n_4832),
.B2(n_4827),
.Y(n_8330)
);

INVxp67_ASAP7_75t_L g8331 ( 
.A(n_8154),
.Y(n_8331)
);

NOR2x1p5_ASAP7_75t_L g8332 ( 
.A(n_8094),
.B(n_4834),
.Y(n_8332)
);

NAND2xp5_ASAP7_75t_L g8333 ( 
.A(n_7777),
.B(n_4835),
.Y(n_8333)
);

INVx1_ASAP7_75t_L g8334 ( 
.A(n_7779),
.Y(n_8334)
);

NOR2xp33_ASAP7_75t_L g8335 ( 
.A(n_7662),
.B(n_7712),
.Y(n_8335)
);

INVx1_ASAP7_75t_L g8336 ( 
.A(n_7781),
.Y(n_8336)
);

INVx2_ASAP7_75t_L g8337 ( 
.A(n_7792),
.Y(n_8337)
);

INVx2_ASAP7_75t_SL g8338 ( 
.A(n_7975),
.Y(n_8338)
);

INVx1_ASAP7_75t_L g8339 ( 
.A(n_7784),
.Y(n_8339)
);

OAI22xp33_ASAP7_75t_L g8340 ( 
.A1(n_8038),
.A2(n_4844),
.B1(n_4851),
.B2(n_4838),
.Y(n_8340)
);

NOR2xp33_ASAP7_75t_L g8341 ( 
.A(n_7728),
.B(n_4852),
.Y(n_8341)
);

INVx1_ASAP7_75t_L g8342 ( 
.A(n_7785),
.Y(n_8342)
);

HB1xp67_ASAP7_75t_L g8343 ( 
.A(n_7872),
.Y(n_8343)
);

NAND2xp5_ASAP7_75t_L g8344 ( 
.A(n_7790),
.B(n_4855),
.Y(n_8344)
);

INVx1_ASAP7_75t_L g8345 ( 
.A(n_7803),
.Y(n_8345)
);

INVx1_ASAP7_75t_L g8346 ( 
.A(n_7806),
.Y(n_8346)
);

BUFx4f_ASAP7_75t_L g8347 ( 
.A(n_8163),
.Y(n_8347)
);

INVxp33_ASAP7_75t_L g8348 ( 
.A(n_7810),
.Y(n_8348)
);

INVx2_ASAP7_75t_L g8349 ( 
.A(n_7799),
.Y(n_8349)
);

NAND2xp5_ASAP7_75t_SL g8350 ( 
.A(n_7694),
.B(n_4857),
.Y(n_8350)
);

OAI22xp5_ASAP7_75t_SL g8351 ( 
.A1(n_8181),
.A2(n_4859),
.B1(n_4860),
.B2(n_4858),
.Y(n_8351)
);

AOI22xp33_ASAP7_75t_L g8352 ( 
.A1(n_7807),
.A2(n_5501),
.B1(n_5496),
.B2(n_4476),
.Y(n_8352)
);

INVx2_ASAP7_75t_SL g8353 ( 
.A(n_8022),
.Y(n_8353)
);

INVx4_ASAP7_75t_L g8354 ( 
.A(n_7926),
.Y(n_8354)
);

HB1xp67_ASAP7_75t_L g8355 ( 
.A(n_7926),
.Y(n_8355)
);

INVx4_ASAP7_75t_L g8356 ( 
.A(n_8040),
.Y(n_8356)
);

NOR2xp33_ASAP7_75t_L g8357 ( 
.A(n_8029),
.B(n_4861),
.Y(n_8357)
);

NOR2xp33_ASAP7_75t_L g8358 ( 
.A(n_7724),
.B(n_4863),
.Y(n_8358)
);

INVx3_ASAP7_75t_L g8359 ( 
.A(n_8040),
.Y(n_8359)
);

OAI22xp33_ASAP7_75t_L g8360 ( 
.A1(n_7987),
.A2(n_4869),
.B1(n_4870),
.B2(n_4864),
.Y(n_8360)
);

NAND2xp5_ASAP7_75t_L g8361 ( 
.A(n_7815),
.B(n_4872),
.Y(n_8361)
);

INVx3_ASAP7_75t_L g8362 ( 
.A(n_8092),
.Y(n_8362)
);

INVx1_ASAP7_75t_L g8363 ( 
.A(n_7817),
.Y(n_8363)
);

INVxp67_ASAP7_75t_L g8364 ( 
.A(n_8128),
.Y(n_8364)
);

NOR2xp33_ASAP7_75t_L g8365 ( 
.A(n_7869),
.B(n_4875),
.Y(n_8365)
);

INVx2_ASAP7_75t_L g8366 ( 
.A(n_7808),
.Y(n_8366)
);

INVx1_ASAP7_75t_L g8367 ( 
.A(n_7819),
.Y(n_8367)
);

BUFx2_ASAP7_75t_L g8368 ( 
.A(n_7936),
.Y(n_8368)
);

NAND2xp5_ASAP7_75t_SL g8369 ( 
.A(n_7811),
.B(n_4880),
.Y(n_8369)
);

AND2x4_ASAP7_75t_L g8370 ( 
.A(n_7888),
.B(n_4474),
.Y(n_8370)
);

INVx1_ASAP7_75t_L g8371 ( 
.A(n_7820),
.Y(n_8371)
);

OAI221xp5_ASAP7_75t_L g8372 ( 
.A1(n_8147),
.A2(n_4885),
.B1(n_4886),
.B2(n_4884),
.C(n_4882),
.Y(n_8372)
);

BUFx10_ASAP7_75t_L g8373 ( 
.A(n_7903),
.Y(n_8373)
);

AND2x6_ASAP7_75t_L g8374 ( 
.A(n_8138),
.B(n_4477),
.Y(n_8374)
);

NOR2xp33_ASAP7_75t_L g8375 ( 
.A(n_8075),
.B(n_4887),
.Y(n_8375)
);

AOI22xp33_ASAP7_75t_L g8376 ( 
.A1(n_7814),
.A2(n_4491),
.B1(n_4492),
.B2(n_4487),
.Y(n_8376)
);

INVx3_ASAP7_75t_L g8377 ( 
.A(n_8092),
.Y(n_8377)
);

INVx1_ASAP7_75t_SL g8378 ( 
.A(n_7812),
.Y(n_8378)
);

BUFx2_ASAP7_75t_L g8379 ( 
.A(n_8046),
.Y(n_8379)
);

BUFx4f_ASAP7_75t_L g8380 ( 
.A(n_8163),
.Y(n_8380)
);

INVx1_ASAP7_75t_L g8381 ( 
.A(n_7828),
.Y(n_8381)
);

NAND2xp5_ASAP7_75t_L g8382 ( 
.A(n_7823),
.B(n_4889),
.Y(n_8382)
);

NOR2xp33_ASAP7_75t_L g8383 ( 
.A(n_7824),
.B(n_4890),
.Y(n_8383)
);

INVx3_ASAP7_75t_L g8384 ( 
.A(n_7805),
.Y(n_8384)
);

AND2x6_ASAP7_75t_L g8385 ( 
.A(n_8131),
.B(n_4506),
.Y(n_8385)
);

NAND2xp5_ASAP7_75t_SL g8386 ( 
.A(n_7825),
.B(n_4893),
.Y(n_8386)
);

INVx1_ASAP7_75t_L g8387 ( 
.A(n_7826),
.Y(n_8387)
);

INVx1_ASAP7_75t_L g8388 ( 
.A(n_7838),
.Y(n_8388)
);

NAND2xp5_ASAP7_75t_L g8389 ( 
.A(n_7972),
.B(n_4896),
.Y(n_8389)
);

INVx1_ASAP7_75t_L g8390 ( 
.A(n_7840),
.Y(n_8390)
);

AO22x2_ASAP7_75t_L g8391 ( 
.A1(n_7699),
.A2(n_4510),
.B1(n_4513),
.B2(n_4509),
.Y(n_8391)
);

INVx4_ASAP7_75t_SL g8392 ( 
.A(n_8051),
.Y(n_8392)
);

INVx2_ASAP7_75t_L g8393 ( 
.A(n_7628),
.Y(n_8393)
);

INVx1_ASAP7_75t_L g8394 ( 
.A(n_7842),
.Y(n_8394)
);

NOR2xp33_ASAP7_75t_L g8395 ( 
.A(n_8145),
.B(n_4897),
.Y(n_8395)
);

INVx1_ASAP7_75t_L g8396 ( 
.A(n_7843),
.Y(n_8396)
);

INVx2_ASAP7_75t_L g8397 ( 
.A(n_7638),
.Y(n_8397)
);

NAND2xp33_ASAP7_75t_L g8398 ( 
.A(n_7931),
.B(n_4898),
.Y(n_8398)
);

INVx3_ASAP7_75t_L g8399 ( 
.A(n_7942),
.Y(n_8399)
);

INVx1_ASAP7_75t_L g8400 ( 
.A(n_7845),
.Y(n_8400)
);

INVx1_ASAP7_75t_L g8401 ( 
.A(n_7847),
.Y(n_8401)
);

INVx1_ASAP7_75t_L g8402 ( 
.A(n_7848),
.Y(n_8402)
);

AO22x2_ASAP7_75t_L g8403 ( 
.A1(n_8090),
.A2(n_4524),
.B1(n_4528),
.B2(n_4521),
.Y(n_8403)
);

NAND2xp5_ASAP7_75t_L g8404 ( 
.A(n_7809),
.B(n_4899),
.Y(n_8404)
);

OR2x6_ASAP7_75t_L g8405 ( 
.A(n_8167),
.B(n_4529),
.Y(n_8405)
);

INVx1_ASAP7_75t_L g8406 ( 
.A(n_7849),
.Y(n_8406)
);

NAND3xp33_ASAP7_75t_L g8407 ( 
.A(n_7932),
.B(n_4901),
.C(n_4900),
.Y(n_8407)
);

NOR2x1p5_ASAP7_75t_L g8408 ( 
.A(n_8133),
.B(n_4902),
.Y(n_8408)
);

INVx1_ASAP7_75t_SL g8409 ( 
.A(n_8103),
.Y(n_8409)
);

NAND3x1_ASAP7_75t_L g8410 ( 
.A(n_8158),
.B(n_4542),
.C(n_4539),
.Y(n_8410)
);

INVx2_ASAP7_75t_L g8411 ( 
.A(n_7641),
.Y(n_8411)
);

NOR2xp33_ASAP7_75t_L g8412 ( 
.A(n_7940),
.B(n_7646),
.Y(n_8412)
);

INVx1_ASAP7_75t_L g8413 ( 
.A(n_7856),
.Y(n_8413)
);

BUFx10_ASAP7_75t_L g8414 ( 
.A(n_8174),
.Y(n_8414)
);

NAND2xp5_ASAP7_75t_L g8415 ( 
.A(n_7857),
.B(n_4903),
.Y(n_8415)
);

AOI21x1_ASAP7_75t_L g8416 ( 
.A1(n_7944),
.A2(n_4564),
.B(n_4556),
.Y(n_8416)
);

INVx1_ASAP7_75t_L g8417 ( 
.A(n_7860),
.Y(n_8417)
);

AND2x2_ASAP7_75t_L g8418 ( 
.A(n_7786),
.B(n_4905),
.Y(n_8418)
);

AO22x2_ASAP7_75t_L g8419 ( 
.A1(n_7681),
.A2(n_4573),
.B1(n_4574),
.B2(n_4566),
.Y(n_8419)
);

AND2x6_ASAP7_75t_L g8420 ( 
.A(n_8149),
.B(n_4575),
.Y(n_8420)
);

INVx4_ASAP7_75t_L g8421 ( 
.A(n_8084),
.Y(n_8421)
);

INVxp67_ASAP7_75t_SL g8422 ( 
.A(n_7921),
.Y(n_8422)
);

INVxp67_ASAP7_75t_L g8423 ( 
.A(n_7802),
.Y(n_8423)
);

NOR2xp33_ASAP7_75t_L g8424 ( 
.A(n_7827),
.B(n_4912),
.Y(n_8424)
);

INVx3_ASAP7_75t_L g8425 ( 
.A(n_8039),
.Y(n_8425)
);

INVx4_ASAP7_75t_SL g8426 ( 
.A(n_8051),
.Y(n_8426)
);

INVx3_ASAP7_75t_L g8427 ( 
.A(n_8071),
.Y(n_8427)
);

OAI22xp5_ASAP7_75t_L g8428 ( 
.A1(n_7922),
.A2(n_4916),
.B1(n_4918),
.B2(n_4915),
.Y(n_8428)
);

INVx3_ASAP7_75t_L g8429 ( 
.A(n_7853),
.Y(n_8429)
);

INVx2_ASAP7_75t_L g8430 ( 
.A(n_7644),
.Y(n_8430)
);

NAND2xp5_ASAP7_75t_L g8431 ( 
.A(n_7695),
.B(n_4919),
.Y(n_8431)
);

INVx2_ASAP7_75t_L g8432 ( 
.A(n_7647),
.Y(n_8432)
);

INVx1_ASAP7_75t_L g8433 ( 
.A(n_7861),
.Y(n_8433)
);

BUFx3_ASAP7_75t_L g8434 ( 
.A(n_8146),
.Y(n_8434)
);

AND2x6_ASAP7_75t_L g8435 ( 
.A(n_8142),
.B(n_4582),
.Y(n_8435)
);

AND2x2_ASAP7_75t_L g8436 ( 
.A(n_7760),
.B(n_4920),
.Y(n_8436)
);

INVx2_ASAP7_75t_L g8437 ( 
.A(n_7650),
.Y(n_8437)
);

NOR2xp33_ASAP7_75t_L g8438 ( 
.A(n_7729),
.B(n_4921),
.Y(n_8438)
);

INVx2_ASAP7_75t_L g8439 ( 
.A(n_7651),
.Y(n_8439)
);

INVx1_ASAP7_75t_L g8440 ( 
.A(n_7863),
.Y(n_8440)
);

INVx2_ASAP7_75t_L g8441 ( 
.A(n_7660),
.Y(n_8441)
);

NAND2xp5_ASAP7_75t_L g8442 ( 
.A(n_7708),
.B(n_4923),
.Y(n_8442)
);

NAND3xp33_ASAP7_75t_L g8443 ( 
.A(n_7736),
.B(n_4927),
.C(n_4926),
.Y(n_8443)
);

INVx1_ASAP7_75t_SL g8444 ( 
.A(n_8160),
.Y(n_8444)
);

CKINVDCx5p33_ASAP7_75t_R g8445 ( 
.A(n_7652),
.Y(n_8445)
);

INVx2_ASAP7_75t_SL g8446 ( 
.A(n_7997),
.Y(n_8446)
);

INVx1_ASAP7_75t_L g8447 ( 
.A(n_7864),
.Y(n_8447)
);

INVx1_ASAP7_75t_L g8448 ( 
.A(n_7867),
.Y(n_8448)
);

NOR2xp33_ASAP7_75t_L g8449 ( 
.A(n_7761),
.B(n_4930),
.Y(n_8449)
);

NOR2xp33_ASAP7_75t_L g8450 ( 
.A(n_8067),
.B(n_4935),
.Y(n_8450)
);

AND2x4_ASAP7_75t_L g8451 ( 
.A(n_7813),
.B(n_4583),
.Y(n_8451)
);

INVx1_ASAP7_75t_L g8452 ( 
.A(n_7868),
.Y(n_8452)
);

INVx1_ASAP7_75t_L g8453 ( 
.A(n_7880),
.Y(n_8453)
);

AOI22xp5_ASAP7_75t_L g8454 ( 
.A1(n_8050),
.A2(n_4939),
.B1(n_4940),
.B2(n_4938),
.Y(n_8454)
);

INVx2_ASAP7_75t_L g8455 ( 
.A(n_7670),
.Y(n_8455)
);

INVx1_ASAP7_75t_L g8456 ( 
.A(n_7901),
.Y(n_8456)
);

INVx2_ASAP7_75t_L g8457 ( 
.A(n_7675),
.Y(n_8457)
);

INVx1_ASAP7_75t_L g8458 ( 
.A(n_7906),
.Y(n_8458)
);

INVx2_ASAP7_75t_L g8459 ( 
.A(n_7684),
.Y(n_8459)
);

NAND2xp5_ASAP7_75t_L g8460 ( 
.A(n_7718),
.B(n_4944),
.Y(n_8460)
);

INVx2_ASAP7_75t_L g8461 ( 
.A(n_7692),
.Y(n_8461)
);

NAND2xp5_ASAP7_75t_L g8462 ( 
.A(n_7723),
.B(n_7730),
.Y(n_8462)
);

AND2x4_ASAP7_75t_L g8463 ( 
.A(n_7846),
.B(n_4586),
.Y(n_8463)
);

INVx1_ASAP7_75t_SL g8464 ( 
.A(n_8168),
.Y(n_8464)
);

INVx1_ASAP7_75t_L g8465 ( 
.A(n_7907),
.Y(n_8465)
);

AO22x2_ASAP7_75t_L g8466 ( 
.A1(n_8012),
.A2(n_4598),
.B1(n_4599),
.B2(n_4597),
.Y(n_8466)
);

INVx1_ASAP7_75t_L g8467 ( 
.A(n_7908),
.Y(n_8467)
);

INVx1_ASAP7_75t_SL g8468 ( 
.A(n_7971),
.Y(n_8468)
);

NOR2xp33_ASAP7_75t_L g8469 ( 
.A(n_7965),
.B(n_8143),
.Y(n_8469)
);

INVx2_ASAP7_75t_L g8470 ( 
.A(n_7698),
.Y(n_8470)
);

INVx3_ASAP7_75t_L g8471 ( 
.A(n_8059),
.Y(n_8471)
);

INVx1_ASAP7_75t_L g8472 ( 
.A(n_7902),
.Y(n_8472)
);

NAND2xp5_ASAP7_75t_L g8473 ( 
.A(n_7738),
.B(n_4945),
.Y(n_8473)
);

INVx1_ASAP7_75t_L g8474 ( 
.A(n_7905),
.Y(n_8474)
);

AND2x2_ASAP7_75t_L g8475 ( 
.A(n_8153),
.B(n_4946),
.Y(n_8475)
);

NAND2xp33_ASAP7_75t_L g8476 ( 
.A(n_7931),
.B(n_4947),
.Y(n_8476)
);

INVx4_ASAP7_75t_SL g8477 ( 
.A(n_8051),
.Y(n_8477)
);

INVx2_ASAP7_75t_L g8478 ( 
.A(n_7701),
.Y(n_8478)
);

INVx2_ASAP7_75t_L g8479 ( 
.A(n_7702),
.Y(n_8479)
);

INVx5_ASAP7_75t_L g8480 ( 
.A(n_7711),
.Y(n_8480)
);

INVx1_ASAP7_75t_L g8481 ( 
.A(n_7912),
.Y(n_8481)
);

INVx1_ASAP7_75t_SL g8482 ( 
.A(n_7971),
.Y(n_8482)
);

INVx2_ASAP7_75t_L g8483 ( 
.A(n_7703),
.Y(n_8483)
);

INVx2_ASAP7_75t_L g8484 ( 
.A(n_7704),
.Y(n_8484)
);

INVx1_ASAP7_75t_L g8485 ( 
.A(n_7710),
.Y(n_8485)
);

AO21x2_ASAP7_75t_L g8486 ( 
.A1(n_7964),
.A2(n_4619),
.B(n_4606),
.Y(n_8486)
);

AOI22xp33_ASAP7_75t_L g8487 ( 
.A1(n_8026),
.A2(n_4621),
.B1(n_4626),
.B2(n_4620),
.Y(n_8487)
);

NAND3xp33_ASAP7_75t_L g8488 ( 
.A(n_8021),
.B(n_4953),
.C(n_4951),
.Y(n_8488)
);

INVx2_ASAP7_75t_SL g8489 ( 
.A(n_8003),
.Y(n_8489)
);

AND2x2_ASAP7_75t_L g8490 ( 
.A(n_8134),
.B(n_4954),
.Y(n_8490)
);

NOR2xp33_ASAP7_75t_L g8491 ( 
.A(n_7643),
.B(n_4956),
.Y(n_8491)
);

INVx2_ASAP7_75t_L g8492 ( 
.A(n_7714),
.Y(n_8492)
);

INVx6_ASAP7_75t_L g8493 ( 
.A(n_7721),
.Y(n_8493)
);

NAND2xp5_ASAP7_75t_L g8494 ( 
.A(n_7743),
.B(n_4958),
.Y(n_8494)
);

INVx1_ASAP7_75t_L g8495 ( 
.A(n_7715),
.Y(n_8495)
);

INVx2_ASAP7_75t_L g8496 ( 
.A(n_7717),
.Y(n_8496)
);

CKINVDCx5p33_ASAP7_75t_R g8497 ( 
.A(n_8175),
.Y(n_8497)
);

AND2x2_ASAP7_75t_L g8498 ( 
.A(n_8152),
.B(n_4963),
.Y(n_8498)
);

BUFx3_ASAP7_75t_L g8499 ( 
.A(n_8062),
.Y(n_8499)
);

NOR2xp33_ASAP7_75t_L g8500 ( 
.A(n_7870),
.B(n_4964),
.Y(n_8500)
);

INVx1_ASAP7_75t_L g8501 ( 
.A(n_7719),
.Y(n_8501)
);

INVx1_ASAP7_75t_L g8502 ( 
.A(n_7720),
.Y(n_8502)
);

BUFx10_ASAP7_75t_L g8503 ( 
.A(n_8105),
.Y(n_8503)
);

INVx1_ASAP7_75t_L g8504 ( 
.A(n_7733),
.Y(n_8504)
);

NAND2xp5_ASAP7_75t_SL g8505 ( 
.A(n_8120),
.B(n_4965),
.Y(n_8505)
);

INVx6_ASAP7_75t_L g8506 ( 
.A(n_7920),
.Y(n_8506)
);

INVx1_ASAP7_75t_L g8507 ( 
.A(n_7735),
.Y(n_8507)
);

INVx2_ASAP7_75t_L g8508 ( 
.A(n_7739),
.Y(n_8508)
);

INVx1_ASAP7_75t_L g8509 ( 
.A(n_7746),
.Y(n_8509)
);

BUFx3_ASAP7_75t_L g8510 ( 
.A(n_7821),
.Y(n_8510)
);

INVx2_ASAP7_75t_L g8511 ( 
.A(n_7831),
.Y(n_8511)
);

NOR2xp33_ASAP7_75t_L g8512 ( 
.A(n_8169),
.B(n_4968),
.Y(n_8512)
);

BUFx3_ASAP7_75t_L g8513 ( 
.A(n_7661),
.Y(n_8513)
);

AND2x4_ASAP7_75t_L g8514 ( 
.A(n_7897),
.B(n_4629),
.Y(n_8514)
);

INVx2_ASAP7_75t_L g8515 ( 
.A(n_7832),
.Y(n_8515)
);

OR2x6_ASAP7_75t_L g8516 ( 
.A(n_8167),
.B(n_4631),
.Y(n_8516)
);

AND3x4_ASAP7_75t_L g8517 ( 
.A(n_8170),
.B(n_4971),
.C(n_4970),
.Y(n_8517)
);

BUFx2_ASAP7_75t_L g8518 ( 
.A(n_8171),
.Y(n_8518)
);

AND2x4_ASAP7_75t_L g8519 ( 
.A(n_7955),
.B(n_4633),
.Y(n_8519)
);

BUFx3_ASAP7_75t_L g8520 ( 
.A(n_7707),
.Y(n_8520)
);

INVx4_ASAP7_75t_L g8521 ( 
.A(n_7920),
.Y(n_8521)
);

INVx1_ASAP7_75t_L g8522 ( 
.A(n_7833),
.Y(n_8522)
);

INVx1_ASAP7_75t_SL g8523 ( 
.A(n_8048),
.Y(n_8523)
);

INVx3_ASAP7_75t_L g8524 ( 
.A(n_7740),
.Y(n_8524)
);

INVx3_ASAP7_75t_L g8525 ( 
.A(n_7742),
.Y(n_8525)
);

NAND2xp5_ASAP7_75t_L g8526 ( 
.A(n_7745),
.B(n_4973),
.Y(n_8526)
);

AND2x6_ASAP7_75t_L g8527 ( 
.A(n_8136),
.B(n_4636),
.Y(n_8527)
);

INVx2_ASAP7_75t_L g8528 ( 
.A(n_7835),
.Y(n_8528)
);

AO22x2_ASAP7_75t_L g8529 ( 
.A1(n_8155),
.A2(n_8137),
.B1(n_8028),
.B2(n_8031),
.Y(n_8529)
);

INVx2_ASAP7_75t_L g8530 ( 
.A(n_7839),
.Y(n_8530)
);

INVx2_ASAP7_75t_SL g8531 ( 
.A(n_8043),
.Y(n_8531)
);

INVx2_ASAP7_75t_L g8532 ( 
.A(n_7841),
.Y(n_8532)
);

INVx1_ASAP7_75t_L g8533 ( 
.A(n_7850),
.Y(n_8533)
);

INVx4_ASAP7_75t_L g8534 ( 
.A(n_7763),
.Y(n_8534)
);

NOR2xp33_ASAP7_75t_SL g8535 ( 
.A(n_8161),
.B(n_4977),
.Y(n_8535)
);

NAND2xp5_ASAP7_75t_L g8536 ( 
.A(n_7759),
.B(n_4978),
.Y(n_8536)
);

INVx3_ASAP7_75t_L g8537 ( 
.A(n_7776),
.Y(n_8537)
);

INVx3_ASAP7_75t_L g8538 ( 
.A(n_7789),
.Y(n_8538)
);

INVx1_ASAP7_75t_L g8539 ( 
.A(n_7855),
.Y(n_8539)
);

INVx1_ASAP7_75t_L g8540 ( 
.A(n_7858),
.Y(n_8540)
);

BUFx6f_ASAP7_75t_L g8541 ( 
.A(n_7793),
.Y(n_8541)
);

NAND2xp5_ASAP7_75t_L g8542 ( 
.A(n_7768),
.B(n_4980),
.Y(n_8542)
);

AND2x6_ASAP7_75t_L g8543 ( 
.A(n_8088),
.B(n_8089),
.Y(n_8543)
);

INVx1_ASAP7_75t_L g8544 ( 
.A(n_7862),
.Y(n_8544)
);

INVx1_ASAP7_75t_L g8545 ( 
.A(n_7866),
.Y(n_8545)
);

BUFx6f_ASAP7_75t_L g8546 ( 
.A(n_7795),
.Y(n_8546)
);

AND2x4_ASAP7_75t_L g8547 ( 
.A(n_7958),
.B(n_4638),
.Y(n_8547)
);

NAND2xp5_ASAP7_75t_L g8548 ( 
.A(n_7794),
.B(n_4986),
.Y(n_8548)
);

INVx2_ASAP7_75t_L g8549 ( 
.A(n_7871),
.Y(n_8549)
);

INVx2_ASAP7_75t_L g8550 ( 
.A(n_7873),
.Y(n_8550)
);

OR2x2_ASAP7_75t_L g8551 ( 
.A(n_7816),
.B(n_4988),
.Y(n_8551)
);

INVx1_ASAP7_75t_L g8552 ( 
.A(n_7875),
.Y(n_8552)
);

NOR2xp33_ASAP7_75t_L g8553 ( 
.A(n_8053),
.B(n_4991),
.Y(n_8553)
);

BUFx2_ASAP7_75t_L g8554 ( 
.A(n_8177),
.Y(n_8554)
);

BUFx6f_ASAP7_75t_L g8555 ( 
.A(n_7801),
.Y(n_8555)
);

INVx3_ASAP7_75t_L g8556 ( 
.A(n_7836),
.Y(n_8556)
);

INVx1_ASAP7_75t_L g8557 ( 
.A(n_7877),
.Y(n_8557)
);

NAND2xp5_ASAP7_75t_SL g8558 ( 
.A(n_8068),
.B(n_5000),
.Y(n_8558)
);

BUFx2_ASAP7_75t_L g8559 ( 
.A(n_8178),
.Y(n_8559)
);

INVx4_ASAP7_75t_L g8560 ( 
.A(n_7874),
.Y(n_8560)
);

INVx1_ASAP7_75t_L g8561 ( 
.A(n_7878),
.Y(n_8561)
);

NAND2xp5_ASAP7_75t_L g8562 ( 
.A(n_7804),
.B(n_5002),
.Y(n_8562)
);

BUFx6f_ASAP7_75t_L g8563 ( 
.A(n_7890),
.Y(n_8563)
);

NAND2xp5_ASAP7_75t_SL g8564 ( 
.A(n_8072),
.B(n_5003),
.Y(n_8564)
);

NAND2xp5_ASAP7_75t_SL g8565 ( 
.A(n_8082),
.B(n_5006),
.Y(n_8565)
);

INVx1_ASAP7_75t_L g8566 ( 
.A(n_7881),
.Y(n_8566)
);

INVx1_ASAP7_75t_L g8567 ( 
.A(n_7882),
.Y(n_8567)
);

INVx1_ASAP7_75t_L g8568 ( 
.A(n_7884),
.Y(n_8568)
);

INVx2_ASAP7_75t_SL g8569 ( 
.A(n_7924),
.Y(n_8569)
);

NAND2xp5_ASAP7_75t_L g8570 ( 
.A(n_7829),
.B(n_7895),
.Y(n_8570)
);

NAND2xp5_ASAP7_75t_SL g8571 ( 
.A(n_8095),
.B(n_5007),
.Y(n_8571)
);

NAND2xp5_ASAP7_75t_L g8572 ( 
.A(n_7899),
.B(n_5008),
.Y(n_8572)
);

NAND2xp5_ASAP7_75t_L g8573 ( 
.A(n_7913),
.B(n_5009),
.Y(n_8573)
);

NOR2xp33_ASAP7_75t_SL g8574 ( 
.A(n_8180),
.B(n_5011),
.Y(n_8574)
);

BUFx6f_ASAP7_75t_L g8575 ( 
.A(n_7939),
.Y(n_8575)
);

NAND2xp5_ASAP7_75t_L g8576 ( 
.A(n_7929),
.B(n_5016),
.Y(n_8576)
);

INVx1_ASAP7_75t_L g8577 ( 
.A(n_7887),
.Y(n_8577)
);

INVx1_ASAP7_75t_L g8578 ( 
.A(n_7889),
.Y(n_8578)
);

INVx2_ASAP7_75t_L g8579 ( 
.A(n_7892),
.Y(n_8579)
);

NAND2xp5_ASAP7_75t_L g8580 ( 
.A(n_7894),
.B(n_5020),
.Y(n_8580)
);

AND2x2_ASAP7_75t_L g8581 ( 
.A(n_7797),
.B(n_5021),
.Y(n_8581)
);

AOI22xp5_ASAP7_75t_L g8582 ( 
.A1(n_7642),
.A2(n_5028),
.B1(n_5034),
.B2(n_5027),
.Y(n_8582)
);

BUFx4f_ASAP7_75t_L g8583 ( 
.A(n_8036),
.Y(n_8583)
);

INVx2_ASAP7_75t_L g8584 ( 
.A(n_7900),
.Y(n_8584)
);

AND2x2_ASAP7_75t_L g8585 ( 
.A(n_8009),
.B(n_5035),
.Y(n_8585)
);

NAND2xp5_ASAP7_75t_SL g8586 ( 
.A(n_7941),
.B(n_5036),
.Y(n_8586)
);

AND2x6_ASAP7_75t_L g8587 ( 
.A(n_8034),
.B(n_4640),
.Y(n_8587)
);

INVx3_ASAP7_75t_L g8588 ( 
.A(n_7947),
.Y(n_8588)
);

NAND2xp5_ASAP7_75t_SL g8589 ( 
.A(n_7949),
.B(n_5037),
.Y(n_8589)
);

INVx3_ASAP7_75t_L g8590 ( 
.A(n_7953),
.Y(n_8590)
);

INVxp33_ASAP7_75t_L g8591 ( 
.A(n_8058),
.Y(n_8591)
);

INVx1_ASAP7_75t_L g8592 ( 
.A(n_8001),
.Y(n_8592)
);

INVx3_ASAP7_75t_L g8593 ( 
.A(n_8018),
.Y(n_8593)
);

BUFx6f_ASAP7_75t_L g8594 ( 
.A(n_8030),
.Y(n_8594)
);

NAND2xp5_ASAP7_75t_L g8595 ( 
.A(n_7923),
.B(n_5038),
.Y(n_8595)
);

INVx2_ASAP7_75t_L g8596 ( 
.A(n_7935),
.Y(n_8596)
);

NOR2xp33_ASAP7_75t_L g8597 ( 
.A(n_7741),
.B(n_5039),
.Y(n_8597)
);

INVx3_ASAP7_75t_L g8598 ( 
.A(n_8122),
.Y(n_8598)
);

NOR2xp33_ASAP7_75t_L g8599 ( 
.A(n_7754),
.B(n_5040),
.Y(n_8599)
);

AND2x6_ASAP7_75t_L g8600 ( 
.A(n_8061),
.B(n_4651),
.Y(n_8600)
);

INVx2_ASAP7_75t_L g8601 ( 
.A(n_7938),
.Y(n_8601)
);

BUFx3_ASAP7_75t_L g8602 ( 
.A(n_8119),
.Y(n_8602)
);

AOI22xp33_ASAP7_75t_L g8603 ( 
.A1(n_8017),
.A2(n_4657),
.B1(n_4663),
.B2(n_4652),
.Y(n_8603)
);

INVx3_ASAP7_75t_L g8604 ( 
.A(n_8124),
.Y(n_8604)
);

INVx1_ASAP7_75t_L g8605 ( 
.A(n_8002),
.Y(n_8605)
);

NOR2xp33_ASAP7_75t_L g8606 ( 
.A(n_8112),
.B(n_7930),
.Y(n_8606)
);

BUFx3_ASAP7_75t_L g8607 ( 
.A(n_8121),
.Y(n_8607)
);

INVx2_ASAP7_75t_L g8608 ( 
.A(n_7954),
.Y(n_8608)
);

INVx1_ASAP7_75t_L g8609 ( 
.A(n_8004),
.Y(n_8609)
);

INVx2_ASAP7_75t_SL g8610 ( 
.A(n_8054),
.Y(n_8610)
);

INVx2_ASAP7_75t_L g8611 ( 
.A(n_7961),
.Y(n_8611)
);

INVx2_ASAP7_75t_L g8612 ( 
.A(n_7914),
.Y(n_8612)
);

INVx1_ASAP7_75t_L g8613 ( 
.A(n_8006),
.Y(n_8613)
);

NOR2xp33_ASAP7_75t_L g8614 ( 
.A(n_7950),
.B(n_5044),
.Y(n_8614)
);

BUFx6f_ASAP7_75t_L g8615 ( 
.A(n_8093),
.Y(n_8615)
);

BUFx6f_ASAP7_75t_L g8616 ( 
.A(n_8129),
.Y(n_8616)
);

INVx1_ASAP7_75t_L g8617 ( 
.A(n_8007),
.Y(n_8617)
);

INVx1_ASAP7_75t_L g8618 ( 
.A(n_8010),
.Y(n_8618)
);

BUFx3_ASAP7_75t_L g8619 ( 
.A(n_8126),
.Y(n_8619)
);

INVx2_ASAP7_75t_L g8620 ( 
.A(n_7918),
.Y(n_8620)
);

BUFx6f_ASAP7_75t_L g8621 ( 
.A(n_8096),
.Y(n_8621)
);

INVx1_ASAP7_75t_L g8622 ( 
.A(n_7928),
.Y(n_8622)
);

NOR2xp33_ASAP7_75t_L g8623 ( 
.A(n_7956),
.B(n_5046),
.Y(n_8623)
);

NAND2xp5_ASAP7_75t_L g8624 ( 
.A(n_7934),
.B(n_5049),
.Y(n_8624)
);

HB1xp67_ASAP7_75t_L g8625 ( 
.A(n_7879),
.Y(n_8625)
);

AND2x4_ASAP7_75t_L g8626 ( 
.A(n_8091),
.B(n_4664),
.Y(n_8626)
);

AND2x6_ASAP7_75t_L g8627 ( 
.A(n_8117),
.B(n_4665),
.Y(n_8627)
);

AND2x4_ASAP7_75t_L g8628 ( 
.A(n_8125),
.B(n_4669),
.Y(n_8628)
);

INVx1_ASAP7_75t_L g8629 ( 
.A(n_7943),
.Y(n_8629)
);

OR2x2_ASAP7_75t_L g8630 ( 
.A(n_8063),
.B(n_5051),
.Y(n_8630)
);

BUFx6f_ASAP7_75t_L g8631 ( 
.A(n_8130),
.Y(n_8631)
);

OR2x2_ASAP7_75t_SL g8632 ( 
.A(n_8166),
.B(n_4670),
.Y(n_8632)
);

INVx1_ASAP7_75t_L g8633 ( 
.A(n_7948),
.Y(n_8633)
);

OR2x6_ASAP7_75t_L g8634 ( 
.A(n_8036),
.B(n_4672),
.Y(n_8634)
);

INVx2_ASAP7_75t_L g8635 ( 
.A(n_7951),
.Y(n_8635)
);

AND3x1_ASAP7_75t_L g8636 ( 
.A(n_8108),
.B(n_4676),
.C(n_4675),
.Y(n_8636)
);

INVx1_ASAP7_75t_L g8637 ( 
.A(n_7957),
.Y(n_8637)
);

INVx2_ASAP7_75t_L g8638 ( 
.A(n_7970),
.Y(n_8638)
);

OR2x2_ASAP7_75t_L g8639 ( 
.A(n_7981),
.B(n_5055),
.Y(n_8639)
);

INVx4_ASAP7_75t_L g8640 ( 
.A(n_8118),
.Y(n_8640)
);

AND2x2_ASAP7_75t_L g8641 ( 
.A(n_7773),
.B(n_5056),
.Y(n_8641)
);

INVx2_ASAP7_75t_L g8642 ( 
.A(n_7991),
.Y(n_8642)
);

INVx2_ASAP7_75t_SL g8643 ( 
.A(n_7896),
.Y(n_8643)
);

AND2x2_ASAP7_75t_L g8644 ( 
.A(n_7854),
.B(n_5058),
.Y(n_8644)
);

INVx2_ASAP7_75t_L g8645 ( 
.A(n_7992),
.Y(n_8645)
);

OR2x2_ASAP7_75t_L g8646 ( 
.A(n_7767),
.B(n_5059),
.Y(n_8646)
);

NAND2xp5_ASAP7_75t_SL g8647 ( 
.A(n_7689),
.B(n_5060),
.Y(n_8647)
);

BUFx6f_ASAP7_75t_L g8648 ( 
.A(n_8073),
.Y(n_8648)
);

NOR2xp33_ASAP7_75t_L g8649 ( 
.A(n_7966),
.B(n_5061),
.Y(n_8649)
);

INVx2_ASAP7_75t_L g8650 ( 
.A(n_7993),
.Y(n_8650)
);

INVx1_ASAP7_75t_L g8651 ( 
.A(n_7994),
.Y(n_8651)
);

NOR2xp33_ASAP7_75t_L g8652 ( 
.A(n_7968),
.B(n_5064),
.Y(n_8652)
);

OR2x2_ASAP7_75t_L g8653 ( 
.A(n_7830),
.B(n_5065),
.Y(n_8653)
);

INVx1_ASAP7_75t_L g8654 ( 
.A(n_7995),
.Y(n_8654)
);

INVx1_ASAP7_75t_L g8655 ( 
.A(n_7996),
.Y(n_8655)
);

AND2x4_ASAP7_75t_L g8656 ( 
.A(n_8078),
.B(n_4678),
.Y(n_8656)
);

NOR2xp33_ASAP7_75t_L g8657 ( 
.A(n_8151),
.B(n_5072),
.Y(n_8657)
);

AND2x4_ASAP7_75t_L g8658 ( 
.A(n_8102),
.B(n_4684),
.Y(n_8658)
);

INVx6_ASAP7_75t_L g8659 ( 
.A(n_7963),
.Y(n_8659)
);

INVx2_ASAP7_75t_L g8660 ( 
.A(n_8008),
.Y(n_8660)
);

INVx2_ASAP7_75t_L g8661 ( 
.A(n_8011),
.Y(n_8661)
);

INVx1_ASAP7_75t_L g8662 ( 
.A(n_8014),
.Y(n_8662)
);

AND2x6_ASAP7_75t_L g8663 ( 
.A(n_8027),
.B(n_4685),
.Y(n_8663)
);

AND2x6_ASAP7_75t_L g8664 ( 
.A(n_8032),
.B(n_4688),
.Y(n_8664)
);

INVx3_ASAP7_75t_L g8665 ( 
.A(n_8107),
.Y(n_8665)
);

BUFx10_ASAP7_75t_L g8666 ( 
.A(n_7979),
.Y(n_8666)
);

NAND2xp33_ASAP7_75t_SL g8667 ( 
.A(n_7998),
.B(n_5075),
.Y(n_8667)
);

CKINVDCx5p33_ASAP7_75t_R g8668 ( 
.A(n_7682),
.Y(n_8668)
);

NOR2xp33_ASAP7_75t_L g8669 ( 
.A(n_8141),
.B(n_5076),
.Y(n_8669)
);

NAND2x1p5_ASAP7_75t_L g8670 ( 
.A(n_8035),
.B(n_4689),
.Y(n_8670)
);

INVx3_ASAP7_75t_L g8671 ( 
.A(n_8109),
.Y(n_8671)
);

INVx1_ASAP7_75t_L g8672 ( 
.A(n_8015),
.Y(n_8672)
);

INVx1_ASAP7_75t_L g8673 ( 
.A(n_8016),
.Y(n_8673)
);

INVx5_ASAP7_75t_L g8674 ( 
.A(n_8017),
.Y(n_8674)
);

INVx2_ASAP7_75t_L g8675 ( 
.A(n_8060),
.Y(n_8675)
);

NAND2xp5_ASAP7_75t_L g8676 ( 
.A(n_7883),
.B(n_5078),
.Y(n_8676)
);

NOR2xp33_ASAP7_75t_L g8677 ( 
.A(n_7788),
.B(n_5079),
.Y(n_8677)
);

NOR2xp33_ASAP7_75t_L g8678 ( 
.A(n_8064),
.B(n_5080),
.Y(n_8678)
);

INVx4_ASAP7_75t_L g8679 ( 
.A(n_7931),
.Y(n_8679)
);

AND2x6_ASAP7_75t_L g8680 ( 
.A(n_8037),
.B(n_8079),
.Y(n_8680)
);

BUFx4f_ASAP7_75t_L g8681 ( 
.A(n_8017),
.Y(n_8681)
);

NAND2xp5_ASAP7_75t_SL g8682 ( 
.A(n_7911),
.B(n_5081),
.Y(n_8682)
);

NOR2xp33_ASAP7_75t_L g8683 ( 
.A(n_8065),
.B(n_8069),
.Y(n_8683)
);

INVx2_ASAP7_75t_L g8684 ( 
.A(n_7962),
.Y(n_8684)
);

BUFx6f_ASAP7_75t_L g8685 ( 
.A(n_8110),
.Y(n_8685)
);

OAI22xp5_ASAP7_75t_L g8686 ( 
.A1(n_7737),
.A2(n_5085),
.B1(n_5086),
.B2(n_5082),
.Y(n_8686)
);

INVx1_ASAP7_75t_L g8687 ( 
.A(n_8045),
.Y(n_8687)
);

NAND2xp5_ASAP7_75t_SL g8688 ( 
.A(n_8023),
.B(n_5092),
.Y(n_8688)
);

INVx1_ASAP7_75t_SL g8689 ( 
.A(n_8057),
.Y(n_8689)
);

INVx1_ASAP7_75t_L g8690 ( 
.A(n_8081),
.Y(n_8690)
);

NAND2xp5_ASAP7_75t_SL g8691 ( 
.A(n_8140),
.B(n_8085),
.Y(n_8691)
);

NAND3x1_ASAP7_75t_L g8692 ( 
.A(n_8000),
.B(n_4698),
.C(n_4697),
.Y(n_8692)
);

NAND2xp5_ASAP7_75t_SL g8693 ( 
.A(n_8220),
.B(n_8083),
.Y(n_8693)
);

NAND2xp5_ASAP7_75t_L g8694 ( 
.A(n_8462),
.B(n_8570),
.Y(n_8694)
);

NAND2xp5_ASAP7_75t_L g8695 ( 
.A(n_8412),
.B(n_7978),
.Y(n_8695)
);

AND2x6_ASAP7_75t_L g8696 ( 
.A(n_8689),
.B(n_8086),
.Y(n_8696)
);

INVx1_ASAP7_75t_L g8697 ( 
.A(n_8183),
.Y(n_8697)
);

AOI22xp5_ASAP7_75t_L g8698 ( 
.A1(n_8365),
.A2(n_8156),
.B1(n_7676),
.B2(n_7885),
.Y(n_8698)
);

INVx3_ASAP7_75t_L g8699 ( 
.A(n_8493),
.Y(n_8699)
);

INVx1_ASAP7_75t_L g8700 ( 
.A(n_8191),
.Y(n_8700)
);

AND2x2_ASAP7_75t_L g8701 ( 
.A(n_8301),
.B(n_8229),
.Y(n_8701)
);

INVx2_ASAP7_75t_L g8702 ( 
.A(n_8196),
.Y(n_8702)
);

NAND2xp5_ASAP7_75t_L g8703 ( 
.A(n_8204),
.B(n_7891),
.Y(n_8703)
);

AOI22xp33_ASAP7_75t_L g8704 ( 
.A1(n_8449),
.A2(n_7999),
.B1(n_7960),
.B2(n_7865),
.Y(n_8704)
);

INVx2_ASAP7_75t_L g8705 ( 
.A(n_8212),
.Y(n_8705)
);

NOR3xp33_ASAP7_75t_L g8706 ( 
.A(n_8383),
.B(n_8172),
.C(n_8164),
.Y(n_8706)
);

INVx2_ASAP7_75t_L g8707 ( 
.A(n_8222),
.Y(n_8707)
);

AOI22xp5_ASAP7_75t_L g8708 ( 
.A1(n_8335),
.A2(n_8077),
.B1(n_8076),
.B2(n_8070),
.Y(n_8708)
);

NAND2xp5_ASAP7_75t_L g8709 ( 
.A(n_8585),
.B(n_7898),
.Y(n_8709)
);

NAND2xp5_ASAP7_75t_L g8710 ( 
.A(n_8389),
.B(n_7852),
.Y(n_8710)
);

AOI22xp5_ASAP7_75t_L g8711 ( 
.A1(n_8201),
.A2(n_8358),
.B1(n_8424),
.B2(n_8491),
.Y(n_8711)
);

INVx1_ASAP7_75t_L g8712 ( 
.A(n_8227),
.Y(n_8712)
);

INVx1_ASAP7_75t_L g8713 ( 
.A(n_8228),
.Y(n_8713)
);

NOR2xp33_ASAP7_75t_L g8714 ( 
.A(n_8378),
.B(n_8159),
.Y(n_8714)
);

INVx1_ASAP7_75t_L g8715 ( 
.A(n_8230),
.Y(n_8715)
);

NAND2xp5_ASAP7_75t_SL g8716 ( 
.A(n_8373),
.B(n_8503),
.Y(n_8716)
);

NAND2xp5_ASAP7_75t_L g8717 ( 
.A(n_8395),
.B(n_7959),
.Y(n_8717)
);

NAND2xp5_ASAP7_75t_L g8718 ( 
.A(n_8436),
.B(n_8139),
.Y(n_8718)
);

INVx1_ASAP7_75t_L g8719 ( 
.A(n_8234),
.Y(n_8719)
);

NAND2xp5_ASAP7_75t_SL g8720 ( 
.A(n_8469),
.B(n_8116),
.Y(n_8720)
);

NAND2xp5_ASAP7_75t_SL g8721 ( 
.A(n_8423),
.B(n_8099),
.Y(n_8721)
);

INVx1_ASAP7_75t_L g8722 ( 
.A(n_8240),
.Y(n_8722)
);

NAND2xp5_ASAP7_75t_SL g8723 ( 
.A(n_8262),
.B(n_8100),
.Y(n_8723)
);

NAND2xp5_ASAP7_75t_L g8724 ( 
.A(n_8581),
.B(n_8162),
.Y(n_8724)
);

INVx3_ASAP7_75t_L g8725 ( 
.A(n_8506),
.Y(n_8725)
);

INVx2_ASAP7_75t_L g8726 ( 
.A(n_8245),
.Y(n_8726)
);

INVx1_ASAP7_75t_L g8727 ( 
.A(n_8258),
.Y(n_8727)
);

NOR2xp33_ASAP7_75t_L g8728 ( 
.A(n_8247),
.B(n_8176),
.Y(n_8728)
);

INVx2_ASAP7_75t_SL g8729 ( 
.A(n_8510),
.Y(n_8729)
);

NAND2xp5_ASAP7_75t_L g8730 ( 
.A(n_8404),
.B(n_7925),
.Y(n_8730)
);

INVxp67_ASAP7_75t_SL g8731 ( 
.A(n_8303),
.Y(n_8731)
);

NAND2xp5_ASAP7_75t_L g8732 ( 
.A(n_8187),
.B(n_8418),
.Y(n_8732)
);

NAND2xp5_ASAP7_75t_L g8733 ( 
.A(n_8323),
.B(n_8106),
.Y(n_8733)
);

NOR2xp33_ASAP7_75t_L g8734 ( 
.A(n_8251),
.B(n_8179),
.Y(n_8734)
);

NOR2xp67_ASAP7_75t_L g8735 ( 
.A(n_8208),
.B(n_8111),
.Y(n_8735)
);

OR2x2_ASAP7_75t_L g8736 ( 
.A(n_8409),
.B(n_8114),
.Y(n_8736)
);

NAND2xp5_ASAP7_75t_L g8737 ( 
.A(n_8324),
.B(n_7667),
.Y(n_8737)
);

OR2x6_ASAP7_75t_L g8738 ( 
.A(n_8279),
.B(n_8052),
.Y(n_8738)
);

INVx2_ASAP7_75t_L g8739 ( 
.A(n_8259),
.Y(n_8739)
);

NOR2xp33_ASAP7_75t_SL g8740 ( 
.A(n_8185),
.B(n_5099),
.Y(n_8740)
);

INVx2_ASAP7_75t_L g8741 ( 
.A(n_8263),
.Y(n_8741)
);

NAND2xp5_ASAP7_75t_L g8742 ( 
.A(n_8328),
.B(n_7977),
.Y(n_8742)
);

NAND2xp5_ASAP7_75t_SL g8743 ( 
.A(n_8414),
.B(n_7748),
.Y(n_8743)
);

NAND2xp5_ASAP7_75t_L g8744 ( 
.A(n_8211),
.B(n_7980),
.Y(n_8744)
);

AOI22xp5_ASAP7_75t_L g8745 ( 
.A1(n_8375),
.A2(n_7818),
.B1(n_7984),
.B2(n_7983),
.Y(n_8745)
);

INVx2_ASAP7_75t_L g8746 ( 
.A(n_8264),
.Y(n_8746)
);

INVx2_ASAP7_75t_L g8747 ( 
.A(n_8273),
.Y(n_8747)
);

NOR2x1p5_ASAP7_75t_L g8748 ( 
.A(n_8421),
.B(n_8144),
.Y(n_8748)
);

INVx2_ASAP7_75t_L g8749 ( 
.A(n_8278),
.Y(n_8749)
);

INVx1_ASAP7_75t_L g8750 ( 
.A(n_8286),
.Y(n_8750)
);

NAND2xp33_ASAP7_75t_L g8751 ( 
.A(n_8680),
.B(n_7985),
.Y(n_8751)
);

NAND2xp5_ASAP7_75t_L g8752 ( 
.A(n_8431),
.B(n_7904),
.Y(n_8752)
);

INVx3_ASAP7_75t_L g8753 ( 
.A(n_8480),
.Y(n_8753)
);

NAND2xp5_ASAP7_75t_SL g8754 ( 
.A(n_8523),
.B(n_7933),
.Y(n_8754)
);

INVx1_ASAP7_75t_L g8755 ( 
.A(n_8291),
.Y(n_8755)
);

AND2x2_ASAP7_75t_L g8756 ( 
.A(n_8300),
.B(n_5100),
.Y(n_8756)
);

AND2x2_ASAP7_75t_L g8757 ( 
.A(n_8475),
.B(n_5102),
.Y(n_8757)
);

INVx2_ASAP7_75t_L g8758 ( 
.A(n_8297),
.Y(n_8758)
);

INVx1_ASAP7_75t_L g8759 ( 
.A(n_8307),
.Y(n_8759)
);

NAND2xp5_ASAP7_75t_SL g8760 ( 
.A(n_8607),
.B(n_5107),
.Y(n_8760)
);

BUFx8_ASAP7_75t_L g8761 ( 
.A(n_8226),
.Y(n_8761)
);

AND2x2_ASAP7_75t_L g8762 ( 
.A(n_8641),
.B(n_5109),
.Y(n_8762)
);

NAND2xp5_ASAP7_75t_SL g8763 ( 
.A(n_8619),
.B(n_5113),
.Y(n_8763)
);

O2A1O1Ixp33_ASAP7_75t_L g8764 ( 
.A1(n_8677),
.A2(n_4704),
.B(n_4706),
.C(n_4703),
.Y(n_8764)
);

NAND2xp5_ASAP7_75t_L g8765 ( 
.A(n_8442),
.B(n_4708),
.Y(n_8765)
);

NAND2x1p5_ASAP7_75t_L g8766 ( 
.A(n_8480),
.B(n_8055),
.Y(n_8766)
);

AND2x2_ASAP7_75t_L g8767 ( 
.A(n_8644),
.B(n_5114),
.Y(n_8767)
);

AND2x6_ASAP7_75t_L g8768 ( 
.A(n_8309),
.B(n_8020),
.Y(n_8768)
);

NAND2xp5_ASAP7_75t_L g8769 ( 
.A(n_8460),
.B(n_4717),
.Y(n_8769)
);

NAND2xp5_ASAP7_75t_SL g8770 ( 
.A(n_8518),
.B(n_5117),
.Y(n_8770)
);

INVx2_ASAP7_75t_L g8771 ( 
.A(n_8318),
.Y(n_8771)
);

INVx2_ASAP7_75t_L g8772 ( 
.A(n_8334),
.Y(n_8772)
);

OAI22xp5_ASAP7_75t_L g8773 ( 
.A1(n_8336),
.A2(n_8033),
.B1(n_8024),
.B2(n_5124),
.Y(n_8773)
);

INVx1_ASAP7_75t_L g8774 ( 
.A(n_8339),
.Y(n_8774)
);

NOR2xp33_ASAP7_75t_L g8775 ( 
.A(n_8473),
.B(n_5122),
.Y(n_8775)
);

NAND2xp5_ASAP7_75t_L g8776 ( 
.A(n_8494),
.B(n_8526),
.Y(n_8776)
);

BUFx8_ASAP7_75t_L g8777 ( 
.A(n_8239),
.Y(n_8777)
);

NAND2xp5_ASAP7_75t_L g8778 ( 
.A(n_8536),
.B(n_4730),
.Y(n_8778)
);

NAND2xp5_ASAP7_75t_SL g8779 ( 
.A(n_8331),
.B(n_8261),
.Y(n_8779)
);

NAND2xp5_ASAP7_75t_SL g8780 ( 
.A(n_8266),
.B(n_5125),
.Y(n_8780)
);

NAND2xp5_ASAP7_75t_L g8781 ( 
.A(n_8542),
.B(n_4737),
.Y(n_8781)
);

NAND2xp5_ASAP7_75t_L g8782 ( 
.A(n_8548),
.B(n_4740),
.Y(n_8782)
);

AND2x4_ASAP7_75t_L g8783 ( 
.A(n_8362),
.B(n_7945),
.Y(n_8783)
);

NAND2xp5_ASAP7_75t_L g8784 ( 
.A(n_8562),
.B(n_4741),
.Y(n_8784)
);

AOI22xp5_ASAP7_75t_L g8785 ( 
.A1(n_8357),
.A2(n_8047),
.B1(n_8042),
.B2(n_5129),
.Y(n_8785)
);

INVx2_ASAP7_75t_L g8786 ( 
.A(n_8342),
.Y(n_8786)
);

CKINVDCx20_ASAP7_75t_R g8787 ( 
.A(n_8238),
.Y(n_8787)
);

NAND2xp5_ASAP7_75t_SL g8788 ( 
.A(n_8270),
.B(n_5128),
.Y(n_8788)
);

NAND2xp33_ASAP7_75t_L g8789 ( 
.A(n_8680),
.B(n_5130),
.Y(n_8789)
);

AOI22xp5_ASAP7_75t_L g8790 ( 
.A1(n_8450),
.A2(n_5137),
.B1(n_5140),
.B2(n_5136),
.Y(n_8790)
);

INVx1_ASAP7_75t_L g8791 ( 
.A(n_8345),
.Y(n_8791)
);

NAND2xp5_ASAP7_75t_L g8792 ( 
.A(n_8572),
.B(n_4745),
.Y(n_8792)
);

OAI22xp5_ASAP7_75t_L g8793 ( 
.A1(n_8346),
.A2(n_5145),
.B1(n_5146),
.B2(n_5142),
.Y(n_8793)
);

NAND2xp5_ASAP7_75t_SL g8794 ( 
.A(n_8290),
.B(n_5147),
.Y(n_8794)
);

NOR2xp33_ASAP7_75t_L g8795 ( 
.A(n_8573),
.B(n_5151),
.Y(n_8795)
);

NAND3xp33_ASAP7_75t_L g8796 ( 
.A(n_8669),
.B(n_5154),
.C(n_5153),
.Y(n_8796)
);

NOR2xp33_ASAP7_75t_L g8797 ( 
.A(n_8415),
.B(n_5155),
.Y(n_8797)
);

INVx2_ASAP7_75t_L g8798 ( 
.A(n_8363),
.Y(n_8798)
);

NAND2xp5_ASAP7_75t_L g8799 ( 
.A(n_8576),
.B(n_4747),
.Y(n_8799)
);

NAND2x1_ASAP7_75t_L g8800 ( 
.A(n_8679),
.B(n_4749),
.Y(n_8800)
);

NOR2xp33_ASAP7_75t_L g8801 ( 
.A(n_8304),
.B(n_5156),
.Y(n_8801)
);

NAND2xp5_ASAP7_75t_SL g8802 ( 
.A(n_8320),
.B(n_5157),
.Y(n_8802)
);

NOR2xp33_ASAP7_75t_L g8803 ( 
.A(n_8315),
.B(n_5158),
.Y(n_8803)
);

NAND2xp5_ASAP7_75t_L g8804 ( 
.A(n_8367),
.B(n_4762),
.Y(n_8804)
);

INVx1_ASAP7_75t_SL g8805 ( 
.A(n_8368),
.Y(n_8805)
);

INVx1_ASAP7_75t_L g8806 ( 
.A(n_8371),
.Y(n_8806)
);

NAND2xp5_ASAP7_75t_L g8807 ( 
.A(n_8381),
.B(n_4763),
.Y(n_8807)
);

INVx2_ASAP7_75t_SL g8808 ( 
.A(n_8195),
.Y(n_8808)
);

NAND2xp5_ASAP7_75t_SL g8809 ( 
.A(n_8208),
.B(n_5160),
.Y(n_8809)
);

INVx1_ASAP7_75t_L g8810 ( 
.A(n_8388),
.Y(n_8810)
);

NOR2xp33_ASAP7_75t_L g8811 ( 
.A(n_8321),
.B(n_5166),
.Y(n_8811)
);

INVx2_ASAP7_75t_L g8812 ( 
.A(n_8622),
.Y(n_8812)
);

NAND2xp5_ASAP7_75t_SL g8813 ( 
.A(n_8621),
.B(n_5167),
.Y(n_8813)
);

NOR2xp33_ASAP7_75t_L g8814 ( 
.A(n_8341),
.B(n_5168),
.Y(n_8814)
);

INVx2_ASAP7_75t_L g8815 ( 
.A(n_8629),
.Y(n_8815)
);

NAND2xp5_ASAP7_75t_L g8816 ( 
.A(n_8231),
.B(n_4765),
.Y(n_8816)
);

NAND2xp5_ASAP7_75t_SL g8817 ( 
.A(n_8621),
.B(n_5170),
.Y(n_8817)
);

INVx3_ASAP7_75t_L g8818 ( 
.A(n_8289),
.Y(n_8818)
);

BUFx6f_ASAP7_75t_L g8819 ( 
.A(n_8195),
.Y(n_8819)
);

NAND2xp5_ASAP7_75t_L g8820 ( 
.A(n_8243),
.B(n_4766),
.Y(n_8820)
);

NAND2xp5_ASAP7_75t_SL g8821 ( 
.A(n_8668),
.B(n_5173),
.Y(n_8821)
);

NOR3xp33_ASAP7_75t_L g8822 ( 
.A(n_8438),
.B(n_4775),
.C(n_4767),
.Y(n_8822)
);

NAND2xp5_ASAP7_75t_SL g8823 ( 
.A(n_8190),
.B(n_5174),
.Y(n_8823)
);

CKINVDCx20_ASAP7_75t_R g8824 ( 
.A(n_8253),
.Y(n_8824)
);

NAND2xp5_ASAP7_75t_L g8825 ( 
.A(n_8254),
.B(n_4776),
.Y(n_8825)
);

NAND2xp5_ASAP7_75t_L g8826 ( 
.A(n_8271),
.B(n_4777),
.Y(n_8826)
);

NOR2xp33_ASAP7_75t_L g8827 ( 
.A(n_8444),
.B(n_5175),
.Y(n_8827)
);

NAND2xp5_ASAP7_75t_L g8828 ( 
.A(n_8287),
.B(n_4782),
.Y(n_8828)
);

INVxp67_ASAP7_75t_L g8829 ( 
.A(n_8554),
.Y(n_8829)
);

OAI22xp33_ASAP7_75t_L g8830 ( 
.A1(n_8268),
.A2(n_5179),
.B1(n_5181),
.B2(n_5177),
.Y(n_8830)
);

INVx1_ASAP7_75t_L g8831 ( 
.A(n_8390),
.Y(n_8831)
);

INVx1_ASAP7_75t_L g8832 ( 
.A(n_8394),
.Y(n_8832)
);

NAND2xp5_ASAP7_75t_L g8833 ( 
.A(n_8288),
.B(n_4785),
.Y(n_8833)
);

INVx1_ASAP7_75t_L g8834 ( 
.A(n_8396),
.Y(n_8834)
);

INVx1_ASAP7_75t_L g8835 ( 
.A(n_8400),
.Y(n_8835)
);

NAND2xp5_ASAP7_75t_L g8836 ( 
.A(n_8319),
.B(n_4786),
.Y(n_8836)
);

INVx2_ASAP7_75t_L g8837 ( 
.A(n_8633),
.Y(n_8837)
);

NAND2xp5_ASAP7_75t_L g8838 ( 
.A(n_8606),
.B(n_4787),
.Y(n_8838)
);

NAND2xp5_ASAP7_75t_L g8839 ( 
.A(n_8592),
.B(n_4797),
.Y(n_8839)
);

NAND2xp5_ASAP7_75t_L g8840 ( 
.A(n_8605),
.B(n_4805),
.Y(n_8840)
);

NAND2xp5_ASAP7_75t_SL g8841 ( 
.A(n_8615),
.B(n_5182),
.Y(n_8841)
);

NAND2x1p5_ASAP7_75t_L g8842 ( 
.A(n_8218),
.B(n_4808),
.Y(n_8842)
);

NOR2x1p5_ASAP7_75t_L g8843 ( 
.A(n_8246),
.B(n_5183),
.Y(n_8843)
);

INVx1_ASAP7_75t_L g8844 ( 
.A(n_8401),
.Y(n_8844)
);

NAND2xp5_ASAP7_75t_L g8845 ( 
.A(n_8609),
.B(n_4821),
.Y(n_8845)
);

NAND2xp5_ASAP7_75t_SL g8846 ( 
.A(n_8615),
.B(n_5191),
.Y(n_8846)
);

O2A1O1Ixp33_ASAP7_75t_L g8847 ( 
.A1(n_8330),
.A2(n_8340),
.B(n_8688),
.C(n_8682),
.Y(n_8847)
);

INVx2_ASAP7_75t_L g8848 ( 
.A(n_8637),
.Y(n_8848)
);

INVx2_ASAP7_75t_L g8849 ( 
.A(n_8612),
.Y(n_8849)
);

NAND2xp5_ASAP7_75t_L g8850 ( 
.A(n_8613),
.B(n_4837),
.Y(n_8850)
);

NAND2xp5_ASAP7_75t_SL g8851 ( 
.A(n_8574),
.B(n_5193),
.Y(n_8851)
);

NAND2xp5_ASAP7_75t_L g8852 ( 
.A(n_8617),
.B(n_4841),
.Y(n_8852)
);

NOR3xp33_ASAP7_75t_L g8853 ( 
.A(n_8488),
.B(n_4845),
.C(n_4842),
.Y(n_8853)
);

INVx4_ASAP7_75t_L g8854 ( 
.A(n_8206),
.Y(n_8854)
);

BUFx3_ASAP7_75t_L g8855 ( 
.A(n_8194),
.Y(n_8855)
);

NAND2xp5_ASAP7_75t_L g8856 ( 
.A(n_8618),
.B(n_4867),
.Y(n_8856)
);

NAND2xp5_ASAP7_75t_SL g8857 ( 
.A(n_8559),
.B(n_5194),
.Y(n_8857)
);

INVxp33_ASAP7_75t_L g8858 ( 
.A(n_8512),
.Y(n_8858)
);

AND2x2_ASAP7_75t_L g8859 ( 
.A(n_8490),
.B(n_5195),
.Y(n_8859)
);

NAND2xp5_ASAP7_75t_SL g8860 ( 
.A(n_8364),
.B(n_5197),
.Y(n_8860)
);

NAND2xp5_ASAP7_75t_L g8861 ( 
.A(n_8387),
.B(n_8683),
.Y(n_8861)
);

NOR2xp33_ASAP7_75t_L g8862 ( 
.A(n_8464),
.B(n_5198),
.Y(n_8862)
);

NAND2xp5_ASAP7_75t_SL g8863 ( 
.A(n_8244),
.B(n_5200),
.Y(n_8863)
);

BUFx3_ASAP7_75t_L g8864 ( 
.A(n_8206),
.Y(n_8864)
);

NOR2xp33_ASAP7_75t_L g8865 ( 
.A(n_8591),
.B(n_8348),
.Y(n_8865)
);

OR2x2_ASAP7_75t_L g8866 ( 
.A(n_8298),
.B(n_5202),
.Y(n_8866)
);

NAND2xp5_ASAP7_75t_L g8867 ( 
.A(n_8402),
.B(n_4868),
.Y(n_8867)
);

INVx1_ASAP7_75t_L g8868 ( 
.A(n_8406),
.Y(n_8868)
);

OAI22xp33_ASAP7_75t_L g8869 ( 
.A1(n_8535),
.A2(n_8582),
.B1(n_8216),
.B2(n_8551),
.Y(n_8869)
);

INVx8_ASAP7_75t_L g8870 ( 
.A(n_8302),
.Y(n_8870)
);

INVx1_ASAP7_75t_L g8871 ( 
.A(n_8413),
.Y(n_8871)
);

NAND2xp5_ASAP7_75t_SL g8872 ( 
.A(n_8184),
.B(n_5203),
.Y(n_8872)
);

INVx2_ASAP7_75t_L g8873 ( 
.A(n_8620),
.Y(n_8873)
);

NAND2xp5_ASAP7_75t_L g8874 ( 
.A(n_8417),
.B(n_8433),
.Y(n_8874)
);

OAI22xp33_ASAP7_75t_L g8875 ( 
.A1(n_8583),
.A2(n_5206),
.B1(n_5207),
.B2(n_5204),
.Y(n_8875)
);

NAND2xp5_ASAP7_75t_L g8876 ( 
.A(n_8440),
.B(n_4874),
.Y(n_8876)
);

NOR2xp33_ASAP7_75t_L g8877 ( 
.A(n_8276),
.B(n_5208),
.Y(n_8877)
);

NAND2xp5_ASAP7_75t_L g8878 ( 
.A(n_8447),
.B(n_4876),
.Y(n_8878)
);

INVx2_ASAP7_75t_L g8879 ( 
.A(n_8635),
.Y(n_8879)
);

NAND2xp5_ASAP7_75t_L g8880 ( 
.A(n_8448),
.B(n_4907),
.Y(n_8880)
);

NAND2xp5_ASAP7_75t_L g8881 ( 
.A(n_8452),
.B(n_4909),
.Y(n_8881)
);

BUFx3_ASAP7_75t_L g8882 ( 
.A(n_8219),
.Y(n_8882)
);

O2A1O1Ixp33_ASAP7_75t_L g8883 ( 
.A1(n_8360),
.A2(n_4914),
.B(n_4928),
.C(n_4913),
.Y(n_8883)
);

NAND2xp5_ASAP7_75t_L g8884 ( 
.A(n_8453),
.B(n_4936),
.Y(n_8884)
);

INVx1_ASAP7_75t_L g8885 ( 
.A(n_8456),
.Y(n_8885)
);

INVx2_ASAP7_75t_SL g8886 ( 
.A(n_8219),
.Y(n_8886)
);

INVx1_ASAP7_75t_L g8887 ( 
.A(n_8458),
.Y(n_8887)
);

NOR2xp33_ASAP7_75t_L g8888 ( 
.A(n_8225),
.B(n_5211),
.Y(n_8888)
);

NAND2xp5_ASAP7_75t_L g8889 ( 
.A(n_8465),
.B(n_4937),
.Y(n_8889)
);

NAND2xp33_ASAP7_75t_L g8890 ( 
.A(n_8445),
.B(n_5213),
.Y(n_8890)
);

INVx2_ASAP7_75t_L g8891 ( 
.A(n_8467),
.Y(n_8891)
);

NAND2xp5_ASAP7_75t_L g8892 ( 
.A(n_8182),
.B(n_4948),
.Y(n_8892)
);

NAND2xp5_ASAP7_75t_L g8893 ( 
.A(n_8192),
.B(n_4952),
.Y(n_8893)
);

NAND2x1p5_ASAP7_75t_L g8894 ( 
.A(n_8233),
.B(n_4961),
.Y(n_8894)
);

INVxp67_ASAP7_75t_SL g8895 ( 
.A(n_8422),
.Y(n_8895)
);

A2O1A1Ixp33_ASAP7_75t_L g8896 ( 
.A1(n_8597),
.A2(n_4966),
.B(n_4979),
.C(n_4962),
.Y(n_8896)
);

INVx2_ASAP7_75t_L g8897 ( 
.A(n_8684),
.Y(n_8897)
);

AND2x2_ASAP7_75t_L g8898 ( 
.A(n_8498),
.B(n_5215),
.Y(n_8898)
);

INVxp67_ASAP7_75t_L g8899 ( 
.A(n_8343),
.Y(n_8899)
);

AOI221xp5_ASAP7_75t_L g8900 ( 
.A1(n_8403),
.A2(n_4984),
.B1(n_4985),
.B2(n_4983),
.C(n_4982),
.Y(n_8900)
);

NAND2xp5_ASAP7_75t_L g8901 ( 
.A(n_8193),
.B(n_4987),
.Y(n_8901)
);

INVx1_ASAP7_75t_L g8902 ( 
.A(n_8199),
.Y(n_8902)
);

INVx1_ASAP7_75t_L g8903 ( 
.A(n_8200),
.Y(n_8903)
);

OR2x2_ASAP7_75t_L g8904 ( 
.A(n_8379),
.B(n_5219),
.Y(n_8904)
);

BUFx6f_ASAP7_75t_L g8905 ( 
.A(n_8255),
.Y(n_8905)
);

NAND2xp5_ASAP7_75t_L g8906 ( 
.A(n_8215),
.B(n_4990),
.Y(n_8906)
);

INVx1_ASAP7_75t_L g8907 ( 
.A(n_8217),
.Y(n_8907)
);

INVx2_ASAP7_75t_L g8908 ( 
.A(n_8248),
.Y(n_8908)
);

AOI21xp5_ASAP7_75t_L g8909 ( 
.A1(n_8691),
.A2(n_8505),
.B(n_8558),
.Y(n_8909)
);

BUFx3_ASAP7_75t_L g8910 ( 
.A(n_8255),
.Y(n_8910)
);

INVx8_ASAP7_75t_L g8911 ( 
.A(n_8260),
.Y(n_8911)
);

NOR2xp33_ASAP7_75t_L g8912 ( 
.A(n_8236),
.B(n_5230),
.Y(n_8912)
);

INVx1_ASAP7_75t_L g8913 ( 
.A(n_8267),
.Y(n_8913)
);

INVx2_ASAP7_75t_L g8914 ( 
.A(n_8280),
.Y(n_8914)
);

NAND2xp33_ASAP7_75t_L g8915 ( 
.A(n_8543),
.B(n_5232),
.Y(n_8915)
);

NAND2xp5_ASAP7_75t_L g8916 ( 
.A(n_8281),
.B(n_4992),
.Y(n_8916)
);

INVx2_ASAP7_75t_SL g8917 ( 
.A(n_8260),
.Y(n_8917)
);

NOR2x1p5_ASAP7_75t_L g8918 ( 
.A(n_8269),
.B(n_5241),
.Y(n_8918)
);

NAND2xp5_ASAP7_75t_SL g8919 ( 
.A(n_8186),
.B(n_5242),
.Y(n_8919)
);

NAND2xp5_ASAP7_75t_SL g8920 ( 
.A(n_8237),
.B(n_5246),
.Y(n_8920)
);

AOI22xp5_ASAP7_75t_L g8921 ( 
.A1(n_8657),
.A2(n_5251),
.B1(n_5252),
.B2(n_5247),
.Y(n_8921)
);

INVx1_ASAP7_75t_L g8922 ( 
.A(n_8285),
.Y(n_8922)
);

NAND2xp5_ASAP7_75t_L g8923 ( 
.A(n_8292),
.B(n_4996),
.Y(n_8923)
);

INVx1_ASAP7_75t_L g8924 ( 
.A(n_8306),
.Y(n_8924)
);

AOI21xp5_ASAP7_75t_L g8925 ( 
.A1(n_8564),
.A2(n_5004),
.B(n_4998),
.Y(n_8925)
);

NAND2xp5_ASAP7_75t_L g8926 ( 
.A(n_8322),
.B(n_5018),
.Y(n_8926)
);

BUFx2_ASAP7_75t_L g8927 ( 
.A(n_8295),
.Y(n_8927)
);

NAND2xp5_ASAP7_75t_L g8928 ( 
.A(n_8329),
.B(n_5025),
.Y(n_8928)
);

NOR2xp33_ASAP7_75t_L g8929 ( 
.A(n_8630),
.B(n_5256),
.Y(n_8929)
);

BUFx5_ASAP7_75t_L g8930 ( 
.A(n_8472),
.Y(n_8930)
);

NAND2xp5_ASAP7_75t_SL g8931 ( 
.A(n_8213),
.B(n_8429),
.Y(n_8931)
);

NAND2xp5_ASAP7_75t_SL g8932 ( 
.A(n_8283),
.B(n_5258),
.Y(n_8932)
);

INVx2_ASAP7_75t_SL g8933 ( 
.A(n_8295),
.Y(n_8933)
);

NAND2xp5_ASAP7_75t_SL g8934 ( 
.A(n_8674),
.B(n_5259),
.Y(n_8934)
);

NAND2xp5_ASAP7_75t_L g8935 ( 
.A(n_8337),
.B(n_8349),
.Y(n_8935)
);

NAND2xp5_ASAP7_75t_L g8936 ( 
.A(n_8366),
.B(n_5026),
.Y(n_8936)
);

INVx2_ASAP7_75t_SL g8937 ( 
.A(n_8316),
.Y(n_8937)
);

NOR2xp33_ASAP7_75t_L g8938 ( 
.A(n_8299),
.B(n_5262),
.Y(n_8938)
);

NAND2xp33_ASAP7_75t_SL g8939 ( 
.A(n_8521),
.B(n_5263),
.Y(n_8939)
);

NOR2xp33_ASAP7_75t_L g8940 ( 
.A(n_8500),
.B(n_5264),
.Y(n_8940)
);

INVx2_ASAP7_75t_SL g8941 ( 
.A(n_8316),
.Y(n_8941)
);

BUFx3_ASAP7_75t_L g8942 ( 
.A(n_8257),
.Y(n_8942)
);

INVx2_ASAP7_75t_L g8943 ( 
.A(n_8393),
.Y(n_8943)
);

NAND2xp5_ASAP7_75t_L g8944 ( 
.A(n_8474),
.B(n_5041),
.Y(n_8944)
);

CKINVDCx20_ASAP7_75t_R g8945 ( 
.A(n_8202),
.Y(n_8945)
);

NAND2xp5_ASAP7_75t_L g8946 ( 
.A(n_8481),
.B(n_8553),
.Y(n_8946)
);

NOR3xp33_ASAP7_75t_L g8947 ( 
.A(n_8407),
.B(n_5047),
.C(n_5043),
.Y(n_8947)
);

NOR2xp33_ASAP7_75t_L g8948 ( 
.A(n_8599),
.B(n_5265),
.Y(n_8948)
);

INVx2_ASAP7_75t_L g8949 ( 
.A(n_8397),
.Y(n_8949)
);

INVx1_ASAP7_75t_L g8950 ( 
.A(n_8485),
.Y(n_8950)
);

NAND2xp5_ASAP7_75t_L g8951 ( 
.A(n_8614),
.B(n_5048),
.Y(n_8951)
);

NAND2xp5_ASAP7_75t_L g8952 ( 
.A(n_8623),
.B(n_5052),
.Y(n_8952)
);

AOI22xp5_ASAP7_75t_L g8953 ( 
.A1(n_8221),
.A2(n_5269),
.B1(n_5274),
.B2(n_5266),
.Y(n_8953)
);

NOR2xp67_ASAP7_75t_L g8954 ( 
.A(n_8443),
.B(n_5),
.Y(n_8954)
);

NAND2xp5_ASAP7_75t_L g8955 ( 
.A(n_8649),
.B(n_5054),
.Y(n_8955)
);

NOR2x1p5_ASAP7_75t_L g8956 ( 
.A(n_8377),
.B(n_5276),
.Y(n_8956)
);

OAI22x1_ASAP7_75t_SL g8957 ( 
.A1(n_8497),
.A2(n_5280),
.B1(n_5282),
.B2(n_5277),
.Y(n_8957)
);

INVx2_ASAP7_75t_L g8958 ( 
.A(n_8411),
.Y(n_8958)
);

INVxp33_ASAP7_75t_SL g8959 ( 
.A(n_8355),
.Y(n_8959)
);

NAND2xp5_ASAP7_75t_L g8960 ( 
.A(n_8652),
.B(n_5057),
.Y(n_8960)
);

INVx2_ASAP7_75t_L g8961 ( 
.A(n_8430),
.Y(n_8961)
);

NAND2xp5_ASAP7_75t_SL g8962 ( 
.A(n_8674),
.B(n_5283),
.Y(n_8962)
);

INVx2_ASAP7_75t_SL g8963 ( 
.A(n_8282),
.Y(n_8963)
);

INVx2_ASAP7_75t_SL g8964 ( 
.A(n_8338),
.Y(n_8964)
);

INVx1_ASAP7_75t_L g8965 ( 
.A(n_8495),
.Y(n_8965)
);

NOR2xp33_ASAP7_75t_L g8966 ( 
.A(n_8209),
.B(n_5285),
.Y(n_8966)
);

NAND2xp5_ASAP7_75t_L g8967 ( 
.A(n_8608),
.B(n_5062),
.Y(n_8967)
);

NAND2xp5_ASAP7_75t_L g8968 ( 
.A(n_8611),
.B(n_5068),
.Y(n_8968)
);

INVx2_ASAP7_75t_L g8969 ( 
.A(n_8432),
.Y(n_8969)
);

NAND2xp5_ASAP7_75t_L g8970 ( 
.A(n_8529),
.B(n_5069),
.Y(n_8970)
);

AND2x6_ASAP7_75t_SL g8971 ( 
.A(n_8224),
.B(n_5073),
.Y(n_8971)
);

AND2x4_ASAP7_75t_L g8972 ( 
.A(n_8434),
.B(n_5077),
.Y(n_8972)
);

INVx1_ASAP7_75t_L g8973 ( 
.A(n_8501),
.Y(n_8973)
);

OAI22xp33_ASAP7_75t_L g8974 ( 
.A1(n_8670),
.A2(n_5289),
.B1(n_5292),
.B2(n_5288),
.Y(n_8974)
);

NAND2xp5_ASAP7_75t_SL g8975 ( 
.A(n_8631),
.B(n_5294),
.Y(n_8975)
);

NAND2xp5_ASAP7_75t_SL g8976 ( 
.A(n_8631),
.B(n_5298),
.Y(n_8976)
);

INVx1_ASAP7_75t_SL g8977 ( 
.A(n_8249),
.Y(n_8977)
);

NAND2xp5_ASAP7_75t_L g8978 ( 
.A(n_8595),
.B(n_5084),
.Y(n_8978)
);

INVx3_ASAP7_75t_L g8979 ( 
.A(n_8294),
.Y(n_8979)
);

INVx1_ASAP7_75t_SL g8980 ( 
.A(n_8384),
.Y(n_8980)
);

NOR3xp33_ASAP7_75t_L g8981 ( 
.A(n_8678),
.B(n_8571),
.C(n_8565),
.Y(n_8981)
);

INVx1_ASAP7_75t_L g8982 ( 
.A(n_8502),
.Y(n_8982)
);

INVx1_ASAP7_75t_L g8983 ( 
.A(n_8504),
.Y(n_8983)
);

NAND2xp33_ASAP7_75t_L g8984 ( 
.A(n_8543),
.B(n_5299),
.Y(n_8984)
);

NAND2xp5_ASAP7_75t_L g8985 ( 
.A(n_8333),
.B(n_5090),
.Y(n_8985)
);

INVx1_ASAP7_75t_L g8986 ( 
.A(n_8507),
.Y(n_8986)
);

NAND2xp5_ASAP7_75t_L g8987 ( 
.A(n_8344),
.B(n_5091),
.Y(n_8987)
);

NOR2xp33_ASAP7_75t_L g8988 ( 
.A(n_8646),
.B(n_8653),
.Y(n_8988)
);

NOR2xp33_ASAP7_75t_L g8989 ( 
.A(n_8639),
.B(n_5300),
.Y(n_8989)
);

AOI22xp5_ASAP7_75t_SL g8990 ( 
.A1(n_8420),
.A2(n_5304),
.B1(n_5310),
.B2(n_5302),
.Y(n_8990)
);

AOI22xp5_ASAP7_75t_L g8991 ( 
.A1(n_8517),
.A2(n_5312),
.B1(n_5314),
.B2(n_5311),
.Y(n_8991)
);

INVx2_ASAP7_75t_L g8992 ( 
.A(n_8437),
.Y(n_8992)
);

AND2x4_ASAP7_75t_L g8993 ( 
.A(n_8602),
.B(n_5093),
.Y(n_8993)
);

INVx1_ASAP7_75t_L g8994 ( 
.A(n_8509),
.Y(n_8994)
);

NAND2xp5_ASAP7_75t_SL g8995 ( 
.A(n_8648),
.B(n_5317),
.Y(n_8995)
);

NAND2xp5_ASAP7_75t_SL g8996 ( 
.A(n_8648),
.B(n_5318),
.Y(n_8996)
);

INVx1_ASAP7_75t_L g8997 ( 
.A(n_8522),
.Y(n_8997)
);

AOI21xp5_ASAP7_75t_L g8998 ( 
.A1(n_8241),
.A2(n_5096),
.B(n_5095),
.Y(n_8998)
);

INVx1_ASAP7_75t_L g8999 ( 
.A(n_8533),
.Y(n_8999)
);

INVx2_ASAP7_75t_L g9000 ( 
.A(n_8439),
.Y(n_9000)
);

NOR2xp33_ASAP7_75t_L g9001 ( 
.A(n_8311),
.B(n_5319),
.Y(n_9001)
);

AOI22xp33_ASAP7_75t_L g9002 ( 
.A1(n_8391),
.A2(n_5104),
.B1(n_5105),
.B2(n_5097),
.Y(n_9002)
);

NAND2xp5_ASAP7_75t_SL g9003 ( 
.A(n_8685),
.B(n_5322),
.Y(n_9003)
);

BUFx6f_ASAP7_75t_L g9004 ( 
.A(n_8347),
.Y(n_9004)
);

NOR3xp33_ASAP7_75t_L g9005 ( 
.A(n_8265),
.B(n_8667),
.C(n_8372),
.Y(n_9005)
);

INVx1_ASAP7_75t_L g9006 ( 
.A(n_8539),
.Y(n_9006)
);

INVx2_ASAP7_75t_L g9007 ( 
.A(n_8441),
.Y(n_9007)
);

INVx1_ASAP7_75t_L g9008 ( 
.A(n_8540),
.Y(n_9008)
);

INVx1_ASAP7_75t_L g9009 ( 
.A(n_8544),
.Y(n_9009)
);

NAND2xp5_ASAP7_75t_L g9010 ( 
.A(n_8361),
.B(n_8687),
.Y(n_9010)
);

NAND2xp5_ASAP7_75t_L g9011 ( 
.A(n_8690),
.B(n_5106),
.Y(n_9011)
);

INVx1_ASAP7_75t_L g9012 ( 
.A(n_8545),
.Y(n_9012)
);

NAND2xp5_ASAP7_75t_SL g9013 ( 
.A(n_8685),
.B(n_8399),
.Y(n_9013)
);

INVx2_ASAP7_75t_L g9014 ( 
.A(n_8455),
.Y(n_9014)
);

INVx4_ASAP7_75t_L g9015 ( 
.A(n_8380),
.Y(n_9015)
);

INVx2_ASAP7_75t_L g9016 ( 
.A(n_8457),
.Y(n_9016)
);

INVx3_ASAP7_75t_L g9017 ( 
.A(n_8310),
.Y(n_9017)
);

INVx2_ASAP7_75t_L g9018 ( 
.A(n_8459),
.Y(n_9018)
);

INVx3_ASAP7_75t_L g9019 ( 
.A(n_8327),
.Y(n_9019)
);

INVx1_ASAP7_75t_L g9020 ( 
.A(n_8552),
.Y(n_9020)
);

AOI21xp5_ASAP7_75t_L g9021 ( 
.A1(n_8350),
.A2(n_5111),
.B(n_5110),
.Y(n_9021)
);

NOR2xp33_ASAP7_75t_L g9022 ( 
.A(n_8326),
.B(n_5323),
.Y(n_9022)
);

NAND2xp5_ASAP7_75t_L g9023 ( 
.A(n_8382),
.B(n_5112),
.Y(n_9023)
);

AOI22xp5_ASAP7_75t_L g9024 ( 
.A1(n_8232),
.A2(n_5330),
.B1(n_5331),
.B2(n_5326),
.Y(n_9024)
);

NAND2xp5_ASAP7_75t_L g9025 ( 
.A(n_8557),
.B(n_5118),
.Y(n_9025)
);

NAND2xp5_ASAP7_75t_SL g9026 ( 
.A(n_8425),
.B(n_8427),
.Y(n_9026)
);

NAND2xp5_ASAP7_75t_L g9027 ( 
.A(n_8561),
.B(n_5119),
.Y(n_9027)
);

NAND2xp5_ASAP7_75t_L g9028 ( 
.A(n_8566),
.B(n_5127),
.Y(n_9028)
);

INVx2_ASAP7_75t_L g9029 ( 
.A(n_8461),
.Y(n_9029)
);

AOI22xp5_ASAP7_75t_L g9030 ( 
.A1(n_8610),
.A2(n_5335),
.B1(n_5336),
.B2(n_5334),
.Y(n_9030)
);

INVx3_ASAP7_75t_L g9031 ( 
.A(n_8354),
.Y(n_9031)
);

INVx1_ASAP7_75t_L g9032 ( 
.A(n_8567),
.Y(n_9032)
);

NOR2xp33_ASAP7_75t_L g9033 ( 
.A(n_8369),
.B(n_5340),
.Y(n_9033)
);

INVx2_ASAP7_75t_L g9034 ( 
.A(n_8470),
.Y(n_9034)
);

OAI21xp5_ASAP7_75t_L g9035 ( 
.A1(n_8676),
.A2(n_5134),
.B(n_5133),
.Y(n_9035)
);

INVx1_ASAP7_75t_L g9036 ( 
.A(n_8568),
.Y(n_9036)
);

NAND2xp33_ASAP7_75t_L g9037 ( 
.A(n_8312),
.B(n_5343),
.Y(n_9037)
);

AOI22xp33_ASAP7_75t_L g9038 ( 
.A1(n_8626),
.A2(n_5138),
.B1(n_5139),
.B2(n_5135),
.Y(n_9038)
);

NOR3xp33_ASAP7_75t_L g9039 ( 
.A(n_8351),
.B(n_5162),
.C(n_5161),
.Y(n_9039)
);

INVx2_ASAP7_75t_L g9040 ( 
.A(n_8478),
.Y(n_9040)
);

INVx1_ASAP7_75t_L g9041 ( 
.A(n_8577),
.Y(n_9041)
);

BUFx6f_ASAP7_75t_SL g9042 ( 
.A(n_8235),
.Y(n_9042)
);

NAND2xp5_ASAP7_75t_L g9043 ( 
.A(n_8578),
.B(n_5172),
.Y(n_9043)
);

INVxp67_ASAP7_75t_L g9044 ( 
.A(n_8625),
.Y(n_9044)
);

NAND2xp5_ASAP7_75t_L g9045 ( 
.A(n_8479),
.B(n_5178),
.Y(n_9045)
);

NAND2xp5_ASAP7_75t_L g9046 ( 
.A(n_8483),
.B(n_5180),
.Y(n_9046)
);

INVx1_ASAP7_75t_L g9047 ( 
.A(n_8484),
.Y(n_9047)
);

INVx2_ASAP7_75t_L g9048 ( 
.A(n_8492),
.Y(n_9048)
);

AND2x2_ASAP7_75t_L g9049 ( 
.A(n_8628),
.B(n_5344),
.Y(n_9049)
);

INVx1_ASAP7_75t_L g9050 ( 
.A(n_8496),
.Y(n_9050)
);

INVx2_ASAP7_75t_SL g9051 ( 
.A(n_8353),
.Y(n_9051)
);

AOI22xp33_ASAP7_75t_L g9052 ( 
.A1(n_8374),
.A2(n_5186),
.B1(n_5189),
.B2(n_5185),
.Y(n_9052)
);

NAND2xp5_ASAP7_75t_L g9053 ( 
.A(n_8508),
.B(n_5209),
.Y(n_9053)
);

OR2x2_ASAP7_75t_SL g9054 ( 
.A(n_8188),
.B(n_5210),
.Y(n_9054)
);

NAND2xp5_ASAP7_75t_L g9055 ( 
.A(n_8511),
.B(n_5217),
.Y(n_9055)
);

NAND2x1_ASAP7_75t_L g9056 ( 
.A(n_8515),
.B(n_5218),
.Y(n_9056)
);

NAND2xp33_ASAP7_75t_L g9057 ( 
.A(n_8312),
.B(n_5347),
.Y(n_9057)
);

AND2x2_ASAP7_75t_L g9058 ( 
.A(n_8656),
.B(n_5349),
.Y(n_9058)
);

NOR2xp33_ASAP7_75t_L g9059 ( 
.A(n_8386),
.B(n_5350),
.Y(n_9059)
);

INVx1_ASAP7_75t_L g9060 ( 
.A(n_8528),
.Y(n_9060)
);

INVx2_ASAP7_75t_L g9061 ( 
.A(n_8530),
.Y(n_9061)
);

NOR2xp33_ASAP7_75t_L g9062 ( 
.A(n_8313),
.B(n_5351),
.Y(n_9062)
);

NAND2xp5_ASAP7_75t_L g9063 ( 
.A(n_8532),
.B(n_5220),
.Y(n_9063)
);

NAND2xp5_ASAP7_75t_L g9064 ( 
.A(n_8549),
.B(n_5222),
.Y(n_9064)
);

NAND2xp5_ASAP7_75t_L g9065 ( 
.A(n_8550),
.B(n_5223),
.Y(n_9065)
);

NOR2xp67_ASAP7_75t_L g9066 ( 
.A(n_8598),
.B(n_5),
.Y(n_9066)
);

NOR2xp33_ASAP7_75t_L g9067 ( 
.A(n_8325),
.B(n_5354),
.Y(n_9067)
);

AOI221xp5_ASAP7_75t_SL g9068 ( 
.A1(n_8686),
.A2(n_5245),
.B1(n_5249),
.B2(n_5240),
.C(n_5227),
.Y(n_9068)
);

INVx1_ASAP7_75t_L g9069 ( 
.A(n_8579),
.Y(n_9069)
);

NOR2xp67_ASAP7_75t_SL g9070 ( 
.A(n_8616),
.B(n_5355),
.Y(n_9070)
);

BUFx3_ASAP7_75t_L g9071 ( 
.A(n_8189),
.Y(n_9071)
);

INVx1_ASAP7_75t_L g9072 ( 
.A(n_8584),
.Y(n_9072)
);

INVx1_ASAP7_75t_L g9073 ( 
.A(n_8596),
.Y(n_9073)
);

INVxp67_ASAP7_75t_L g9074 ( 
.A(n_8541),
.Y(n_9074)
);

NAND2xp5_ASAP7_75t_SL g9075 ( 
.A(n_8468),
.B(n_5358),
.Y(n_9075)
);

OAI22xp5_ASAP7_75t_L g9076 ( 
.A1(n_8651),
.A2(n_5360),
.B1(n_5362),
.B2(n_5359),
.Y(n_9076)
);

INVx1_ASAP7_75t_L g9077 ( 
.A(n_8601),
.Y(n_9077)
);

NOR2xp67_ASAP7_75t_L g9078 ( 
.A(n_8604),
.B(n_6),
.Y(n_9078)
);

AND2x2_ASAP7_75t_L g9079 ( 
.A(n_8658),
.B(n_5363),
.Y(n_9079)
);

BUFx5_ASAP7_75t_L g9080 ( 
.A(n_8654),
.Y(n_9080)
);

OAI22xp5_ASAP7_75t_SL g9081 ( 
.A1(n_8632),
.A2(n_5370),
.B1(n_5373),
.B2(n_5365),
.Y(n_9081)
);

NAND2xp5_ASAP7_75t_SL g9082 ( 
.A(n_8482),
.B(n_5377),
.Y(n_9082)
);

NOR2xp33_ASAP7_75t_L g9083 ( 
.A(n_8296),
.B(n_5378),
.Y(n_9083)
);

NAND2xp5_ASAP7_75t_L g9084 ( 
.A(n_8580),
.B(n_5250),
.Y(n_9084)
);

INVx1_ASAP7_75t_L g9085 ( 
.A(n_8655),
.Y(n_9085)
);

INVx2_ASAP7_75t_L g9086 ( 
.A(n_8638),
.Y(n_9086)
);

INVx1_ASAP7_75t_L g9087 ( 
.A(n_8662),
.Y(n_9087)
);

INVx1_ASAP7_75t_L g9088 ( 
.A(n_8672),
.Y(n_9088)
);

INVx1_ASAP7_75t_L g9089 ( 
.A(n_8673),
.Y(n_9089)
);

INVx1_ASAP7_75t_L g9090 ( 
.A(n_8642),
.Y(n_9090)
);

AOI22xp5_ASAP7_75t_L g9091 ( 
.A1(n_8274),
.A2(n_5380),
.B1(n_5382),
.B2(n_5379),
.Y(n_9091)
);

INVx2_ASAP7_75t_L g9092 ( 
.A(n_8645),
.Y(n_9092)
);

INVx2_ASAP7_75t_L g9093 ( 
.A(n_8650),
.Y(n_9093)
);

NAND2xp5_ASAP7_75t_L g9094 ( 
.A(n_8487),
.B(n_5253),
.Y(n_9094)
);

INVx2_ASAP7_75t_SL g9095 ( 
.A(n_8541),
.Y(n_9095)
);

NAND2xp5_ASAP7_75t_SL g9096 ( 
.A(n_8665),
.B(n_5383),
.Y(n_9096)
);

INVx1_ASAP7_75t_L g9097 ( 
.A(n_8660),
.Y(n_9097)
);

NOR2xp67_ASAP7_75t_L g9098 ( 
.A(n_8671),
.B(n_6),
.Y(n_9098)
);

INVx1_ASAP7_75t_L g9099 ( 
.A(n_8661),
.Y(n_9099)
);

NOR2xp33_ASAP7_75t_L g9100 ( 
.A(n_8277),
.B(n_5385),
.Y(n_9100)
);

BUFx3_ASAP7_75t_L g9101 ( 
.A(n_8203),
.Y(n_9101)
);

NOR2xp33_ASAP7_75t_L g9102 ( 
.A(n_8293),
.B(n_5387),
.Y(n_9102)
);

INVx2_ASAP7_75t_L g9103 ( 
.A(n_8675),
.Y(n_9103)
);

INVxp67_ASAP7_75t_L g9104 ( 
.A(n_8546),
.Y(n_9104)
);

INVx1_ASAP7_75t_L g9105 ( 
.A(n_8486),
.Y(n_9105)
);

NAND2xp5_ASAP7_75t_L g9106 ( 
.A(n_8624),
.B(n_5255),
.Y(n_9106)
);

NAND2xp5_ASAP7_75t_SL g9107 ( 
.A(n_8534),
.B(n_5388),
.Y(n_9107)
);

AND2x2_ASAP7_75t_L g9108 ( 
.A(n_8451),
.B(n_5390),
.Y(n_9108)
);

INVx1_ASAP7_75t_L g9109 ( 
.A(n_8463),
.Y(n_9109)
);

NAND2xp5_ASAP7_75t_SL g9110 ( 
.A(n_8560),
.B(n_5391),
.Y(n_9110)
);

NAND2xp5_ASAP7_75t_L g9111 ( 
.A(n_8374),
.B(n_8527),
.Y(n_9111)
);

INVxp33_ASAP7_75t_L g9112 ( 
.A(n_8546),
.Y(n_9112)
);

NAND2xp33_ASAP7_75t_L g9113 ( 
.A(n_8527),
.B(n_5393),
.Y(n_9113)
);

INVx2_ASAP7_75t_L g9114 ( 
.A(n_8416),
.Y(n_9114)
);

NAND2xp5_ASAP7_75t_L g9115 ( 
.A(n_8376),
.B(n_8663),
.Y(n_9115)
);

NOR2xp33_ASAP7_75t_SL g9116 ( 
.A(n_8198),
.B(n_5397),
.Y(n_9116)
);

NAND2xp5_ASAP7_75t_SL g9117 ( 
.A(n_8555),
.B(n_5398),
.Y(n_9117)
);

INVx2_ASAP7_75t_L g9118 ( 
.A(n_8370),
.Y(n_9118)
);

INVx2_ASAP7_75t_L g9119 ( 
.A(n_8514),
.Y(n_9119)
);

NAND2xp5_ASAP7_75t_L g9120 ( 
.A(n_8663),
.B(n_5260),
.Y(n_9120)
);

AND2x2_ASAP7_75t_L g9121 ( 
.A(n_8519),
.B(n_5401),
.Y(n_9121)
);

AOI22xp5_ASAP7_75t_L g9122 ( 
.A1(n_8223),
.A2(n_5407),
.B1(n_5409),
.B2(n_5406),
.Y(n_9122)
);

OAI22xp5_ASAP7_75t_L g9123 ( 
.A1(n_8471),
.A2(n_8524),
.B1(n_8537),
.B2(n_8525),
.Y(n_9123)
);

NAND2xp5_ASAP7_75t_SL g9124 ( 
.A(n_8555),
.B(n_5413),
.Y(n_9124)
);

OAI22xp33_ASAP7_75t_L g9125 ( 
.A1(n_8634),
.A2(n_5419),
.B1(n_5420),
.B2(n_5418),
.Y(n_9125)
);

AOI22xp5_ASAP7_75t_L g9126 ( 
.A1(n_8664),
.A2(n_8643),
.B1(n_8419),
.B2(n_8647),
.Y(n_9126)
);

OR2x6_ASAP7_75t_L g9127 ( 
.A(n_8250),
.B(n_5261),
.Y(n_9127)
);

AOI22xp33_ASAP7_75t_SL g9128 ( 
.A1(n_8420),
.A2(n_5425),
.B1(n_5426),
.B2(n_5421),
.Y(n_9128)
);

INVx2_ASAP7_75t_L g9129 ( 
.A(n_8547),
.Y(n_9129)
);

NAND2xp5_ASAP7_75t_SL g9130 ( 
.A(n_8563),
.B(n_5428),
.Y(n_9130)
);

NAND2xp5_ASAP7_75t_L g9131 ( 
.A(n_8664),
.B(n_5267),
.Y(n_9131)
);

INVx1_ASAP7_75t_L g9132 ( 
.A(n_8466),
.Y(n_9132)
);

INVx2_ASAP7_75t_L g9133 ( 
.A(n_8538),
.Y(n_9133)
);

INVx1_ASAP7_75t_L g9134 ( 
.A(n_8556),
.Y(n_9134)
);

NOR2xp33_ASAP7_75t_L g9135 ( 
.A(n_8428),
.B(n_5432),
.Y(n_9135)
);

INVx1_ASAP7_75t_L g9136 ( 
.A(n_8588),
.Y(n_9136)
);

NAND2xp5_ASAP7_75t_L g9137 ( 
.A(n_8352),
.B(n_5270),
.Y(n_9137)
);

AOI22xp33_ASAP7_75t_L g9138 ( 
.A1(n_8587),
.A2(n_5273),
.B1(n_5275),
.B2(n_5272),
.Y(n_9138)
);

NAND2xp5_ASAP7_75t_L g9139 ( 
.A(n_8284),
.B(n_5278),
.Y(n_9139)
);

O2A1O1Ixp5_ASAP7_75t_L g9140 ( 
.A1(n_8586),
.A2(n_5284),
.B(n_5287),
.C(n_5279),
.Y(n_9140)
);

NAND2xp33_ASAP7_75t_L g9141 ( 
.A(n_8332),
.B(n_8563),
.Y(n_9141)
);

NAND2xp5_ASAP7_75t_L g9142 ( 
.A(n_8590),
.B(n_8593),
.Y(n_9142)
);

NAND2xp5_ASAP7_75t_SL g9143 ( 
.A(n_8575),
.B(n_5435),
.Y(n_9143)
);

NOR2x1_ASAP7_75t_L g9144 ( 
.A(n_8356),
.B(n_5291),
.Y(n_9144)
);

NAND2xp5_ASAP7_75t_L g9145 ( 
.A(n_8589),
.B(n_5293),
.Y(n_9145)
);

INVxp33_ASAP7_75t_L g9146 ( 
.A(n_8575),
.Y(n_9146)
);

INVx2_ASAP7_75t_L g9147 ( 
.A(n_8569),
.Y(n_9147)
);

AND2x4_ASAP7_75t_SL g9148 ( 
.A(n_8252),
.B(n_5308),
.Y(n_9148)
);

NOR2xp33_ASAP7_75t_SL g9149 ( 
.A(n_8681),
.B(n_8640),
.Y(n_9149)
);

AND2x2_ASAP7_75t_L g9150 ( 
.A(n_8272),
.B(n_5437),
.Y(n_9150)
);

INVx3_ASAP7_75t_L g9151 ( 
.A(n_8499),
.Y(n_9151)
);

INVxp67_ASAP7_75t_L g9152 ( 
.A(n_8594),
.Y(n_9152)
);

INVx2_ASAP7_75t_L g9153 ( 
.A(n_8594),
.Y(n_9153)
);

NAND2xp5_ASAP7_75t_L g9154 ( 
.A(n_8454),
.B(n_5309),
.Y(n_9154)
);

CKINVDCx5p33_ASAP7_75t_R g9155 ( 
.A(n_8659),
.Y(n_9155)
);

NAND2xp5_ASAP7_75t_SL g9156 ( 
.A(n_8616),
.B(n_5439),
.Y(n_9156)
);

NAND2xp5_ASAP7_75t_L g9157 ( 
.A(n_8636),
.B(n_5313),
.Y(n_9157)
);

INVx1_ASAP7_75t_L g9158 ( 
.A(n_8446),
.Y(n_9158)
);

NAND2xp5_ASAP7_75t_L g9159 ( 
.A(n_8603),
.B(n_5316),
.Y(n_9159)
);

INVx2_ASAP7_75t_L g9160 ( 
.A(n_8489),
.Y(n_9160)
);

INVx2_ASAP7_75t_SL g9161 ( 
.A(n_8513),
.Y(n_9161)
);

INVx1_ASAP7_75t_L g9162 ( 
.A(n_8531),
.Y(n_9162)
);

AOI21xp5_ASAP7_75t_L g9163 ( 
.A1(n_8398),
.A2(n_5327),
.B(n_5321),
.Y(n_9163)
);

INVx3_ASAP7_75t_L g9164 ( 
.A(n_8520),
.Y(n_9164)
);

NAND2xp5_ASAP7_75t_L g9165 ( 
.A(n_8476),
.B(n_8314),
.Y(n_9165)
);

NAND2xp5_ASAP7_75t_L g9166 ( 
.A(n_8359),
.B(n_8692),
.Y(n_9166)
);

NAND2xp5_ASAP7_75t_SL g9167 ( 
.A(n_8275),
.B(n_5440),
.Y(n_9167)
);

NAND2xp5_ASAP7_75t_L g9168 ( 
.A(n_8627),
.B(n_5328),
.Y(n_9168)
);

AOI221xp5_ASAP7_75t_L g9169 ( 
.A1(n_8197),
.A2(n_5353),
.B1(n_5356),
.B2(n_5346),
.C(n_5342),
.Y(n_9169)
);

INVx1_ASAP7_75t_L g9170 ( 
.A(n_8205),
.Y(n_9170)
);

NOR2xp33_ASAP7_75t_L g9171 ( 
.A(n_8207),
.B(n_5443),
.Y(n_9171)
);

NAND2xp5_ASAP7_75t_SL g9172 ( 
.A(n_8392),
.B(n_5444),
.Y(n_9172)
);

NAND2xp5_ASAP7_75t_L g9173 ( 
.A(n_8627),
.B(n_5357),
.Y(n_9173)
);

INVx1_ASAP7_75t_L g9174 ( 
.A(n_8587),
.Y(n_9174)
);

AOI22xp33_ASAP7_75t_L g9175 ( 
.A1(n_8600),
.A2(n_8408),
.B1(n_8385),
.B2(n_8435),
.Y(n_9175)
);

INVx4_ASAP7_75t_L g9176 ( 
.A(n_8210),
.Y(n_9176)
);

NAND2xp5_ASAP7_75t_SL g9177 ( 
.A(n_8426),
.B(n_5445),
.Y(n_9177)
);

NAND2xp5_ASAP7_75t_L g9178 ( 
.A(n_8600),
.B(n_5361),
.Y(n_9178)
);

INVx2_ASAP7_75t_L g9179 ( 
.A(n_8385),
.Y(n_9179)
);

AOI22xp5_ASAP7_75t_L g9180 ( 
.A1(n_8435),
.A2(n_5447),
.B1(n_5448),
.B2(n_5446),
.Y(n_9180)
);

NAND2xp5_ASAP7_75t_L g9181 ( 
.A(n_8477),
.B(n_5366),
.Y(n_9181)
);

INVx1_ASAP7_75t_L g9182 ( 
.A(n_8305),
.Y(n_9182)
);

BUFx3_ASAP7_75t_L g9183 ( 
.A(n_8214),
.Y(n_9183)
);

NAND2xp5_ASAP7_75t_L g9184 ( 
.A(n_8214),
.B(n_5375),
.Y(n_9184)
);

NAND2xp5_ASAP7_75t_L g9185 ( 
.A(n_8256),
.B(n_5381),
.Y(n_9185)
);

OAI22xp33_ASAP7_75t_L g9186 ( 
.A1(n_8308),
.A2(n_5453),
.B1(n_5456),
.B2(n_5451),
.Y(n_9186)
);

NAND2xp5_ASAP7_75t_L g9187 ( 
.A(n_8256),
.B(n_5384),
.Y(n_9187)
);

NAND2xp5_ASAP7_75t_L g9188 ( 
.A(n_8410),
.B(n_5386),
.Y(n_9188)
);

AND2x2_ASAP7_75t_L g9189 ( 
.A(n_8405),
.B(n_5462),
.Y(n_9189)
);

AOI22xp33_ASAP7_75t_L g9190 ( 
.A1(n_8516),
.A2(n_5402),
.B1(n_5411),
.B2(n_5389),
.Y(n_9190)
);

NAND2xp5_ASAP7_75t_L g9191 ( 
.A(n_8666),
.B(n_5422),
.Y(n_9191)
);

NAND2xp5_ASAP7_75t_SL g9192 ( 
.A(n_8242),
.B(n_5463),
.Y(n_9192)
);

NAND2xp5_ASAP7_75t_L g9193 ( 
.A(n_8317),
.B(n_5427),
.Y(n_9193)
);

BUFx6f_ASAP7_75t_L g9194 ( 
.A(n_8195),
.Y(n_9194)
);

OAI21xp5_ASAP7_75t_L g9195 ( 
.A1(n_8462),
.A2(n_5431),
.B(n_5430),
.Y(n_9195)
);

INVx1_ASAP7_75t_L g9196 ( 
.A(n_8183),
.Y(n_9196)
);

BUFx3_ASAP7_75t_L g9197 ( 
.A(n_8493),
.Y(n_9197)
);

NOR2xp33_ASAP7_75t_L g9198 ( 
.A(n_8204),
.B(n_5464),
.Y(n_9198)
);

NAND2xp5_ASAP7_75t_SL g9199 ( 
.A(n_8220),
.B(n_5465),
.Y(n_9199)
);

NAND2xp5_ASAP7_75t_L g9200 ( 
.A(n_8220),
.B(n_5433),
.Y(n_9200)
);

NAND2xp5_ASAP7_75t_L g9201 ( 
.A(n_8220),
.B(n_5449),
.Y(n_9201)
);

NOR2xp33_ASAP7_75t_SL g9202 ( 
.A(n_8185),
.B(n_5468),
.Y(n_9202)
);

AND2x4_ASAP7_75t_L g9203 ( 
.A(n_8362),
.B(n_5454),
.Y(n_9203)
);

INVx1_ASAP7_75t_L g9204 ( 
.A(n_8183),
.Y(n_9204)
);

AND2x2_ASAP7_75t_L g9205 ( 
.A(n_8301),
.B(n_5471),
.Y(n_9205)
);

INVx1_ASAP7_75t_L g9206 ( 
.A(n_8183),
.Y(n_9206)
);

NAND2xp5_ASAP7_75t_L g9207 ( 
.A(n_8220),
.B(n_5455),
.Y(n_9207)
);

NAND2xp5_ASAP7_75t_SL g9208 ( 
.A(n_8220),
.B(n_5472),
.Y(n_9208)
);

INVx1_ASAP7_75t_L g9209 ( 
.A(n_8183),
.Y(n_9209)
);

INVxp67_ASAP7_75t_L g9210 ( 
.A(n_8226),
.Y(n_9210)
);

INVx1_ASAP7_75t_L g9211 ( 
.A(n_8874),
.Y(n_9211)
);

BUFx3_ASAP7_75t_L g9212 ( 
.A(n_9197),
.Y(n_9212)
);

INVxp67_ASAP7_75t_L g9213 ( 
.A(n_8731),
.Y(n_9213)
);

AND2x2_ASAP7_75t_L g9214 ( 
.A(n_8701),
.B(n_5460),
.Y(n_9214)
);

NAND2xp5_ASAP7_75t_L g9215 ( 
.A(n_8694),
.B(n_5476),
.Y(n_9215)
);

AND2x4_ASAP7_75t_L g9216 ( 
.A(n_8699),
.B(n_5461),
.Y(n_9216)
);

INVx2_ASAP7_75t_L g9217 ( 
.A(n_8702),
.Y(n_9217)
);

BUFx6f_ASAP7_75t_L g9218 ( 
.A(n_9004),
.Y(n_9218)
);

INVx1_ASAP7_75t_L g9219 ( 
.A(n_8705),
.Y(n_9219)
);

INVx2_ASAP7_75t_L g9220 ( 
.A(n_8707),
.Y(n_9220)
);

AND2x2_ASAP7_75t_L g9221 ( 
.A(n_8767),
.B(n_5470),
.Y(n_9221)
);

AND2x2_ASAP7_75t_L g9222 ( 
.A(n_8757),
.B(n_5478),
.Y(n_9222)
);

INVx4_ASAP7_75t_L g9223 ( 
.A(n_9004),
.Y(n_9223)
);

BUFx6f_ASAP7_75t_L g9224 ( 
.A(n_8819),
.Y(n_9224)
);

BUFx3_ASAP7_75t_L g9225 ( 
.A(n_8911),
.Y(n_9225)
);

AND2x2_ASAP7_75t_L g9226 ( 
.A(n_9205),
.B(n_5480),
.Y(n_9226)
);

NAND2x1p5_ASAP7_75t_L g9227 ( 
.A(n_9015),
.B(n_8753),
.Y(n_9227)
);

BUFx2_ASAP7_75t_L g9228 ( 
.A(n_8761),
.Y(n_9228)
);

AND2x2_ASAP7_75t_L g9229 ( 
.A(n_8762),
.B(n_5485),
.Y(n_9229)
);

NAND2xp5_ASAP7_75t_L g9230 ( 
.A(n_8711),
.B(n_5479),
.Y(n_9230)
);

INVx3_ASAP7_75t_L g9231 ( 
.A(n_8855),
.Y(n_9231)
);

INVx1_ASAP7_75t_L g9232 ( 
.A(n_8726),
.Y(n_9232)
);

AND2x2_ASAP7_75t_L g9233 ( 
.A(n_8756),
.B(n_5487),
.Y(n_9233)
);

INVx3_ASAP7_75t_SL g9234 ( 
.A(n_9155),
.Y(n_9234)
);

AND2x6_ASAP7_75t_L g9235 ( 
.A(n_8698),
.B(n_5489),
.Y(n_9235)
);

BUFx3_ASAP7_75t_L g9236 ( 
.A(n_8911),
.Y(n_9236)
);

AND2x4_ASAP7_75t_L g9237 ( 
.A(n_8942),
.B(n_5491),
.Y(n_9237)
);

NAND2xp5_ASAP7_75t_SL g9238 ( 
.A(n_8858),
.B(n_5481),
.Y(n_9238)
);

BUFx6f_ASAP7_75t_L g9239 ( 
.A(n_8819),
.Y(n_9239)
);

BUFx6f_ASAP7_75t_L g9240 ( 
.A(n_8905),
.Y(n_9240)
);

NAND2xp5_ASAP7_75t_L g9241 ( 
.A(n_9198),
.B(n_5482),
.Y(n_9241)
);

AND2x4_ASAP7_75t_L g9242 ( 
.A(n_8725),
.B(n_5494),
.Y(n_9242)
);

INVx1_ASAP7_75t_L g9243 ( 
.A(n_8739),
.Y(n_9243)
);

NAND2xp5_ASAP7_75t_L g9244 ( 
.A(n_8776),
.B(n_5483),
.Y(n_9244)
);

BUFx6f_ASAP7_75t_L g9245 ( 
.A(n_8905),
.Y(n_9245)
);

INVx1_ASAP7_75t_L g9246 ( 
.A(n_8741),
.Y(n_9246)
);

INVxp67_ASAP7_75t_SL g9247 ( 
.A(n_8895),
.Y(n_9247)
);

INVx2_ASAP7_75t_L g9248 ( 
.A(n_8746),
.Y(n_9248)
);

INVx2_ASAP7_75t_SL g9249 ( 
.A(n_8870),
.Y(n_9249)
);

INVx1_ASAP7_75t_L g9250 ( 
.A(n_8747),
.Y(n_9250)
);

INVx3_ASAP7_75t_L g9251 ( 
.A(n_9151),
.Y(n_9251)
);

OR2x2_ASAP7_75t_L g9252 ( 
.A(n_8946),
.B(n_5500),
.Y(n_9252)
);

NAND2xp5_ASAP7_75t_L g9253 ( 
.A(n_8732),
.B(n_5492),
.Y(n_9253)
);

INVx2_ASAP7_75t_L g9254 ( 
.A(n_8749),
.Y(n_9254)
);

INVx2_ASAP7_75t_SL g9255 ( 
.A(n_8870),
.Y(n_9255)
);

NAND2xp5_ASAP7_75t_L g9256 ( 
.A(n_8988),
.B(n_5493),
.Y(n_9256)
);

NAND2xp5_ASAP7_75t_L g9257 ( 
.A(n_8801),
.B(n_5505),
.Y(n_9257)
);

AND2x2_ASAP7_75t_SL g9258 ( 
.A(n_8940),
.B(n_5514),
.Y(n_9258)
);

NAND2xp5_ASAP7_75t_L g9259 ( 
.A(n_8803),
.B(n_5516),
.Y(n_9259)
);

NAND2x1p5_ASAP7_75t_L g9260 ( 
.A(n_8805),
.B(n_5518),
.Y(n_9260)
);

BUFx6f_ASAP7_75t_L g9261 ( 
.A(n_9194),
.Y(n_9261)
);

OAI21xp5_ASAP7_75t_L g9262 ( 
.A1(n_8948),
.A2(n_5524),
.B(n_5521),
.Y(n_9262)
);

AND2x2_ASAP7_75t_L g9263 ( 
.A(n_8859),
.B(n_6),
.Y(n_9263)
);

AND2x4_ASAP7_75t_L g9264 ( 
.A(n_9164),
.B(n_303),
.Y(n_9264)
);

INVx1_ASAP7_75t_L g9265 ( 
.A(n_8758),
.Y(n_9265)
);

NAND2xp5_ASAP7_75t_SL g9266 ( 
.A(n_8869),
.B(n_303),
.Y(n_9266)
);

AND2x2_ASAP7_75t_L g9267 ( 
.A(n_8898),
.B(n_7),
.Y(n_9267)
);

AND2x4_ASAP7_75t_L g9268 ( 
.A(n_9161),
.B(n_304),
.Y(n_9268)
);

INVx1_ASAP7_75t_L g9269 ( 
.A(n_8771),
.Y(n_9269)
);

AND2x2_ASAP7_75t_L g9270 ( 
.A(n_9118),
.B(n_7),
.Y(n_9270)
);

INVx1_ASAP7_75t_L g9271 ( 
.A(n_8772),
.Y(n_9271)
);

BUFx3_ASAP7_75t_L g9272 ( 
.A(n_8864),
.Y(n_9272)
);

AND2x2_ASAP7_75t_L g9273 ( 
.A(n_9119),
.B(n_8),
.Y(n_9273)
);

AND2x2_ASAP7_75t_L g9274 ( 
.A(n_9129),
.B(n_8),
.Y(n_9274)
);

HB1xp67_ASAP7_75t_L g9275 ( 
.A(n_8829),
.Y(n_9275)
);

INVx1_ASAP7_75t_L g9276 ( 
.A(n_8786),
.Y(n_9276)
);

NAND2xp5_ASAP7_75t_SL g9277 ( 
.A(n_8695),
.B(n_305),
.Y(n_9277)
);

INVx2_ASAP7_75t_L g9278 ( 
.A(n_8798),
.Y(n_9278)
);

AND2x2_ASAP7_75t_L g9279 ( 
.A(n_9132),
.B(n_8),
.Y(n_9279)
);

HB1xp67_ASAP7_75t_L g9280 ( 
.A(n_9210),
.Y(n_9280)
);

NOR2xp33_ASAP7_75t_L g9281 ( 
.A(n_8811),
.B(n_305),
.Y(n_9281)
);

NAND2xp5_ASAP7_75t_L g9282 ( 
.A(n_8814),
.B(n_9),
.Y(n_9282)
);

AND2x2_ASAP7_75t_L g9283 ( 
.A(n_9108),
.B(n_9),
.Y(n_9283)
);

NAND2xp5_ASAP7_75t_L g9284 ( 
.A(n_8861),
.B(n_10),
.Y(n_9284)
);

INVx3_ASAP7_75t_L g9285 ( 
.A(n_9071),
.Y(n_9285)
);

AND2x2_ASAP7_75t_L g9286 ( 
.A(n_9121),
.B(n_9049),
.Y(n_9286)
);

HB1xp67_ASAP7_75t_L g9287 ( 
.A(n_9044),
.Y(n_9287)
);

AND2x2_ASAP7_75t_L g9288 ( 
.A(n_9058),
.B(n_10),
.Y(n_9288)
);

INVx3_ASAP7_75t_L g9289 ( 
.A(n_9101),
.Y(n_9289)
);

AND2x2_ASAP7_75t_L g9290 ( 
.A(n_9079),
.B(n_11),
.Y(n_9290)
);

NAND2xp5_ASAP7_75t_L g9291 ( 
.A(n_8912),
.B(n_11),
.Y(n_9291)
);

INVx1_ASAP7_75t_L g9292 ( 
.A(n_8812),
.Y(n_9292)
);

INVx3_ASAP7_75t_L g9293 ( 
.A(n_8854),
.Y(n_9293)
);

AND2x2_ASAP7_75t_L g9294 ( 
.A(n_9109),
.B(n_8849),
.Y(n_9294)
);

NAND2xp5_ASAP7_75t_L g9295 ( 
.A(n_8938),
.B(n_12),
.Y(n_9295)
);

INVxp67_ASAP7_75t_SL g9296 ( 
.A(n_8736),
.Y(n_9296)
);

HB1xp67_ASAP7_75t_L g9297 ( 
.A(n_8779),
.Y(n_9297)
);

BUFx3_ASAP7_75t_L g9298 ( 
.A(n_8882),
.Y(n_9298)
);

AND2x2_ASAP7_75t_L g9299 ( 
.A(n_8873),
.B(n_12),
.Y(n_9299)
);

INVx3_ASAP7_75t_SL g9300 ( 
.A(n_8787),
.Y(n_9300)
);

AND2x2_ASAP7_75t_L g9301 ( 
.A(n_8879),
.B(n_13),
.Y(n_9301)
);

NAND2xp5_ASAP7_75t_L g9302 ( 
.A(n_8703),
.B(n_13),
.Y(n_9302)
);

INVx2_ASAP7_75t_L g9303 ( 
.A(n_8815),
.Y(n_9303)
);

AND2x6_ASAP7_75t_L g9304 ( 
.A(n_9111),
.B(n_306),
.Y(n_9304)
);

INVx1_ASAP7_75t_L g9305 ( 
.A(n_8837),
.Y(n_9305)
);

OR2x2_ASAP7_75t_L g9306 ( 
.A(n_8838),
.B(n_307),
.Y(n_9306)
);

INVx1_ASAP7_75t_L g9307 ( 
.A(n_8848),
.Y(n_9307)
);

AND2x2_ASAP7_75t_L g9308 ( 
.A(n_8822),
.B(n_13),
.Y(n_9308)
);

INVx4_ASAP7_75t_L g9309 ( 
.A(n_9194),
.Y(n_9309)
);

HB1xp67_ASAP7_75t_L g9310 ( 
.A(n_8927),
.Y(n_9310)
);

INVx1_ASAP7_75t_L g9311 ( 
.A(n_8891),
.Y(n_9311)
);

AND2x2_ASAP7_75t_L g9312 ( 
.A(n_8908),
.B(n_14),
.Y(n_9312)
);

HB1xp67_ASAP7_75t_L g9313 ( 
.A(n_8980),
.Y(n_9313)
);

AND2x2_ASAP7_75t_L g9314 ( 
.A(n_8914),
.B(n_8951),
.Y(n_9314)
);

INVx1_ASAP7_75t_L g9315 ( 
.A(n_8697),
.Y(n_9315)
);

INVx1_ASAP7_75t_L g9316 ( 
.A(n_8700),
.Y(n_9316)
);

INVx3_ASAP7_75t_L g9317 ( 
.A(n_8979),
.Y(n_9317)
);

AND2x4_ASAP7_75t_L g9318 ( 
.A(n_8729),
.B(n_307),
.Y(n_9318)
);

INVx3_ASAP7_75t_L g9319 ( 
.A(n_9017),
.Y(n_9319)
);

INVx1_ASAP7_75t_SL g9320 ( 
.A(n_8959),
.Y(n_9320)
);

NAND2xp5_ASAP7_75t_L g9321 ( 
.A(n_8797),
.B(n_14),
.Y(n_9321)
);

INVx1_ASAP7_75t_L g9322 ( 
.A(n_8712),
.Y(n_9322)
);

AND2x2_ASAP7_75t_L g9323 ( 
.A(n_8952),
.B(n_14),
.Y(n_9323)
);

AND2x2_ASAP7_75t_L g9324 ( 
.A(n_8955),
.B(n_15),
.Y(n_9324)
);

NOR2xp33_ASAP7_75t_L g9325 ( 
.A(n_8717),
.B(n_308),
.Y(n_9325)
);

HB1xp67_ASAP7_75t_L g9326 ( 
.A(n_8899),
.Y(n_9326)
);

AND2x2_ASAP7_75t_L g9327 ( 
.A(n_8960),
.B(n_15),
.Y(n_9327)
);

AND2x2_ASAP7_75t_L g9328 ( 
.A(n_8943),
.B(n_15),
.Y(n_9328)
);

INVx1_ASAP7_75t_L g9329 ( 
.A(n_8713),
.Y(n_9329)
);

AND2x2_ASAP7_75t_L g9330 ( 
.A(n_8949),
.B(n_16),
.Y(n_9330)
);

NAND2xp5_ASAP7_75t_L g9331 ( 
.A(n_8775),
.B(n_16),
.Y(n_9331)
);

INVx1_ASAP7_75t_L g9332 ( 
.A(n_8715),
.Y(n_9332)
);

BUFx3_ASAP7_75t_L g9333 ( 
.A(n_8910),
.Y(n_9333)
);

INVx2_ASAP7_75t_SL g9334 ( 
.A(n_8777),
.Y(n_9334)
);

OAI21xp33_ASAP7_75t_L g9335 ( 
.A1(n_9195),
.A2(n_16),
.B(n_17),
.Y(n_9335)
);

NAND2xp5_ASAP7_75t_L g9336 ( 
.A(n_8795),
.B(n_17),
.Y(n_9336)
);

INVx3_ASAP7_75t_L g9337 ( 
.A(n_9019),
.Y(n_9337)
);

NAND2xp5_ASAP7_75t_L g9338 ( 
.A(n_9010),
.B(n_17),
.Y(n_9338)
);

NOR2x1p5_ASAP7_75t_L g9339 ( 
.A(n_9115),
.B(n_308),
.Y(n_9339)
);

NAND2xp5_ASAP7_75t_L g9340 ( 
.A(n_8989),
.B(n_18),
.Y(n_9340)
);

BUFx3_ASAP7_75t_L g9341 ( 
.A(n_8824),
.Y(n_9341)
);

INVxp67_ASAP7_75t_L g9342 ( 
.A(n_8734),
.Y(n_9342)
);

INVx1_ASAP7_75t_L g9343 ( 
.A(n_8719),
.Y(n_9343)
);

AND2x4_ASAP7_75t_L g9344 ( 
.A(n_9095),
.B(n_309),
.Y(n_9344)
);

AND2x2_ASAP7_75t_L g9345 ( 
.A(n_8958),
.B(n_18),
.Y(n_9345)
);

INVx2_ASAP7_75t_L g9346 ( 
.A(n_8961),
.Y(n_9346)
);

AND2x2_ASAP7_75t_L g9347 ( 
.A(n_8969),
.B(n_18),
.Y(n_9347)
);

HB1xp67_ASAP7_75t_L g9348 ( 
.A(n_9160),
.Y(n_9348)
);

INVx1_ASAP7_75t_L g9349 ( 
.A(n_8722),
.Y(n_9349)
);

NAND2xp5_ASAP7_75t_L g9350 ( 
.A(n_8929),
.B(n_19),
.Y(n_9350)
);

AND2x2_ASAP7_75t_L g9351 ( 
.A(n_8992),
.B(n_9000),
.Y(n_9351)
);

AND2x2_ASAP7_75t_L g9352 ( 
.A(n_9007),
.B(n_19),
.Y(n_9352)
);

OAI21xp5_ASAP7_75t_L g9353 ( 
.A1(n_9035),
.A2(n_19),
.B(n_20),
.Y(n_9353)
);

AND2x2_ASAP7_75t_L g9354 ( 
.A(n_9014),
.B(n_9016),
.Y(n_9354)
);

AND2x6_ASAP7_75t_L g9355 ( 
.A(n_9126),
.B(n_309),
.Y(n_9355)
);

AND2x2_ASAP7_75t_L g9356 ( 
.A(n_9018),
.B(n_20),
.Y(n_9356)
);

NAND2xp5_ASAP7_75t_SL g9357 ( 
.A(n_8708),
.B(n_310),
.Y(n_9357)
);

NAND2xp5_ASAP7_75t_L g9358 ( 
.A(n_8877),
.B(n_20),
.Y(n_9358)
);

INVx3_ASAP7_75t_L g9359 ( 
.A(n_9031),
.Y(n_9359)
);

NAND2xp5_ASAP7_75t_SL g9360 ( 
.A(n_8724),
.B(n_310),
.Y(n_9360)
);

INVx2_ASAP7_75t_L g9361 ( 
.A(n_9029),
.Y(n_9361)
);

NAND2xp5_ASAP7_75t_SL g9362 ( 
.A(n_8718),
.B(n_311),
.Y(n_9362)
);

AND2x4_ASAP7_75t_L g9363 ( 
.A(n_9074),
.B(n_311),
.Y(n_9363)
);

NOR2xp33_ASAP7_75t_SL g9364 ( 
.A(n_9176),
.B(n_21),
.Y(n_9364)
);

INVxp67_ASAP7_75t_L g9365 ( 
.A(n_8866),
.Y(n_9365)
);

INVx2_ASAP7_75t_L g9366 ( 
.A(n_9034),
.Y(n_9366)
);

INVx1_ASAP7_75t_L g9367 ( 
.A(n_8727),
.Y(n_9367)
);

INVx1_ASAP7_75t_L g9368 ( 
.A(n_8750),
.Y(n_9368)
);

NAND2xp5_ASAP7_75t_L g9369 ( 
.A(n_9001),
.B(n_21),
.Y(n_9369)
);

AOI22xp5_ASAP7_75t_L g9370 ( 
.A1(n_9005),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_9370)
);

INVx2_ASAP7_75t_SL g9371 ( 
.A(n_8808),
.Y(n_9371)
);

HB1xp67_ASAP7_75t_L g9372 ( 
.A(n_8886),
.Y(n_9372)
);

INVx1_ASAP7_75t_L g9373 ( 
.A(n_8755),
.Y(n_9373)
);

NAND2xp5_ASAP7_75t_L g9374 ( 
.A(n_9022),
.B(n_22),
.Y(n_9374)
);

INVx2_ASAP7_75t_L g9375 ( 
.A(n_9040),
.Y(n_9375)
);

CKINVDCx5p33_ASAP7_75t_R g9376 ( 
.A(n_8945),
.Y(n_9376)
);

NAND2xp5_ASAP7_75t_L g9377 ( 
.A(n_8714),
.B(n_22),
.Y(n_9377)
);

AND2x4_ASAP7_75t_SL g9378 ( 
.A(n_8818),
.B(n_312),
.Y(n_9378)
);

AND2x2_ASAP7_75t_L g9379 ( 
.A(n_9048),
.B(n_23),
.Y(n_9379)
);

NOR2xp33_ASAP7_75t_L g9380 ( 
.A(n_8865),
.B(n_312),
.Y(n_9380)
);

AND2x2_ASAP7_75t_L g9381 ( 
.A(n_9061),
.B(n_23),
.Y(n_9381)
);

NAND2xp5_ASAP7_75t_L g9382 ( 
.A(n_8799),
.B(n_24),
.Y(n_9382)
);

NAND2xp5_ASAP7_75t_L g9383 ( 
.A(n_8765),
.B(n_24),
.Y(n_9383)
);

INVx2_ASAP7_75t_L g9384 ( 
.A(n_9086),
.Y(n_9384)
);

INVx2_ASAP7_75t_L g9385 ( 
.A(n_9092),
.Y(n_9385)
);

INVx2_ASAP7_75t_L g9386 ( 
.A(n_9093),
.Y(n_9386)
);

BUFx6f_ASAP7_75t_L g9387 ( 
.A(n_8917),
.Y(n_9387)
);

INVx2_ASAP7_75t_L g9388 ( 
.A(n_9103),
.Y(n_9388)
);

BUFx6f_ASAP7_75t_L g9389 ( 
.A(n_8933),
.Y(n_9389)
);

INVx2_ASAP7_75t_SL g9390 ( 
.A(n_8937),
.Y(n_9390)
);

AND2x2_ASAP7_75t_L g9391 ( 
.A(n_8954),
.B(n_25),
.Y(n_9391)
);

NOR2xp33_ASAP7_75t_L g9392 ( 
.A(n_8710),
.B(n_313),
.Y(n_9392)
);

BUFx6f_ASAP7_75t_L g9393 ( 
.A(n_8941),
.Y(n_9393)
);

INVx1_ASAP7_75t_L g9394 ( 
.A(n_8759),
.Y(n_9394)
);

AND2x2_ASAP7_75t_L g9395 ( 
.A(n_9150),
.B(n_25),
.Y(n_9395)
);

AND2x2_ASAP7_75t_L g9396 ( 
.A(n_8902),
.B(n_25),
.Y(n_9396)
);

INVx1_ASAP7_75t_L g9397 ( 
.A(n_8774),
.Y(n_9397)
);

INVx2_ASAP7_75t_L g9398 ( 
.A(n_8791),
.Y(n_9398)
);

NAND2xp5_ASAP7_75t_L g9399 ( 
.A(n_8769),
.B(n_26),
.Y(n_9399)
);

AND2x2_ASAP7_75t_L g9400 ( 
.A(n_8903),
.B(n_26),
.Y(n_9400)
);

BUFx6f_ASAP7_75t_L g9401 ( 
.A(n_9153),
.Y(n_9401)
);

INVx1_ASAP7_75t_L g9402 ( 
.A(n_8806),
.Y(n_9402)
);

NAND2xp5_ASAP7_75t_L g9403 ( 
.A(n_8778),
.B(n_26),
.Y(n_9403)
);

NAND2xp5_ASAP7_75t_L g9404 ( 
.A(n_8781),
.B(n_27),
.Y(n_9404)
);

AND2x2_ASAP7_75t_L g9405 ( 
.A(n_8907),
.B(n_28),
.Y(n_9405)
);

INVxp67_ASAP7_75t_SL g9406 ( 
.A(n_8751),
.Y(n_9406)
);

INVx2_ASAP7_75t_L g9407 ( 
.A(n_8810),
.Y(n_9407)
);

AND2x2_ASAP7_75t_L g9408 ( 
.A(n_8913),
.B(n_28),
.Y(n_9408)
);

BUFx4_ASAP7_75t_SL g9409 ( 
.A(n_8971),
.Y(n_9409)
);

INVx1_ASAP7_75t_L g9410 ( 
.A(n_8831),
.Y(n_9410)
);

BUFx2_ASAP7_75t_L g9411 ( 
.A(n_9104),
.Y(n_9411)
);

AND2x2_ASAP7_75t_L g9412 ( 
.A(n_8922),
.B(n_28),
.Y(n_9412)
);

AND2x2_ASAP7_75t_L g9413 ( 
.A(n_8924),
.B(n_30),
.Y(n_9413)
);

INVx1_ASAP7_75t_L g9414 ( 
.A(n_8832),
.Y(n_9414)
);

NAND2xp5_ASAP7_75t_L g9415 ( 
.A(n_8782),
.B(n_30),
.Y(n_9415)
);

AND2x2_ASAP7_75t_SL g9416 ( 
.A(n_8981),
.B(n_313),
.Y(n_9416)
);

NAND2xp5_ASAP7_75t_SL g9417 ( 
.A(n_8709),
.B(n_314),
.Y(n_9417)
);

AND2x4_ASAP7_75t_L g9418 ( 
.A(n_9152),
.B(n_315),
.Y(n_9418)
);

INVx2_ASAP7_75t_L g9419 ( 
.A(n_8834),
.Y(n_9419)
);

NAND2xp5_ASAP7_75t_L g9420 ( 
.A(n_8784),
.B(n_30),
.Y(n_9420)
);

NAND2xp5_ASAP7_75t_L g9421 ( 
.A(n_8792),
.B(n_31),
.Y(n_9421)
);

OR2x2_ASAP7_75t_L g9422 ( 
.A(n_9200),
.B(n_316),
.Y(n_9422)
);

OAI21xp5_ASAP7_75t_L g9423 ( 
.A1(n_9199),
.A2(n_31),
.B(n_32),
.Y(n_9423)
);

NAND2xp5_ASAP7_75t_L g9424 ( 
.A(n_8816),
.B(n_31),
.Y(n_9424)
);

AND2x2_ASAP7_75t_L g9425 ( 
.A(n_9067),
.B(n_32),
.Y(n_9425)
);

HB1xp67_ASAP7_75t_L g9426 ( 
.A(n_9158),
.Y(n_9426)
);

AND2x2_ASAP7_75t_SL g9427 ( 
.A(n_8706),
.B(n_316),
.Y(n_9427)
);

AND2x2_ASAP7_75t_L g9428 ( 
.A(n_9083),
.B(n_32),
.Y(n_9428)
);

INVx1_ASAP7_75t_L g9429 ( 
.A(n_8835),
.Y(n_9429)
);

INVx1_ASAP7_75t_L g9430 ( 
.A(n_8844),
.Y(n_9430)
);

INVx1_ASAP7_75t_L g9431 ( 
.A(n_8868),
.Y(n_9431)
);

AND2x2_ASAP7_75t_L g9432 ( 
.A(n_9047),
.B(n_33),
.Y(n_9432)
);

INVx2_ASAP7_75t_L g9433 ( 
.A(n_8871),
.Y(n_9433)
);

AND2x2_ASAP7_75t_L g9434 ( 
.A(n_9050),
.B(n_9060),
.Y(n_9434)
);

HB1xp67_ASAP7_75t_L g9435 ( 
.A(n_9162),
.Y(n_9435)
);

BUFx3_ASAP7_75t_L g9436 ( 
.A(n_8963),
.Y(n_9436)
);

AND2x2_ASAP7_75t_L g9437 ( 
.A(n_9069),
.B(n_33),
.Y(n_9437)
);

NAND2xp5_ASAP7_75t_L g9438 ( 
.A(n_8820),
.B(n_33),
.Y(n_9438)
);

INVx2_ASAP7_75t_L g9439 ( 
.A(n_8885),
.Y(n_9439)
);

HB1xp67_ASAP7_75t_L g9440 ( 
.A(n_9170),
.Y(n_9440)
);

NAND2x1p5_ASAP7_75t_L g9441 ( 
.A(n_9013),
.B(n_317),
.Y(n_9441)
);

HB1xp67_ASAP7_75t_L g9442 ( 
.A(n_8964),
.Y(n_9442)
);

OAI21xp5_ASAP7_75t_L g9443 ( 
.A1(n_9208),
.A2(n_34),
.B(n_35),
.Y(n_9443)
);

BUFx6f_ASAP7_75t_L g9444 ( 
.A(n_9051),
.Y(n_9444)
);

AND2x2_ASAP7_75t_L g9445 ( 
.A(n_9072),
.B(n_34),
.Y(n_9445)
);

INVx2_ASAP7_75t_L g9446 ( 
.A(n_8887),
.Y(n_9446)
);

INVx1_ASAP7_75t_L g9447 ( 
.A(n_9196),
.Y(n_9447)
);

INVx2_ASAP7_75t_L g9448 ( 
.A(n_9204),
.Y(n_9448)
);

OR2x2_ASAP7_75t_L g9449 ( 
.A(n_9201),
.B(n_9207),
.Y(n_9449)
);

CKINVDCx5p33_ASAP7_75t_R g9450 ( 
.A(n_9042),
.Y(n_9450)
);

NAND2xp5_ASAP7_75t_L g9451 ( 
.A(n_8825),
.B(n_34),
.Y(n_9451)
);

INVx1_ASAP7_75t_L g9452 ( 
.A(n_9206),
.Y(n_9452)
);

AND2x2_ASAP7_75t_L g9453 ( 
.A(n_9073),
.B(n_35),
.Y(n_9453)
);

NAND2xp5_ASAP7_75t_L g9454 ( 
.A(n_8826),
.B(n_35),
.Y(n_9454)
);

AND2x2_ASAP7_75t_L g9455 ( 
.A(n_9077),
.B(n_9090),
.Y(n_9455)
);

INVx2_ASAP7_75t_L g9456 ( 
.A(n_9209),
.Y(n_9456)
);

BUFx3_ASAP7_75t_L g9457 ( 
.A(n_9147),
.Y(n_9457)
);

AND2x2_ASAP7_75t_L g9458 ( 
.A(n_9097),
.B(n_36),
.Y(n_9458)
);

INVx4_ASAP7_75t_L g9459 ( 
.A(n_8696),
.Y(n_9459)
);

INVx1_ASAP7_75t_L g9460 ( 
.A(n_8950),
.Y(n_9460)
);

NOR2xp67_ASAP7_75t_L g9461 ( 
.A(n_9142),
.B(n_36),
.Y(n_9461)
);

OAI21xp5_ASAP7_75t_L g9462 ( 
.A1(n_8693),
.A2(n_36),
.B(n_37),
.Y(n_9462)
);

NAND2xp5_ASAP7_75t_L g9463 ( 
.A(n_8828),
.B(n_37),
.Y(n_9463)
);

BUFx3_ASAP7_75t_L g9464 ( 
.A(n_9133),
.Y(n_9464)
);

NAND2xp5_ASAP7_75t_L g9465 ( 
.A(n_8833),
.B(n_37),
.Y(n_9465)
);

INVx2_ASAP7_75t_L g9466 ( 
.A(n_9099),
.Y(n_9466)
);

HB1xp67_ASAP7_75t_L g9467 ( 
.A(n_9026),
.Y(n_9467)
);

INVx1_ASAP7_75t_L g9468 ( 
.A(n_8965),
.Y(n_9468)
);

BUFx6f_ASAP7_75t_L g9469 ( 
.A(n_9203),
.Y(n_9469)
);

INVx1_ASAP7_75t_SL g9470 ( 
.A(n_8904),
.Y(n_9470)
);

OR2x2_ASAP7_75t_L g9471 ( 
.A(n_8836),
.B(n_317),
.Y(n_9471)
);

BUFx2_ASAP7_75t_L g9472 ( 
.A(n_8696),
.Y(n_9472)
);

AND2x4_ASAP7_75t_L g9473 ( 
.A(n_8735),
.B(n_318),
.Y(n_9473)
);

AND2x2_ASAP7_75t_L g9474 ( 
.A(n_9078),
.B(n_38),
.Y(n_9474)
);

BUFx4f_ASAP7_75t_L g9475 ( 
.A(n_8696),
.Y(n_9475)
);

INVx2_ASAP7_75t_L g9476 ( 
.A(n_8897),
.Y(n_9476)
);

AND2x2_ASAP7_75t_L g9477 ( 
.A(n_9098),
.B(n_8947),
.Y(n_9477)
);

INVx1_ASAP7_75t_SL g9478 ( 
.A(n_8977),
.Y(n_9478)
);

INVx2_ASAP7_75t_L g9479 ( 
.A(n_8973),
.Y(n_9479)
);

INVx4_ASAP7_75t_L g9480 ( 
.A(n_8783),
.Y(n_9480)
);

BUFx3_ASAP7_75t_L g9481 ( 
.A(n_9134),
.Y(n_9481)
);

AND2x2_ASAP7_75t_L g9482 ( 
.A(n_8827),
.B(n_38),
.Y(n_9482)
);

BUFx3_ASAP7_75t_L g9483 ( 
.A(n_9136),
.Y(n_9483)
);

INVx2_ASAP7_75t_L g9484 ( 
.A(n_8982),
.Y(n_9484)
);

AND3x1_ASAP7_75t_SL g9485 ( 
.A(n_8900),
.B(n_38),
.C(n_39),
.Y(n_9485)
);

INVx1_ASAP7_75t_L g9486 ( 
.A(n_8983),
.Y(n_9486)
);

AND2x2_ASAP7_75t_L g9487 ( 
.A(n_8862),
.B(n_39),
.Y(n_9487)
);

NAND2xp5_ASAP7_75t_L g9488 ( 
.A(n_8733),
.B(n_39),
.Y(n_9488)
);

NAND2xp5_ASAP7_75t_L g9489 ( 
.A(n_8985),
.B(n_40),
.Y(n_9489)
);

AND2x2_ASAP7_75t_L g9490 ( 
.A(n_9033),
.B(n_41),
.Y(n_9490)
);

NAND2xp5_ASAP7_75t_L g9491 ( 
.A(n_8987),
.B(n_41),
.Y(n_9491)
);

BUFx3_ASAP7_75t_L g9492 ( 
.A(n_9174),
.Y(n_9492)
);

AND2x4_ASAP7_75t_L g9493 ( 
.A(n_8843),
.B(n_318),
.Y(n_9493)
);

NAND2xp5_ASAP7_75t_L g9494 ( 
.A(n_9106),
.B(n_41),
.Y(n_9494)
);

INVx2_ASAP7_75t_L g9495 ( 
.A(n_8986),
.Y(n_9495)
);

NAND2xp5_ASAP7_75t_L g9496 ( 
.A(n_8742),
.B(n_42),
.Y(n_9496)
);

AND2x2_ASAP7_75t_L g9497 ( 
.A(n_9059),
.B(n_42),
.Y(n_9497)
);

INVx1_ASAP7_75t_L g9498 ( 
.A(n_8994),
.Y(n_9498)
);

INVx2_ASAP7_75t_L g9499 ( 
.A(n_8997),
.Y(n_9499)
);

INVxp33_ASAP7_75t_L g9500 ( 
.A(n_8728),
.Y(n_9500)
);

AND2x2_ASAP7_75t_L g9501 ( 
.A(n_9066),
.B(n_42),
.Y(n_9501)
);

AND2x2_ASAP7_75t_L g9502 ( 
.A(n_8853),
.B(n_43),
.Y(n_9502)
);

INVx1_ASAP7_75t_L g9503 ( 
.A(n_8999),
.Y(n_9503)
);

BUFx6f_ASAP7_75t_L g9504 ( 
.A(n_9183),
.Y(n_9504)
);

INVx3_ASAP7_75t_L g9505 ( 
.A(n_8766),
.Y(n_9505)
);

NAND2xp5_ASAP7_75t_L g9506 ( 
.A(n_9023),
.B(n_43),
.Y(n_9506)
);

AND2x2_ASAP7_75t_L g9507 ( 
.A(n_9062),
.B(n_44),
.Y(n_9507)
);

AND2x2_ASAP7_75t_L g9508 ( 
.A(n_8966),
.B(n_44),
.Y(n_9508)
);

INVxp67_ASAP7_75t_L g9509 ( 
.A(n_9171),
.Y(n_9509)
);

NAND2xp5_ASAP7_75t_L g9510 ( 
.A(n_9084),
.B(n_44),
.Y(n_9510)
);

INVx1_ASAP7_75t_L g9511 ( 
.A(n_9006),
.Y(n_9511)
);

BUFx3_ASAP7_75t_L g9512 ( 
.A(n_9179),
.Y(n_9512)
);

BUFx2_ASAP7_75t_L g9513 ( 
.A(n_9166),
.Y(n_9513)
);

CKINVDCx5p33_ASAP7_75t_R g9514 ( 
.A(n_8716),
.Y(n_9514)
);

INVx2_ASAP7_75t_L g9515 ( 
.A(n_9008),
.Y(n_9515)
);

AND2x2_ASAP7_75t_L g9516 ( 
.A(n_8888),
.B(n_45),
.Y(n_9516)
);

CKINVDCx5p33_ASAP7_75t_R g9517 ( 
.A(n_8957),
.Y(n_9517)
);

AND2x2_ASAP7_75t_L g9518 ( 
.A(n_9157),
.B(n_45),
.Y(n_9518)
);

INVx2_ASAP7_75t_L g9519 ( 
.A(n_9009),
.Y(n_9519)
);

INVx3_ASAP7_75t_L g9520 ( 
.A(n_8993),
.Y(n_9520)
);

AND2x2_ASAP7_75t_L g9521 ( 
.A(n_9002),
.B(n_45),
.Y(n_9521)
);

INVx2_ASAP7_75t_L g9522 ( 
.A(n_9012),
.Y(n_9522)
);

AND2x2_ASAP7_75t_L g9523 ( 
.A(n_9100),
.B(n_46),
.Y(n_9523)
);

AND2x2_ASAP7_75t_L g9524 ( 
.A(n_9102),
.B(n_46),
.Y(n_9524)
);

NAND2xp5_ASAP7_75t_L g9525 ( 
.A(n_8978),
.B(n_46),
.Y(n_9525)
);

INVx4_ASAP7_75t_L g9526 ( 
.A(n_8738),
.Y(n_9526)
);

AND2x2_ASAP7_75t_SL g9527 ( 
.A(n_9039),
.B(n_319),
.Y(n_9527)
);

INVx3_ASAP7_75t_L g9528 ( 
.A(n_8972),
.Y(n_9528)
);

AND2x6_ASAP7_75t_L g9529 ( 
.A(n_8745),
.B(n_320),
.Y(n_9529)
);

INVx1_ASAP7_75t_L g9530 ( 
.A(n_9020),
.Y(n_9530)
);

NAND2xp5_ASAP7_75t_L g9531 ( 
.A(n_8720),
.B(n_47),
.Y(n_9531)
);

NOR2xp33_ASAP7_75t_L g9532 ( 
.A(n_8823),
.B(n_321),
.Y(n_9532)
);

INVx4_ASAP7_75t_L g9533 ( 
.A(n_8738),
.Y(n_9533)
);

BUFx3_ASAP7_75t_L g9534 ( 
.A(n_9182),
.Y(n_9534)
);

HB1xp67_ASAP7_75t_L g9535 ( 
.A(n_9112),
.Y(n_9535)
);

INVx3_ASAP7_75t_L g9536 ( 
.A(n_9056),
.Y(n_9536)
);

NAND2xp5_ASAP7_75t_L g9537 ( 
.A(n_9135),
.B(n_47),
.Y(n_9537)
);

AND2x2_ASAP7_75t_SL g9538 ( 
.A(n_8704),
.B(n_322),
.Y(n_9538)
);

NAND2xp5_ASAP7_75t_L g9539 ( 
.A(n_8935),
.B(n_48),
.Y(n_9539)
);

AND2x2_ASAP7_75t_L g9540 ( 
.A(n_9052),
.B(n_8990),
.Y(n_9540)
);

INVx1_ASAP7_75t_L g9541 ( 
.A(n_9032),
.Y(n_9541)
);

NAND2xp5_ASAP7_75t_L g9542 ( 
.A(n_8744),
.B(n_48),
.Y(n_9542)
);

INVx2_ASAP7_75t_L g9543 ( 
.A(n_9036),
.Y(n_9543)
);

INVx2_ASAP7_75t_L g9544 ( 
.A(n_9041),
.Y(n_9544)
);

INVx1_ASAP7_75t_SL g9545 ( 
.A(n_9146),
.Y(n_9545)
);

NOR2xp67_ASAP7_75t_L g9546 ( 
.A(n_8909),
.B(n_8796),
.Y(n_9546)
);

NAND2xp5_ASAP7_75t_SL g9547 ( 
.A(n_8847),
.B(n_322),
.Y(n_9547)
);

INVx4_ASAP7_75t_L g9548 ( 
.A(n_9127),
.Y(n_9548)
);

AND2x4_ASAP7_75t_SL g9549 ( 
.A(n_9127),
.B(n_323),
.Y(n_9549)
);

INVx2_ASAP7_75t_L g9550 ( 
.A(n_9085),
.Y(n_9550)
);

INVx2_ASAP7_75t_SL g9551 ( 
.A(n_8956),
.Y(n_9551)
);

INVx1_ASAP7_75t_L g9552 ( 
.A(n_9087),
.Y(n_9552)
);

NAND2xp5_ASAP7_75t_L g9553 ( 
.A(n_9154),
.B(n_48),
.Y(n_9553)
);

HB1xp67_ASAP7_75t_L g9554 ( 
.A(n_8721),
.Y(n_9554)
);

AND2x2_ASAP7_75t_L g9555 ( 
.A(n_9038),
.B(n_49),
.Y(n_9555)
);

AND2x2_ASAP7_75t_L g9556 ( 
.A(n_9120),
.B(n_49),
.Y(n_9556)
);

INVx2_ASAP7_75t_L g9557 ( 
.A(n_9088),
.Y(n_9557)
);

NOR2xp33_ASAP7_75t_L g9558 ( 
.A(n_8863),
.B(n_8740),
.Y(n_9558)
);

INVx1_ASAP7_75t_L g9559 ( 
.A(n_9089),
.Y(n_9559)
);

INVx1_ASAP7_75t_L g9560 ( 
.A(n_9025),
.Y(n_9560)
);

AND2x2_ASAP7_75t_L g9561 ( 
.A(n_9131),
.B(n_49),
.Y(n_9561)
);

AND2x2_ASAP7_75t_L g9562 ( 
.A(n_8970),
.B(n_50),
.Y(n_9562)
);

AND2x2_ASAP7_75t_L g9563 ( 
.A(n_9138),
.B(n_50),
.Y(n_9563)
);

AND2x4_ASAP7_75t_SL g9564 ( 
.A(n_9175),
.B(n_323),
.Y(n_9564)
);

HB1xp67_ASAP7_75t_L g9565 ( 
.A(n_9165),
.Y(n_9565)
);

NAND2xp5_ASAP7_75t_L g9566 ( 
.A(n_8921),
.B(n_50),
.Y(n_9566)
);

INVx2_ASAP7_75t_L g9567 ( 
.A(n_8930),
.Y(n_9567)
);

INVx1_ASAP7_75t_L g9568 ( 
.A(n_9027),
.Y(n_9568)
);

INVx3_ASAP7_75t_L g9569 ( 
.A(n_8842),
.Y(n_9569)
);

NAND2xp5_ASAP7_75t_L g9570 ( 
.A(n_8790),
.B(n_51),
.Y(n_9570)
);

AND2x2_ASAP7_75t_L g9571 ( 
.A(n_9168),
.B(n_51),
.Y(n_9571)
);

INVx1_ASAP7_75t_L g9572 ( 
.A(n_9028),
.Y(n_9572)
);

NAND2xp5_ASAP7_75t_L g9573 ( 
.A(n_8730),
.B(n_51),
.Y(n_9573)
);

INVx1_ASAP7_75t_L g9574 ( 
.A(n_9043),
.Y(n_9574)
);

AND2x2_ASAP7_75t_L g9575 ( 
.A(n_9173),
.B(n_52),
.Y(n_9575)
);

AND2x2_ASAP7_75t_L g9576 ( 
.A(n_9128),
.B(n_52),
.Y(n_9576)
);

INVx3_ASAP7_75t_L g9577 ( 
.A(n_8894),
.Y(n_9577)
);

INVxp67_ASAP7_75t_L g9578 ( 
.A(n_9202),
.Y(n_9578)
);

NAND2xp5_ASAP7_75t_L g9579 ( 
.A(n_9139),
.B(n_52),
.Y(n_9579)
);

NAND2x1p5_ASAP7_75t_L g9580 ( 
.A(n_8931),
.B(n_324),
.Y(n_9580)
);

INVx2_ASAP7_75t_L g9581 ( 
.A(n_8930),
.Y(n_9581)
);

NAND2xp5_ASAP7_75t_L g9582 ( 
.A(n_8804),
.B(n_53),
.Y(n_9582)
);

INVx1_ASAP7_75t_L g9583 ( 
.A(n_9045),
.Y(n_9583)
);

INVx1_ASAP7_75t_L g9584 ( 
.A(n_9046),
.Y(n_9584)
);

NOR2xp67_ASAP7_75t_L g9585 ( 
.A(n_8743),
.B(n_53),
.Y(n_9585)
);

OR2x2_ASAP7_75t_L g9586 ( 
.A(n_8944),
.B(n_9011),
.Y(n_9586)
);

NOR2xp33_ASAP7_75t_L g9587 ( 
.A(n_8932),
.B(n_324),
.Y(n_9587)
);

NAND2xp5_ASAP7_75t_L g9588 ( 
.A(n_8807),
.B(n_54),
.Y(n_9588)
);

OAI21x1_ASAP7_75t_L g9589 ( 
.A1(n_9114),
.A2(n_54),
.B(n_55),
.Y(n_9589)
);

INVx3_ASAP7_75t_L g9590 ( 
.A(n_8800),
.Y(n_9590)
);

OAI21x1_ASAP7_75t_L g9591 ( 
.A1(n_9105),
.A2(n_55),
.B(n_56),
.Y(n_9591)
);

HB1xp67_ASAP7_75t_L g9592 ( 
.A(n_9123),
.Y(n_9592)
);

AND2x2_ASAP7_75t_L g9593 ( 
.A(n_9178),
.B(n_55),
.Y(n_9593)
);

AND2x2_ASAP7_75t_L g9594 ( 
.A(n_8872),
.B(n_56),
.Y(n_9594)
);

AND2x2_ASAP7_75t_L g9595 ( 
.A(n_8896),
.B(n_56),
.Y(n_9595)
);

BUFx6f_ASAP7_75t_L g9596 ( 
.A(n_8813),
.Y(n_9596)
);

INVx2_ASAP7_75t_L g9597 ( 
.A(n_8930),
.Y(n_9597)
);

NAND2xp5_ASAP7_75t_L g9598 ( 
.A(n_8839),
.B(n_57),
.Y(n_9598)
);

AND2x2_ASAP7_75t_L g9599 ( 
.A(n_9188),
.B(n_57),
.Y(n_9599)
);

INVx2_ASAP7_75t_L g9600 ( 
.A(n_8930),
.Y(n_9600)
);

NAND2xp5_ASAP7_75t_L g9601 ( 
.A(n_8840),
.B(n_57),
.Y(n_9601)
);

AND2x2_ASAP7_75t_L g9602 ( 
.A(n_8919),
.B(n_58),
.Y(n_9602)
);

AND2x2_ASAP7_75t_L g9603 ( 
.A(n_8920),
.B(n_58),
.Y(n_9603)
);

INVx2_ASAP7_75t_SL g9604 ( 
.A(n_8918),
.Y(n_9604)
);

INVx2_ASAP7_75t_SL g9605 ( 
.A(n_9117),
.Y(n_9605)
);

AND2x6_ASAP7_75t_L g9606 ( 
.A(n_8737),
.B(n_325),
.Y(n_9606)
);

INVx1_ASAP7_75t_L g9607 ( 
.A(n_9053),
.Y(n_9607)
);

INVx2_ASAP7_75t_L g9608 ( 
.A(n_9080),
.Y(n_9608)
);

AND2x2_ASAP7_75t_L g9609 ( 
.A(n_9145),
.B(n_59),
.Y(n_9609)
);

INVx3_ASAP7_75t_L g9610 ( 
.A(n_9148),
.Y(n_9610)
);

AND2x2_ASAP7_75t_L g9611 ( 
.A(n_8860),
.B(n_59),
.Y(n_9611)
);

INVx4_ASAP7_75t_L g9612 ( 
.A(n_8768),
.Y(n_9612)
);

OR2x2_ASAP7_75t_L g9613 ( 
.A(n_8845),
.B(n_325),
.Y(n_9613)
);

NAND2xp5_ASAP7_75t_L g9614 ( 
.A(n_8850),
.B(n_59),
.Y(n_9614)
);

INVx2_ASAP7_75t_L g9615 ( 
.A(n_9080),
.Y(n_9615)
);

BUFx6f_ASAP7_75t_L g9616 ( 
.A(n_8817),
.Y(n_9616)
);

AND2x2_ASAP7_75t_L g9617 ( 
.A(n_8821),
.B(n_60),
.Y(n_9617)
);

AND2x2_ASAP7_75t_L g9618 ( 
.A(n_9144),
.B(n_60),
.Y(n_9618)
);

AND2x2_ASAP7_75t_L g9619 ( 
.A(n_9094),
.B(n_60),
.Y(n_9619)
);

AND2x2_ASAP7_75t_L g9620 ( 
.A(n_8770),
.B(n_61),
.Y(n_9620)
);

INVx3_ASAP7_75t_L g9621 ( 
.A(n_9080),
.Y(n_9621)
);

INVx1_ASAP7_75t_SL g9622 ( 
.A(n_8890),
.Y(n_9622)
);

NAND2xp5_ASAP7_75t_L g9623 ( 
.A(n_8852),
.B(n_61),
.Y(n_9623)
);

AND2x4_ASAP7_75t_SL g9624 ( 
.A(n_9189),
.B(n_326),
.Y(n_9624)
);

OAI21xp5_ASAP7_75t_L g9625 ( 
.A1(n_8752),
.A2(n_61),
.B(n_62),
.Y(n_9625)
);

HB1xp67_ASAP7_75t_L g9626 ( 
.A(n_8892),
.Y(n_9626)
);

INVx1_ASAP7_75t_L g9627 ( 
.A(n_9055),
.Y(n_9627)
);

AND2x4_ASAP7_75t_L g9628 ( 
.A(n_8748),
.B(n_326),
.Y(n_9628)
);

NAND2xp5_ASAP7_75t_L g9629 ( 
.A(n_8856),
.B(n_62),
.Y(n_9629)
);

INVx2_ASAP7_75t_L g9630 ( 
.A(n_9080),
.Y(n_9630)
);

NAND2xp5_ASAP7_75t_L g9631 ( 
.A(n_8867),
.B(n_62),
.Y(n_9631)
);

AND2x2_ASAP7_75t_L g9632 ( 
.A(n_8857),
.B(n_63),
.Y(n_9632)
);

NAND2xp5_ASAP7_75t_L g9633 ( 
.A(n_8876),
.B(n_63),
.Y(n_9633)
);

INVx3_ASAP7_75t_L g9634 ( 
.A(n_8768),
.Y(n_9634)
);

INVx1_ASAP7_75t_L g9635 ( 
.A(n_9063),
.Y(n_9635)
);

INVx1_ASAP7_75t_L g9636 ( 
.A(n_9064),
.Y(n_9636)
);

INVx2_ASAP7_75t_L g9637 ( 
.A(n_9065),
.Y(n_9637)
);

INVx2_ASAP7_75t_L g9638 ( 
.A(n_8893),
.Y(n_9638)
);

AND2x2_ASAP7_75t_L g9639 ( 
.A(n_9159),
.B(n_63),
.Y(n_9639)
);

BUFx3_ASAP7_75t_L g9640 ( 
.A(n_9054),
.Y(n_9640)
);

AND2x2_ASAP7_75t_SL g9641 ( 
.A(n_9113),
.B(n_327),
.Y(n_9641)
);

AND2x2_ASAP7_75t_L g9642 ( 
.A(n_9184),
.B(n_64),
.Y(n_9642)
);

INVx1_ASAP7_75t_L g9643 ( 
.A(n_8901),
.Y(n_9643)
);

INVx1_ASAP7_75t_L g9644 ( 
.A(n_8906),
.Y(n_9644)
);

AOI22xp5_ASAP7_75t_L g9645 ( 
.A1(n_8851),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_9645)
);

INVx1_ASAP7_75t_L g9646 ( 
.A(n_8916),
.Y(n_9646)
);

NAND2xp5_ASAP7_75t_L g9647 ( 
.A(n_8878),
.B(n_8880),
.Y(n_9647)
);

HB1xp67_ASAP7_75t_L g9648 ( 
.A(n_8923),
.Y(n_9648)
);

AND2x2_ASAP7_75t_L g9649 ( 
.A(n_9185),
.B(n_64),
.Y(n_9649)
);

INVx2_ASAP7_75t_L g9650 ( 
.A(n_8926),
.Y(n_9650)
);

INVx1_ASAP7_75t_L g9651 ( 
.A(n_8928),
.Y(n_9651)
);

INVx3_ASAP7_75t_L g9652 ( 
.A(n_8768),
.Y(n_9652)
);

INVx3_ASAP7_75t_L g9653 ( 
.A(n_8936),
.Y(n_9653)
);

INVx1_ASAP7_75t_L g9654 ( 
.A(n_8967),
.Y(n_9654)
);

INVx1_ASAP7_75t_L g9655 ( 
.A(n_8968),
.Y(n_9655)
);

OAI21xp5_ASAP7_75t_L g9656 ( 
.A1(n_8830),
.A2(n_65),
.B(n_66),
.Y(n_9656)
);

NAND2xp5_ASAP7_75t_L g9657 ( 
.A(n_8881),
.B(n_65),
.Y(n_9657)
);

NAND2xp5_ASAP7_75t_L g9658 ( 
.A(n_8884),
.B(n_66),
.Y(n_9658)
);

BUFx3_ASAP7_75t_L g9659 ( 
.A(n_9181),
.Y(n_9659)
);

INVx3_ASAP7_75t_L g9660 ( 
.A(n_8889),
.Y(n_9660)
);

HB1xp67_ASAP7_75t_L g9661 ( 
.A(n_8760),
.Y(n_9661)
);

INVx1_ASAP7_75t_L g9662 ( 
.A(n_8998),
.Y(n_9662)
);

AND2x2_ASAP7_75t_L g9663 ( 
.A(n_9187),
.B(n_9030),
.Y(n_9663)
);

NAND2xp5_ASAP7_75t_L g9664 ( 
.A(n_8953),
.B(n_67),
.Y(n_9664)
);

INVx1_ASAP7_75t_L g9665 ( 
.A(n_8754),
.Y(n_9665)
);

BUFx6f_ASAP7_75t_L g9666 ( 
.A(n_9124),
.Y(n_9666)
);

NAND2xp5_ASAP7_75t_L g9667 ( 
.A(n_9068),
.B(n_8974),
.Y(n_9667)
);

AND2x2_ASAP7_75t_L g9668 ( 
.A(n_8763),
.B(n_67),
.Y(n_9668)
);

INVx2_ASAP7_75t_L g9669 ( 
.A(n_9140),
.Y(n_9669)
);

NAND2xp5_ASAP7_75t_L g9670 ( 
.A(n_8723),
.B(n_9167),
.Y(n_9670)
);

INVx3_ASAP7_75t_SL g9671 ( 
.A(n_9156),
.Y(n_9671)
);

NAND2xp5_ASAP7_75t_L g9672 ( 
.A(n_9091),
.B(n_68),
.Y(n_9672)
);

NAND2xp5_ASAP7_75t_L g9673 ( 
.A(n_9125),
.B(n_68),
.Y(n_9673)
);

NAND2xp5_ASAP7_75t_SL g9674 ( 
.A(n_8875),
.B(n_327),
.Y(n_9674)
);

INVx1_ASAP7_75t_L g9675 ( 
.A(n_9021),
.Y(n_9675)
);

NAND2xp5_ASAP7_75t_L g9676 ( 
.A(n_9137),
.B(n_68),
.Y(n_9676)
);

AND2x2_ASAP7_75t_L g9677 ( 
.A(n_8780),
.B(n_69),
.Y(n_9677)
);

INVx2_ASAP7_75t_L g9678 ( 
.A(n_9096),
.Y(n_9678)
);

INVxp67_ASAP7_75t_L g9679 ( 
.A(n_9191),
.Y(n_9679)
);

INVx1_ASAP7_75t_L g9680 ( 
.A(n_9163),
.Y(n_9680)
);

INVx2_ASAP7_75t_SL g9681 ( 
.A(n_9130),
.Y(n_9681)
);

BUFx2_ASAP7_75t_L g9682 ( 
.A(n_8939),
.Y(n_9682)
);

AND2x4_ASAP7_75t_L g9683 ( 
.A(n_9143),
.B(n_328),
.Y(n_9683)
);

NAND2xp5_ASAP7_75t_L g9684 ( 
.A(n_8793),
.B(n_9122),
.Y(n_9684)
);

INVx2_ASAP7_75t_L g9685 ( 
.A(n_8975),
.Y(n_9685)
);

NAND2xp5_ASAP7_75t_L g9686 ( 
.A(n_9076),
.B(n_70),
.Y(n_9686)
);

NAND2xp5_ASAP7_75t_L g9687 ( 
.A(n_8764),
.B(n_70),
.Y(n_9687)
);

NOR2xp33_ASAP7_75t_L g9688 ( 
.A(n_8788),
.B(n_328),
.Y(n_9688)
);

OAI21xp5_ASAP7_75t_L g9689 ( 
.A1(n_8785),
.A2(n_70),
.B(n_71),
.Y(n_9689)
);

AND2x2_ASAP7_75t_L g9690 ( 
.A(n_8794),
.B(n_71),
.Y(n_9690)
);

INVx2_ASAP7_75t_L g9691 ( 
.A(n_8976),
.Y(n_9691)
);

BUFx6f_ASAP7_75t_L g9692 ( 
.A(n_8995),
.Y(n_9692)
);

AND2x4_ASAP7_75t_L g9693 ( 
.A(n_8996),
.B(n_329),
.Y(n_9693)
);

INVx1_ASAP7_75t_L g9694 ( 
.A(n_8883),
.Y(n_9694)
);

INVx1_ASAP7_75t_L g9695 ( 
.A(n_8925),
.Y(n_9695)
);

AND2x2_ASAP7_75t_L g9696 ( 
.A(n_8802),
.B(n_8841),
.Y(n_9696)
);

NAND2xp5_ASAP7_75t_L g9697 ( 
.A(n_8991),
.B(n_71),
.Y(n_9697)
);

AND2x2_ASAP7_75t_L g9698 ( 
.A(n_8846),
.B(n_72),
.Y(n_9698)
);

NAND2xp5_ASAP7_75t_L g9699 ( 
.A(n_9003),
.B(n_72),
.Y(n_9699)
);

AND2x2_ASAP7_75t_L g9700 ( 
.A(n_9193),
.B(n_73),
.Y(n_9700)
);

AND2x2_ASAP7_75t_L g9701 ( 
.A(n_9024),
.B(n_73),
.Y(n_9701)
);

NAND2xp5_ASAP7_75t_L g9702 ( 
.A(n_9186),
.B(n_74),
.Y(n_9702)
);

AND2x2_ASAP7_75t_L g9703 ( 
.A(n_9180),
.B(n_74),
.Y(n_9703)
);

HB1xp67_ASAP7_75t_L g9704 ( 
.A(n_9075),
.Y(n_9704)
);

NAND2xp5_ASAP7_75t_L g9705 ( 
.A(n_9149),
.B(n_74),
.Y(n_9705)
);

INVxp67_ASAP7_75t_L g9706 ( 
.A(n_9082),
.Y(n_9706)
);

INVx1_ASAP7_75t_L g9707 ( 
.A(n_8773),
.Y(n_9707)
);

NAND2xp5_ASAP7_75t_L g9708 ( 
.A(n_8789),
.B(n_75),
.Y(n_9708)
);

AND2x4_ASAP7_75t_L g9709 ( 
.A(n_8934),
.B(n_329),
.Y(n_9709)
);

NOR2xp33_ASAP7_75t_L g9710 ( 
.A(n_9081),
.B(n_330),
.Y(n_9710)
);

OAI21xp5_ASAP7_75t_L g9711 ( 
.A1(n_8915),
.A2(n_8984),
.B(n_9107),
.Y(n_9711)
);

AND2x2_ASAP7_75t_L g9712 ( 
.A(n_8962),
.B(n_75),
.Y(n_9712)
);

BUFx6f_ASAP7_75t_L g9713 ( 
.A(n_8809),
.Y(n_9713)
);

NAND2xp5_ASAP7_75t_L g9714 ( 
.A(n_9141),
.B(n_75),
.Y(n_9714)
);

HB1xp67_ASAP7_75t_L g9715 ( 
.A(n_9110),
.Y(n_9715)
);

NOR2xp33_ASAP7_75t_L g9716 ( 
.A(n_9037),
.B(n_330),
.Y(n_9716)
);

NAND2xp5_ASAP7_75t_L g9717 ( 
.A(n_9057),
.B(n_9070),
.Y(n_9717)
);

INVx2_ASAP7_75t_SL g9718 ( 
.A(n_9172),
.Y(n_9718)
);

NAND2xp5_ASAP7_75t_L g9719 ( 
.A(n_9190),
.B(n_76),
.Y(n_9719)
);

OAI21xp5_ASAP7_75t_L g9720 ( 
.A1(n_9177),
.A2(n_76),
.B(n_77),
.Y(n_9720)
);

INVx1_ASAP7_75t_L g9721 ( 
.A(n_9169),
.Y(n_9721)
);

INVx1_ASAP7_75t_L g9722 ( 
.A(n_9192),
.Y(n_9722)
);

INVx1_ASAP7_75t_L g9723 ( 
.A(n_9116),
.Y(n_9723)
);

AND2x2_ASAP7_75t_L g9724 ( 
.A(n_8701),
.B(n_76),
.Y(n_9724)
);

INVx2_ASAP7_75t_L g9725 ( 
.A(n_8702),
.Y(n_9725)
);

INVx3_ASAP7_75t_L g9726 ( 
.A(n_9197),
.Y(n_9726)
);

INVx3_ASAP7_75t_L g9727 ( 
.A(n_9197),
.Y(n_9727)
);

INVx2_ASAP7_75t_L g9728 ( 
.A(n_8702),
.Y(n_9728)
);

INVx1_ASAP7_75t_L g9729 ( 
.A(n_8874),
.Y(n_9729)
);

INVx4_ASAP7_75t_L g9730 ( 
.A(n_9004),
.Y(n_9730)
);

INVx1_ASAP7_75t_SL g9731 ( 
.A(n_8805),
.Y(n_9731)
);

INVxp67_ASAP7_75t_SL g9732 ( 
.A(n_8895),
.Y(n_9732)
);

NOR2xp33_ASAP7_75t_L g9733 ( 
.A(n_8711),
.B(n_331),
.Y(n_9733)
);

AND2x4_ASAP7_75t_L g9734 ( 
.A(n_9197),
.B(n_331),
.Y(n_9734)
);

INVx3_ASAP7_75t_L g9735 ( 
.A(n_9197),
.Y(n_9735)
);

INVx1_ASAP7_75t_L g9736 ( 
.A(n_8874),
.Y(n_9736)
);

NAND2xp5_ASAP7_75t_SL g9737 ( 
.A(n_8711),
.B(n_332),
.Y(n_9737)
);

INVx2_ASAP7_75t_L g9738 ( 
.A(n_8702),
.Y(n_9738)
);

AND2x2_ASAP7_75t_L g9739 ( 
.A(n_8701),
.B(n_77),
.Y(n_9739)
);

INVx2_ASAP7_75t_L g9740 ( 
.A(n_8702),
.Y(n_9740)
);

HB1xp67_ASAP7_75t_L g9741 ( 
.A(n_8829),
.Y(n_9741)
);

AND2x2_ASAP7_75t_L g9742 ( 
.A(n_8701),
.B(n_77),
.Y(n_9742)
);

INVx1_ASAP7_75t_L g9743 ( 
.A(n_8874),
.Y(n_9743)
);

INVx2_ASAP7_75t_L g9744 ( 
.A(n_8702),
.Y(n_9744)
);

INVx1_ASAP7_75t_L g9745 ( 
.A(n_8874),
.Y(n_9745)
);

NOR2xp33_ASAP7_75t_L g9746 ( 
.A(n_8711),
.B(n_332),
.Y(n_9746)
);

BUFx8_ASAP7_75t_L g9747 ( 
.A(n_9042),
.Y(n_9747)
);

INVx2_ASAP7_75t_L g9748 ( 
.A(n_8702),
.Y(n_9748)
);

NAND2xp5_ASAP7_75t_L g9749 ( 
.A(n_8694),
.B(n_78),
.Y(n_9749)
);

INVxp67_ASAP7_75t_L g9750 ( 
.A(n_8731),
.Y(n_9750)
);

NAND2xp5_ASAP7_75t_L g9751 ( 
.A(n_8694),
.B(n_78),
.Y(n_9751)
);

BUFx3_ASAP7_75t_L g9752 ( 
.A(n_9197),
.Y(n_9752)
);

INVx2_ASAP7_75t_L g9753 ( 
.A(n_8702),
.Y(n_9753)
);

INVx1_ASAP7_75t_L g9754 ( 
.A(n_8874),
.Y(n_9754)
);

BUFx3_ASAP7_75t_L g9755 ( 
.A(n_9197),
.Y(n_9755)
);

NAND2xp5_ASAP7_75t_L g9756 ( 
.A(n_8694),
.B(n_79),
.Y(n_9756)
);

NOR2xp33_ASAP7_75t_L g9757 ( 
.A(n_8711),
.B(n_333),
.Y(n_9757)
);

HB1xp67_ASAP7_75t_L g9758 ( 
.A(n_8829),
.Y(n_9758)
);

NAND2xp5_ASAP7_75t_L g9759 ( 
.A(n_8694),
.B(n_80),
.Y(n_9759)
);

NAND2xp5_ASAP7_75t_L g9760 ( 
.A(n_8694),
.B(n_80),
.Y(n_9760)
);

INVx3_ASAP7_75t_L g9761 ( 
.A(n_9197),
.Y(n_9761)
);

AND2x4_ASAP7_75t_L g9762 ( 
.A(n_9197),
.B(n_333),
.Y(n_9762)
);

BUFx4f_ASAP7_75t_L g9763 ( 
.A(n_9004),
.Y(n_9763)
);

INVx2_ASAP7_75t_L g9764 ( 
.A(n_8702),
.Y(n_9764)
);

AND2x2_ASAP7_75t_L g9765 ( 
.A(n_8701),
.B(n_80),
.Y(n_9765)
);

AND2x2_ASAP7_75t_L g9766 ( 
.A(n_8701),
.B(n_81),
.Y(n_9766)
);

INVx4_ASAP7_75t_L g9767 ( 
.A(n_9004),
.Y(n_9767)
);

NAND2xp5_ASAP7_75t_L g9768 ( 
.A(n_8694),
.B(n_81),
.Y(n_9768)
);

NAND2xp5_ASAP7_75t_L g9769 ( 
.A(n_8694),
.B(n_81),
.Y(n_9769)
);

INVx2_ASAP7_75t_L g9770 ( 
.A(n_8702),
.Y(n_9770)
);

INVx1_ASAP7_75t_L g9771 ( 
.A(n_8874),
.Y(n_9771)
);

NOR2xp33_ASAP7_75t_L g9772 ( 
.A(n_8711),
.B(n_334),
.Y(n_9772)
);

AND2x2_ASAP7_75t_L g9773 ( 
.A(n_8701),
.B(n_82),
.Y(n_9773)
);

NAND2xp5_ASAP7_75t_SL g9774 ( 
.A(n_8711),
.B(n_334),
.Y(n_9774)
);

AND2x4_ASAP7_75t_L g9775 ( 
.A(n_9197),
.B(n_335),
.Y(n_9775)
);

INVx1_ASAP7_75t_SL g9776 ( 
.A(n_8805),
.Y(n_9776)
);

HB1xp67_ASAP7_75t_L g9777 ( 
.A(n_8829),
.Y(n_9777)
);

NOR2xp33_ASAP7_75t_L g9778 ( 
.A(n_8711),
.B(n_335),
.Y(n_9778)
);

AND2x2_ASAP7_75t_L g9779 ( 
.A(n_8701),
.B(n_82),
.Y(n_9779)
);

INVx2_ASAP7_75t_L g9780 ( 
.A(n_8702),
.Y(n_9780)
);

HB1xp67_ASAP7_75t_L g9781 ( 
.A(n_8829),
.Y(n_9781)
);

BUFx3_ASAP7_75t_L g9782 ( 
.A(n_9197),
.Y(n_9782)
);

AND2x2_ASAP7_75t_L g9783 ( 
.A(n_8701),
.B(n_82),
.Y(n_9783)
);

NAND2xp5_ASAP7_75t_L g9784 ( 
.A(n_8694),
.B(n_83),
.Y(n_9784)
);

AOI22xp5_ASAP7_75t_L g9785 ( 
.A1(n_8711),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_9785)
);

INVx1_ASAP7_75t_L g9786 ( 
.A(n_8874),
.Y(n_9786)
);

INVx2_ASAP7_75t_L g9787 ( 
.A(n_8702),
.Y(n_9787)
);

NAND2xp5_ASAP7_75t_L g9788 ( 
.A(n_8694),
.B(n_83),
.Y(n_9788)
);

INVx3_ASAP7_75t_L g9789 ( 
.A(n_9197),
.Y(n_9789)
);

AND2x2_ASAP7_75t_L g9790 ( 
.A(n_8701),
.B(n_84),
.Y(n_9790)
);

INVx2_ASAP7_75t_L g9791 ( 
.A(n_8702),
.Y(n_9791)
);

BUFx3_ASAP7_75t_L g9792 ( 
.A(n_9197),
.Y(n_9792)
);

HB1xp67_ASAP7_75t_L g9793 ( 
.A(n_8829),
.Y(n_9793)
);

BUFx3_ASAP7_75t_L g9794 ( 
.A(n_9197),
.Y(n_9794)
);

INVx1_ASAP7_75t_L g9795 ( 
.A(n_8874),
.Y(n_9795)
);

BUFx3_ASAP7_75t_L g9796 ( 
.A(n_9197),
.Y(n_9796)
);

NAND2xp5_ASAP7_75t_L g9797 ( 
.A(n_8694),
.B(n_84),
.Y(n_9797)
);

INVx2_ASAP7_75t_SL g9798 ( 
.A(n_8911),
.Y(n_9798)
);

AND2x2_ASAP7_75t_L g9799 ( 
.A(n_8701),
.B(n_85),
.Y(n_9799)
);

NOR2xp33_ASAP7_75t_L g9800 ( 
.A(n_8711),
.B(n_336),
.Y(n_9800)
);

AND2x2_ASAP7_75t_SL g9801 ( 
.A(n_8711),
.B(n_336),
.Y(n_9801)
);

INVx1_ASAP7_75t_L g9802 ( 
.A(n_8874),
.Y(n_9802)
);

NAND2xp5_ASAP7_75t_SL g9803 ( 
.A(n_8711),
.B(n_337),
.Y(n_9803)
);

INVx1_ASAP7_75t_L g9804 ( 
.A(n_8874),
.Y(n_9804)
);

INVx2_ASAP7_75t_L g9805 ( 
.A(n_8702),
.Y(n_9805)
);

INVx2_ASAP7_75t_L g9806 ( 
.A(n_8702),
.Y(n_9806)
);

AND2x2_ASAP7_75t_L g9807 ( 
.A(n_8701),
.B(n_86),
.Y(n_9807)
);

AND2x2_ASAP7_75t_L g9808 ( 
.A(n_8701),
.B(n_86),
.Y(n_9808)
);

INVx1_ASAP7_75t_L g9809 ( 
.A(n_8874),
.Y(n_9809)
);

NAND2xp5_ASAP7_75t_L g9810 ( 
.A(n_8694),
.B(n_86),
.Y(n_9810)
);

AOI21xp5_ASAP7_75t_L g9811 ( 
.A1(n_9406),
.A2(n_338),
.B(n_337),
.Y(n_9811)
);

NOR3xp33_ASAP7_75t_L g9812 ( 
.A(n_9266),
.B(n_87),
.C(n_88),
.Y(n_9812)
);

BUFx12f_ASAP7_75t_L g9813 ( 
.A(n_9376),
.Y(n_9813)
);

AOI21xp5_ASAP7_75t_L g9814 ( 
.A1(n_9680),
.A2(n_339),
.B(n_338),
.Y(n_9814)
);

INVx1_ASAP7_75t_L g9815 ( 
.A(n_9315),
.Y(n_9815)
);

AOI21xp5_ASAP7_75t_L g9816 ( 
.A1(n_9353),
.A2(n_340),
.B(n_339),
.Y(n_9816)
);

NAND2xp5_ASAP7_75t_L g9817 ( 
.A(n_9296),
.B(n_341),
.Y(n_9817)
);

NAND2xp5_ASAP7_75t_L g9818 ( 
.A(n_9211),
.B(n_341),
.Y(n_9818)
);

BUFx12f_ASAP7_75t_L g9819 ( 
.A(n_9747),
.Y(n_9819)
);

AOI21xp5_ASAP7_75t_L g9820 ( 
.A1(n_9546),
.A2(n_344),
.B(n_342),
.Y(n_9820)
);

BUFx4f_ASAP7_75t_L g9821 ( 
.A(n_9218),
.Y(n_9821)
);

OAI22xp5_ASAP7_75t_L g9822 ( 
.A1(n_9258),
.A2(n_9281),
.B1(n_9801),
.B2(n_9509),
.Y(n_9822)
);

AOI21x1_ASAP7_75t_L g9823 ( 
.A1(n_9547),
.A2(n_87),
.B(n_88),
.Y(n_9823)
);

INVx1_ASAP7_75t_L g9824 ( 
.A(n_9316),
.Y(n_9824)
);

AND2x2_ASAP7_75t_L g9825 ( 
.A(n_9314),
.B(n_342),
.Y(n_9825)
);

NOR2xp33_ASAP7_75t_L g9826 ( 
.A(n_9500),
.B(n_344),
.Y(n_9826)
);

NAND2xp5_ASAP7_75t_L g9827 ( 
.A(n_9729),
.B(n_9736),
.Y(n_9827)
);

BUFx6f_ASAP7_75t_L g9828 ( 
.A(n_9763),
.Y(n_9828)
);

AND2x2_ASAP7_75t_L g9829 ( 
.A(n_9562),
.B(n_345),
.Y(n_9829)
);

NAND2xp5_ASAP7_75t_SL g9830 ( 
.A(n_9449),
.B(n_346),
.Y(n_9830)
);

NAND2xp5_ASAP7_75t_L g9831 ( 
.A(n_9743),
.B(n_347),
.Y(n_9831)
);

BUFx6f_ASAP7_75t_L g9832 ( 
.A(n_9218),
.Y(n_9832)
);

O2A1O1Ixp33_ASAP7_75t_L g9833 ( 
.A1(n_9537),
.A2(n_91),
.B(n_89),
.C(n_90),
.Y(n_9833)
);

BUFx6f_ASAP7_75t_L g9834 ( 
.A(n_9224),
.Y(n_9834)
);

NOR3xp33_ASAP7_75t_L g9835 ( 
.A(n_9262),
.B(n_89),
.C(n_91),
.Y(n_9835)
);

AND2x4_ASAP7_75t_L g9836 ( 
.A(n_9480),
.B(n_347),
.Y(n_9836)
);

AOI22xp5_ASAP7_75t_L g9837 ( 
.A1(n_9733),
.A2(n_9746),
.B1(n_9772),
.B2(n_9757),
.Y(n_9837)
);

NAND2xp5_ASAP7_75t_L g9838 ( 
.A(n_9745),
.B(n_348),
.Y(n_9838)
);

AOI21xp5_ASAP7_75t_L g9839 ( 
.A1(n_9662),
.A2(n_349),
.B(n_348),
.Y(n_9839)
);

OAI22xp5_ASAP7_75t_L g9840 ( 
.A1(n_9342),
.A2(n_93),
.B1(n_89),
.B2(n_92),
.Y(n_9840)
);

O2A1O1Ixp33_ASAP7_75t_L g9841 ( 
.A1(n_9778),
.A2(n_95),
.B(n_92),
.C(n_94),
.Y(n_9841)
);

NOR2xp33_ASAP7_75t_L g9842 ( 
.A(n_9320),
.B(n_350),
.Y(n_9842)
);

NOR2xp33_ASAP7_75t_L g9843 ( 
.A(n_9731),
.B(n_350),
.Y(n_9843)
);

AOI21x1_ASAP7_75t_L g9844 ( 
.A1(n_9667),
.A2(n_92),
.B(n_94),
.Y(n_9844)
);

NOR2xp33_ASAP7_75t_L g9845 ( 
.A(n_9776),
.B(n_351),
.Y(n_9845)
);

BUFx4f_ASAP7_75t_L g9846 ( 
.A(n_9224),
.Y(n_9846)
);

BUFx2_ASAP7_75t_L g9847 ( 
.A(n_9313),
.Y(n_9847)
);

BUFx2_ASAP7_75t_L g9848 ( 
.A(n_9310),
.Y(n_9848)
);

NAND2xp5_ASAP7_75t_L g9849 ( 
.A(n_9754),
.B(n_351),
.Y(n_9849)
);

NAND2xp5_ASAP7_75t_L g9850 ( 
.A(n_9771),
.B(n_352),
.Y(n_9850)
);

INVx1_ASAP7_75t_L g9851 ( 
.A(n_9322),
.Y(n_9851)
);

INVx2_ASAP7_75t_L g9852 ( 
.A(n_9217),
.Y(n_9852)
);

AOI21xp5_ASAP7_75t_L g9853 ( 
.A1(n_9247),
.A2(n_353),
.B(n_352),
.Y(n_9853)
);

AOI22xp5_ASAP7_75t_L g9854 ( 
.A1(n_9800),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_9854)
);

AOI21xp5_ASAP7_75t_L g9855 ( 
.A1(n_9732),
.A2(n_357),
.B(n_355),
.Y(n_9855)
);

AOI21xp5_ASAP7_75t_L g9856 ( 
.A1(n_9689),
.A2(n_358),
.B(n_357),
.Y(n_9856)
);

OAI321xp33_ASAP7_75t_L g9857 ( 
.A1(n_9656),
.A2(n_98),
.A3(n_100),
.B1(n_96),
.B2(n_97),
.C(n_99),
.Y(n_9857)
);

NAND2xp5_ASAP7_75t_SL g9858 ( 
.A(n_9475),
.B(n_358),
.Y(n_9858)
);

NOR3xp33_ASAP7_75t_L g9859 ( 
.A(n_9257),
.B(n_97),
.C(n_98),
.Y(n_9859)
);

AOI21xp5_ASAP7_75t_L g9860 ( 
.A1(n_9711),
.A2(n_360),
.B(n_359),
.Y(n_9860)
);

AOI21xp5_ASAP7_75t_L g9861 ( 
.A1(n_9647),
.A2(n_360),
.B(n_359),
.Y(n_9861)
);

AOI222xp33_ASAP7_75t_L g9862 ( 
.A1(n_9538),
.A2(n_100),
.B1(n_102),
.B2(n_98),
.C1(n_99),
.C2(n_101),
.Y(n_9862)
);

O2A1O1Ixp5_ASAP7_75t_L g9863 ( 
.A1(n_9625),
.A2(n_103),
.B(n_101),
.C(n_102),
.Y(n_9863)
);

O2A1O1Ixp5_ASAP7_75t_L g9864 ( 
.A1(n_9357),
.A2(n_103),
.B(n_101),
.C(n_102),
.Y(n_9864)
);

INVx2_ASAP7_75t_L g9865 ( 
.A(n_9220),
.Y(n_9865)
);

AOI21xp5_ASAP7_75t_L g9866 ( 
.A1(n_9335),
.A2(n_363),
.B(n_361),
.Y(n_9866)
);

INVx1_ASAP7_75t_L g9867 ( 
.A(n_9329),
.Y(n_9867)
);

AOI21xp5_ASAP7_75t_L g9868 ( 
.A1(n_9675),
.A2(n_363),
.B(n_361),
.Y(n_9868)
);

BUFx6f_ASAP7_75t_L g9869 ( 
.A(n_9239),
.Y(n_9869)
);

AOI21xp5_ASAP7_75t_L g9870 ( 
.A1(n_9695),
.A2(n_365),
.B(n_364),
.Y(n_9870)
);

AOI21x1_ASAP7_75t_L g9871 ( 
.A1(n_9707),
.A2(n_9573),
.B(n_9665),
.Y(n_9871)
);

AOI21x1_ASAP7_75t_L g9872 ( 
.A1(n_9362),
.A2(n_104),
.B(n_105),
.Y(n_9872)
);

INVx1_ASAP7_75t_L g9873 ( 
.A(n_9332),
.Y(n_9873)
);

NAND2xp5_ASAP7_75t_L g9874 ( 
.A(n_9786),
.B(n_364),
.Y(n_9874)
);

AOI21x1_ASAP7_75t_L g9875 ( 
.A1(n_9669),
.A2(n_104),
.B(n_105),
.Y(n_9875)
);

NAND2xp5_ASAP7_75t_L g9876 ( 
.A(n_9795),
.B(n_366),
.Y(n_9876)
);

AOI21xp5_ASAP7_75t_L g9877 ( 
.A1(n_9462),
.A2(n_367),
.B(n_366),
.Y(n_9877)
);

NAND2xp5_ASAP7_75t_L g9878 ( 
.A(n_9802),
.B(n_367),
.Y(n_9878)
);

NAND2xp5_ASAP7_75t_L g9879 ( 
.A(n_9804),
.B(n_368),
.Y(n_9879)
);

INVx1_ASAP7_75t_L g9880 ( 
.A(n_9343),
.Y(n_9880)
);

INVx5_ASAP7_75t_L g9881 ( 
.A(n_9529),
.Y(n_9881)
);

AOI21xp5_ASAP7_75t_L g9882 ( 
.A1(n_9809),
.A2(n_369),
.B(n_368),
.Y(n_9882)
);

NOR2xp33_ASAP7_75t_L g9883 ( 
.A(n_9545),
.B(n_9300),
.Y(n_9883)
);

O2A1O1Ixp33_ASAP7_75t_L g9884 ( 
.A1(n_9282),
.A2(n_106),
.B(n_104),
.C(n_105),
.Y(n_9884)
);

AOI21xp5_ASAP7_75t_L g9885 ( 
.A1(n_9684),
.A2(n_9259),
.B(n_9637),
.Y(n_9885)
);

AOI21xp5_ASAP7_75t_L g9886 ( 
.A1(n_9638),
.A2(n_371),
.B(n_370),
.Y(n_9886)
);

OAI21xp33_ASAP7_75t_L g9887 ( 
.A1(n_9295),
.A2(n_106),
.B(n_107),
.Y(n_9887)
);

AOI21xp5_ASAP7_75t_L g9888 ( 
.A1(n_9650),
.A2(n_9586),
.B(n_9612),
.Y(n_9888)
);

AOI21xp5_ASAP7_75t_L g9889 ( 
.A1(n_9621),
.A2(n_9584),
.B(n_9583),
.Y(n_9889)
);

BUFx4f_ASAP7_75t_L g9890 ( 
.A(n_9239),
.Y(n_9890)
);

INVxp67_ASAP7_75t_L g9891 ( 
.A(n_9275),
.Y(n_9891)
);

INVx1_ASAP7_75t_L g9892 ( 
.A(n_9349),
.Y(n_9892)
);

AOI21xp5_ASAP7_75t_L g9893 ( 
.A1(n_9607),
.A2(n_372),
.B(n_370),
.Y(n_9893)
);

CKINVDCx8_ASAP7_75t_R g9894 ( 
.A(n_9450),
.Y(n_9894)
);

NAND2xp5_ASAP7_75t_SL g9895 ( 
.A(n_9660),
.B(n_372),
.Y(n_9895)
);

NAND2xp5_ASAP7_75t_L g9896 ( 
.A(n_9560),
.B(n_373),
.Y(n_9896)
);

O2A1O1Ixp5_ASAP7_75t_L g9897 ( 
.A1(n_9423),
.A2(n_108),
.B(n_106),
.C(n_107),
.Y(n_9897)
);

NAND2xp5_ASAP7_75t_L g9898 ( 
.A(n_9568),
.B(n_374),
.Y(n_9898)
);

CKINVDCx20_ASAP7_75t_R g9899 ( 
.A(n_9234),
.Y(n_9899)
);

NOR2x1p5_ASAP7_75t_SL g9900 ( 
.A(n_9567),
.B(n_374),
.Y(n_9900)
);

NAND2xp5_ASAP7_75t_L g9901 ( 
.A(n_9572),
.B(n_375),
.Y(n_9901)
);

AND2x4_ASAP7_75t_L g9902 ( 
.A(n_9341),
.B(n_9231),
.Y(n_9902)
);

NAND2xp5_ASAP7_75t_L g9903 ( 
.A(n_9574),
.B(n_375),
.Y(n_9903)
);

OAI21xp5_ASAP7_75t_L g9904 ( 
.A1(n_9241),
.A2(n_108),
.B(n_109),
.Y(n_9904)
);

INVx1_ASAP7_75t_L g9905 ( 
.A(n_9367),
.Y(n_9905)
);

NOR2xp33_ASAP7_75t_L g9906 ( 
.A(n_9659),
.B(n_376),
.Y(n_9906)
);

AOI21x1_ASAP7_75t_L g9907 ( 
.A1(n_9694),
.A2(n_108),
.B(n_109),
.Y(n_9907)
);

HB1xp67_ASAP7_75t_L g9908 ( 
.A(n_9426),
.Y(n_9908)
);

OAI321xp33_ASAP7_75t_L g9909 ( 
.A1(n_9370),
.A2(n_9443),
.A3(n_9785),
.B1(n_9710),
.B2(n_9340),
.C(n_9291),
.Y(n_9909)
);

INVx2_ASAP7_75t_L g9910 ( 
.A(n_9248),
.Y(n_9910)
);

INVx11_ASAP7_75t_L g9911 ( 
.A(n_9304),
.Y(n_9911)
);

INVx1_ASAP7_75t_L g9912 ( 
.A(n_9368),
.Y(n_9912)
);

O2A1O1Ixp33_ASAP7_75t_L g9913 ( 
.A1(n_9737),
.A2(n_9803),
.B(n_9774),
.C(n_9374),
.Y(n_9913)
);

OAI21x1_ASAP7_75t_L g9914 ( 
.A1(n_9581),
.A2(n_109),
.B(n_110),
.Y(n_9914)
);

AOI21xp5_ASAP7_75t_L g9915 ( 
.A1(n_9627),
.A2(n_377),
.B(n_376),
.Y(n_9915)
);

AOI21xp5_ASAP7_75t_L g9916 ( 
.A1(n_9635),
.A2(n_379),
.B(n_378),
.Y(n_9916)
);

NOR3xp33_ASAP7_75t_L g9917 ( 
.A(n_9674),
.B(n_9230),
.C(n_9321),
.Y(n_9917)
);

AOI21xp5_ASAP7_75t_L g9918 ( 
.A1(n_9636),
.A2(n_381),
.B(n_380),
.Y(n_9918)
);

AOI21xp5_ASAP7_75t_L g9919 ( 
.A1(n_9643),
.A2(n_382),
.B(n_381),
.Y(n_9919)
);

INVx3_ASAP7_75t_L g9920 ( 
.A(n_9212),
.Y(n_9920)
);

AOI21xp33_ASAP7_75t_L g9921 ( 
.A1(n_9369),
.A2(n_110),
.B(n_111),
.Y(n_9921)
);

NOR2x1_ASAP7_75t_L g9922 ( 
.A(n_9459),
.B(n_383),
.Y(n_9922)
);

HB1xp67_ASAP7_75t_L g9923 ( 
.A(n_9435),
.Y(n_9923)
);

OAI21xp5_ASAP7_75t_L g9924 ( 
.A1(n_9331),
.A2(n_110),
.B(n_111),
.Y(n_9924)
);

NAND2xp5_ASAP7_75t_L g9925 ( 
.A(n_9626),
.B(n_383),
.Y(n_9925)
);

AOI21xp5_ASAP7_75t_L g9926 ( 
.A1(n_9644),
.A2(n_9651),
.B(n_9646),
.Y(n_9926)
);

NAND2xp5_ASAP7_75t_SL g9927 ( 
.A(n_9653),
.B(n_384),
.Y(n_9927)
);

O2A1O1Ixp33_ASAP7_75t_L g9928 ( 
.A1(n_9336),
.A2(n_113),
.B(n_111),
.C(n_112),
.Y(n_9928)
);

INVx2_ASAP7_75t_L g9929 ( 
.A(n_9254),
.Y(n_9929)
);

NAND2xp5_ASAP7_75t_L g9930 ( 
.A(n_9648),
.B(n_384),
.Y(n_9930)
);

INVx3_ASAP7_75t_L g9931 ( 
.A(n_9752),
.Y(n_9931)
);

OAI21xp5_ASAP7_75t_L g9932 ( 
.A1(n_9256),
.A2(n_112),
.B(n_113),
.Y(n_9932)
);

A2O1A1Ixp33_ASAP7_75t_L g9933 ( 
.A1(n_9716),
.A2(n_386),
.B(n_387),
.C(n_385),
.Y(n_9933)
);

INVx1_ASAP7_75t_L g9934 ( 
.A(n_9373),
.Y(n_9934)
);

AND2x2_ASAP7_75t_SL g9935 ( 
.A(n_9427),
.B(n_9416),
.Y(n_9935)
);

INVx1_ASAP7_75t_L g9936 ( 
.A(n_9394),
.Y(n_9936)
);

OAI21x1_ASAP7_75t_L g9937 ( 
.A1(n_9597),
.A2(n_113),
.B(n_114),
.Y(n_9937)
);

AOI21xp5_ASAP7_75t_L g9938 ( 
.A1(n_9654),
.A2(n_386),
.B(n_385),
.Y(n_9938)
);

HB1xp67_ASAP7_75t_L g9939 ( 
.A(n_9297),
.Y(n_9939)
);

AND2x4_ASAP7_75t_L g9940 ( 
.A(n_9272),
.B(n_9298),
.Y(n_9940)
);

AOI22xp5_ASAP7_75t_L g9941 ( 
.A1(n_9532),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_9941)
);

INVx2_ASAP7_75t_L g9942 ( 
.A(n_9278),
.Y(n_9942)
);

AOI21x1_ASAP7_75t_L g9943 ( 
.A1(n_9472),
.A2(n_114),
.B(n_115),
.Y(n_9943)
);

AOI21xp5_ASAP7_75t_L g9944 ( 
.A1(n_9655),
.A2(n_389),
.B(n_388),
.Y(n_9944)
);

HB1xp67_ASAP7_75t_L g9945 ( 
.A(n_9565),
.Y(n_9945)
);

NOR2xp33_ASAP7_75t_L g9946 ( 
.A(n_9470),
.B(n_388),
.Y(n_9946)
);

AND2x2_ASAP7_75t_L g9947 ( 
.A(n_9724),
.B(n_389),
.Y(n_9947)
);

NAND2xp5_ASAP7_75t_L g9948 ( 
.A(n_9392),
.B(n_9542),
.Y(n_9948)
);

AOI21xp5_ASAP7_75t_L g9949 ( 
.A1(n_9600),
.A2(n_391),
.B(n_390),
.Y(n_9949)
);

AND2x4_ASAP7_75t_L g9950 ( 
.A(n_9333),
.B(n_390),
.Y(n_9950)
);

OAI22xp5_ASAP7_75t_L g9951 ( 
.A1(n_9721),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_9951)
);

NOR2xp33_ASAP7_75t_L g9952 ( 
.A(n_9679),
.B(n_392),
.Y(n_9952)
);

OAI22xp5_ASAP7_75t_L g9953 ( 
.A1(n_9513),
.A2(n_9350),
.B1(n_9358),
.B2(n_9365),
.Y(n_9953)
);

CKINVDCx6p67_ASAP7_75t_R g9954 ( 
.A(n_9755),
.Y(n_9954)
);

NAND2xp5_ASAP7_75t_L g9955 ( 
.A(n_9488),
.B(n_9496),
.Y(n_9955)
);

INVx1_ASAP7_75t_L g9956 ( 
.A(n_9397),
.Y(n_9956)
);

AOI21xp5_ASAP7_75t_L g9957 ( 
.A1(n_9608),
.A2(n_393),
.B(n_392),
.Y(n_9957)
);

O2A1O1Ixp5_ASAP7_75t_L g9958 ( 
.A1(n_9687),
.A2(n_118),
.B(n_116),
.C(n_117),
.Y(n_9958)
);

AOI21xp5_ASAP7_75t_L g9959 ( 
.A1(n_9615),
.A2(n_394),
.B(n_393),
.Y(n_9959)
);

NOR2xp33_ASAP7_75t_L g9960 ( 
.A(n_9622),
.B(n_394),
.Y(n_9960)
);

NAND2xp5_ASAP7_75t_L g9961 ( 
.A(n_9325),
.B(n_395),
.Y(n_9961)
);

NAND2xp5_ASAP7_75t_L g9962 ( 
.A(n_9235),
.B(n_9360),
.Y(n_9962)
);

AOI21x1_ASAP7_75t_L g9963 ( 
.A1(n_9417),
.A2(n_117),
.B(n_119),
.Y(n_9963)
);

AOI21xp5_ASAP7_75t_L g9964 ( 
.A1(n_9630),
.A2(n_396),
.B(n_395),
.Y(n_9964)
);

INVx1_ASAP7_75t_L g9965 ( 
.A(n_9402),
.Y(n_9965)
);

OAI21xp5_ASAP7_75t_L g9966 ( 
.A1(n_9244),
.A2(n_119),
.B(n_120),
.Y(n_9966)
);

AOI21xp5_ASAP7_75t_L g9967 ( 
.A1(n_9670),
.A2(n_398),
.B(n_397),
.Y(n_9967)
);

AOI21xp5_ASAP7_75t_L g9968 ( 
.A1(n_9253),
.A2(n_398),
.B(n_397),
.Y(n_9968)
);

OAI22xp5_ASAP7_75t_L g9969 ( 
.A1(n_9527),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_9969)
);

BUFx4f_ASAP7_75t_L g9970 ( 
.A(n_9240),
.Y(n_9970)
);

NAND2xp5_ASAP7_75t_L g9971 ( 
.A(n_9235),
.B(n_399),
.Y(n_9971)
);

AOI21xp5_ASAP7_75t_L g9972 ( 
.A1(n_9215),
.A2(n_400),
.B(n_399),
.Y(n_9972)
);

NAND2xp5_ASAP7_75t_L g9973 ( 
.A(n_9235),
.B(n_400),
.Y(n_9973)
);

NAND3xp33_ASAP7_75t_SL g9974 ( 
.A(n_9364),
.B(n_120),
.C(n_121),
.Y(n_9974)
);

AOI21xp5_ASAP7_75t_L g9975 ( 
.A1(n_9717),
.A2(n_402),
.B(n_401),
.Y(n_9975)
);

OAI21xp5_ASAP7_75t_L g9976 ( 
.A1(n_9553),
.A2(n_9566),
.B(n_9477),
.Y(n_9976)
);

NAND2xp5_ASAP7_75t_L g9977 ( 
.A(n_9302),
.B(n_401),
.Y(n_9977)
);

NAND2xp5_ASAP7_75t_L g9978 ( 
.A(n_9749),
.B(n_402),
.Y(n_9978)
);

NAND2xp5_ASAP7_75t_L g9979 ( 
.A(n_9751),
.B(n_403),
.Y(n_9979)
);

AOI21xp5_ASAP7_75t_L g9980 ( 
.A1(n_9634),
.A2(n_404),
.B(n_403),
.Y(n_9980)
);

NOR3xp33_ASAP7_75t_L g9981 ( 
.A(n_9587),
.B(n_121),
.C(n_123),
.Y(n_9981)
);

AND2x4_ASAP7_75t_L g9982 ( 
.A(n_9534),
.B(n_405),
.Y(n_9982)
);

NOR2xp33_ASAP7_75t_L g9983 ( 
.A(n_9286),
.B(n_9578),
.Y(n_9983)
);

NAND2xp5_ASAP7_75t_L g9984 ( 
.A(n_9756),
.B(n_405),
.Y(n_9984)
);

O2A1O1Ixp33_ASAP7_75t_L g9985 ( 
.A1(n_9697),
.A2(n_125),
.B(n_123),
.C(n_124),
.Y(n_9985)
);

AOI21xp5_ASAP7_75t_L g9986 ( 
.A1(n_9652),
.A2(n_407),
.B(n_406),
.Y(n_9986)
);

INVx2_ASAP7_75t_L g9987 ( 
.A(n_9303),
.Y(n_9987)
);

BUFx6f_ASAP7_75t_L g9988 ( 
.A(n_9240),
.Y(n_9988)
);

INVx4_ASAP7_75t_L g9989 ( 
.A(n_9245),
.Y(n_9989)
);

AOI21xp5_ASAP7_75t_L g9990 ( 
.A1(n_9759),
.A2(n_407),
.B(n_406),
.Y(n_9990)
);

INVx2_ASAP7_75t_L g9991 ( 
.A(n_9725),
.Y(n_9991)
);

OAI21xp5_ASAP7_75t_L g9992 ( 
.A1(n_9672),
.A2(n_123),
.B(n_124),
.Y(n_9992)
);

OAI22xp5_ASAP7_75t_L g9993 ( 
.A1(n_9641),
.A2(n_9750),
.B1(n_9213),
.B2(n_9570),
.Y(n_9993)
);

AOI21xp5_ASAP7_75t_L g9994 ( 
.A1(n_9760),
.A2(n_409),
.B(n_408),
.Y(n_9994)
);

INVx2_ASAP7_75t_SL g9995 ( 
.A(n_9782),
.Y(n_9995)
);

BUFx6f_ASAP7_75t_L g9996 ( 
.A(n_9245),
.Y(n_9996)
);

NOR2xp33_ASAP7_75t_SL g9997 ( 
.A(n_9223),
.B(n_124),
.Y(n_9997)
);

NOR2xp33_ASAP7_75t_SL g9998 ( 
.A(n_9730),
.B(n_125),
.Y(n_9998)
);

NOR2xp67_ASAP7_75t_L g9999 ( 
.A(n_9317),
.B(n_9319),
.Y(n_9999)
);

A2O1A1Ixp33_ASAP7_75t_L g10000 ( 
.A1(n_9558),
.A2(n_409),
.B(n_410),
.C(n_408),
.Y(n_10000)
);

NAND2xp5_ASAP7_75t_L g10001 ( 
.A(n_9768),
.B(n_410),
.Y(n_10001)
);

AOI21xp5_ASAP7_75t_L g10002 ( 
.A1(n_9769),
.A2(n_412),
.B(n_411),
.Y(n_10002)
);

CKINVDCx5p33_ASAP7_75t_R g10003 ( 
.A(n_9792),
.Y(n_10003)
);

INVx1_ASAP7_75t_L g10004 ( 
.A(n_9410),
.Y(n_10004)
);

AOI21xp5_ASAP7_75t_L g10005 ( 
.A1(n_9784),
.A2(n_413),
.B(n_412),
.Y(n_10005)
);

AOI21xp5_ASAP7_75t_L g10006 ( 
.A1(n_9788),
.A2(n_414),
.B(n_413),
.Y(n_10006)
);

O2A1O1Ixp33_ASAP7_75t_L g10007 ( 
.A1(n_9673),
.A2(n_127),
.B(n_125),
.C(n_126),
.Y(n_10007)
);

NAND2xp5_ASAP7_75t_L g10008 ( 
.A(n_9797),
.B(n_414),
.Y(n_10008)
);

NOR3xp33_ASAP7_75t_L g10009 ( 
.A(n_9720),
.B(n_126),
.C(n_127),
.Y(n_10009)
);

AOI21xp5_ASAP7_75t_L g10010 ( 
.A1(n_9810),
.A2(n_416),
.B(n_415),
.Y(n_10010)
);

INVx2_ASAP7_75t_L g10011 ( 
.A(n_9728),
.Y(n_10011)
);

INVx2_ASAP7_75t_L g10012 ( 
.A(n_9738),
.Y(n_10012)
);

BUFx6f_ASAP7_75t_L g10013 ( 
.A(n_9261),
.Y(n_10013)
);

AOI21xp5_ASAP7_75t_L g10014 ( 
.A1(n_9678),
.A2(n_416),
.B(n_415),
.Y(n_10014)
);

OAI21xp5_ASAP7_75t_L g10015 ( 
.A1(n_9664),
.A2(n_126),
.B(n_127),
.Y(n_10015)
);

NAND2xp5_ASAP7_75t_L g10016 ( 
.A(n_9351),
.B(n_417),
.Y(n_10016)
);

AOI21x1_ASAP7_75t_L g10017 ( 
.A1(n_9277),
.A2(n_128),
.B(n_129),
.Y(n_10017)
);

NAND2xp5_ASAP7_75t_L g10018 ( 
.A(n_9354),
.B(n_417),
.Y(n_10018)
);

AOI21x1_ASAP7_75t_L g10019 ( 
.A1(n_9592),
.A2(n_128),
.B(n_129),
.Y(n_10019)
);

INVx2_ASAP7_75t_L g10020 ( 
.A(n_9740),
.Y(n_10020)
);

INVx1_ASAP7_75t_L g10021 ( 
.A(n_9414),
.Y(n_10021)
);

INVxp67_ASAP7_75t_SL g10022 ( 
.A(n_9554),
.Y(n_10022)
);

AOI21xp5_ASAP7_75t_L g10023 ( 
.A1(n_9744),
.A2(n_419),
.B(n_418),
.Y(n_10023)
);

O2A1O1Ixp33_ASAP7_75t_SL g10024 ( 
.A1(n_9702),
.A2(n_131),
.B(n_128),
.C(n_130),
.Y(n_10024)
);

NOR2x1p5_ASAP7_75t_SL g10025 ( 
.A(n_9346),
.B(n_418),
.Y(n_10025)
);

AND2x2_ASAP7_75t_L g10026 ( 
.A(n_9739),
.B(n_420),
.Y(n_10026)
);

AND2x4_ASAP7_75t_L g10027 ( 
.A(n_9249),
.B(n_420),
.Y(n_10027)
);

BUFx3_ASAP7_75t_L g10028 ( 
.A(n_9794),
.Y(n_10028)
);

OAI21xp5_ASAP7_75t_L g10029 ( 
.A1(n_9663),
.A2(n_130),
.B(n_131),
.Y(n_10029)
);

AOI22xp5_ASAP7_75t_L g10030 ( 
.A1(n_9355),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.Y(n_10030)
);

AO21x1_ASAP7_75t_L g10031 ( 
.A1(n_9708),
.A2(n_132),
.B(n_133),
.Y(n_10031)
);

NAND2xp5_ASAP7_75t_SL g10032 ( 
.A(n_9682),
.B(n_421),
.Y(n_10032)
);

NAND2xp5_ASAP7_75t_SL g10033 ( 
.A(n_9596),
.B(n_421),
.Y(n_10033)
);

AOI21xp5_ASAP7_75t_L g10034 ( 
.A1(n_9748),
.A2(n_423),
.B(n_422),
.Y(n_10034)
);

AOI21xp5_ASAP7_75t_L g10035 ( 
.A1(n_9753),
.A2(n_423),
.B(n_422),
.Y(n_10035)
);

AOI21xp5_ASAP7_75t_L g10036 ( 
.A1(n_9764),
.A2(n_425),
.B(n_424),
.Y(n_10036)
);

BUFx5_ASAP7_75t_L g10037 ( 
.A(n_9529),
.Y(n_10037)
);

AOI21xp5_ASAP7_75t_L g10038 ( 
.A1(n_9770),
.A2(n_425),
.B(n_424),
.Y(n_10038)
);

INVx1_ASAP7_75t_SL g10039 ( 
.A(n_9411),
.Y(n_10039)
);

NAND3xp33_ASAP7_75t_L g10040 ( 
.A(n_9688),
.B(n_132),
.C(n_133),
.Y(n_10040)
);

NAND2xp5_ASAP7_75t_L g10041 ( 
.A(n_9780),
.B(n_426),
.Y(n_10041)
);

INVx2_ASAP7_75t_L g10042 ( 
.A(n_9787),
.Y(n_10042)
);

AOI21xp5_ASAP7_75t_L g10043 ( 
.A1(n_9791),
.A2(n_9806),
.B(n_9805),
.Y(n_10043)
);

AOI22xp5_ASAP7_75t_L g10044 ( 
.A1(n_9355),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.Y(n_10044)
);

INVx1_ASAP7_75t_L g10045 ( 
.A(n_9429),
.Y(n_10045)
);

AOI21xp5_ASAP7_75t_L g10046 ( 
.A1(n_9479),
.A2(n_428),
.B(n_427),
.Y(n_10046)
);

INVxp67_ASAP7_75t_L g10047 ( 
.A(n_9741),
.Y(n_10047)
);

BUFx6f_ASAP7_75t_L g10048 ( 
.A(n_9261),
.Y(n_10048)
);

NAND2xp5_ASAP7_75t_L g10049 ( 
.A(n_9434),
.B(n_427),
.Y(n_10049)
);

AOI21xp5_ASAP7_75t_L g10050 ( 
.A1(n_9484),
.A2(n_430),
.B(n_429),
.Y(n_10050)
);

INVx2_ASAP7_75t_SL g10051 ( 
.A(n_9796),
.Y(n_10051)
);

O2A1O1Ixp33_ASAP7_75t_L g10052 ( 
.A1(n_9686),
.A2(n_136),
.B(n_134),
.C(n_135),
.Y(n_10052)
);

INVx3_ASAP7_75t_L g10053 ( 
.A(n_9726),
.Y(n_10053)
);

CKINVDCx5p33_ASAP7_75t_R g10054 ( 
.A(n_9409),
.Y(n_10054)
);

AOI21xp5_ASAP7_75t_L g10055 ( 
.A1(n_9495),
.A2(n_430),
.B(n_429),
.Y(n_10055)
);

NAND2xp5_ASAP7_75t_L g10056 ( 
.A(n_9455),
.B(n_431),
.Y(n_10056)
);

NAND2xp5_ASAP7_75t_L g10057 ( 
.A(n_9338),
.B(n_432),
.Y(n_10057)
);

OAI21xp5_ASAP7_75t_L g10058 ( 
.A1(n_9382),
.A2(n_136),
.B(n_137),
.Y(n_10058)
);

NAND2xp5_ASAP7_75t_SL g10059 ( 
.A(n_9596),
.B(n_432),
.Y(n_10059)
);

OAI22x1_ASAP7_75t_L g10060 ( 
.A1(n_9339),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.Y(n_10060)
);

BUFx6f_ASAP7_75t_L g10061 ( 
.A(n_9225),
.Y(n_10061)
);

AND2x4_ASAP7_75t_L g10062 ( 
.A(n_9255),
.B(n_433),
.Y(n_10062)
);

OAI21xp33_ASAP7_75t_L g10063 ( 
.A1(n_9645),
.A2(n_138),
.B(n_139),
.Y(n_10063)
);

CKINVDCx10_ASAP7_75t_R g10064 ( 
.A(n_9517),
.Y(n_10064)
);

NOR2xp33_ASAP7_75t_L g10065 ( 
.A(n_9478),
.B(n_433),
.Y(n_10065)
);

A2O1A1Ixp33_ASAP7_75t_L g10066 ( 
.A1(n_9383),
.A2(n_435),
.B(n_436),
.C(n_434),
.Y(n_10066)
);

OAI21xp5_ASAP7_75t_L g10067 ( 
.A1(n_9399),
.A2(n_138),
.B(n_139),
.Y(n_10067)
);

AOI21xp5_ASAP7_75t_L g10068 ( 
.A1(n_9499),
.A2(n_435),
.B(n_434),
.Y(n_10068)
);

AND2x2_ASAP7_75t_L g10069 ( 
.A(n_9742),
.B(n_9765),
.Y(n_10069)
);

INVx2_ASAP7_75t_SL g10070 ( 
.A(n_9444),
.Y(n_10070)
);

AOI21xp5_ASAP7_75t_L g10071 ( 
.A1(n_9515),
.A2(n_438),
.B(n_437),
.Y(n_10071)
);

AOI21xp5_ASAP7_75t_L g10072 ( 
.A1(n_9519),
.A2(n_439),
.B(n_437),
.Y(n_10072)
);

NAND2xp5_ASAP7_75t_L g10073 ( 
.A(n_9280),
.B(n_439),
.Y(n_10073)
);

OAI22xp5_ASAP7_75t_L g10074 ( 
.A1(n_9706),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.Y(n_10074)
);

OAI22xp5_ASAP7_75t_L g10075 ( 
.A1(n_9661),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.Y(n_10075)
);

NAND2xp5_ASAP7_75t_L g10076 ( 
.A(n_9758),
.B(n_440),
.Y(n_10076)
);

A2O1A1Ixp33_ASAP7_75t_L g10077 ( 
.A1(n_9403),
.A2(n_441),
.B(n_442),
.C(n_440),
.Y(n_10077)
);

INVx1_ASAP7_75t_L g10078 ( 
.A(n_9430),
.Y(n_10078)
);

OAI21xp5_ASAP7_75t_L g10079 ( 
.A1(n_9404),
.A2(n_140),
.B(n_141),
.Y(n_10079)
);

O2A1O1Ixp5_ASAP7_75t_L g10080 ( 
.A1(n_9628),
.A2(n_9284),
.B(n_9533),
.C(n_9526),
.Y(n_10080)
);

O2A1O1Ixp33_ASAP7_75t_L g10081 ( 
.A1(n_9377),
.A2(n_144),
.B(n_142),
.C(n_143),
.Y(n_10081)
);

AOI22xp5_ASAP7_75t_L g10082 ( 
.A1(n_9355),
.A2(n_144),
.B1(n_142),
.B2(n_143),
.Y(n_10082)
);

AOI22xp5_ASAP7_75t_L g10083 ( 
.A1(n_9540),
.A2(n_146),
.B1(n_144),
.B2(n_145),
.Y(n_10083)
);

NAND2xp5_ASAP7_75t_L g10084 ( 
.A(n_9777),
.B(n_441),
.Y(n_10084)
);

INVx1_ASAP7_75t_L g10085 ( 
.A(n_9431),
.Y(n_10085)
);

AOI21x1_ASAP7_75t_L g10086 ( 
.A1(n_9591),
.A2(n_145),
.B(n_146),
.Y(n_10086)
);

INVx1_ASAP7_75t_L g10087 ( 
.A(n_9447),
.Y(n_10087)
);

INVx2_ASAP7_75t_L g10088 ( 
.A(n_9398),
.Y(n_10088)
);

A2O1A1Ixp33_ASAP7_75t_L g10089 ( 
.A1(n_9415),
.A2(n_444),
.B(n_445),
.C(n_443),
.Y(n_10089)
);

AOI21x1_ASAP7_75t_L g10090 ( 
.A1(n_9531),
.A2(n_145),
.B(n_146),
.Y(n_10090)
);

A2O1A1Ixp33_ASAP7_75t_L g10091 ( 
.A1(n_9420),
.A2(n_445),
.B(n_446),
.C(n_443),
.Y(n_10091)
);

O2A1O1Ixp33_ASAP7_75t_L g10092 ( 
.A1(n_9705),
.A2(n_149),
.B(n_147),
.C(n_148),
.Y(n_10092)
);

INVx1_ASAP7_75t_L g10093 ( 
.A(n_9452),
.Y(n_10093)
);

O2A1O1Ixp33_ASAP7_75t_L g10094 ( 
.A1(n_9424),
.A2(n_149),
.B(n_147),
.C(n_148),
.Y(n_10094)
);

BUFx2_ASAP7_75t_L g10095 ( 
.A(n_9781),
.Y(n_10095)
);

AOI21xp5_ASAP7_75t_L g10096 ( 
.A1(n_9522),
.A2(n_448),
.B(n_446),
.Y(n_10096)
);

AOI21xp5_ASAP7_75t_L g10097 ( 
.A1(n_9543),
.A2(n_450),
.B(n_449),
.Y(n_10097)
);

NOR2xp33_ASAP7_75t_L g10098 ( 
.A(n_9535),
.B(n_449),
.Y(n_10098)
);

AOI21xp5_ASAP7_75t_L g10099 ( 
.A1(n_9544),
.A2(n_452),
.B(n_450),
.Y(n_10099)
);

OAI22xp5_ASAP7_75t_L g10100 ( 
.A1(n_9585),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.Y(n_10100)
);

INVx2_ASAP7_75t_L g10101 ( 
.A(n_9407),
.Y(n_10101)
);

NAND2xp5_ASAP7_75t_L g10102 ( 
.A(n_9793),
.B(n_9287),
.Y(n_10102)
);

NAND2xp5_ASAP7_75t_L g10103 ( 
.A(n_9219),
.B(n_452),
.Y(n_10103)
);

NOR2xp33_ASAP7_75t_L g10104 ( 
.A(n_9671),
.B(n_453),
.Y(n_10104)
);

AOI21xp5_ASAP7_75t_L g10105 ( 
.A1(n_9550),
.A2(n_454),
.B(n_453),
.Y(n_10105)
);

INVx1_ASAP7_75t_SL g10106 ( 
.A(n_9457),
.Y(n_10106)
);

OAI21xp5_ASAP7_75t_L g10107 ( 
.A1(n_9421),
.A2(n_150),
.B(n_151),
.Y(n_10107)
);

BUFx12f_ASAP7_75t_L g10108 ( 
.A(n_9228),
.Y(n_10108)
);

AOI22xp33_ASAP7_75t_L g10109 ( 
.A1(n_9529),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.Y(n_10109)
);

INVxp67_ASAP7_75t_L g10110 ( 
.A(n_9326),
.Y(n_10110)
);

INVx1_ASAP7_75t_L g10111 ( 
.A(n_9460),
.Y(n_10111)
);

NAND2xp5_ASAP7_75t_L g10112 ( 
.A(n_9232),
.B(n_454),
.Y(n_10112)
);

INVx1_ASAP7_75t_SL g10113 ( 
.A(n_9442),
.Y(n_10113)
);

NOR3xp33_ASAP7_75t_L g10114 ( 
.A(n_9490),
.B(n_152),
.C(n_154),
.Y(n_10114)
);

OAI22xp5_ASAP7_75t_L g10115 ( 
.A1(n_9605),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_10115)
);

AOI21xp5_ASAP7_75t_L g10116 ( 
.A1(n_9557),
.A2(n_9433),
.B(n_9419),
.Y(n_10116)
);

O2A1O1Ixp33_ASAP7_75t_L g10117 ( 
.A1(n_9438),
.A2(n_157),
.B(n_155),
.C(n_156),
.Y(n_10117)
);

INVx1_ASAP7_75t_L g10118 ( 
.A(n_9468),
.Y(n_10118)
);

NOR2xp33_ASAP7_75t_L g10119 ( 
.A(n_9727),
.B(n_455),
.Y(n_10119)
);

OAI21xp5_ASAP7_75t_L g10120 ( 
.A1(n_9451),
.A2(n_9463),
.B(n_9454),
.Y(n_10120)
);

AOI21xp5_ASAP7_75t_L g10121 ( 
.A1(n_9439),
.A2(n_9448),
.B(n_9446),
.Y(n_10121)
);

NAND2xp5_ASAP7_75t_L g10122 ( 
.A(n_9243),
.B(n_455),
.Y(n_10122)
);

AOI21xp5_ASAP7_75t_L g10123 ( 
.A1(n_9456),
.A2(n_457),
.B(n_456),
.Y(n_10123)
);

NAND3xp33_ASAP7_75t_L g10124 ( 
.A(n_9497),
.B(n_155),
.C(n_156),
.Y(n_10124)
);

INVx1_ASAP7_75t_L g10125 ( 
.A(n_9486),
.Y(n_10125)
);

AOI21xp5_ASAP7_75t_L g10126 ( 
.A1(n_9466),
.A2(n_457),
.B(n_456),
.Y(n_10126)
);

OAI22xp33_ASAP7_75t_L g10127 ( 
.A1(n_9422),
.A2(n_459),
.B1(n_460),
.B2(n_458),
.Y(n_10127)
);

NAND2xp5_ASAP7_75t_L g10128 ( 
.A(n_9246),
.B(n_458),
.Y(n_10128)
);

AOI22xp5_ASAP7_75t_L g10129 ( 
.A1(n_9508),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.Y(n_10129)
);

INVx1_ASAP7_75t_L g10130 ( 
.A(n_9498),
.Y(n_10130)
);

A2O1A1Ixp33_ASAP7_75t_L g10131 ( 
.A1(n_9465),
.A2(n_460),
.B(n_461),
.C(n_459),
.Y(n_10131)
);

NOR2xp33_ASAP7_75t_L g10132 ( 
.A(n_9735),
.B(n_461),
.Y(n_10132)
);

NAND2xp5_ASAP7_75t_L g10133 ( 
.A(n_9250),
.B(n_462),
.Y(n_10133)
);

OAI21xp5_ASAP7_75t_L g10134 ( 
.A1(n_9489),
.A2(n_157),
.B(n_158),
.Y(n_10134)
);

OAI22xp5_ASAP7_75t_L g10135 ( 
.A1(n_9681),
.A2(n_161),
.B1(n_159),
.B2(n_160),
.Y(n_10135)
);

NOR2x1_ASAP7_75t_L g10136 ( 
.A(n_9505),
.B(n_462),
.Y(n_10136)
);

A2O1A1Ixp33_ASAP7_75t_L g10137 ( 
.A1(n_9491),
.A2(n_464),
.B(n_465),
.C(n_463),
.Y(n_10137)
);

AOI21xp5_ASAP7_75t_L g10138 ( 
.A1(n_9265),
.A2(n_464),
.B(n_463),
.Y(n_10138)
);

NAND2xp5_ASAP7_75t_L g10139 ( 
.A(n_9269),
.B(n_465),
.Y(n_10139)
);

OAI21xp33_ASAP7_75t_L g10140 ( 
.A1(n_9516),
.A2(n_159),
.B(n_160),
.Y(n_10140)
);

AOI21xp5_ASAP7_75t_L g10141 ( 
.A1(n_9271),
.A2(n_467),
.B(n_466),
.Y(n_10141)
);

NAND2xp5_ASAP7_75t_L g10142 ( 
.A(n_9276),
.B(n_466),
.Y(n_10142)
);

NAND2xp5_ASAP7_75t_L g10143 ( 
.A(n_9292),
.B(n_9305),
.Y(n_10143)
);

INVx1_ASAP7_75t_L g10144 ( 
.A(n_9503),
.Y(n_10144)
);

AOI21xp5_ASAP7_75t_L g10145 ( 
.A1(n_9307),
.A2(n_469),
.B(n_468),
.Y(n_10145)
);

O2A1O1Ixp33_ASAP7_75t_L g10146 ( 
.A1(n_9494),
.A2(n_163),
.B(n_161),
.C(n_162),
.Y(n_10146)
);

OAI321xp33_ASAP7_75t_L g10147 ( 
.A1(n_9580),
.A2(n_164),
.A3(n_166),
.B1(n_162),
.B2(n_163),
.C(n_165),
.Y(n_10147)
);

NAND2xp5_ASAP7_75t_SL g10148 ( 
.A(n_9616),
.B(n_468),
.Y(n_10148)
);

AOI21xp5_ASAP7_75t_L g10149 ( 
.A1(n_9311),
.A2(n_9691),
.B(n_9685),
.Y(n_10149)
);

A2O1A1Ixp33_ASAP7_75t_L g10150 ( 
.A1(n_9506),
.A2(n_471),
.B(n_472),
.C(n_469),
.Y(n_10150)
);

BUFx4f_ASAP7_75t_L g10151 ( 
.A(n_9504),
.Y(n_10151)
);

AOI21xp5_ASAP7_75t_L g10152 ( 
.A1(n_9511),
.A2(n_473),
.B(n_472),
.Y(n_10152)
);

NAND2xp5_ASAP7_75t_L g10153 ( 
.A(n_9323),
.B(n_473),
.Y(n_10153)
);

AOI21xp5_ASAP7_75t_L g10154 ( 
.A1(n_9530),
.A2(n_475),
.B(n_474),
.Y(n_10154)
);

NAND2xp5_ASAP7_75t_L g10155 ( 
.A(n_9324),
.B(n_474),
.Y(n_10155)
);

AND2x2_ASAP7_75t_L g10156 ( 
.A(n_9766),
.B(n_9773),
.Y(n_10156)
);

AOI21xp5_ASAP7_75t_L g10157 ( 
.A1(n_9541),
.A2(n_476),
.B(n_475),
.Y(n_10157)
);

INVx2_ASAP7_75t_L g10158 ( 
.A(n_9361),
.Y(n_10158)
);

AOI21xp5_ASAP7_75t_L g10159 ( 
.A1(n_9552),
.A2(n_478),
.B(n_477),
.Y(n_10159)
);

CKINVDCx10_ASAP7_75t_R g10160 ( 
.A(n_9334),
.Y(n_10160)
);

OAI21xp5_ASAP7_75t_L g10161 ( 
.A1(n_9510),
.A2(n_162),
.B(n_163),
.Y(n_10161)
);

NAND2xp5_ASAP7_75t_L g10162 ( 
.A(n_9327),
.B(n_477),
.Y(n_10162)
);

NAND2xp5_ASAP7_75t_L g10163 ( 
.A(n_9366),
.B(n_9375),
.Y(n_10163)
);

INVx8_ASAP7_75t_L g10164 ( 
.A(n_9387),
.Y(n_10164)
);

AOI21xp5_ASAP7_75t_L g10165 ( 
.A1(n_9559),
.A2(n_480),
.B(n_478),
.Y(n_10165)
);

O2A1O1Ixp33_ASAP7_75t_L g10166 ( 
.A1(n_9714),
.A2(n_166),
.B(n_164),
.C(n_165),
.Y(n_10166)
);

NOR2xp33_ASAP7_75t_L g10167 ( 
.A(n_9761),
.B(n_480),
.Y(n_10167)
);

INVx1_ASAP7_75t_L g10168 ( 
.A(n_9384),
.Y(n_10168)
);

AOI21x1_ASAP7_75t_L g10169 ( 
.A1(n_9589),
.A2(n_9539),
.B(n_9579),
.Y(n_10169)
);

AOI21xp5_ASAP7_75t_L g10170 ( 
.A1(n_9536),
.A2(n_482),
.B(n_481),
.Y(n_10170)
);

AOI22xp5_ASAP7_75t_L g10171 ( 
.A1(n_9425),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.Y(n_10171)
);

INVx1_ASAP7_75t_L g10172 ( 
.A(n_9385),
.Y(n_10172)
);

BUFx3_ASAP7_75t_L g10173 ( 
.A(n_9789),
.Y(n_10173)
);

NOR2xp33_ASAP7_75t_L g10174 ( 
.A(n_9238),
.B(n_481),
.Y(n_10174)
);

AOI21xp5_ASAP7_75t_L g10175 ( 
.A1(n_9525),
.A2(n_483),
.B(n_482),
.Y(n_10175)
);

NOR2xp33_ASAP7_75t_L g10176 ( 
.A(n_9520),
.B(n_483),
.Y(n_10176)
);

AND2x2_ASAP7_75t_L g10177 ( 
.A(n_9779),
.B(n_484),
.Y(n_10177)
);

NAND2xp5_ASAP7_75t_L g10178 ( 
.A(n_9386),
.B(n_485),
.Y(n_10178)
);

BUFx4f_ASAP7_75t_L g10179 ( 
.A(n_9504),
.Y(n_10179)
);

BUFx2_ASAP7_75t_L g10180 ( 
.A(n_9440),
.Y(n_10180)
);

A2O1A1Ixp33_ASAP7_75t_L g10181 ( 
.A1(n_9428),
.A2(n_486),
.B(n_487),
.C(n_485),
.Y(n_10181)
);

NOR2x1_ASAP7_75t_L g10182 ( 
.A(n_9481),
.B(n_486),
.Y(n_10182)
);

NAND2xp5_ASAP7_75t_L g10183 ( 
.A(n_9388),
.B(n_488),
.Y(n_10183)
);

AOI21xp33_ASAP7_75t_L g10184 ( 
.A1(n_9676),
.A2(n_167),
.B(n_168),
.Y(n_10184)
);

NAND2xp5_ASAP7_75t_L g10185 ( 
.A(n_9476),
.B(n_489),
.Y(n_10185)
);

AOI21xp5_ASAP7_75t_L g10186 ( 
.A1(n_9590),
.A2(n_490),
.B(n_489),
.Y(n_10186)
);

OAI22xp5_ASAP7_75t_L g10187 ( 
.A1(n_9514),
.A2(n_9715),
.B1(n_9704),
.B2(n_9723),
.Y(n_10187)
);

INVx3_ASAP7_75t_L g10188 ( 
.A(n_9444),
.Y(n_10188)
);

O2A1O1Ixp33_ASAP7_75t_L g10189 ( 
.A1(n_9308),
.A2(n_9507),
.B(n_9524),
.C(n_9523),
.Y(n_10189)
);

OAI21xp5_ASAP7_75t_L g10190 ( 
.A1(n_9252),
.A2(n_167),
.B(n_168),
.Y(n_10190)
);

INVx1_ASAP7_75t_L g10191 ( 
.A(n_9294),
.Y(n_10191)
);

OAI21xp5_ASAP7_75t_L g10192 ( 
.A1(n_9582),
.A2(n_168),
.B(n_169),
.Y(n_10192)
);

BUFx2_ASAP7_75t_L g10193 ( 
.A(n_9467),
.Y(n_10193)
);

INVx2_ASAP7_75t_L g10194 ( 
.A(n_9348),
.Y(n_10194)
);

NAND2xp5_ASAP7_75t_SL g10195 ( 
.A(n_9616),
.B(n_491),
.Y(n_10195)
);

NAND2xp5_ASAP7_75t_L g10196 ( 
.A(n_9606),
.B(n_492),
.Y(n_10196)
);

AND2x4_ASAP7_75t_L g10197 ( 
.A(n_9512),
.B(n_492),
.Y(n_10197)
);

AOI21xp5_ASAP7_75t_L g10198 ( 
.A1(n_9588),
.A2(n_9601),
.B(n_9598),
.Y(n_10198)
);

NAND2xp5_ASAP7_75t_SL g10199 ( 
.A(n_9692),
.B(n_493),
.Y(n_10199)
);

AOI21xp33_ASAP7_75t_L g10200 ( 
.A1(n_9306),
.A2(n_169),
.B(n_170),
.Y(n_10200)
);

AOI21xp5_ASAP7_75t_L g10201 ( 
.A1(n_9614),
.A2(n_494),
.B(n_493),
.Y(n_10201)
);

NAND2xp5_ASAP7_75t_L g10202 ( 
.A(n_9606),
.B(n_494),
.Y(n_10202)
);

AOI22xp5_ASAP7_75t_L g10203 ( 
.A1(n_9722),
.A2(n_171),
.B1(n_169),
.B2(n_170),
.Y(n_10203)
);

AND2x4_ASAP7_75t_L g10204 ( 
.A(n_9492),
.B(n_495),
.Y(n_10204)
);

INVx2_ASAP7_75t_L g10205 ( 
.A(n_9483),
.Y(n_10205)
);

AOI22xp33_ASAP7_75t_L g10206 ( 
.A1(n_9606),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.Y(n_10206)
);

BUFx6f_ASAP7_75t_L g10207 ( 
.A(n_9387),
.Y(n_10207)
);

NAND2xp5_ASAP7_75t_L g10208 ( 
.A(n_9214),
.B(n_497),
.Y(n_10208)
);

AOI21xp5_ASAP7_75t_L g10209 ( 
.A1(n_9623),
.A2(n_498),
.B(n_497),
.Y(n_10209)
);

AOI21xp5_ASAP7_75t_L g10210 ( 
.A1(n_9629),
.A2(n_500),
.B(n_499),
.Y(n_10210)
);

A2O1A1Ixp33_ASAP7_75t_L g10211 ( 
.A1(n_9631),
.A2(n_501),
.B(n_502),
.C(n_499),
.Y(n_10211)
);

AOI21xp5_ASAP7_75t_L g10212 ( 
.A1(n_9633),
.A2(n_503),
.B(n_502),
.Y(n_10212)
);

NAND2xp5_ASAP7_75t_L g10213 ( 
.A(n_9521),
.B(n_503),
.Y(n_10213)
);

INVx1_ASAP7_75t_L g10214 ( 
.A(n_9312),
.Y(n_10214)
);

AOI21x1_ASAP7_75t_L g10215 ( 
.A1(n_9657),
.A2(n_9658),
.B(n_9699),
.Y(n_10215)
);

OAI22xp5_ASAP7_75t_L g10216 ( 
.A1(n_9718),
.A2(n_173),
.B1(n_171),
.B2(n_172),
.Y(n_10216)
);

NOR2xp33_ASAP7_75t_L g10217 ( 
.A(n_9692),
.B(n_504),
.Y(n_10217)
);

NOR2xp33_ASAP7_75t_L g10218 ( 
.A(n_9528),
.B(n_504),
.Y(n_10218)
);

NAND2xp5_ASAP7_75t_L g10219 ( 
.A(n_9518),
.B(n_505),
.Y(n_10219)
);

NAND2xp5_ASAP7_75t_SL g10220 ( 
.A(n_9666),
.B(n_505),
.Y(n_10220)
);

NAND2xp5_ASAP7_75t_L g10221 ( 
.A(n_9555),
.B(n_506),
.Y(n_10221)
);

OAI21xp33_ASAP7_75t_L g10222 ( 
.A1(n_9502),
.A2(n_173),
.B(n_174),
.Y(n_10222)
);

OAI22xp5_ASAP7_75t_L g10223 ( 
.A1(n_9380),
.A2(n_9548),
.B1(n_9471),
.B2(n_9436),
.Y(n_10223)
);

NAND2xp5_ASAP7_75t_L g10224 ( 
.A(n_9639),
.B(n_506),
.Y(n_10224)
);

AND2x4_ASAP7_75t_SL g10225 ( 
.A(n_9767),
.B(n_507),
.Y(n_10225)
);

AOI22xp5_ASAP7_75t_L g10226 ( 
.A1(n_9696),
.A2(n_176),
.B1(n_173),
.B2(n_175),
.Y(n_10226)
);

AOI21xp5_ASAP7_75t_L g10227 ( 
.A1(n_9719),
.A2(n_509),
.B(n_508),
.Y(n_10227)
);

NAND2xp5_ASAP7_75t_SL g10228 ( 
.A(n_9666),
.B(n_509),
.Y(n_10228)
);

BUFx2_ASAP7_75t_L g10229 ( 
.A(n_9372),
.Y(n_10229)
);

BUFx6f_ASAP7_75t_L g10230 ( 
.A(n_9236),
.Y(n_10230)
);

A2O1A1Ixp33_ASAP7_75t_L g10231 ( 
.A1(n_9701),
.A2(n_9595),
.B(n_9703),
.C(n_9609),
.Y(n_10231)
);

NOR3xp33_ASAP7_75t_L g10232 ( 
.A(n_9569),
.B(n_175),
.C(n_176),
.Y(n_10232)
);

CKINVDCx10_ASAP7_75t_R g10233 ( 
.A(n_9640),
.Y(n_10233)
);

INVx2_ASAP7_75t_L g10234 ( 
.A(n_9328),
.Y(n_10234)
);

AOI21xp5_ASAP7_75t_L g10235 ( 
.A1(n_9613),
.A2(n_511),
.B(n_510),
.Y(n_10235)
);

AND2x2_ASAP7_75t_L g10236 ( 
.A(n_9783),
.B(n_510),
.Y(n_10236)
);

AND2x2_ASAP7_75t_L g10237 ( 
.A(n_9790),
.B(n_511),
.Y(n_10237)
);

NAND2xp5_ASAP7_75t_L g10238 ( 
.A(n_9619),
.B(n_512),
.Y(n_10238)
);

NAND2xp5_ASAP7_75t_L g10239 ( 
.A(n_9563),
.B(n_512),
.Y(n_10239)
);

AOI21x1_ASAP7_75t_L g10240 ( 
.A1(n_9229),
.A2(n_175),
.B(n_176),
.Y(n_10240)
);

AOI22xp5_ASAP7_75t_L g10241 ( 
.A1(n_9693),
.A2(n_179),
.B1(n_177),
.B2(n_178),
.Y(n_10241)
);

NOR2xp33_ASAP7_75t_SL g10242 ( 
.A(n_9610),
.B(n_177),
.Y(n_10242)
);

O2A1O1Ixp33_ASAP7_75t_SL g10243 ( 
.A1(n_9604),
.A2(n_9551),
.B(n_9798),
.C(n_9371),
.Y(n_10243)
);

NOR2xp33_ASAP7_75t_L g10244 ( 
.A(n_9251),
.B(n_513),
.Y(n_10244)
);

OAI21xp5_ASAP7_75t_L g10245 ( 
.A1(n_9221),
.A2(n_178),
.B(n_179),
.Y(n_10245)
);

AOI22xp33_ASAP7_75t_L g10246 ( 
.A1(n_9576),
.A2(n_180),
.B1(n_178),
.B2(n_179),
.Y(n_10246)
);

AOI21xp5_ASAP7_75t_L g10247 ( 
.A1(n_9441),
.A2(n_514),
.B(n_513),
.Y(n_10247)
);

NAND2xp5_ASAP7_75t_L g10248 ( 
.A(n_9594),
.B(n_514),
.Y(n_10248)
);

AOI21x1_ASAP7_75t_L g10249 ( 
.A1(n_9461),
.A2(n_180),
.B(n_181),
.Y(n_10249)
);

OAI21xp5_ASAP7_75t_L g10250 ( 
.A1(n_9222),
.A2(n_180),
.B(n_181),
.Y(n_10250)
);

NAND2xp5_ASAP7_75t_L g10251 ( 
.A(n_9599),
.B(n_516),
.Y(n_10251)
);

OAI22xp5_ASAP7_75t_L g10252 ( 
.A1(n_9564),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.Y(n_10252)
);

AND2x2_ASAP7_75t_L g10253 ( 
.A(n_9799),
.B(n_517),
.Y(n_10253)
);

NAND2xp5_ASAP7_75t_L g10254 ( 
.A(n_9226),
.B(n_517),
.Y(n_10254)
);

OAI21xp5_ASAP7_75t_L g10255 ( 
.A1(n_9233),
.A2(n_182),
.B(n_183),
.Y(n_10255)
);

AOI21xp5_ASAP7_75t_L g10256 ( 
.A1(n_9474),
.A2(n_520),
.B(n_518),
.Y(n_10256)
);

OAI21xp5_ASAP7_75t_L g10257 ( 
.A1(n_9482),
.A2(n_182),
.B(n_183),
.Y(n_10257)
);

NAND2xp5_ASAP7_75t_L g10258 ( 
.A(n_9330),
.B(n_518),
.Y(n_10258)
);

BUFx12f_ASAP7_75t_L g10259 ( 
.A(n_9469),
.Y(n_10259)
);

AOI21x1_ASAP7_75t_L g10260 ( 
.A1(n_9501),
.A2(n_184),
.B(n_185),
.Y(n_10260)
);

NAND2xp5_ASAP7_75t_SL g10261 ( 
.A(n_9713),
.B(n_520),
.Y(n_10261)
);

HB1xp67_ASAP7_75t_L g10262 ( 
.A(n_9464),
.Y(n_10262)
);

A2O1A1Ixp33_ASAP7_75t_L g10263 ( 
.A1(n_9602),
.A2(n_522),
.B(n_523),
.C(n_521),
.Y(n_10263)
);

OAI22xp5_ASAP7_75t_L g10264 ( 
.A1(n_9260),
.A2(n_187),
.B1(n_184),
.B2(n_186),
.Y(n_10264)
);

AOI21xp5_ASAP7_75t_L g10265 ( 
.A1(n_9603),
.A2(n_522),
.B(n_521),
.Y(n_10265)
);

AO21x1_ASAP7_75t_L g10266 ( 
.A1(n_9391),
.A2(n_9279),
.B(n_9487),
.Y(n_10266)
);

NAND2xp5_ASAP7_75t_SL g10267 ( 
.A(n_9713),
.B(n_524),
.Y(n_10267)
);

OAI22xp5_ASAP7_75t_L g10268 ( 
.A1(n_9577),
.A2(n_188),
.B1(n_186),
.B2(n_187),
.Y(n_10268)
);

AOI22xp5_ASAP7_75t_L g10269 ( 
.A1(n_9709),
.A2(n_188),
.B1(n_186),
.B2(n_187),
.Y(n_10269)
);

AOI21xp5_ASAP7_75t_L g10270 ( 
.A1(n_9683),
.A2(n_526),
.B(n_525),
.Y(n_10270)
);

AOI21xp5_ASAP7_75t_L g10271 ( 
.A1(n_9345),
.A2(n_526),
.B(n_525),
.Y(n_10271)
);

AOI21xp5_ASAP7_75t_L g10272 ( 
.A1(n_9347),
.A2(n_9356),
.B(n_9352),
.Y(n_10272)
);

INVx1_ASAP7_75t_L g10273 ( 
.A(n_9379),
.Y(n_10273)
);

NAND2xp5_ASAP7_75t_L g10274 ( 
.A(n_9381),
.B(n_9299),
.Y(n_10274)
);

AOI21xp5_ASAP7_75t_L g10275 ( 
.A1(n_9698),
.A2(n_528),
.B(n_527),
.Y(n_10275)
);

BUFx6f_ASAP7_75t_L g10276 ( 
.A(n_9389),
.Y(n_10276)
);

NAND2xp5_ASAP7_75t_L g10277 ( 
.A(n_9301),
.B(n_527),
.Y(n_10277)
);

BUFx2_ASAP7_75t_L g10278 ( 
.A(n_9285),
.Y(n_10278)
);

AOI21xp5_ASAP7_75t_L g10279 ( 
.A1(n_9263),
.A2(n_529),
.B(n_528),
.Y(n_10279)
);

NAND2xp5_ASAP7_75t_L g10280 ( 
.A(n_9396),
.B(n_530),
.Y(n_10280)
);

OAI22xp5_ASAP7_75t_L g10281 ( 
.A1(n_9227),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.Y(n_10281)
);

NAND2xp5_ASAP7_75t_L g10282 ( 
.A(n_9400),
.B(n_531),
.Y(n_10282)
);

INVx3_ASAP7_75t_L g10283 ( 
.A(n_9289),
.Y(n_10283)
);

OAI321xp33_ASAP7_75t_L g10284 ( 
.A1(n_9618),
.A2(n_191),
.A3(n_193),
.B1(n_189),
.B2(n_190),
.C(n_192),
.Y(n_10284)
);

NAND2xp5_ASAP7_75t_L g10285 ( 
.A(n_9405),
.B(n_531),
.Y(n_10285)
);

AOI21xp5_ASAP7_75t_L g10286 ( 
.A1(n_9267),
.A2(n_533),
.B(n_532),
.Y(n_10286)
);

O2A1O1Ixp33_ASAP7_75t_L g10287 ( 
.A1(n_9700),
.A2(n_192),
.B(n_190),
.C(n_191),
.Y(n_10287)
);

AOI21x1_ASAP7_75t_L g10288 ( 
.A1(n_9408),
.A2(n_191),
.B(n_192),
.Y(n_10288)
);

BUFx6f_ASAP7_75t_L g10289 ( 
.A(n_9389),
.Y(n_10289)
);

A2O1A1Ixp33_ASAP7_75t_L g10290 ( 
.A1(n_9611),
.A2(n_533),
.B(n_534),
.C(n_532),
.Y(n_10290)
);

NOR2xp33_ASAP7_75t_L g10291 ( 
.A(n_9469),
.B(n_534),
.Y(n_10291)
);

AOI21xp5_ASAP7_75t_L g10292 ( 
.A1(n_9337),
.A2(n_536),
.B(n_535),
.Y(n_10292)
);

NOR2x1_ASAP7_75t_L g10293 ( 
.A(n_9359),
.B(n_535),
.Y(n_10293)
);

NOR3xp33_ASAP7_75t_L g10294 ( 
.A(n_9556),
.B(n_9561),
.C(n_9642),
.Y(n_10294)
);

NAND2xp5_ASAP7_75t_L g10295 ( 
.A(n_9412),
.B(n_536),
.Y(n_10295)
);

NAND2xp5_ASAP7_75t_L g10296 ( 
.A(n_9413),
.B(n_537),
.Y(n_10296)
);

AOI21xp5_ASAP7_75t_L g10297 ( 
.A1(n_9432),
.A2(n_539),
.B(n_538),
.Y(n_10297)
);

O2A1O1Ixp33_ASAP7_75t_SL g10298 ( 
.A1(n_9390),
.A2(n_195),
.B(n_193),
.C(n_194),
.Y(n_10298)
);

O2A1O1Ixp33_ASAP7_75t_L g10299 ( 
.A1(n_9649),
.A2(n_195),
.B(n_193),
.C(n_194),
.Y(n_10299)
);

INVx2_ASAP7_75t_L g10300 ( 
.A(n_9401),
.Y(n_10300)
);

AND2x2_ASAP7_75t_L g10301 ( 
.A(n_9807),
.B(n_538),
.Y(n_10301)
);

AOI21x1_ASAP7_75t_L g10302 ( 
.A1(n_9437),
.A2(n_195),
.B(n_196),
.Y(n_10302)
);

NOR2xp33_ASAP7_75t_L g10303 ( 
.A(n_9401),
.B(n_540),
.Y(n_10303)
);

AOI21xp5_ASAP7_75t_L g10304 ( 
.A1(n_9445),
.A2(n_541),
.B(n_540),
.Y(n_10304)
);

NAND2xp5_ASAP7_75t_L g10305 ( 
.A(n_9453),
.B(n_541),
.Y(n_10305)
);

NAND2xp5_ASAP7_75t_L g10306 ( 
.A(n_9458),
.B(n_542),
.Y(n_10306)
);

AOI21xp5_ASAP7_75t_L g10307 ( 
.A1(n_9668),
.A2(n_543),
.B(n_542),
.Y(n_10307)
);

AOI21xp5_ASAP7_75t_L g10308 ( 
.A1(n_9712),
.A2(n_544),
.B(n_543),
.Y(n_10308)
);

NAND2xp5_ASAP7_75t_L g10309 ( 
.A(n_9808),
.B(n_544),
.Y(n_10309)
);

OAI21xp5_ASAP7_75t_L g10310 ( 
.A1(n_9620),
.A2(n_9632),
.B(n_9575),
.Y(n_10310)
);

AOI21xp5_ASAP7_75t_L g10311 ( 
.A1(n_9473),
.A2(n_546),
.B(n_545),
.Y(n_10311)
);

AND2x2_ASAP7_75t_L g10312 ( 
.A(n_9571),
.B(n_545),
.Y(n_10312)
);

NAND3xp33_ASAP7_75t_L g10313 ( 
.A(n_9593),
.B(n_196),
.C(n_197),
.Y(n_10313)
);

NAND2xp5_ASAP7_75t_L g10314 ( 
.A(n_9617),
.B(n_546),
.Y(n_10314)
);

AND2x2_ASAP7_75t_L g10315 ( 
.A(n_9677),
.B(n_9690),
.Y(n_10315)
);

AOI21xp5_ASAP7_75t_L g10316 ( 
.A1(n_9378),
.A2(n_548),
.B(n_547),
.Y(n_10316)
);

AOI21xp5_ASAP7_75t_L g10317 ( 
.A1(n_9493),
.A2(n_548),
.B(n_547),
.Y(n_10317)
);

OAI21xp5_ASAP7_75t_L g10318 ( 
.A1(n_9283),
.A2(n_196),
.B(n_197),
.Y(n_10318)
);

NOR2xp33_ASAP7_75t_L g10319 ( 
.A(n_9395),
.B(n_549),
.Y(n_10319)
);

OAI21xp5_ASAP7_75t_L g10320 ( 
.A1(n_9288),
.A2(n_197),
.B(n_198),
.Y(n_10320)
);

AOI21xp5_ASAP7_75t_L g10321 ( 
.A1(n_9264),
.A2(n_551),
.B(n_550),
.Y(n_10321)
);

AND2x2_ASAP7_75t_L g10322 ( 
.A(n_9270),
.B(n_550),
.Y(n_10322)
);

NAND2xp5_ASAP7_75t_L g10323 ( 
.A(n_9273),
.B(n_551),
.Y(n_10323)
);

OAI21x1_ASAP7_75t_L g10324 ( 
.A1(n_9293),
.A2(n_198),
.B(n_199),
.Y(n_10324)
);

BUFx8_ASAP7_75t_L g10325 ( 
.A(n_9393),
.Y(n_10325)
);

AOI22xp5_ASAP7_75t_L g10326 ( 
.A1(n_9485),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_10326)
);

NAND2xp5_ASAP7_75t_L g10327 ( 
.A(n_9274),
.B(n_552),
.Y(n_10327)
);

INVx1_ASAP7_75t_L g10328 ( 
.A(n_9344),
.Y(n_10328)
);

NAND2xp5_ASAP7_75t_L g10329 ( 
.A(n_9290),
.B(n_552),
.Y(n_10329)
);

OAI22xp5_ASAP7_75t_L g10330 ( 
.A1(n_9549),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.Y(n_10330)
);

NAND2xp5_ASAP7_75t_L g10331 ( 
.A(n_9304),
.B(n_554),
.Y(n_10331)
);

AOI21x1_ASAP7_75t_L g10332 ( 
.A1(n_9237),
.A2(n_9216),
.B(n_9242),
.Y(n_10332)
);

INVx2_ASAP7_75t_L g10333 ( 
.A(n_9393),
.Y(n_10333)
);

AOI21x1_ASAP7_75t_L g10334 ( 
.A1(n_9268),
.A2(n_9318),
.B(n_9363),
.Y(n_10334)
);

OAI21x1_ASAP7_75t_L g10335 ( 
.A1(n_9304),
.A2(n_201),
.B(n_202),
.Y(n_10335)
);

NOR3xp33_ASAP7_75t_L g10336 ( 
.A(n_9734),
.B(n_203),
.C(n_204),
.Y(n_10336)
);

O2A1O1Ixp5_ASAP7_75t_L g10337 ( 
.A1(n_9418),
.A2(n_206),
.B(n_204),
.C(n_205),
.Y(n_10337)
);

A2O1A1Ixp33_ASAP7_75t_L g10338 ( 
.A1(n_9624),
.A2(n_555),
.B(n_556),
.C(n_554),
.Y(n_10338)
);

AOI21xp5_ASAP7_75t_L g10339 ( 
.A1(n_9762),
.A2(n_557),
.B(n_556),
.Y(n_10339)
);

O2A1O1Ixp33_ASAP7_75t_L g10340 ( 
.A1(n_9775),
.A2(n_206),
.B(n_204),
.C(n_205),
.Y(n_10340)
);

OAI22xp5_ASAP7_75t_L g10341 ( 
.A1(n_9309),
.A2(n_208),
.B1(n_206),
.B2(n_207),
.Y(n_10341)
);

O2A1O1Ixp33_ASAP7_75t_L g10342 ( 
.A1(n_9281),
.A2(n_209),
.B(n_207),
.C(n_208),
.Y(n_10342)
);

NAND2xp5_ASAP7_75t_L g10343 ( 
.A(n_9296),
.B(n_558),
.Y(n_10343)
);

INVx3_ASAP7_75t_L g10344 ( 
.A(n_9212),
.Y(n_10344)
);

CKINVDCx10_ASAP7_75t_R g10345 ( 
.A(n_9409),
.Y(n_10345)
);

AOI21xp5_ASAP7_75t_L g10346 ( 
.A1(n_9406),
.A2(n_560),
.B(n_559),
.Y(n_10346)
);

INVx2_ASAP7_75t_SL g10347 ( 
.A(n_9763),
.Y(n_10347)
);

NAND2xp5_ASAP7_75t_SL g10348 ( 
.A(n_9258),
.B(n_559),
.Y(n_10348)
);

AOI21xp5_ASAP7_75t_L g10349 ( 
.A1(n_9406),
.A2(n_561),
.B(n_560),
.Y(n_10349)
);

INVx1_ASAP7_75t_L g10350 ( 
.A(n_9315),
.Y(n_10350)
);

INVx2_ASAP7_75t_L g10351 ( 
.A(n_9217),
.Y(n_10351)
);

OAI21xp33_ASAP7_75t_L g10352 ( 
.A1(n_9258),
.A2(n_208),
.B(n_209),
.Y(n_10352)
);

NAND2xp5_ASAP7_75t_L g10353 ( 
.A(n_9296),
.B(n_561),
.Y(n_10353)
);

AOI21xp5_ASAP7_75t_L g10354 ( 
.A1(n_9406),
.A2(n_563),
.B(n_562),
.Y(n_10354)
);

AOI21xp5_ASAP7_75t_L g10355 ( 
.A1(n_9406),
.A2(n_563),
.B(n_562),
.Y(n_10355)
);

NOR2xp33_ASAP7_75t_SL g10356 ( 
.A(n_9258),
.B(n_210),
.Y(n_10356)
);

A2O1A1Ixp33_ASAP7_75t_L g10357 ( 
.A1(n_9281),
.A2(n_565),
.B(n_566),
.C(n_564),
.Y(n_10357)
);

INVx3_ASAP7_75t_L g10358 ( 
.A(n_9212),
.Y(n_10358)
);

NAND2xp5_ASAP7_75t_L g10359 ( 
.A(n_9296),
.B(n_564),
.Y(n_10359)
);

NAND2xp5_ASAP7_75t_L g10360 ( 
.A(n_9296),
.B(n_565),
.Y(n_10360)
);

NAND2xp5_ASAP7_75t_L g10361 ( 
.A(n_9296),
.B(n_566),
.Y(n_10361)
);

O2A1O1Ixp5_ASAP7_75t_L g10362 ( 
.A1(n_9547),
.A2(n_213),
.B(n_211),
.C(n_212),
.Y(n_10362)
);

OAI21xp5_ASAP7_75t_L g10363 ( 
.A1(n_9258),
.A2(n_211),
.B(n_212),
.Y(n_10363)
);

NAND2xp5_ASAP7_75t_L g10364 ( 
.A(n_9296),
.B(n_567),
.Y(n_10364)
);

AOI21xp5_ASAP7_75t_L g10365 ( 
.A1(n_9406),
.A2(n_568),
.B(n_567),
.Y(n_10365)
);

OAI21xp5_ASAP7_75t_L g10366 ( 
.A1(n_9258),
.A2(n_211),
.B(n_212),
.Y(n_10366)
);

NAND2xp5_ASAP7_75t_L g10367 ( 
.A(n_9296),
.B(n_568),
.Y(n_10367)
);

NAND2xp5_ASAP7_75t_L g10368 ( 
.A(n_9296),
.B(n_569),
.Y(n_10368)
);

NAND2xp5_ASAP7_75t_SL g10369 ( 
.A(n_9258),
.B(n_569),
.Y(n_10369)
);

OAI21xp5_ASAP7_75t_L g10370 ( 
.A1(n_9258),
.A2(n_213),
.B(n_214),
.Y(n_10370)
);

NAND2xp5_ASAP7_75t_SL g10371 ( 
.A(n_9258),
.B(n_570),
.Y(n_10371)
);

NAND2xp5_ASAP7_75t_L g10372 ( 
.A(n_9296),
.B(n_571),
.Y(n_10372)
);

INVx2_ASAP7_75t_L g10373 ( 
.A(n_9217),
.Y(n_10373)
);

NAND2xp5_ASAP7_75t_L g10374 ( 
.A(n_9296),
.B(n_571),
.Y(n_10374)
);

AOI22xp5_ASAP7_75t_L g10375 ( 
.A1(n_9258),
.A2(n_215),
.B1(n_213),
.B2(n_214),
.Y(n_10375)
);

BUFx4f_ASAP7_75t_L g10376 ( 
.A(n_9218),
.Y(n_10376)
);

OAI21xp33_ASAP7_75t_L g10377 ( 
.A1(n_9258),
.A2(n_214),
.B(n_215),
.Y(n_10377)
);

NOR2xp33_ASAP7_75t_L g10378 ( 
.A(n_9500),
.B(n_572),
.Y(n_10378)
);

NAND2xp5_ASAP7_75t_L g10379 ( 
.A(n_9296),
.B(n_573),
.Y(n_10379)
);

INVx1_ASAP7_75t_L g10380 ( 
.A(n_9315),
.Y(n_10380)
);

NAND2xp5_ASAP7_75t_L g10381 ( 
.A(n_9296),
.B(n_574),
.Y(n_10381)
);

AOI22xp5_ASAP7_75t_L g10382 ( 
.A1(n_9258),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_10382)
);

BUFx4f_ASAP7_75t_L g10383 ( 
.A(n_9218),
.Y(n_10383)
);

AND2x2_ASAP7_75t_L g10384 ( 
.A(n_9314),
.B(n_575),
.Y(n_10384)
);

INVx1_ASAP7_75t_L g10385 ( 
.A(n_9315),
.Y(n_10385)
);

AOI21xp5_ASAP7_75t_L g10386 ( 
.A1(n_9406),
.A2(n_576),
.B(n_575),
.Y(n_10386)
);

AOI22xp5_ASAP7_75t_L g10387 ( 
.A1(n_9258),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_10387)
);

OAI22xp5_ASAP7_75t_L g10388 ( 
.A1(n_9258),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_10388)
);

INVx8_ASAP7_75t_L g10389 ( 
.A(n_9218),
.Y(n_10389)
);

AOI21xp5_ASAP7_75t_L g10390 ( 
.A1(n_9406),
.A2(n_578),
.B(n_577),
.Y(n_10390)
);

OAI21xp5_ASAP7_75t_L g10391 ( 
.A1(n_9258),
.A2(n_219),
.B(n_220),
.Y(n_10391)
);

NAND2xp5_ASAP7_75t_SL g10392 ( 
.A(n_9258),
.B(n_578),
.Y(n_10392)
);

AOI21xp5_ASAP7_75t_L g10393 ( 
.A1(n_9406),
.A2(n_580),
.B(n_579),
.Y(n_10393)
);

AOI22xp5_ASAP7_75t_L g10394 ( 
.A1(n_9258),
.A2(n_221),
.B1(n_219),
.B2(n_220),
.Y(n_10394)
);

O2A1O1Ixp5_ASAP7_75t_L g10395 ( 
.A1(n_9547),
.A2(n_221),
.B(n_219),
.C(n_220),
.Y(n_10395)
);

OAI21xp5_ASAP7_75t_L g10396 ( 
.A1(n_9258),
.A2(n_222),
.B(n_223),
.Y(n_10396)
);

NOR2xp33_ASAP7_75t_L g10397 ( 
.A(n_9500),
.B(n_579),
.Y(n_10397)
);

NAND2xp5_ASAP7_75t_L g10398 ( 
.A(n_9296),
.B(n_581),
.Y(n_10398)
);

OAI21xp33_ASAP7_75t_L g10399 ( 
.A1(n_9258),
.A2(n_222),
.B(n_223),
.Y(n_10399)
);

AOI21xp5_ASAP7_75t_L g10400 ( 
.A1(n_9406),
.A2(n_582),
.B(n_581),
.Y(n_10400)
);

AOI21xp5_ASAP7_75t_L g10401 ( 
.A1(n_9406),
.A2(n_583),
.B(n_582),
.Y(n_10401)
);

AOI22xp5_ASAP7_75t_L g10402 ( 
.A1(n_9258),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.Y(n_10402)
);

INVx2_ASAP7_75t_L g10403 ( 
.A(n_9217),
.Y(n_10403)
);

AO32x2_ASAP7_75t_L g10404 ( 
.A1(n_9526),
.A2(n_226),
.A3(n_224),
.B1(n_225),
.B2(n_227),
.Y(n_10404)
);

O2A1O1Ixp33_ASAP7_75t_L g10405 ( 
.A1(n_9281),
.A2(n_226),
.B(n_224),
.C(n_225),
.Y(n_10405)
);

NAND2xp5_ASAP7_75t_L g10406 ( 
.A(n_9296),
.B(n_583),
.Y(n_10406)
);

NAND3xp33_ASAP7_75t_L g10407 ( 
.A(n_9281),
.B(n_226),
.C(n_227),
.Y(n_10407)
);

AOI21xp5_ASAP7_75t_L g10408 ( 
.A1(n_9406),
.A2(n_585),
.B(n_584),
.Y(n_10408)
);

AOI21xp5_ASAP7_75t_L g10409 ( 
.A1(n_9406),
.A2(n_585),
.B(n_584),
.Y(n_10409)
);

AOI21x1_ASAP7_75t_L g10410 ( 
.A1(n_9547),
.A2(n_227),
.B(n_228),
.Y(n_10410)
);

INVx1_ASAP7_75t_L g10411 ( 
.A(n_9315),
.Y(n_10411)
);

NAND2xp5_ASAP7_75t_L g10412 ( 
.A(n_9296),
.B(n_586),
.Y(n_10412)
);

NAND2xp5_ASAP7_75t_SL g10413 ( 
.A(n_9258),
.B(n_586),
.Y(n_10413)
);

AOI21xp5_ASAP7_75t_L g10414 ( 
.A1(n_9406),
.A2(n_588),
.B(n_587),
.Y(n_10414)
);

O2A1O1Ixp33_ASAP7_75t_L g10415 ( 
.A1(n_9281),
.A2(n_230),
.B(n_228),
.C(n_229),
.Y(n_10415)
);

CKINVDCx5p33_ASAP7_75t_R g10416 ( 
.A(n_9376),
.Y(n_10416)
);

NOR3xp33_ASAP7_75t_L g10417 ( 
.A(n_9266),
.B(n_228),
.C(n_229),
.Y(n_10417)
);

CKINVDCx20_ASAP7_75t_R g10418 ( 
.A(n_9376),
.Y(n_10418)
);

O2A1O1Ixp33_ASAP7_75t_L g10419 ( 
.A1(n_9281),
.A2(n_231),
.B(n_229),
.C(n_230),
.Y(n_10419)
);

BUFx4f_ASAP7_75t_L g10420 ( 
.A(n_9218),
.Y(n_10420)
);

OAI21x1_ASAP7_75t_L g10421 ( 
.A1(n_9662),
.A2(n_231),
.B(n_232),
.Y(n_10421)
);

NAND2xp5_ASAP7_75t_L g10422 ( 
.A(n_9296),
.B(n_587),
.Y(n_10422)
);

NAND2xp5_ASAP7_75t_L g10423 ( 
.A(n_9296),
.B(n_589),
.Y(n_10423)
);

AOI21xp5_ASAP7_75t_L g10424 ( 
.A1(n_9406),
.A2(n_590),
.B(n_589),
.Y(n_10424)
);

AOI21xp5_ASAP7_75t_L g10425 ( 
.A1(n_9406),
.A2(n_592),
.B(n_591),
.Y(n_10425)
);

NAND2xp5_ASAP7_75t_L g10426 ( 
.A(n_9296),
.B(n_591),
.Y(n_10426)
);

INVx1_ASAP7_75t_L g10427 ( 
.A(n_9315),
.Y(n_10427)
);

NOR3xp33_ASAP7_75t_L g10428 ( 
.A(n_9266),
.B(n_231),
.C(n_232),
.Y(n_10428)
);

AOI21xp5_ASAP7_75t_L g10429 ( 
.A1(n_9406),
.A2(n_593),
.B(n_592),
.Y(n_10429)
);

AND2x2_ASAP7_75t_L g10430 ( 
.A(n_9314),
.B(n_593),
.Y(n_10430)
);

AND2x2_ASAP7_75t_L g10431 ( 
.A(n_9314),
.B(n_594),
.Y(n_10431)
);

AOI21x1_ASAP7_75t_L g10432 ( 
.A1(n_9547),
.A2(n_232),
.B(n_233),
.Y(n_10432)
);

OAI321xp33_ASAP7_75t_L g10433 ( 
.A1(n_9656),
.A2(n_235),
.A3(n_237),
.B1(n_233),
.B2(n_234),
.C(n_236),
.Y(n_10433)
);

A2O1A1Ixp33_ASAP7_75t_L g10434 ( 
.A1(n_9281),
.A2(n_595),
.B(n_596),
.C(n_594),
.Y(n_10434)
);

O2A1O1Ixp33_ASAP7_75t_L g10435 ( 
.A1(n_9281),
.A2(n_235),
.B(n_233),
.C(n_234),
.Y(n_10435)
);

CKINVDCx5p33_ASAP7_75t_R g10436 ( 
.A(n_9376),
.Y(n_10436)
);

AOI21xp5_ASAP7_75t_L g10437 ( 
.A1(n_9406),
.A2(n_598),
.B(n_597),
.Y(n_10437)
);

AOI21xp5_ASAP7_75t_L g10438 ( 
.A1(n_9406),
.A2(n_598),
.B(n_597),
.Y(n_10438)
);

AO21x1_ASAP7_75t_L g10439 ( 
.A1(n_9547),
.A2(n_234),
.B(n_235),
.Y(n_10439)
);

AND2x4_ASAP7_75t_L g10440 ( 
.A(n_9480),
.B(n_600),
.Y(n_10440)
);

AOI22xp5_ASAP7_75t_L g10441 ( 
.A1(n_9258),
.A2(n_238),
.B1(n_236),
.B2(n_237),
.Y(n_10441)
);

NAND2xp5_ASAP7_75t_SL g10442 ( 
.A(n_9258),
.B(n_600),
.Y(n_10442)
);

NOR2xp33_ASAP7_75t_L g10443 ( 
.A(n_9500),
.B(n_601),
.Y(n_10443)
);

NAND2xp5_ASAP7_75t_L g10444 ( 
.A(n_9296),
.B(n_601),
.Y(n_10444)
);

AOI21xp5_ASAP7_75t_L g10445 ( 
.A1(n_9406),
.A2(n_603),
.B(n_602),
.Y(n_10445)
);

INVx1_ASAP7_75t_L g10446 ( 
.A(n_9315),
.Y(n_10446)
);

O2A1O1Ixp5_ASAP7_75t_L g10447 ( 
.A1(n_9547),
.A2(n_238),
.B(n_236),
.C(n_237),
.Y(n_10447)
);

NAND2xp5_ASAP7_75t_L g10448 ( 
.A(n_9296),
.B(n_602),
.Y(n_10448)
);

O2A1O1Ixp5_ASAP7_75t_L g10449 ( 
.A1(n_9547),
.A2(n_240),
.B(n_238),
.C(n_239),
.Y(n_10449)
);

AOI21xp5_ASAP7_75t_L g10450 ( 
.A1(n_9406),
.A2(n_604),
.B(n_603),
.Y(n_10450)
);

BUFx6f_ASAP7_75t_L g10451 ( 
.A(n_9763),
.Y(n_10451)
);

NAND2xp5_ASAP7_75t_L g10452 ( 
.A(n_9296),
.B(n_604),
.Y(n_10452)
);

AO22x1_ASAP7_75t_L g10453 ( 
.A1(n_9281),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.Y(n_10453)
);

NAND2xp5_ASAP7_75t_SL g10454 ( 
.A(n_9258),
.B(n_605),
.Y(n_10454)
);

AOI22xp33_ASAP7_75t_L g10455 ( 
.A1(n_9258),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.Y(n_10455)
);

BUFx6f_ASAP7_75t_L g10456 ( 
.A(n_9763),
.Y(n_10456)
);

NAND2xp5_ASAP7_75t_L g10457 ( 
.A(n_9296),
.B(n_605),
.Y(n_10457)
);

HB1xp67_ASAP7_75t_L g10458 ( 
.A(n_9296),
.Y(n_10458)
);

AOI22xp33_ASAP7_75t_L g10459 ( 
.A1(n_9258),
.A2(n_243),
.B1(n_241),
.B2(n_242),
.Y(n_10459)
);

AOI21xp5_ASAP7_75t_L g10460 ( 
.A1(n_9406),
.A2(n_607),
.B(n_606),
.Y(n_10460)
);

AND2x2_ASAP7_75t_L g10461 ( 
.A(n_9314),
.B(n_606),
.Y(n_10461)
);

BUFx3_ASAP7_75t_L g10462 ( 
.A(n_9763),
.Y(n_10462)
);

NOR2xp33_ASAP7_75t_L g10463 ( 
.A(n_9500),
.B(n_608),
.Y(n_10463)
);

AND2x2_ASAP7_75t_L g10464 ( 
.A(n_9314),
.B(n_608),
.Y(n_10464)
);

NAND2xp5_ASAP7_75t_SL g10465 ( 
.A(n_9258),
.B(n_609),
.Y(n_10465)
);

BUFx6f_ASAP7_75t_L g10466 ( 
.A(n_9763),
.Y(n_10466)
);

INVx2_ASAP7_75t_SL g10467 ( 
.A(n_9763),
.Y(n_10467)
);

AOI21xp5_ASAP7_75t_L g10468 ( 
.A1(n_9406),
.A2(n_610),
.B(n_609),
.Y(n_10468)
);

AOI22xp5_ASAP7_75t_L g10469 ( 
.A1(n_9258),
.A2(n_244),
.B1(n_242),
.B2(n_243),
.Y(n_10469)
);

NAND2xp5_ASAP7_75t_L g10470 ( 
.A(n_9296),
.B(n_610),
.Y(n_10470)
);

NOR2xp33_ASAP7_75t_L g10471 ( 
.A(n_9500),
.B(n_611),
.Y(n_10471)
);

AOI21xp5_ASAP7_75t_L g10472 ( 
.A1(n_9406),
.A2(n_612),
.B(n_611),
.Y(n_10472)
);

NOR2xp33_ASAP7_75t_L g10473 ( 
.A(n_9500),
.B(n_612),
.Y(n_10473)
);

NOR2xp33_ASAP7_75t_L g10474 ( 
.A(n_9500),
.B(n_613),
.Y(n_10474)
);

BUFx2_ASAP7_75t_L g10475 ( 
.A(n_9296),
.Y(n_10475)
);

OAI321xp33_ASAP7_75t_L g10476 ( 
.A1(n_9656),
.A2(n_245),
.A3(n_247),
.B1(n_242),
.B2(n_244),
.C(n_246),
.Y(n_10476)
);

AND2x2_ASAP7_75t_L g10477 ( 
.A(n_9314),
.B(n_614),
.Y(n_10477)
);

INVx1_ASAP7_75t_L g10478 ( 
.A(n_9315),
.Y(n_10478)
);

INVx1_ASAP7_75t_SL g10479 ( 
.A(n_9731),
.Y(n_10479)
);

AOI21xp5_ASAP7_75t_L g10480 ( 
.A1(n_9406),
.A2(n_615),
.B(n_614),
.Y(n_10480)
);

OAI21xp5_ASAP7_75t_L g10481 ( 
.A1(n_9258),
.A2(n_245),
.B(n_246),
.Y(n_10481)
);

NOR2xp67_ASAP7_75t_L g10482 ( 
.A(n_9342),
.B(n_246),
.Y(n_10482)
);

O2A1O1Ixp5_ASAP7_75t_L g10483 ( 
.A1(n_9547),
.A2(n_249),
.B(n_247),
.C(n_248),
.Y(n_10483)
);

A2O1A1Ixp33_ASAP7_75t_L g10484 ( 
.A1(n_9281),
.A2(n_616),
.B(n_617),
.C(n_615),
.Y(n_10484)
);

AOI21x1_ASAP7_75t_L g10485 ( 
.A1(n_9547),
.A2(n_247),
.B(n_249),
.Y(n_10485)
);

AOI22xp5_ASAP7_75t_L g10486 ( 
.A1(n_9258),
.A2(n_251),
.B1(n_249),
.B2(n_250),
.Y(n_10486)
);

INVx4_ASAP7_75t_L g10487 ( 
.A(n_9763),
.Y(n_10487)
);

NOR2xp67_ASAP7_75t_L g10488 ( 
.A(n_9342),
.B(n_250),
.Y(n_10488)
);

AOI22xp33_ASAP7_75t_L g10489 ( 
.A1(n_9258),
.A2(n_252),
.B1(n_250),
.B2(n_251),
.Y(n_10489)
);

OAI21xp5_ASAP7_75t_L g10490 ( 
.A1(n_9258),
.A2(n_251),
.B(n_252),
.Y(n_10490)
);

NAND2xp5_ASAP7_75t_L g10491 ( 
.A(n_9296),
.B(n_616),
.Y(n_10491)
);

INVx1_ASAP7_75t_L g10492 ( 
.A(n_9315),
.Y(n_10492)
);

AOI21xp5_ASAP7_75t_L g10493 ( 
.A1(n_9406),
.A2(n_619),
.B(n_618),
.Y(n_10493)
);

NOR2xp33_ASAP7_75t_L g10494 ( 
.A(n_9500),
.B(n_618),
.Y(n_10494)
);

O2A1O1Ixp33_ASAP7_75t_L g10495 ( 
.A1(n_9281),
.A2(n_254),
.B(n_252),
.C(n_253),
.Y(n_10495)
);

BUFx6f_ASAP7_75t_L g10496 ( 
.A(n_9763),
.Y(n_10496)
);

A2O1A1Ixp33_ASAP7_75t_L g10497 ( 
.A1(n_9281),
.A2(n_621),
.B(n_622),
.C(n_620),
.Y(n_10497)
);

BUFx6f_ASAP7_75t_L g10498 ( 
.A(n_9763),
.Y(n_10498)
);

OAI21xp5_ASAP7_75t_L g10499 ( 
.A1(n_9258),
.A2(n_253),
.B(n_254),
.Y(n_10499)
);

NOR2xp33_ASAP7_75t_L g10500 ( 
.A(n_9500),
.B(n_620),
.Y(n_10500)
);

BUFx3_ASAP7_75t_L g10501 ( 
.A(n_9763),
.Y(n_10501)
);

NAND2xp5_ASAP7_75t_L g10502 ( 
.A(n_9296),
.B(n_621),
.Y(n_10502)
);

A2O1A1Ixp33_ASAP7_75t_L g10503 ( 
.A1(n_9281),
.A2(n_624),
.B(n_625),
.C(n_622),
.Y(n_10503)
);

NAND2xp5_ASAP7_75t_L g10504 ( 
.A(n_9296),
.B(n_624),
.Y(n_10504)
);

INVx2_ASAP7_75t_L g10505 ( 
.A(n_9217),
.Y(n_10505)
);

NAND2xp5_ASAP7_75t_L g10506 ( 
.A(n_9296),
.B(n_625),
.Y(n_10506)
);

NOR2xp33_ASAP7_75t_L g10507 ( 
.A(n_9500),
.B(n_626),
.Y(n_10507)
);

INVx11_ASAP7_75t_L g10508 ( 
.A(n_9747),
.Y(n_10508)
);

NOR2x1p5_ASAP7_75t_SL g10509 ( 
.A(n_9662),
.B(n_626),
.Y(n_10509)
);

INVx1_ASAP7_75t_L g10510 ( 
.A(n_9315),
.Y(n_10510)
);

NAND2xp5_ASAP7_75t_L g10511 ( 
.A(n_9296),
.B(n_627),
.Y(n_10511)
);

AOI22xp33_ASAP7_75t_L g10512 ( 
.A1(n_9258),
.A2(n_256),
.B1(n_254),
.B2(n_255),
.Y(n_10512)
);

AOI21xp5_ASAP7_75t_L g10513 ( 
.A1(n_9406),
.A2(n_628),
.B(n_627),
.Y(n_10513)
);

O2A1O1Ixp5_ASAP7_75t_L g10514 ( 
.A1(n_9547),
.A2(n_257),
.B(n_255),
.C(n_256),
.Y(n_10514)
);

OAI21xp5_ASAP7_75t_L g10515 ( 
.A1(n_9258),
.A2(n_255),
.B(n_257),
.Y(n_10515)
);

AND2x2_ASAP7_75t_L g10516 ( 
.A(n_9314),
.B(n_629),
.Y(n_10516)
);

AOI21xp5_ASAP7_75t_L g10517 ( 
.A1(n_9406),
.A2(n_631),
.B(n_630),
.Y(n_10517)
);

AOI21xp5_ASAP7_75t_L g10518 ( 
.A1(n_9406),
.A2(n_632),
.B(n_631),
.Y(n_10518)
);

BUFx6f_ASAP7_75t_L g10519 ( 
.A(n_9763),
.Y(n_10519)
);

O2A1O1Ixp33_ASAP7_75t_L g10520 ( 
.A1(n_9281),
.A2(n_259),
.B(n_257),
.C(n_258),
.Y(n_10520)
);

NAND2xp5_ASAP7_75t_L g10521 ( 
.A(n_9296),
.B(n_632),
.Y(n_10521)
);

NOR2xp33_ASAP7_75t_L g10522 ( 
.A(n_9500),
.B(n_633),
.Y(n_10522)
);

OAI21xp5_ASAP7_75t_L g10523 ( 
.A1(n_9258),
.A2(n_258),
.B(n_259),
.Y(n_10523)
);

AOI21xp5_ASAP7_75t_L g10524 ( 
.A1(n_9406),
.A2(n_634),
.B(n_633),
.Y(n_10524)
);

OAI21xp5_ASAP7_75t_L g10525 ( 
.A1(n_9258),
.A2(n_259),
.B(n_260),
.Y(n_10525)
);

OAI22xp5_ASAP7_75t_L g10526 ( 
.A1(n_9258),
.A2(n_262),
.B1(n_260),
.B2(n_261),
.Y(n_10526)
);

AOI21xp5_ASAP7_75t_L g10527 ( 
.A1(n_9406),
.A2(n_635),
.B(n_634),
.Y(n_10527)
);

OAI22xp5_ASAP7_75t_L g10528 ( 
.A1(n_9258),
.A2(n_262),
.B1(n_260),
.B2(n_261),
.Y(n_10528)
);

AOI21xp5_ASAP7_75t_L g10529 ( 
.A1(n_9406),
.A2(n_636),
.B(n_635),
.Y(n_10529)
);

AOI21xp5_ASAP7_75t_L g10530 ( 
.A1(n_9406),
.A2(n_638),
.B(n_637),
.Y(n_10530)
);

INVx1_ASAP7_75t_L g10531 ( 
.A(n_9315),
.Y(n_10531)
);

OR2x6_ASAP7_75t_L g10532 ( 
.A(n_9459),
.B(n_637),
.Y(n_10532)
);

AOI21xp5_ASAP7_75t_L g10533 ( 
.A1(n_9406),
.A2(n_640),
.B(n_639),
.Y(n_10533)
);

A2O1A1Ixp33_ASAP7_75t_L g10534 ( 
.A1(n_9281),
.A2(n_642),
.B(n_643),
.C(n_641),
.Y(n_10534)
);

INVx1_ASAP7_75t_L g10535 ( 
.A(n_9315),
.Y(n_10535)
);

OAI21xp5_ASAP7_75t_L g10536 ( 
.A1(n_9258),
.A2(n_261),
.B(n_262),
.Y(n_10536)
);

NAND2xp5_ASAP7_75t_SL g10537 ( 
.A(n_9258),
.B(n_642),
.Y(n_10537)
);

AOI22xp5_ASAP7_75t_L g10538 ( 
.A1(n_9258),
.A2(n_265),
.B1(n_263),
.B2(n_264),
.Y(n_10538)
);

INVx3_ASAP7_75t_L g10539 ( 
.A(n_9940),
.Y(n_10539)
);

AND2x4_ASAP7_75t_L g10540 ( 
.A(n_9848),
.B(n_643),
.Y(n_10540)
);

OAI22xp5_ASAP7_75t_SL g10541 ( 
.A1(n_9837),
.A2(n_265),
.B1(n_263),
.B2(n_264),
.Y(n_10541)
);

AOI21xp5_ASAP7_75t_L g10542 ( 
.A1(n_9885),
.A2(n_9856),
.B(n_9816),
.Y(n_10542)
);

NAND2xp5_ASAP7_75t_L g10543 ( 
.A(n_10458),
.B(n_644),
.Y(n_10543)
);

INVx3_ASAP7_75t_L g10544 ( 
.A(n_10028),
.Y(n_10544)
);

INVx1_ASAP7_75t_L g10545 ( 
.A(n_9815),
.Y(n_10545)
);

CKINVDCx5p33_ASAP7_75t_R g10546 ( 
.A(n_10345),
.Y(n_10546)
);

A2O1A1Ixp33_ASAP7_75t_L g10547 ( 
.A1(n_9913),
.A2(n_645),
.B(n_646),
.C(n_644),
.Y(n_10547)
);

INVx1_ASAP7_75t_L g10548 ( 
.A(n_9824),
.Y(n_10548)
);

OAI22xp5_ASAP7_75t_L g10549 ( 
.A1(n_9881),
.A2(n_266),
.B1(n_263),
.B2(n_264),
.Y(n_10549)
);

NAND2xp5_ASAP7_75t_L g10550 ( 
.A(n_9945),
.B(n_645),
.Y(n_10550)
);

AOI21xp5_ASAP7_75t_L g10551 ( 
.A1(n_9888),
.A2(n_266),
.B(n_267),
.Y(n_10551)
);

O2A1O1Ixp33_ASAP7_75t_L g10552 ( 
.A1(n_10534),
.A2(n_268),
.B(n_266),
.C(n_267),
.Y(n_10552)
);

INVx2_ASAP7_75t_SL g10553 ( 
.A(n_10164),
.Y(n_10553)
);

INVx2_ASAP7_75t_L g10554 ( 
.A(n_10088),
.Y(n_10554)
);

OAI22xp5_ASAP7_75t_L g10555 ( 
.A1(n_9881),
.A2(n_269),
.B1(n_267),
.B2(n_268),
.Y(n_10555)
);

O2A1O1Ixp33_ASAP7_75t_L g10556 ( 
.A1(n_10357),
.A2(n_270),
.B(n_268),
.C(n_269),
.Y(n_10556)
);

NAND2xp5_ASAP7_75t_L g10557 ( 
.A(n_10475),
.B(n_646),
.Y(n_10557)
);

NOR2xp33_ASAP7_75t_L g10558 ( 
.A(n_10479),
.B(n_647),
.Y(n_10558)
);

BUFx6f_ASAP7_75t_L g10559 ( 
.A(n_10451),
.Y(n_10559)
);

NAND2xp5_ASAP7_75t_L g10560 ( 
.A(n_10022),
.B(n_10194),
.Y(n_10560)
);

INVx2_ASAP7_75t_L g10561 ( 
.A(n_10101),
.Y(n_10561)
);

NAND2xp5_ASAP7_75t_L g10562 ( 
.A(n_9939),
.B(n_647),
.Y(n_10562)
);

NAND3xp33_ASAP7_75t_SL g10563 ( 
.A(n_10356),
.B(n_269),
.C(n_270),
.Y(n_10563)
);

NAND2xp5_ASAP7_75t_L g10564 ( 
.A(n_9908),
.B(n_648),
.Y(n_10564)
);

AND2x4_ASAP7_75t_L g10565 ( 
.A(n_9847),
.B(n_649),
.Y(n_10565)
);

AOI21xp5_ASAP7_75t_L g10566 ( 
.A1(n_9881),
.A2(n_271),
.B(n_272),
.Y(n_10566)
);

INVx5_ASAP7_75t_L g10567 ( 
.A(n_10532),
.Y(n_10567)
);

BUFx6f_ASAP7_75t_L g10568 ( 
.A(n_10451),
.Y(n_10568)
);

A2O1A1Ixp33_ASAP7_75t_L g10569 ( 
.A1(n_10363),
.A2(n_650),
.B(n_652),
.C(n_649),
.Y(n_10569)
);

BUFx2_ASAP7_75t_L g10570 ( 
.A(n_10095),
.Y(n_10570)
);

BUFx2_ASAP7_75t_L g10571 ( 
.A(n_10180),
.Y(n_10571)
);

NAND2xp5_ASAP7_75t_SL g10572 ( 
.A(n_9935),
.B(n_653),
.Y(n_10572)
);

AND2x2_ASAP7_75t_L g10573 ( 
.A(n_10315),
.B(n_653),
.Y(n_10573)
);

AOI21xp5_ASAP7_75t_L g10574 ( 
.A1(n_9889),
.A2(n_271),
.B(n_272),
.Y(n_10574)
);

HB1xp67_ASAP7_75t_L g10575 ( 
.A(n_9923),
.Y(n_10575)
);

O2A1O1Ixp33_ASAP7_75t_L g10576 ( 
.A1(n_10434),
.A2(n_274),
.B(n_271),
.C(n_273),
.Y(n_10576)
);

INVx2_ASAP7_75t_SL g10577 ( 
.A(n_10164),
.Y(n_10577)
);

AOI22xp33_ASAP7_75t_L g10578 ( 
.A1(n_9835),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.Y(n_10578)
);

NOR2xp67_ASAP7_75t_SL g10579 ( 
.A(n_10407),
.B(n_273),
.Y(n_10579)
);

BUFx6f_ASAP7_75t_L g10580 ( 
.A(n_10451),
.Y(n_10580)
);

INVxp67_ASAP7_75t_L g10581 ( 
.A(n_10262),
.Y(n_10581)
);

AOI21xp5_ASAP7_75t_L g10582 ( 
.A1(n_9926),
.A2(n_9877),
.B(n_9860),
.Y(n_10582)
);

A2O1A1Ixp33_ASAP7_75t_L g10583 ( 
.A1(n_10366),
.A2(n_655),
.B(n_656),
.C(n_654),
.Y(n_10583)
);

BUFx2_ASAP7_75t_L g10584 ( 
.A(n_10193),
.Y(n_10584)
);

A2O1A1Ixp33_ASAP7_75t_L g10585 ( 
.A1(n_10370),
.A2(n_655),
.B(n_657),
.C(n_654),
.Y(n_10585)
);

NAND2xp5_ASAP7_75t_L g10586 ( 
.A(n_9827),
.B(n_657),
.Y(n_10586)
);

INVx1_ASAP7_75t_L g10587 ( 
.A(n_9851),
.Y(n_10587)
);

INVx1_ASAP7_75t_L g10588 ( 
.A(n_9867),
.Y(n_10588)
);

OR2x6_ASAP7_75t_L g10589 ( 
.A(n_10532),
.B(n_658),
.Y(n_10589)
);

AOI21xp5_ASAP7_75t_L g10590 ( 
.A1(n_10198),
.A2(n_9866),
.B(n_10116),
.Y(n_10590)
);

BUFx3_ASAP7_75t_L g10591 ( 
.A(n_10325),
.Y(n_10591)
);

BUFx2_ASAP7_75t_L g10592 ( 
.A(n_10229),
.Y(n_10592)
);

NOR2xp67_ASAP7_75t_L g10593 ( 
.A(n_10149),
.B(n_275),
.Y(n_10593)
);

NOR2xp33_ASAP7_75t_L g10594 ( 
.A(n_9883),
.B(n_659),
.Y(n_10594)
);

NOR3xp33_ASAP7_75t_SL g10595 ( 
.A(n_9974),
.B(n_275),
.C(n_276),
.Y(n_10595)
);

NOR2xp33_ASAP7_75t_R g10596 ( 
.A(n_10418),
.B(n_276),
.Y(n_10596)
);

BUFx8_ASAP7_75t_SL g10597 ( 
.A(n_9819),
.Y(n_10597)
);

NOR2xp33_ASAP7_75t_L g10598 ( 
.A(n_9948),
.B(n_659),
.Y(n_10598)
);

INVx2_ASAP7_75t_L g10599 ( 
.A(n_9873),
.Y(n_10599)
);

OAI22xp5_ASAP7_75t_L g10600 ( 
.A1(n_9822),
.A2(n_278),
.B1(n_276),
.B2(n_277),
.Y(n_10600)
);

CKINVDCx5p33_ASAP7_75t_R g10601 ( 
.A(n_10416),
.Y(n_10601)
);

CKINVDCx20_ASAP7_75t_R g10602 ( 
.A(n_9899),
.Y(n_10602)
);

A2O1A1Ixp33_ASAP7_75t_L g10603 ( 
.A1(n_10391),
.A2(n_661),
.B(n_662),
.C(n_660),
.Y(n_10603)
);

A2O1A1Ixp33_ASAP7_75t_L g10604 ( 
.A1(n_10396),
.A2(n_661),
.B(n_662),
.C(n_660),
.Y(n_10604)
);

AOI21xp5_ASAP7_75t_L g10605 ( 
.A1(n_10121),
.A2(n_277),
.B(n_278),
.Y(n_10605)
);

OAI22xp5_ASAP7_75t_L g10606 ( 
.A1(n_10030),
.A2(n_279),
.B1(n_277),
.B2(n_278),
.Y(n_10606)
);

NAND2xp5_ASAP7_75t_L g10607 ( 
.A(n_10102),
.B(n_663),
.Y(n_10607)
);

NAND2xp5_ASAP7_75t_SL g10608 ( 
.A(n_10080),
.B(n_664),
.Y(n_10608)
);

OAI21xp5_ASAP7_75t_L g10609 ( 
.A1(n_9972),
.A2(n_279),
.B(n_280),
.Y(n_10609)
);

A2O1A1Ixp33_ASAP7_75t_L g10610 ( 
.A1(n_10481),
.A2(n_665),
.B(n_666),
.C(n_664),
.Y(n_10610)
);

INVx1_ASAP7_75t_L g10611 ( 
.A(n_9880),
.Y(n_10611)
);

HB1xp67_ASAP7_75t_L g10612 ( 
.A(n_9892),
.Y(n_10612)
);

NAND2xp5_ASAP7_75t_L g10613 ( 
.A(n_10110),
.B(n_665),
.Y(n_10613)
);

NAND2xp5_ASAP7_75t_L g10614 ( 
.A(n_9891),
.B(n_667),
.Y(n_10614)
);

BUFx2_ASAP7_75t_L g10615 ( 
.A(n_10205),
.Y(n_10615)
);

NAND2xp5_ASAP7_75t_L g10616 ( 
.A(n_10047),
.B(n_667),
.Y(n_10616)
);

AND2x2_ASAP7_75t_L g10617 ( 
.A(n_10069),
.B(n_668),
.Y(n_10617)
);

NAND2xp5_ASAP7_75t_L g10618 ( 
.A(n_9955),
.B(n_668),
.Y(n_10618)
);

BUFx12f_ASAP7_75t_L g10619 ( 
.A(n_10456),
.Y(n_10619)
);

NOR2xp33_ASAP7_75t_L g10620 ( 
.A(n_10436),
.B(n_669),
.Y(n_10620)
);

O2A1O1Ixp33_ASAP7_75t_L g10621 ( 
.A1(n_10484),
.A2(n_281),
.B(n_279),
.C(n_280),
.Y(n_10621)
);

A2O1A1Ixp33_ASAP7_75t_L g10622 ( 
.A1(n_10490),
.A2(n_670),
.B(n_671),
.C(n_669),
.Y(n_10622)
);

INVx1_ASAP7_75t_L g10623 ( 
.A(n_9905),
.Y(n_10623)
);

AOI21xp33_ASAP7_75t_L g10624 ( 
.A1(n_9909),
.A2(n_280),
.B(n_281),
.Y(n_10624)
);

INVx2_ASAP7_75t_L g10625 ( 
.A(n_9912),
.Y(n_10625)
);

NAND2xp5_ASAP7_75t_SL g10626 ( 
.A(n_10037),
.B(n_670),
.Y(n_10626)
);

NOR2xp33_ASAP7_75t_L g10627 ( 
.A(n_9983),
.B(n_671),
.Y(n_10627)
);

AOI21xp5_ASAP7_75t_L g10628 ( 
.A1(n_10009),
.A2(n_281),
.B(n_282),
.Y(n_10628)
);

NAND2xp5_ASAP7_75t_L g10629 ( 
.A(n_10191),
.B(n_672),
.Y(n_10629)
);

INVx3_ASAP7_75t_L g10630 ( 
.A(n_10173),
.Y(n_10630)
);

CKINVDCx5p33_ASAP7_75t_R g10631 ( 
.A(n_9813),
.Y(n_10631)
);

BUFx6f_ASAP7_75t_L g10632 ( 
.A(n_10456),
.Y(n_10632)
);

O2A1O1Ixp33_ASAP7_75t_L g10633 ( 
.A1(n_10497),
.A2(n_284),
.B(n_282),
.C(n_283),
.Y(n_10633)
);

NAND2xp5_ASAP7_75t_L g10634 ( 
.A(n_9976),
.B(n_10168),
.Y(n_10634)
);

OAI22xp5_ASAP7_75t_L g10635 ( 
.A1(n_10044),
.A2(n_10082),
.B1(n_10326),
.B2(n_10109),
.Y(n_10635)
);

BUFx12f_ASAP7_75t_SL g10636 ( 
.A(n_10456),
.Y(n_10636)
);

AND2x2_ASAP7_75t_L g10637 ( 
.A(n_10156),
.B(n_672),
.Y(n_10637)
);

AOI21xp5_ASAP7_75t_L g10638 ( 
.A1(n_9857),
.A2(n_282),
.B(n_283),
.Y(n_10638)
);

O2A1O1Ixp5_ASAP7_75t_SL g10639 ( 
.A1(n_9830),
.A2(n_285),
.B(n_283),
.C(n_284),
.Y(n_10639)
);

NOR2x1_ASAP7_75t_L g10640 ( 
.A(n_10187),
.B(n_673),
.Y(n_10640)
);

NOR2xp33_ASAP7_75t_L g10641 ( 
.A(n_10106),
.B(n_673),
.Y(n_10641)
);

INVx2_ASAP7_75t_L g10642 ( 
.A(n_9934),
.Y(n_10642)
);

NAND2xp5_ASAP7_75t_L g10643 ( 
.A(n_10172),
.B(n_674),
.Y(n_10643)
);

AND2x4_ASAP7_75t_L g10644 ( 
.A(n_10039),
.B(n_675),
.Y(n_10644)
);

O2A1O1Ixp5_ASAP7_75t_L g10645 ( 
.A1(n_10453),
.A2(n_286),
.B(n_284),
.C(n_285),
.Y(n_10645)
);

AOI21xp5_ASAP7_75t_L g10646 ( 
.A1(n_10433),
.A2(n_285),
.B(n_286),
.Y(n_10646)
);

AOI21xp5_ASAP7_75t_L g10647 ( 
.A1(n_10476),
.A2(n_287),
.B(n_288),
.Y(n_10647)
);

INVx3_ASAP7_75t_L g10648 ( 
.A(n_9834),
.Y(n_10648)
);

OR2x4_ASAP7_75t_L g10649 ( 
.A(n_9960),
.B(n_287),
.Y(n_10649)
);

AOI21xp5_ASAP7_75t_L g10650 ( 
.A1(n_9814),
.A2(n_287),
.B(n_288),
.Y(n_10650)
);

NAND2xp5_ASAP7_75t_SL g10651 ( 
.A(n_10037),
.B(n_675),
.Y(n_10651)
);

AOI21xp5_ASAP7_75t_L g10652 ( 
.A1(n_9839),
.A2(n_288),
.B(n_289),
.Y(n_10652)
);

INVx2_ASAP7_75t_L g10653 ( 
.A(n_9936),
.Y(n_10653)
);

INVx1_ASAP7_75t_SL g10654 ( 
.A(n_10278),
.Y(n_10654)
);

AOI21xp5_ASAP7_75t_L g10655 ( 
.A1(n_9863),
.A2(n_289),
.B(n_290),
.Y(n_10655)
);

AOI21xp5_ASAP7_75t_L g10656 ( 
.A1(n_9868),
.A2(n_289),
.B(n_290),
.Y(n_10656)
);

NAND2xp5_ASAP7_75t_SL g10657 ( 
.A(n_10037),
.B(n_676),
.Y(n_10657)
);

NAND2xp5_ASAP7_75t_L g10658 ( 
.A(n_10113),
.B(n_676),
.Y(n_10658)
);

NAND2xp5_ASAP7_75t_L g10659 ( 
.A(n_9852),
.B(n_677),
.Y(n_10659)
);

BUFx6f_ASAP7_75t_L g10660 ( 
.A(n_10466),
.Y(n_10660)
);

BUFx2_ASAP7_75t_SL g10661 ( 
.A(n_9999),
.Y(n_10661)
);

INVx1_ASAP7_75t_SL g10662 ( 
.A(n_9902),
.Y(n_10662)
);

NOR2xp33_ASAP7_75t_L g10663 ( 
.A(n_10053),
.B(n_677),
.Y(n_10663)
);

BUFx2_ASAP7_75t_L g10664 ( 
.A(n_10259),
.Y(n_10664)
);

OAI22xp5_ASAP7_75t_L g10665 ( 
.A1(n_10455),
.A2(n_292),
.B1(n_290),
.B2(n_291),
.Y(n_10665)
);

INVx2_ASAP7_75t_L g10666 ( 
.A(n_9956),
.Y(n_10666)
);

INVxp67_ASAP7_75t_L g10667 ( 
.A(n_10300),
.Y(n_10667)
);

NOR2xp33_ASAP7_75t_L g10668 ( 
.A(n_10003),
.B(n_678),
.Y(n_10668)
);

O2A1O1Ixp33_ASAP7_75t_L g10669 ( 
.A1(n_10503),
.A2(n_293),
.B(n_291),
.C(n_292),
.Y(n_10669)
);

INVx3_ASAP7_75t_L g10670 ( 
.A(n_9834),
.Y(n_10670)
);

NAND2xp5_ASAP7_75t_L g10671 ( 
.A(n_9865),
.B(n_679),
.Y(n_10671)
);

CKINVDCx8_ASAP7_75t_R g10672 ( 
.A(n_10064),
.Y(n_10672)
);

AOI21xp5_ASAP7_75t_L g10673 ( 
.A1(n_9870),
.A2(n_291),
.B(n_292),
.Y(n_10673)
);

AOI21xp5_ASAP7_75t_L g10674 ( 
.A1(n_9820),
.A2(n_293),
.B(n_294),
.Y(n_10674)
);

O2A1O1Ixp33_ASAP7_75t_L g10675 ( 
.A1(n_10342),
.A2(n_295),
.B(n_293),
.C(n_294),
.Y(n_10675)
);

AND2x2_ASAP7_75t_L g10676 ( 
.A(n_10234),
.B(n_680),
.Y(n_10676)
);

BUFx6f_ASAP7_75t_L g10677 ( 
.A(n_10466),
.Y(n_10677)
);

NAND2xp5_ASAP7_75t_L g10678 ( 
.A(n_9910),
.B(n_680),
.Y(n_10678)
);

AOI21xp5_ASAP7_75t_L g10679 ( 
.A1(n_10043),
.A2(n_294),
.B(n_295),
.Y(n_10679)
);

OR2x6_ASAP7_75t_L g10680 ( 
.A(n_10025),
.B(n_681),
.Y(n_10680)
);

INVx2_ASAP7_75t_L g10681 ( 
.A(n_9965),
.Y(n_10681)
);

INVx2_ASAP7_75t_L g10682 ( 
.A(n_10004),
.Y(n_10682)
);

OAI22xp5_ASAP7_75t_L g10683 ( 
.A1(n_10459),
.A2(n_297),
.B1(n_295),
.B2(n_296),
.Y(n_10683)
);

OA21x2_ASAP7_75t_L g10684 ( 
.A1(n_10421),
.A2(n_9958),
.B(n_9937),
.Y(n_10684)
);

O2A1O1Ixp33_ASAP7_75t_L g10685 ( 
.A1(n_10405),
.A2(n_10415),
.B(n_10435),
.C(n_10419),
.Y(n_10685)
);

INVx1_ASAP7_75t_L g10686 ( 
.A(n_10021),
.Y(n_10686)
);

A2O1A1Ixp33_ASAP7_75t_L g10687 ( 
.A1(n_10499),
.A2(n_682),
.B(n_683),
.C(n_681),
.Y(n_10687)
);

INVx1_ASAP7_75t_L g10688 ( 
.A(n_10045),
.Y(n_10688)
);

NAND2xp5_ASAP7_75t_L g10689 ( 
.A(n_9929),
.B(n_682),
.Y(n_10689)
);

INVx1_ASAP7_75t_L g10690 ( 
.A(n_10078),
.Y(n_10690)
);

AOI21xp5_ASAP7_75t_L g10691 ( 
.A1(n_9897),
.A2(n_296),
.B(n_297),
.Y(n_10691)
);

NOR2xp33_ASAP7_75t_SL g10692 ( 
.A(n_10487),
.B(n_296),
.Y(n_10692)
);

NAND2xp5_ASAP7_75t_L g10693 ( 
.A(n_9942),
.B(n_683),
.Y(n_10693)
);

NAND2xp5_ASAP7_75t_L g10694 ( 
.A(n_9987),
.B(n_684),
.Y(n_10694)
);

CKINVDCx5p33_ASAP7_75t_R g10695 ( 
.A(n_10508),
.Y(n_10695)
);

INVx2_ASAP7_75t_L g10696 ( 
.A(n_10085),
.Y(n_10696)
);

INVx5_ASAP7_75t_SL g10697 ( 
.A(n_10466),
.Y(n_10697)
);

INVx1_ASAP7_75t_L g10698 ( 
.A(n_10087),
.Y(n_10698)
);

O2A1O1Ixp33_ASAP7_75t_SL g10699 ( 
.A1(n_9933),
.A2(n_299),
.B(n_297),
.C(n_298),
.Y(n_10699)
);

NAND2x1p5_ASAP7_75t_L g10700 ( 
.A(n_10283),
.B(n_684),
.Y(n_10700)
);

NAND2xp5_ASAP7_75t_SL g10701 ( 
.A(n_10037),
.B(n_685),
.Y(n_10701)
);

NOR2xp33_ASAP7_75t_L g10702 ( 
.A(n_10274),
.B(n_685),
.Y(n_10702)
);

OAI22xp5_ASAP7_75t_L g10703 ( 
.A1(n_10489),
.A2(n_300),
.B1(n_298),
.B2(n_299),
.Y(n_10703)
);

AOI21xp5_ASAP7_75t_L g10704 ( 
.A1(n_9904),
.A2(n_299),
.B(n_300),
.Y(n_10704)
);

OR2x2_ASAP7_75t_L g10705 ( 
.A(n_10093),
.B(n_687),
.Y(n_10705)
);

NOR2xp33_ASAP7_75t_L g10706 ( 
.A(n_10223),
.B(n_687),
.Y(n_10706)
);

AOI21x1_ASAP7_75t_SL g10707 ( 
.A1(n_10196),
.A2(n_689),
.B(n_688),
.Y(n_10707)
);

AND2x4_ASAP7_75t_L g10708 ( 
.A(n_10333),
.B(n_688),
.Y(n_10708)
);

INVx3_ASAP7_75t_L g10709 ( 
.A(n_9869),
.Y(n_10709)
);

AOI21xp5_ASAP7_75t_L g10710 ( 
.A1(n_10120),
.A2(n_300),
.B(n_301),
.Y(n_10710)
);

NAND2xp5_ASAP7_75t_L g10711 ( 
.A(n_9991),
.B(n_689),
.Y(n_10711)
);

INVx1_ASAP7_75t_L g10712 ( 
.A(n_10111),
.Y(n_10712)
);

NAND2xp5_ASAP7_75t_SL g10713 ( 
.A(n_9993),
.B(n_690),
.Y(n_10713)
);

OR2x2_ASAP7_75t_L g10714 ( 
.A(n_10118),
.B(n_691),
.Y(n_10714)
);

AOI21x1_ASAP7_75t_L g10715 ( 
.A1(n_9875),
.A2(n_301),
.B(n_302),
.Y(n_10715)
);

AND2x2_ASAP7_75t_L g10716 ( 
.A(n_10310),
.B(n_691),
.Y(n_10716)
);

AOI21xp5_ASAP7_75t_L g10717 ( 
.A1(n_9966),
.A2(n_301),
.B(n_302),
.Y(n_10717)
);

INVx1_ASAP7_75t_L g10718 ( 
.A(n_10125),
.Y(n_10718)
);

CKINVDCx5p33_ASAP7_75t_R g10719 ( 
.A(n_10160),
.Y(n_10719)
);

NOR2xp33_ASAP7_75t_SL g10720 ( 
.A(n_9894),
.B(n_302),
.Y(n_10720)
);

NAND2xp5_ASAP7_75t_SL g10721 ( 
.A(n_9953),
.B(n_692),
.Y(n_10721)
);

INVx2_ASAP7_75t_L g10722 ( 
.A(n_10130),
.Y(n_10722)
);

O2A1O1Ixp5_ASAP7_75t_L g10723 ( 
.A1(n_10515),
.A2(n_694),
.B(n_692),
.C(n_693),
.Y(n_10723)
);

AOI21xp5_ASAP7_75t_L g10724 ( 
.A1(n_9917),
.A2(n_693),
.B(n_694),
.Y(n_10724)
);

INVxp67_ASAP7_75t_L g10725 ( 
.A(n_10207),
.Y(n_10725)
);

NOR2xp33_ASAP7_75t_L g10726 ( 
.A(n_9920),
.B(n_695),
.Y(n_10726)
);

OAI21xp5_ASAP7_75t_L g10727 ( 
.A1(n_9968),
.A2(n_695),
.B(n_696),
.Y(n_10727)
);

NOR2xp33_ASAP7_75t_L g10728 ( 
.A(n_9931),
.B(n_697),
.Y(n_10728)
);

INVx2_ASAP7_75t_L g10729 ( 
.A(n_10144),
.Y(n_10729)
);

AND2x2_ASAP7_75t_SL g10730 ( 
.A(n_9981),
.B(n_697),
.Y(n_10730)
);

INVx2_ASAP7_75t_L g10731 ( 
.A(n_10350),
.Y(n_10731)
);

AOI21xp5_ASAP7_75t_L g10732 ( 
.A1(n_9932),
.A2(n_698),
.B(n_699),
.Y(n_10732)
);

INVx2_ASAP7_75t_L g10733 ( 
.A(n_10380),
.Y(n_10733)
);

INVxp67_ASAP7_75t_L g10734 ( 
.A(n_10207),
.Y(n_10734)
);

AOI21x1_ASAP7_75t_L g10735 ( 
.A1(n_9871),
.A2(n_698),
.B(n_699),
.Y(n_10735)
);

NAND2xp5_ASAP7_75t_L g10736 ( 
.A(n_10011),
.B(n_700),
.Y(n_10736)
);

INVxp67_ASAP7_75t_SL g10737 ( 
.A(n_10143),
.Y(n_10737)
);

NAND2x1p5_ASAP7_75t_L g10738 ( 
.A(n_10344),
.B(n_701),
.Y(n_10738)
);

AND2x2_ASAP7_75t_L g10739 ( 
.A(n_9825),
.B(n_701),
.Y(n_10739)
);

NOR2x1p5_ASAP7_75t_SL g10740 ( 
.A(n_10086),
.B(n_702),
.Y(n_10740)
);

AO21x1_ASAP7_75t_L g10741 ( 
.A1(n_10348),
.A2(n_703),
.B(n_704),
.Y(n_10741)
);

NAND2xp5_ASAP7_75t_L g10742 ( 
.A(n_10012),
.B(n_703),
.Y(n_10742)
);

BUFx2_ASAP7_75t_SL g10743 ( 
.A(n_9995),
.Y(n_10743)
);

INVx2_ASAP7_75t_L g10744 ( 
.A(n_10385),
.Y(n_10744)
);

NOR2xp33_ASAP7_75t_L g10745 ( 
.A(n_10358),
.B(n_704),
.Y(n_10745)
);

CKINVDCx8_ASAP7_75t_R g10746 ( 
.A(n_9828),
.Y(n_10746)
);

INVx2_ASAP7_75t_L g10747 ( 
.A(n_10411),
.Y(n_10747)
);

INVx1_ASAP7_75t_L g10748 ( 
.A(n_10427),
.Y(n_10748)
);

INVx2_ASAP7_75t_L g10749 ( 
.A(n_10446),
.Y(n_10749)
);

NOR2xp33_ASAP7_75t_L g10750 ( 
.A(n_10051),
.B(n_705),
.Y(n_10750)
);

NAND2xp5_ASAP7_75t_SL g10751 ( 
.A(n_10266),
.B(n_705),
.Y(n_10751)
);

AOI221x1_ASAP7_75t_L g10752 ( 
.A1(n_9859),
.A2(n_10114),
.B1(n_10040),
.B2(n_10525),
.C(n_10523),
.Y(n_10752)
);

OAI22xp5_ASAP7_75t_L g10753 ( 
.A1(n_10512),
.A2(n_708),
.B1(n_706),
.B2(n_707),
.Y(n_10753)
);

AOI21xp5_ASAP7_75t_L g10754 ( 
.A1(n_10029),
.A2(n_706),
.B(n_707),
.Y(n_10754)
);

INVx2_ASAP7_75t_L g10755 ( 
.A(n_10478),
.Y(n_10755)
);

O2A1O1Ixp33_ASAP7_75t_L g10756 ( 
.A1(n_10495),
.A2(n_10520),
.B(n_10000),
.C(n_9841),
.Y(n_10756)
);

AOI21x1_ASAP7_75t_L g10757 ( 
.A1(n_9844),
.A2(n_708),
.B(n_709),
.Y(n_10757)
);

INVx2_ASAP7_75t_L g10758 ( 
.A(n_10492),
.Y(n_10758)
);

NOR2xp33_ASAP7_75t_L g10759 ( 
.A(n_10462),
.B(n_709),
.Y(n_10759)
);

AND2x6_ASAP7_75t_SL g10760 ( 
.A(n_10104),
.B(n_710),
.Y(n_10760)
);

INVx2_ASAP7_75t_L g10761 ( 
.A(n_10510),
.Y(n_10761)
);

AND2x2_ASAP7_75t_L g10762 ( 
.A(n_10384),
.B(n_710),
.Y(n_10762)
);

AOI21xp5_ASAP7_75t_L g10763 ( 
.A1(n_10536),
.A2(n_711),
.B(n_712),
.Y(n_10763)
);

INVx1_ASAP7_75t_L g10764 ( 
.A(n_10531),
.Y(n_10764)
);

INVx1_ASAP7_75t_L g10765 ( 
.A(n_10535),
.Y(n_10765)
);

INVx2_ASAP7_75t_L g10766 ( 
.A(n_10020),
.Y(n_10766)
);

INVx2_ASAP7_75t_L g10767 ( 
.A(n_10042),
.Y(n_10767)
);

AND2x2_ASAP7_75t_L g10768 ( 
.A(n_10430),
.B(n_10431),
.Y(n_10768)
);

AOI21xp5_ASAP7_75t_L g10769 ( 
.A1(n_10063),
.A2(n_712),
.B(n_713),
.Y(n_10769)
);

AOI222xp33_ASAP7_75t_L g10770 ( 
.A1(n_10352),
.A2(n_715),
.B1(n_717),
.B2(n_713),
.C1(n_714),
.C2(n_716),
.Y(n_10770)
);

AOI22xp33_ASAP7_75t_L g10771 ( 
.A1(n_9812),
.A2(n_716),
.B1(n_714),
.B2(n_715),
.Y(n_10771)
);

NOR2xp33_ASAP7_75t_L g10772 ( 
.A(n_10501),
.B(n_717),
.Y(n_10772)
);

AOI21xp5_ASAP7_75t_L g10773 ( 
.A1(n_9811),
.A2(n_10349),
.B(n_10346),
.Y(n_10773)
);

OAI22xp5_ASAP7_75t_L g10774 ( 
.A1(n_10538),
.A2(n_10382),
.B1(n_10387),
.B2(n_10375),
.Y(n_10774)
);

A2O1A1Ixp33_ASAP7_75t_L g10775 ( 
.A1(n_10377),
.A2(n_720),
.B(n_718),
.C(n_719),
.Y(n_10775)
);

BUFx6f_ASAP7_75t_L g10776 ( 
.A(n_9828),
.Y(n_10776)
);

OAI22xp5_ASAP7_75t_L g10777 ( 
.A1(n_10394),
.A2(n_721),
.B1(n_718),
.B2(n_719),
.Y(n_10777)
);

A2O1A1Ixp33_ASAP7_75t_L g10778 ( 
.A1(n_10399),
.A2(n_724),
.B(n_722),
.C(n_723),
.Y(n_10778)
);

NOR2xp33_ASAP7_75t_L g10779 ( 
.A(n_9961),
.B(n_722),
.Y(n_10779)
);

NAND2xp5_ASAP7_75t_L g10780 ( 
.A(n_10351),
.B(n_723),
.Y(n_10780)
);

NAND2xp5_ASAP7_75t_L g10781 ( 
.A(n_10373),
.B(n_726),
.Y(n_10781)
);

OAI22xp5_ASAP7_75t_SL g10782 ( 
.A1(n_10402),
.A2(n_728),
.B1(n_726),
.B2(n_727),
.Y(n_10782)
);

A2O1A1Ixp33_ASAP7_75t_L g10783 ( 
.A1(n_9985),
.A2(n_730),
.B(n_728),
.C(n_729),
.Y(n_10783)
);

OAI22xp5_ASAP7_75t_L g10784 ( 
.A1(n_10441),
.A2(n_10486),
.B1(n_10469),
.B2(n_9854),
.Y(n_10784)
);

OAI22xp5_ASAP7_75t_L g10785 ( 
.A1(n_10206),
.A2(n_731),
.B1(n_729),
.B2(n_730),
.Y(n_10785)
);

INVx2_ASAP7_75t_L g10786 ( 
.A(n_10403),
.Y(n_10786)
);

AOI21xp5_ASAP7_75t_L g10787 ( 
.A1(n_10354),
.A2(n_731),
.B(n_732),
.Y(n_10787)
);

INVx1_ASAP7_75t_SL g10788 ( 
.A(n_10207),
.Y(n_10788)
);

INVx2_ASAP7_75t_L g10789 ( 
.A(n_10505),
.Y(n_10789)
);

NOR2xp33_ASAP7_75t_R g10790 ( 
.A(n_10054),
.B(n_732),
.Y(n_10790)
);

OAI21x1_ASAP7_75t_L g10791 ( 
.A1(n_10169),
.A2(n_733),
.B(n_734),
.Y(n_10791)
);

INVx4_ASAP7_75t_L g10792 ( 
.A(n_10496),
.Y(n_10792)
);

INVx3_ASAP7_75t_L g10793 ( 
.A(n_9869),
.Y(n_10793)
);

NOR2xp33_ASAP7_75t_L g10794 ( 
.A(n_10369),
.B(n_733),
.Y(n_10794)
);

AOI21xp5_ASAP7_75t_L g10795 ( 
.A1(n_10355),
.A2(n_735),
.B(n_736),
.Y(n_10795)
);

AOI22xp5_ASAP7_75t_L g10796 ( 
.A1(n_10417),
.A2(n_737),
.B1(n_735),
.B2(n_736),
.Y(n_10796)
);

INVx2_ASAP7_75t_SL g10797 ( 
.A(n_10276),
.Y(n_10797)
);

OAI21xp5_ASAP7_75t_L g10798 ( 
.A1(n_9975),
.A2(n_737),
.B(n_738),
.Y(n_10798)
);

BUFx6f_ASAP7_75t_L g10799 ( 
.A(n_10496),
.Y(n_10799)
);

O2A1O1Ixp33_ASAP7_75t_L g10800 ( 
.A1(n_10371),
.A2(n_740),
.B(n_738),
.C(n_739),
.Y(n_10800)
);

INVx4_ASAP7_75t_L g10801 ( 
.A(n_10498),
.Y(n_10801)
);

A2O1A1Ixp33_ASAP7_75t_L g10802 ( 
.A1(n_9833),
.A2(n_741),
.B(n_739),
.C(n_740),
.Y(n_10802)
);

AOI21xp5_ASAP7_75t_L g10803 ( 
.A1(n_10365),
.A2(n_741),
.B(n_742),
.Y(n_10803)
);

O2A1O1Ixp33_ASAP7_75t_L g10804 ( 
.A1(n_10392),
.A2(n_744),
.B(n_742),
.C(n_743),
.Y(n_10804)
);

INVx2_ASAP7_75t_SL g10805 ( 
.A(n_10276),
.Y(n_10805)
);

AOI21xp33_ASAP7_75t_L g10806 ( 
.A1(n_10007),
.A2(n_10052),
.B(n_9992),
.Y(n_10806)
);

A2O1A1Ixp33_ASAP7_75t_L g10807 ( 
.A1(n_9884),
.A2(n_746),
.B(n_744),
.C(n_745),
.Y(n_10807)
);

INVx2_ASAP7_75t_L g10808 ( 
.A(n_10158),
.Y(n_10808)
);

NAND2xp5_ASAP7_75t_L g10809 ( 
.A(n_10214),
.B(n_745),
.Y(n_10809)
);

NAND2xp5_ASAP7_75t_L g10810 ( 
.A(n_10273),
.B(n_746),
.Y(n_10810)
);

OAI21x1_ASAP7_75t_L g10811 ( 
.A1(n_9914),
.A2(n_747),
.B(n_748),
.Y(n_10811)
);

AOI21xp5_ASAP7_75t_L g10812 ( 
.A1(n_10386),
.A2(n_747),
.B(n_748),
.Y(n_10812)
);

NAND2xp5_ASAP7_75t_L g10813 ( 
.A(n_10163),
.B(n_751),
.Y(n_10813)
);

CKINVDCx5p33_ASAP7_75t_R g10814 ( 
.A(n_9954),
.Y(n_10814)
);

NAND2xp5_ASAP7_75t_L g10815 ( 
.A(n_10272),
.B(n_10461),
.Y(n_10815)
);

NAND2xp5_ASAP7_75t_L g10816 ( 
.A(n_10464),
.B(n_751),
.Y(n_10816)
);

BUFx6f_ASAP7_75t_L g10817 ( 
.A(n_10498),
.Y(n_10817)
);

INVx3_ASAP7_75t_SL g10818 ( 
.A(n_10519),
.Y(n_10818)
);

INVx1_ASAP7_75t_SL g10819 ( 
.A(n_10276),
.Y(n_10819)
);

OR2x6_ASAP7_75t_L g10820 ( 
.A(n_9900),
.B(n_752),
.Y(n_10820)
);

INVx2_ASAP7_75t_L g10821 ( 
.A(n_10103),
.Y(n_10821)
);

AOI22xp5_ASAP7_75t_L g10822 ( 
.A1(n_10428),
.A2(n_754),
.B1(n_752),
.B2(n_753),
.Y(n_10822)
);

NAND2xp5_ASAP7_75t_L g10823 ( 
.A(n_10477),
.B(n_753),
.Y(n_10823)
);

O2A1O1Ixp33_ASAP7_75t_L g10824 ( 
.A1(n_10413),
.A2(n_756),
.B(n_754),
.C(n_755),
.Y(n_10824)
);

NOR3xp33_ASAP7_75t_SL g10825 ( 
.A(n_10284),
.B(n_755),
.C(n_756),
.Y(n_10825)
);

O2A1O1Ixp33_ASAP7_75t_L g10826 ( 
.A1(n_10442),
.A2(n_759),
.B(n_757),
.C(n_758),
.Y(n_10826)
);

INVx4_ASAP7_75t_L g10827 ( 
.A(n_10519),
.Y(n_10827)
);

HB1xp67_ASAP7_75t_L g10828 ( 
.A(n_10215),
.Y(n_10828)
);

O2A1O1Ixp33_ASAP7_75t_L g10829 ( 
.A1(n_10454),
.A2(n_760),
.B(n_758),
.C(n_759),
.Y(n_10829)
);

AO32x2_ASAP7_75t_L g10830 ( 
.A1(n_9969),
.A2(n_762),
.A3(n_760),
.B1(n_761),
.B2(n_763),
.Y(n_10830)
);

NAND2xp5_ASAP7_75t_L g10831 ( 
.A(n_10516),
.B(n_761),
.Y(n_10831)
);

BUFx12f_ASAP7_75t_L g10832 ( 
.A(n_10108),
.Y(n_10832)
);

NAND2xp5_ASAP7_75t_L g10833 ( 
.A(n_9817),
.B(n_762),
.Y(n_10833)
);

AND2x4_ASAP7_75t_L g10834 ( 
.A(n_10070),
.B(n_763),
.Y(n_10834)
);

INVxp67_ASAP7_75t_SL g10835 ( 
.A(n_10439),
.Y(n_10835)
);

AOI22xp5_ASAP7_75t_L g10836 ( 
.A1(n_10465),
.A2(n_767),
.B1(n_764),
.B2(n_765),
.Y(n_10836)
);

INVx4_ASAP7_75t_L g10837 ( 
.A(n_10151),
.Y(n_10837)
);

BUFx6f_ASAP7_75t_L g10838 ( 
.A(n_9821),
.Y(n_10838)
);

NAND2xp5_ASAP7_75t_L g10839 ( 
.A(n_10343),
.B(n_764),
.Y(n_10839)
);

NAND2xp5_ASAP7_75t_SL g10840 ( 
.A(n_9962),
.B(n_767),
.Y(n_10840)
);

INVx2_ASAP7_75t_L g10841 ( 
.A(n_10112),
.Y(n_10841)
);

NAND2xp5_ASAP7_75t_L g10842 ( 
.A(n_10353),
.B(n_768),
.Y(n_10842)
);

AOI21xp5_ASAP7_75t_L g10843 ( 
.A1(n_10390),
.A2(n_769),
.B(n_770),
.Y(n_10843)
);

OAI22xp5_ASAP7_75t_L g10844 ( 
.A1(n_9941),
.A2(n_771),
.B1(n_769),
.B2(n_770),
.Y(n_10844)
);

O2A1O1Ixp5_ASAP7_75t_L g10845 ( 
.A1(n_10031),
.A2(n_773),
.B(n_771),
.C(n_772),
.Y(n_10845)
);

AOI21xp5_ASAP7_75t_L g10846 ( 
.A1(n_10393),
.A2(n_772),
.B(n_773),
.Y(n_10846)
);

O2A1O1Ixp5_ASAP7_75t_L g10847 ( 
.A1(n_10537),
.A2(n_9924),
.B(n_10015),
.C(n_10058),
.Y(n_10847)
);

INVx3_ASAP7_75t_L g10848 ( 
.A(n_9988),
.Y(n_10848)
);

NAND2xp5_ASAP7_75t_L g10849 ( 
.A(n_10359),
.B(n_774),
.Y(n_10849)
);

A2O1A1Ixp33_ASAP7_75t_L g10850 ( 
.A1(n_9928),
.A2(n_776),
.B(n_774),
.C(n_775),
.Y(n_10850)
);

INVx2_ASAP7_75t_L g10851 ( 
.A(n_10122),
.Y(n_10851)
);

O2A1O1Ixp33_ASAP7_75t_L g10852 ( 
.A1(n_10211),
.A2(n_777),
.B(n_775),
.C(n_776),
.Y(n_10852)
);

NAND2xp5_ASAP7_75t_SL g10853 ( 
.A(n_10189),
.B(n_777),
.Y(n_10853)
);

INVx1_ASAP7_75t_L g10854 ( 
.A(n_10128),
.Y(n_10854)
);

NOR2xp33_ASAP7_75t_L g10855 ( 
.A(n_9826),
.B(n_778),
.Y(n_10855)
);

AOI21xp33_ASAP7_75t_L g10856 ( 
.A1(n_10166),
.A2(n_778),
.B(n_779),
.Y(n_10856)
);

INVx1_ASAP7_75t_SL g10857 ( 
.A(n_10289),
.Y(n_10857)
);

AOI21xp5_ASAP7_75t_L g10858 ( 
.A1(n_10400),
.A2(n_779),
.B(n_780),
.Y(n_10858)
);

INVx2_ASAP7_75t_L g10859 ( 
.A(n_10133),
.Y(n_10859)
);

NOR2xp33_ASAP7_75t_L g10860 ( 
.A(n_10378),
.B(n_780),
.Y(n_10860)
);

NAND2xp33_ASAP7_75t_L g10861 ( 
.A(n_9887),
.B(n_781),
.Y(n_10861)
);

NAND2xp5_ASAP7_75t_SL g10862 ( 
.A(n_9922),
.B(n_10190),
.Y(n_10862)
);

INVx2_ASAP7_75t_L g10863 ( 
.A(n_10139),
.Y(n_10863)
);

NOR2xp33_ASAP7_75t_L g10864 ( 
.A(n_10397),
.B(n_781),
.Y(n_10864)
);

NOR3xp33_ASAP7_75t_L g10865 ( 
.A(n_10067),
.B(n_782),
.C(n_783),
.Y(n_10865)
);

NOR2xp33_ASAP7_75t_SL g10866 ( 
.A(n_10179),
.B(n_782),
.Y(n_10866)
);

BUFx6f_ASAP7_75t_L g10867 ( 
.A(n_10376),
.Y(n_10867)
);

INVx5_ASAP7_75t_L g10868 ( 
.A(n_10013),
.Y(n_10868)
);

NAND2xp5_ASAP7_75t_SL g10869 ( 
.A(n_10182),
.B(n_783),
.Y(n_10869)
);

OAI22xp5_ASAP7_75t_L g10870 ( 
.A1(n_10231),
.A2(n_786),
.B1(n_784),
.B2(n_785),
.Y(n_10870)
);

AOI21x1_ASAP7_75t_L g10871 ( 
.A1(n_10019),
.A2(n_784),
.B(n_785),
.Y(n_10871)
);

AOI21xp5_ASAP7_75t_L g10872 ( 
.A1(n_10401),
.A2(n_786),
.B(n_787),
.Y(n_10872)
);

INVx2_ASAP7_75t_L g10873 ( 
.A(n_10142),
.Y(n_10873)
);

NOR2xp33_ASAP7_75t_R g10874 ( 
.A(n_10383),
.B(n_787),
.Y(n_10874)
);

AOI22xp5_ASAP7_75t_L g10875 ( 
.A1(n_9862),
.A2(n_791),
.B1(n_789),
.B2(n_790),
.Y(n_10875)
);

NAND2xp5_ASAP7_75t_SL g10876 ( 
.A(n_10202),
.B(n_789),
.Y(n_10876)
);

NAND2xp5_ASAP7_75t_L g10877 ( 
.A(n_10360),
.B(n_790),
.Y(n_10877)
);

AOI21xp5_ASAP7_75t_L g10878 ( 
.A1(n_10408),
.A2(n_792),
.B(n_793),
.Y(n_10878)
);

A2O1A1Ixp33_ASAP7_75t_L g10879 ( 
.A1(n_10081),
.A2(n_794),
.B(n_792),
.C(n_793),
.Y(n_10879)
);

O2A1O1Ixp33_ASAP7_75t_L g10880 ( 
.A1(n_10066),
.A2(n_797),
.B(n_795),
.C(n_796),
.Y(n_10880)
);

AND2x6_ASAP7_75t_L g10881 ( 
.A(n_10293),
.B(n_795),
.Y(n_10881)
);

AOI21xp5_ASAP7_75t_L g10882 ( 
.A1(n_10409),
.A2(n_796),
.B(n_797),
.Y(n_10882)
);

NAND2xp5_ASAP7_75t_L g10883 ( 
.A(n_10361),
.B(n_798),
.Y(n_10883)
);

AOI21xp5_ASAP7_75t_L g10884 ( 
.A1(n_10414),
.A2(n_798),
.B(n_799),
.Y(n_10884)
);

HB1xp67_ASAP7_75t_L g10885 ( 
.A(n_10364),
.Y(n_10885)
);

INVx4_ASAP7_75t_L g10886 ( 
.A(n_10420),
.Y(n_10886)
);

NOR2xp33_ASAP7_75t_SL g10887 ( 
.A(n_10347),
.B(n_800),
.Y(n_10887)
);

NAND2xp5_ASAP7_75t_L g10888 ( 
.A(n_10367),
.B(n_800),
.Y(n_10888)
);

AOI21xp5_ASAP7_75t_L g10889 ( 
.A1(n_10424),
.A2(n_801),
.B(n_802),
.Y(n_10889)
);

NAND2xp5_ASAP7_75t_L g10890 ( 
.A(n_10368),
.B(n_801),
.Y(n_10890)
);

AOI22xp5_ASAP7_75t_L g10891 ( 
.A1(n_10222),
.A2(n_10294),
.B1(n_10174),
.B2(n_10388),
.Y(n_10891)
);

INVx1_ASAP7_75t_L g10892 ( 
.A(n_10372),
.Y(n_10892)
);

BUFx2_ASAP7_75t_L g10893 ( 
.A(n_10013),
.Y(n_10893)
);

AOI21xp5_ASAP7_75t_L g10894 ( 
.A1(n_10425),
.A2(n_802),
.B(n_803),
.Y(n_10894)
);

AO22x1_ASAP7_75t_L g10895 ( 
.A1(n_10079),
.A2(n_806),
.B1(n_804),
.B2(n_805),
.Y(n_10895)
);

AOI21xp5_ASAP7_75t_L g10896 ( 
.A1(n_10429),
.A2(n_804),
.B(n_806),
.Y(n_10896)
);

NAND2xp5_ASAP7_75t_L g10897 ( 
.A(n_10374),
.B(n_807),
.Y(n_10897)
);

BUFx2_ASAP7_75t_L g10898 ( 
.A(n_10013),
.Y(n_10898)
);

AOI21xp5_ASAP7_75t_L g10899 ( 
.A1(n_10437),
.A2(n_807),
.B(n_808),
.Y(n_10899)
);

AND2x4_ASAP7_75t_L g10900 ( 
.A(n_10188),
.B(n_808),
.Y(n_10900)
);

BUFx6f_ASAP7_75t_L g10901 ( 
.A(n_9832),
.Y(n_10901)
);

HB1xp67_ASAP7_75t_L g10902 ( 
.A(n_10379),
.Y(n_10902)
);

NAND2xp5_ASAP7_75t_L g10903 ( 
.A(n_10381),
.B(n_809),
.Y(n_10903)
);

AOI21xp5_ASAP7_75t_L g10904 ( 
.A1(n_10438),
.A2(n_809),
.B(n_810),
.Y(n_10904)
);

NOR2xp33_ASAP7_75t_L g10905 ( 
.A(n_10443),
.B(n_10463),
.Y(n_10905)
);

HB1xp67_ASAP7_75t_L g10906 ( 
.A(n_10398),
.Y(n_10906)
);

O2A1O1Ixp33_ASAP7_75t_L g10907 ( 
.A1(n_10077),
.A2(n_812),
.B(n_810),
.C(n_811),
.Y(n_10907)
);

CKINVDCx10_ASAP7_75t_R g10908 ( 
.A(n_10233),
.Y(n_10908)
);

CKINVDCx20_ASAP7_75t_R g10909 ( 
.A(n_10467),
.Y(n_10909)
);

OAI22xp5_ASAP7_75t_L g10910 ( 
.A1(n_10083),
.A2(n_814),
.B1(n_811),
.B2(n_813),
.Y(n_10910)
);

O2A1O1Ixp33_ASAP7_75t_L g10911 ( 
.A1(n_10089),
.A2(n_815),
.B(n_813),
.C(n_814),
.Y(n_10911)
);

NAND2xp5_ASAP7_75t_L g10912 ( 
.A(n_10406),
.B(n_815),
.Y(n_10912)
);

INVx2_ASAP7_75t_L g10913 ( 
.A(n_10041),
.Y(n_10913)
);

INVx2_ASAP7_75t_L g10914 ( 
.A(n_10178),
.Y(n_10914)
);

O2A1O1Ixp5_ASAP7_75t_L g10915 ( 
.A1(n_10107),
.A2(n_819),
.B(n_816),
.C(n_817),
.Y(n_10915)
);

BUFx3_ASAP7_75t_L g10916 ( 
.A(n_9832),
.Y(n_10916)
);

NAND2xp5_ASAP7_75t_SL g10917 ( 
.A(n_10332),
.B(n_10412),
.Y(n_10917)
);

O2A1O1Ixp33_ASAP7_75t_SL g10918 ( 
.A1(n_10338),
.A2(n_819),
.B(n_816),
.C(n_817),
.Y(n_10918)
);

NOR2xp67_ASAP7_75t_SL g10919 ( 
.A(n_10147),
.B(n_820),
.Y(n_10919)
);

AOI21xp5_ASAP7_75t_L g10920 ( 
.A1(n_10445),
.A2(n_821),
.B(n_822),
.Y(n_10920)
);

OAI21xp5_ASAP7_75t_L g10921 ( 
.A1(n_9967),
.A2(n_822),
.B(n_823),
.Y(n_10921)
);

AND2x2_ASAP7_75t_L g10922 ( 
.A(n_10312),
.B(n_823),
.Y(n_10922)
);

A2O1A1Ixp33_ASAP7_75t_L g10923 ( 
.A1(n_10094),
.A2(n_826),
.B(n_824),
.C(n_825),
.Y(n_10923)
);

INVx2_ASAP7_75t_L g10924 ( 
.A(n_10183),
.Y(n_10924)
);

NAND2xp5_ASAP7_75t_SL g10925 ( 
.A(n_10422),
.B(n_824),
.Y(n_10925)
);

NAND2xp5_ASAP7_75t_L g10926 ( 
.A(n_10423),
.B(n_825),
.Y(n_10926)
);

NAND2xp5_ASAP7_75t_SL g10927 ( 
.A(n_10426),
.B(n_826),
.Y(n_10927)
);

NAND2xp5_ASAP7_75t_L g10928 ( 
.A(n_10444),
.B(n_827),
.Y(n_10928)
);

AO21x1_ASAP7_75t_L g10929 ( 
.A1(n_9853),
.A2(n_827),
.B(n_828),
.Y(n_10929)
);

OAI21xp33_ASAP7_75t_SL g10930 ( 
.A1(n_9911),
.A2(n_828),
.B(n_830),
.Y(n_10930)
);

NOR3xp33_ASAP7_75t_SL g10931 ( 
.A(n_10124),
.B(n_10313),
.C(n_10127),
.Y(n_10931)
);

XOR2x2_ASAP7_75t_L g10932 ( 
.A(n_9842),
.B(n_830),
.Y(n_10932)
);

INVx1_ASAP7_75t_L g10933 ( 
.A(n_10448),
.Y(n_10933)
);

NOR2xp33_ASAP7_75t_L g10934 ( 
.A(n_10471),
.B(n_831),
.Y(n_10934)
);

O2A1O1Ixp33_ASAP7_75t_L g10935 ( 
.A1(n_10091),
.A2(n_833),
.B(n_831),
.C(n_832),
.Y(n_10935)
);

OAI21x1_ASAP7_75t_L g10936 ( 
.A1(n_9907),
.A2(n_832),
.B(n_833),
.Y(n_10936)
);

HB1xp67_ASAP7_75t_L g10937 ( 
.A(n_10452),
.Y(n_10937)
);

INVx1_ASAP7_75t_L g10938 ( 
.A(n_10457),
.Y(n_10938)
);

BUFx4f_ASAP7_75t_L g10939 ( 
.A(n_10289),
.Y(n_10939)
);

A2O1A1Ixp33_ASAP7_75t_L g10940 ( 
.A1(n_10117),
.A2(n_837),
.B(n_835),
.C(n_836),
.Y(n_10940)
);

AOI21x1_ASAP7_75t_L g10941 ( 
.A1(n_10090),
.A2(n_835),
.B(n_836),
.Y(n_10941)
);

O2A1O1Ixp5_ASAP7_75t_L g10942 ( 
.A1(n_10134),
.A2(n_839),
.B(n_837),
.C(n_838),
.Y(n_10942)
);

NAND2xp5_ASAP7_75t_L g10943 ( 
.A(n_10470),
.B(n_10491),
.Y(n_10943)
);

NAND2xp5_ASAP7_75t_L g10944 ( 
.A(n_10502),
.B(n_839),
.Y(n_10944)
);

AND2x4_ASAP7_75t_L g10945 ( 
.A(n_10328),
.B(n_840),
.Y(n_10945)
);

NAND2xp5_ASAP7_75t_L g10946 ( 
.A(n_10504),
.B(n_840),
.Y(n_10946)
);

AOI21xp5_ASAP7_75t_L g10947 ( 
.A1(n_10450),
.A2(n_841),
.B(n_842),
.Y(n_10947)
);

BUFx8_ASAP7_75t_SL g10948 ( 
.A(n_9846),
.Y(n_10948)
);

BUFx2_ASAP7_75t_L g10949 ( 
.A(n_9989),
.Y(n_10949)
);

A2O1A1Ixp33_ASAP7_75t_L g10950 ( 
.A1(n_10146),
.A2(n_843),
.B(n_841),
.C(n_842),
.Y(n_10950)
);

INVx1_ASAP7_75t_L g10951 ( 
.A(n_10506),
.Y(n_10951)
);

NAND2xp5_ASAP7_75t_L g10952 ( 
.A(n_10511),
.B(n_844),
.Y(n_10952)
);

AOI21xp5_ASAP7_75t_L g10953 ( 
.A1(n_10460),
.A2(n_844),
.B(n_845),
.Y(n_10953)
);

NAND2xp5_ASAP7_75t_SL g10954 ( 
.A(n_10521),
.B(n_845),
.Y(n_10954)
);

NOR2xp33_ASAP7_75t_L g10955 ( 
.A(n_10473),
.B(n_846),
.Y(n_10955)
);

INVx2_ASAP7_75t_L g10956 ( 
.A(n_10185),
.Y(n_10956)
);

NAND3xp33_ASAP7_75t_SL g10957 ( 
.A(n_10245),
.B(n_847),
.C(n_848),
.Y(n_10957)
);

BUFx6f_ASAP7_75t_L g10958 ( 
.A(n_9890),
.Y(n_10958)
);

AOI21xp5_ASAP7_75t_L g10959 ( 
.A1(n_10468),
.A2(n_847),
.B(n_848),
.Y(n_10959)
);

NOR2xp33_ASAP7_75t_L g10960 ( 
.A(n_10474),
.B(n_849),
.Y(n_10960)
);

NOR2x1_ASAP7_75t_L g10961 ( 
.A(n_9818),
.B(n_850),
.Y(n_10961)
);

NAND2xp5_ASAP7_75t_L g10962 ( 
.A(n_10221),
.B(n_850),
.Y(n_10962)
);

AND2x2_ASAP7_75t_L g10963 ( 
.A(n_9947),
.B(n_851),
.Y(n_10963)
);

NAND2xp5_ASAP7_75t_L g10964 ( 
.A(n_10239),
.B(n_852),
.Y(n_10964)
);

INVx1_ASAP7_75t_L g10965 ( 
.A(n_10404),
.Y(n_10965)
);

NOR2xp33_ASAP7_75t_L g10966 ( 
.A(n_10494),
.B(n_852),
.Y(n_10966)
);

OAI22xp5_ASAP7_75t_L g10967 ( 
.A1(n_10241),
.A2(n_855),
.B1(n_853),
.B2(n_854),
.Y(n_10967)
);

AOI22x1_ASAP7_75t_L g10968 ( 
.A1(n_9861),
.A2(n_857),
.B1(n_853),
.B2(n_856),
.Y(n_10968)
);

NOR3xp33_ASAP7_75t_SL g10969 ( 
.A(n_10140),
.B(n_857),
.C(n_858),
.Y(n_10969)
);

O2A1O1Ixp33_ASAP7_75t_L g10970 ( 
.A1(n_10131),
.A2(n_10137),
.B(n_10150),
.C(n_10181),
.Y(n_10970)
);

OAI22xp5_ASAP7_75t_L g10971 ( 
.A1(n_10269),
.A2(n_860),
.B1(n_858),
.B2(n_859),
.Y(n_10971)
);

INVxp67_ASAP7_75t_SL g10972 ( 
.A(n_10324),
.Y(n_10972)
);

NOR2xp33_ASAP7_75t_L g10973 ( 
.A(n_10500),
.B(n_859),
.Y(n_10973)
);

INVx1_ASAP7_75t_L g10974 ( 
.A(n_10404),
.Y(n_10974)
);

INVx2_ASAP7_75t_L g10975 ( 
.A(n_9831),
.Y(n_10975)
);

AND2x2_ASAP7_75t_L g10976 ( 
.A(n_10026),
.B(n_860),
.Y(n_10976)
);

OAI21xp5_ASAP7_75t_L g10977 ( 
.A1(n_10227),
.A2(n_861),
.B(n_862),
.Y(n_10977)
);

NAND2xp5_ASAP7_75t_L g10978 ( 
.A(n_10213),
.B(n_9838),
.Y(n_10978)
);

AOI21xp5_ASAP7_75t_L g10979 ( 
.A1(n_10472),
.A2(n_10493),
.B(n_10480),
.Y(n_10979)
);

NOR2x1_ASAP7_75t_SL g10980 ( 
.A(n_9943),
.B(n_861),
.Y(n_10980)
);

INVx4_ASAP7_75t_L g10981 ( 
.A(n_10389),
.Y(n_10981)
);

BUFx3_ASAP7_75t_L g10982 ( 
.A(n_10389),
.Y(n_10982)
);

AOI22xp5_ASAP7_75t_L g10983 ( 
.A1(n_10526),
.A2(n_864),
.B1(n_862),
.B2(n_863),
.Y(n_10983)
);

AND2x4_ASAP7_75t_L g10984 ( 
.A(n_10509),
.B(n_863),
.Y(n_10984)
);

NOR3xp33_ASAP7_75t_SL g10985 ( 
.A(n_10528),
.B(n_864),
.C(n_865),
.Y(n_10985)
);

NOR2xp33_ASAP7_75t_L g10986 ( 
.A(n_10507),
.B(n_10522),
.Y(n_10986)
);

AOI22xp5_ASAP7_75t_L g10987 ( 
.A1(n_10161),
.A2(n_867),
.B1(n_865),
.B2(n_866),
.Y(n_10987)
);

NOR2xp33_ASAP7_75t_L g10988 ( 
.A(n_10217),
.B(n_867),
.Y(n_10988)
);

NAND2xp5_ASAP7_75t_L g10989 ( 
.A(n_9849),
.B(n_869),
.Y(n_10989)
);

INVx1_ASAP7_75t_L g10990 ( 
.A(n_10404),
.Y(n_10990)
);

NAND2xp5_ASAP7_75t_L g10991 ( 
.A(n_9850),
.B(n_869),
.Y(n_10991)
);

NAND2xp5_ASAP7_75t_L g10992 ( 
.A(n_9874),
.B(n_870),
.Y(n_10992)
);

A2O1A1Ixp33_ASAP7_75t_L g10993 ( 
.A1(n_10287),
.A2(n_872),
.B(n_870),
.C(n_871),
.Y(n_10993)
);

OR2x6_ASAP7_75t_L g10994 ( 
.A(n_10513),
.B(n_871),
.Y(n_10994)
);

A2O1A1Ixp33_ASAP7_75t_L g10995 ( 
.A1(n_10299),
.A2(n_874),
.B(n_872),
.C(n_873),
.Y(n_10995)
);

A2O1A1Ixp33_ASAP7_75t_L g10996 ( 
.A1(n_10092),
.A2(n_876),
.B(n_874),
.C(n_875),
.Y(n_10996)
);

NAND2xp5_ASAP7_75t_L g10997 ( 
.A(n_9876),
.B(n_875),
.Y(n_10997)
);

O2A1O1Ixp33_ASAP7_75t_L g10998 ( 
.A1(n_10290),
.A2(n_878),
.B(n_876),
.C(n_877),
.Y(n_10998)
);

O2A1O1Ixp5_ASAP7_75t_SL g10999 ( 
.A1(n_9921),
.A2(n_880),
.B(n_878),
.C(n_879),
.Y(n_10999)
);

NAND3xp33_ASAP7_75t_SL g11000 ( 
.A(n_10250),
.B(n_879),
.C(n_880),
.Y(n_11000)
);

OAI22xp5_ASAP7_75t_L g11001 ( 
.A1(n_10226),
.A2(n_883),
.B1(n_881),
.B2(n_882),
.Y(n_11001)
);

AOI21xp5_ASAP7_75t_L g11002 ( 
.A1(n_10517),
.A2(n_881),
.B(n_882),
.Y(n_11002)
);

OAI22xp5_ASAP7_75t_L g11003 ( 
.A1(n_10246),
.A2(n_885),
.B1(n_883),
.B2(n_884),
.Y(n_11003)
);

AOI22xp5_ASAP7_75t_L g11004 ( 
.A1(n_10192),
.A2(n_886),
.B1(n_884),
.B2(n_885),
.Y(n_11004)
);

NAND2xp5_ASAP7_75t_L g11005 ( 
.A(n_9878),
.B(n_886),
.Y(n_11005)
);

A2O1A1Ixp33_ASAP7_75t_L g11006 ( 
.A1(n_10340),
.A2(n_889),
.B(n_887),
.C(n_888),
.Y(n_11006)
);

AOI21xp5_ASAP7_75t_L g11007 ( 
.A1(n_10518),
.A2(n_887),
.B(n_890),
.Y(n_11007)
);

NOR2xp33_ASAP7_75t_SL g11008 ( 
.A(n_9997),
.B(n_890),
.Y(n_11008)
);

O2A1O1Ixp33_ASAP7_75t_L g11009 ( 
.A1(n_10263),
.A2(n_893),
.B(n_891),
.C(n_892),
.Y(n_11009)
);

O2A1O1Ixp33_ASAP7_75t_L g11010 ( 
.A1(n_10255),
.A2(n_10032),
.B(n_10024),
.C(n_9971),
.Y(n_11010)
);

OAI22xp5_ASAP7_75t_SL g11011 ( 
.A1(n_10060),
.A2(n_894),
.B1(n_892),
.B2(n_893),
.Y(n_11011)
);

AOI21xp5_ASAP7_75t_L g11012 ( 
.A1(n_10524),
.A2(n_894),
.B(n_895),
.Y(n_11012)
);

NAND2xp5_ASAP7_75t_L g11013 ( 
.A(n_9879),
.B(n_895),
.Y(n_11013)
);

AND2x4_ASAP7_75t_L g11014 ( 
.A(n_10061),
.B(n_896),
.Y(n_11014)
);

AOI22xp5_ASAP7_75t_L g11015 ( 
.A1(n_9998),
.A2(n_898),
.B1(n_896),
.B2(n_897),
.Y(n_11015)
);

NAND2xp5_ASAP7_75t_L g11016 ( 
.A(n_10016),
.B(n_897),
.Y(n_11016)
);

NAND2xp5_ASAP7_75t_SL g11017 ( 
.A(n_10247),
.B(n_9925),
.Y(n_11017)
);

NAND2xp5_ASAP7_75t_SL g11018 ( 
.A(n_9930),
.B(n_898),
.Y(n_11018)
);

NAND2xp5_ASAP7_75t_L g11019 ( 
.A(n_10018),
.B(n_899),
.Y(n_11019)
);

O2A1O1Ixp33_ASAP7_75t_L g11020 ( 
.A1(n_9973),
.A2(n_902),
.B(n_899),
.C(n_901),
.Y(n_11020)
);

NAND2xp5_ASAP7_75t_L g11021 ( 
.A(n_10049),
.B(n_902),
.Y(n_11021)
);

AOI21xp5_ASAP7_75t_L g11022 ( 
.A1(n_10527),
.A2(n_10530),
.B(n_10529),
.Y(n_11022)
);

NOR3xp33_ASAP7_75t_SL g11023 ( 
.A(n_10257),
.B(n_903),
.C(n_904),
.Y(n_11023)
);

BUFx8_ASAP7_75t_SL g11024 ( 
.A(n_9970),
.Y(n_11024)
);

OAI22xp5_ASAP7_75t_L g11025 ( 
.A1(n_10129),
.A2(n_905),
.B1(n_903),
.B2(n_904),
.Y(n_11025)
);

O2A1O1Ixp33_ASAP7_75t_L g11026 ( 
.A1(n_9858),
.A2(n_908),
.B(n_906),
.C(n_907),
.Y(n_11026)
);

AOI22xp5_ASAP7_75t_L g11027 ( 
.A1(n_10232),
.A2(n_908),
.B1(n_906),
.B2(n_907),
.Y(n_11027)
);

INVx2_ASAP7_75t_L g11028 ( 
.A(n_9896),
.Y(n_11028)
);

NAND2xp5_ASAP7_75t_L g11029 ( 
.A(n_10056),
.B(n_909),
.Y(n_11029)
);

NOR3xp33_ASAP7_75t_SL g11030 ( 
.A(n_10235),
.B(n_909),
.C(n_910),
.Y(n_11030)
);

INVx2_ASAP7_75t_L g11031 ( 
.A(n_9898),
.Y(n_11031)
);

NAND2xp5_ASAP7_75t_L g11032 ( 
.A(n_9901),
.B(n_911),
.Y(n_11032)
);

AOI21xp5_ASAP7_75t_L g11033 ( 
.A1(n_10533),
.A2(n_911),
.B(n_912),
.Y(n_11033)
);

INVx1_ASAP7_75t_L g11034 ( 
.A(n_10260),
.Y(n_11034)
);

NOR2xp33_ASAP7_75t_L g11035 ( 
.A(n_10334),
.B(n_912),
.Y(n_11035)
);

INVx2_ASAP7_75t_L g11036 ( 
.A(n_9903),
.Y(n_11036)
);

AOI21xp5_ASAP7_75t_L g11037 ( 
.A1(n_10046),
.A2(n_913),
.B(n_914),
.Y(n_11037)
);

AOI22xp5_ASAP7_75t_L g11038 ( 
.A1(n_10033),
.A2(n_915),
.B1(n_913),
.B2(n_914),
.Y(n_11038)
);

INVx2_ASAP7_75t_L g11039 ( 
.A(n_10335),
.Y(n_11039)
);

BUFx3_ASAP7_75t_L g11040 ( 
.A(n_9988),
.Y(n_11040)
);

OAI22xp5_ASAP7_75t_L g11041 ( 
.A1(n_10171),
.A2(n_917),
.B1(n_915),
.B2(n_916),
.Y(n_11041)
);

O2A1O1Ixp33_ASAP7_75t_L g11042 ( 
.A1(n_10331),
.A2(n_920),
.B(n_918),
.C(n_919),
.Y(n_11042)
);

INVx2_ASAP7_75t_L g11043 ( 
.A(n_10240),
.Y(n_11043)
);

NOR3xp33_ASAP7_75t_L g11044 ( 
.A(n_9864),
.B(n_918),
.C(n_919),
.Y(n_11044)
);

INVx1_ASAP7_75t_L g11045 ( 
.A(n_10288),
.Y(n_11045)
);

INVx2_ASAP7_75t_L g11046 ( 
.A(n_10302),
.Y(n_11046)
);

NOR2xp33_ASAP7_75t_L g11047 ( 
.A(n_10319),
.B(n_10219),
.Y(n_11047)
);

INVx2_ASAP7_75t_SL g11048 ( 
.A(n_9996),
.Y(n_11048)
);

BUFx6f_ASAP7_75t_L g11049 ( 
.A(n_9996),
.Y(n_11049)
);

INVx6_ASAP7_75t_L g11050 ( 
.A(n_10048),
.Y(n_11050)
);

INVx4_ASAP7_75t_L g11051 ( 
.A(n_10048),
.Y(n_11051)
);

BUFx6f_ASAP7_75t_L g11052 ( 
.A(n_10061),
.Y(n_11052)
);

AOI222xp33_ASAP7_75t_L g11053 ( 
.A1(n_10318),
.A2(n_922),
.B1(n_924),
.B2(n_920),
.C1(n_921),
.C2(n_923),
.Y(n_11053)
);

INVx1_ASAP7_75t_L g11054 ( 
.A(n_9963),
.Y(n_11054)
);

CKINVDCx5p33_ASAP7_75t_R g11055 ( 
.A(n_10230),
.Y(n_11055)
);

BUFx6f_ASAP7_75t_L g11056 ( 
.A(n_10230),
.Y(n_11056)
);

NAND2xp5_ASAP7_75t_SL g11057 ( 
.A(n_10014),
.B(n_921),
.Y(n_11057)
);

INVx1_ASAP7_75t_L g11058 ( 
.A(n_10249),
.Y(n_11058)
);

OAI21xp5_ASAP7_75t_L g11059 ( 
.A1(n_9990),
.A2(n_924),
.B(n_925),
.Y(n_11059)
);

BUFx6f_ASAP7_75t_L g11060 ( 
.A(n_9836),
.Y(n_11060)
);

INVx3_ASAP7_75t_SL g11061 ( 
.A(n_10440),
.Y(n_11061)
);

NAND2xp5_ASAP7_75t_L g11062 ( 
.A(n_9978),
.B(n_925),
.Y(n_11062)
);

AND2x4_ASAP7_75t_L g11063 ( 
.A(n_10204),
.B(n_926),
.Y(n_11063)
);

A2O1A1Ixp33_ASAP7_75t_L g11064 ( 
.A1(n_10175),
.A2(n_928),
.B(n_926),
.C(n_927),
.Y(n_11064)
);

NAND2xp5_ASAP7_75t_SL g11065 ( 
.A(n_9895),
.B(n_927),
.Y(n_11065)
);

NAND2xp5_ASAP7_75t_L g11066 ( 
.A(n_9979),
.B(n_928),
.Y(n_11066)
);

NAND2xp5_ASAP7_75t_SL g11067 ( 
.A(n_9927),
.B(n_929),
.Y(n_11067)
);

NOR2xp33_ASAP7_75t_R g11068 ( 
.A(n_10242),
.B(n_929),
.Y(n_11068)
);

NOR2xp33_ASAP7_75t_L g11069 ( 
.A(n_10254),
.B(n_930),
.Y(n_11069)
);

NOR2xp33_ASAP7_75t_R g11070 ( 
.A(n_10017),
.B(n_930),
.Y(n_11070)
);

AOI21xp5_ASAP7_75t_L g11071 ( 
.A1(n_10050),
.A2(n_931),
.B(n_932),
.Y(n_11071)
);

AND2x4_ASAP7_75t_L g11072 ( 
.A(n_9982),
.B(n_931),
.Y(n_11072)
);

NAND2xp5_ASAP7_75t_L g11073 ( 
.A(n_9984),
.B(n_933),
.Y(n_11073)
);

AOI21xp5_ASAP7_75t_L g11074 ( 
.A1(n_10055),
.A2(n_934),
.B(n_935),
.Y(n_11074)
);

O2A1O1Ixp33_ASAP7_75t_SL g11075 ( 
.A1(n_10261),
.A2(n_937),
.B(n_934),
.C(n_935),
.Y(n_11075)
);

OAI21xp5_ASAP7_75t_L g11076 ( 
.A1(n_9994),
.A2(n_937),
.B(n_938),
.Y(n_11076)
);

INVx2_ASAP7_75t_L g11077 ( 
.A(n_9872),
.Y(n_11077)
);

A2O1A1Ixp33_ASAP7_75t_L g11078 ( 
.A1(n_10201),
.A2(n_940),
.B(n_938),
.C(n_939),
.Y(n_11078)
);

BUFx2_ASAP7_75t_L g11079 ( 
.A(n_10197),
.Y(n_11079)
);

AOI22xp33_ASAP7_75t_L g11080 ( 
.A1(n_10336),
.A2(n_10320),
.B1(n_10210),
.B2(n_10212),
.Y(n_11080)
);

NOR3xp33_ASAP7_75t_SL g11081 ( 
.A(n_10075),
.B(n_939),
.C(n_940),
.Y(n_11081)
);

NAND2xp5_ASAP7_75t_L g11082 ( 
.A(n_10001),
.B(n_941),
.Y(n_11082)
);

CKINVDCx11_ASAP7_75t_R g11083 ( 
.A(n_9950),
.Y(n_11083)
);

NOR2xp33_ASAP7_75t_L g11084 ( 
.A(n_10251),
.B(n_941),
.Y(n_11084)
);

NAND2xp5_ASAP7_75t_SL g11085 ( 
.A(n_9855),
.B(n_942),
.Y(n_11085)
);

AOI21xp5_ASAP7_75t_L g11086 ( 
.A1(n_10068),
.A2(n_943),
.B(n_944),
.Y(n_11086)
);

INVx8_ASAP7_75t_L g11087 ( 
.A(n_10027),
.Y(n_11087)
);

CKINVDCx5p33_ASAP7_75t_R g11088 ( 
.A(n_9946),
.Y(n_11088)
);

NAND2xp5_ASAP7_75t_L g11089 ( 
.A(n_10008),
.B(n_943),
.Y(n_11089)
);

AOI21xp5_ASAP7_75t_L g11090 ( 
.A1(n_10071),
.A2(n_944),
.B(n_945),
.Y(n_11090)
);

BUFx3_ASAP7_75t_L g11091 ( 
.A(n_10062),
.Y(n_11091)
);

AOI21xp5_ASAP7_75t_L g11092 ( 
.A1(n_10072),
.A2(n_946),
.B(n_947),
.Y(n_11092)
);

NAND2xp5_ASAP7_75t_L g11093 ( 
.A(n_10057),
.B(n_947),
.Y(n_11093)
);

A2O1A1Ixp33_ASAP7_75t_L g11094 ( 
.A1(n_10209),
.A2(n_950),
.B(n_948),
.C(n_949),
.Y(n_11094)
);

OAI22x1_ASAP7_75t_L g11095 ( 
.A1(n_10203),
.A2(n_10267),
.B1(n_10059),
.B2(n_10195),
.Y(n_11095)
);

NOR2xp33_ASAP7_75t_L g11096 ( 
.A(n_10248),
.B(n_948),
.Y(n_11096)
);

AOI21xp5_ASAP7_75t_L g11097 ( 
.A1(n_10096),
.A2(n_950),
.B(n_952),
.Y(n_11097)
);

OAI22xp5_ASAP7_75t_L g11098 ( 
.A1(n_9977),
.A2(n_954),
.B1(n_952),
.B2(n_953),
.Y(n_11098)
);

AOI21xp5_ASAP7_75t_L g11099 ( 
.A1(n_10097),
.A2(n_953),
.B(n_954),
.Y(n_11099)
);

AOI22xp33_ASAP7_75t_L g11100 ( 
.A1(n_10002),
.A2(n_957),
.B1(n_955),
.B2(n_956),
.Y(n_11100)
);

NOR2xp33_ASAP7_75t_L g11101 ( 
.A(n_10314),
.B(n_955),
.Y(n_11101)
);

O2A1O1Ixp33_ASAP7_75t_L g11102 ( 
.A1(n_10005),
.A2(n_959),
.B(n_956),
.C(n_957),
.Y(n_11102)
);

INVx2_ASAP7_75t_SL g11103 ( 
.A(n_10073),
.Y(n_11103)
);

INVx1_ASAP7_75t_L g11104 ( 
.A(n_9823),
.Y(n_11104)
);

INVx2_ASAP7_75t_SL g11105 ( 
.A(n_10076),
.Y(n_11105)
);

NAND2xp5_ASAP7_75t_L g11106 ( 
.A(n_9952),
.B(n_960),
.Y(n_11106)
);

AOI21xp5_ASAP7_75t_L g11107 ( 
.A1(n_10099),
.A2(n_960),
.B(n_961),
.Y(n_11107)
);

O2A1O1Ixp33_ASAP7_75t_L g11108 ( 
.A1(n_10006),
.A2(n_963),
.B(n_961),
.C(n_962),
.Y(n_11108)
);

AND2x2_ASAP7_75t_L g11109 ( 
.A(n_10177),
.B(n_10236),
.Y(n_11109)
);

AO32x2_ASAP7_75t_L g11110 ( 
.A1(n_10100),
.A2(n_964),
.A3(n_962),
.B1(n_963),
.B2(n_965),
.Y(n_11110)
);

A2O1A1Ixp33_ASAP7_75t_SL g11111 ( 
.A1(n_10176),
.A2(n_967),
.B(n_965),
.C(n_966),
.Y(n_11111)
);

AND2x2_ASAP7_75t_L g11112 ( 
.A(n_10237),
.B(n_966),
.Y(n_11112)
);

AOI22xp5_ASAP7_75t_L g11113 ( 
.A1(n_10148),
.A2(n_969),
.B1(n_967),
.B2(n_968),
.Y(n_11113)
);

NAND2xp5_ASAP7_75t_SL g11114 ( 
.A(n_9886),
.B(n_968),
.Y(n_11114)
);

AOI21xp5_ASAP7_75t_L g11115 ( 
.A1(n_10105),
.A2(n_969),
.B(n_970),
.Y(n_11115)
);

INVx3_ASAP7_75t_L g11116 ( 
.A(n_10225),
.Y(n_11116)
);

INVx1_ASAP7_75t_L g11117 ( 
.A(n_10410),
.Y(n_11117)
);

NOR2xp33_ASAP7_75t_L g11118 ( 
.A(n_10199),
.B(n_971),
.Y(n_11118)
);

NAND2xp5_ASAP7_75t_L g11119 ( 
.A(n_10010),
.B(n_971),
.Y(n_11119)
);

NAND3xp33_ASAP7_75t_SL g11120 ( 
.A(n_10270),
.B(n_972),
.C(n_973),
.Y(n_11120)
);

A2O1A1Ixp33_ASAP7_75t_L g11121 ( 
.A1(n_10362),
.A2(n_975),
.B(n_973),
.C(n_974),
.Y(n_11121)
);

AOI22xp33_ASAP7_75t_L g11122 ( 
.A1(n_10307),
.A2(n_10265),
.B1(n_10275),
.B2(n_10308),
.Y(n_11122)
);

NAND2xp5_ASAP7_75t_L g11123 ( 
.A(n_10224),
.B(n_974),
.Y(n_11123)
);

A2O1A1Ixp33_ASAP7_75t_L g11124 ( 
.A1(n_10395),
.A2(n_977),
.B(n_975),
.C(n_976),
.Y(n_11124)
);

NOR2x1_ASAP7_75t_R g11125 ( 
.A(n_10220),
.B(n_976),
.Y(n_11125)
);

INVx5_ASAP7_75t_L g11126 ( 
.A(n_10322),
.Y(n_11126)
);

INVx1_ASAP7_75t_L g11127 ( 
.A(n_10432),
.Y(n_11127)
);

AOI21xp5_ASAP7_75t_L g11128 ( 
.A1(n_10123),
.A2(n_978),
.B(n_979),
.Y(n_11128)
);

NAND2xp5_ASAP7_75t_L g11129 ( 
.A(n_10238),
.B(n_978),
.Y(n_11129)
);

NAND2xp5_ASAP7_75t_L g11130 ( 
.A(n_10084),
.B(n_979),
.Y(n_11130)
);

NOR2x1_ASAP7_75t_L g11131 ( 
.A(n_10136),
.B(n_981),
.Y(n_11131)
);

NAND2x1p5_ASAP7_75t_L g11132 ( 
.A(n_10228),
.B(n_981),
.Y(n_11132)
);

AND2x2_ASAP7_75t_L g11133 ( 
.A(n_10253),
.B(n_982),
.Y(n_11133)
);

HB1xp67_ASAP7_75t_SL g11134 ( 
.A(n_9829),
.Y(n_11134)
);

AOI21xp5_ASAP7_75t_L g11135 ( 
.A1(n_10126),
.A2(n_982),
.B(n_983),
.Y(n_11135)
);

NOR2xp33_ASAP7_75t_L g11136 ( 
.A(n_10153),
.B(n_983),
.Y(n_11136)
);

NAND3xp33_ASAP7_75t_SL g11137 ( 
.A(n_10279),
.B(n_984),
.C(n_985),
.Y(n_11137)
);

BUFx2_ASAP7_75t_L g11138 ( 
.A(n_10208),
.Y(n_11138)
);

AOI21xp5_ASAP7_75t_L g11139 ( 
.A1(n_10023),
.A2(n_984),
.B(n_986),
.Y(n_11139)
);

NOR2xp33_ASAP7_75t_R g11140 ( 
.A(n_10485),
.B(n_986),
.Y(n_11140)
);

NAND2xp5_ASAP7_75t_L g11141 ( 
.A(n_10098),
.B(n_987),
.Y(n_11141)
);

NAND2xp5_ASAP7_75t_L g11142 ( 
.A(n_10280),
.B(n_987),
.Y(n_11142)
);

AND2x2_ASAP7_75t_L g11143 ( 
.A(n_10301),
.B(n_988),
.Y(n_11143)
);

NAND2xp5_ASAP7_75t_SL g11144 ( 
.A(n_10337),
.B(n_989),
.Y(n_11144)
);

NAND2xp5_ASAP7_75t_SL g11145 ( 
.A(n_10447),
.B(n_989),
.Y(n_11145)
);

AOI22xp33_ASAP7_75t_L g11146 ( 
.A1(n_10184),
.A2(n_992),
.B1(n_990),
.B2(n_991),
.Y(n_11146)
);

NAND2xp33_ASAP7_75t_L g11147 ( 
.A(n_10264),
.B(n_991),
.Y(n_11147)
);

INVx2_ASAP7_75t_L g11148 ( 
.A(n_10258),
.Y(n_11148)
);

INVx1_ASAP7_75t_L g11149 ( 
.A(n_10298),
.Y(n_11149)
);

AOI22xp5_ASAP7_75t_L g11150 ( 
.A1(n_10317),
.A2(n_994),
.B1(n_992),
.B2(n_993),
.Y(n_11150)
);

AOI21xp5_ASAP7_75t_L g11151 ( 
.A1(n_10034),
.A2(n_993),
.B(n_995),
.Y(n_11151)
);

CKINVDCx5p33_ASAP7_75t_R g11152 ( 
.A(n_9843),
.Y(n_11152)
);

AOI21xp5_ASAP7_75t_L g11153 ( 
.A1(n_10035),
.A2(n_995),
.B(n_996),
.Y(n_11153)
);

AOI22xp33_ASAP7_75t_L g11154 ( 
.A1(n_10200),
.A2(n_998),
.B1(n_996),
.B2(n_997),
.Y(n_11154)
);

INVx2_ASAP7_75t_SL g11155 ( 
.A(n_10277),
.Y(n_11155)
);

INVx3_ASAP7_75t_L g11156 ( 
.A(n_10323),
.Y(n_11156)
);

NAND2xp5_ASAP7_75t_SL g11157 ( 
.A(n_10449),
.B(n_997),
.Y(n_11157)
);

NOR2xp33_ASAP7_75t_L g11158 ( 
.A(n_10155),
.B(n_998),
.Y(n_11158)
);

NOR2xp33_ASAP7_75t_R g11159 ( 
.A(n_10309),
.B(n_999),
.Y(n_11159)
);

INVx1_ASAP7_75t_L g11160 ( 
.A(n_10243),
.Y(n_11160)
);

INVx1_ASAP7_75t_L g11161 ( 
.A(n_10138),
.Y(n_11161)
);

INVx1_ASAP7_75t_L g11162 ( 
.A(n_10141),
.Y(n_11162)
);

O2A1O1Ixp5_ASAP7_75t_L g11163 ( 
.A1(n_9882),
.A2(n_1001),
.B(n_999),
.C(n_1000),
.Y(n_11163)
);

INVx2_ASAP7_75t_L g11164 ( 
.A(n_10282),
.Y(n_11164)
);

INVx2_ASAP7_75t_L g11165 ( 
.A(n_10285),
.Y(n_11165)
);

NOR2x1_ASAP7_75t_L g11166 ( 
.A(n_10482),
.B(n_1000),
.Y(n_11166)
);

OAI22xp5_ASAP7_75t_L g11167 ( 
.A1(n_10488),
.A2(n_1003),
.B1(n_1001),
.B2(n_1002),
.Y(n_11167)
);

AND2x4_ASAP7_75t_L g11168 ( 
.A(n_10303),
.B(n_1002),
.Y(n_11168)
);

NAND2xp5_ASAP7_75t_L g11169 ( 
.A(n_10295),
.B(n_1003),
.Y(n_11169)
);

AO32x1_ASAP7_75t_L g11170 ( 
.A1(n_9951),
.A2(n_9840),
.A3(n_10074),
.B1(n_10341),
.B2(n_10135),
.Y(n_11170)
);

AOI21xp5_ASAP7_75t_L g11171 ( 
.A1(n_10036),
.A2(n_1004),
.B(n_1005),
.Y(n_11171)
);

NAND2xp5_ASAP7_75t_L g11172 ( 
.A(n_10296),
.B(n_1004),
.Y(n_11172)
);

NAND2xp5_ASAP7_75t_L g11173 ( 
.A(n_10305),
.B(n_1005),
.Y(n_11173)
);

AOI21xp5_ASAP7_75t_L g11174 ( 
.A1(n_10038),
.A2(n_1006),
.B(n_1007),
.Y(n_11174)
);

NAND2xp5_ASAP7_75t_L g11175 ( 
.A(n_10306),
.B(n_1008),
.Y(n_11175)
);

AND2x2_ASAP7_75t_L g11176 ( 
.A(n_10244),
.B(n_1009),
.Y(n_11176)
);

A2O1A1Ixp33_ASAP7_75t_L g11177 ( 
.A1(n_10483),
.A2(n_1011),
.B(n_1009),
.C(n_1010),
.Y(n_11177)
);

CKINVDCx5p33_ASAP7_75t_R g11178 ( 
.A(n_9845),
.Y(n_11178)
);

NOR2xp33_ASAP7_75t_L g11179 ( 
.A(n_10162),
.B(n_1011),
.Y(n_11179)
);

INVxp67_ASAP7_75t_L g11180 ( 
.A(n_10065),
.Y(n_11180)
);

BUFx8_ASAP7_75t_L g11181 ( 
.A(n_10291),
.Y(n_11181)
);

NAND2xp5_ASAP7_75t_L g11182 ( 
.A(n_9906),
.B(n_1012),
.Y(n_11182)
);

BUFx6f_ASAP7_75t_L g11183 ( 
.A(n_10327),
.Y(n_11183)
);

AND2x2_ASAP7_75t_L g11184 ( 
.A(n_10119),
.B(n_1012),
.Y(n_11184)
);

NOR2xp33_ASAP7_75t_L g11185 ( 
.A(n_10329),
.B(n_1013),
.Y(n_11185)
);

BUFx6f_ASAP7_75t_L g11186 ( 
.A(n_10218),
.Y(n_11186)
);

BUFx6f_ASAP7_75t_L g11187 ( 
.A(n_10132),
.Y(n_11187)
);

A2O1A1Ixp33_ASAP7_75t_SL g11188 ( 
.A1(n_9893),
.A2(n_1016),
.B(n_1014),
.C(n_1015),
.Y(n_11188)
);

INVx1_ASAP7_75t_L g11189 ( 
.A(n_10145),
.Y(n_11189)
);

NOR3xp33_ASAP7_75t_SL g11190 ( 
.A(n_10281),
.B(n_1014),
.C(n_1015),
.Y(n_11190)
);

OAI22xp33_ASAP7_75t_L g11191 ( 
.A1(n_10286),
.A2(n_1018),
.B1(n_1016),
.B2(n_1017),
.Y(n_11191)
);

AOI21xp5_ASAP7_75t_L g11192 ( 
.A1(n_9949),
.A2(n_1017),
.B(n_1018),
.Y(n_11192)
);

AOI21xp5_ASAP7_75t_L g11193 ( 
.A1(n_9957),
.A2(n_1019),
.B(n_1020),
.Y(n_11193)
);

AOI21xp5_ASAP7_75t_L g11194 ( 
.A1(n_9959),
.A2(n_1019),
.B(n_1020),
.Y(n_11194)
);

NOR2xp33_ASAP7_75t_L g11195 ( 
.A(n_10167),
.B(n_1021),
.Y(n_11195)
);

AND2x2_ASAP7_75t_SL g11196 ( 
.A(n_10514),
.B(n_9915),
.Y(n_11196)
);

INVx1_ASAP7_75t_L g11197 ( 
.A(n_10152),
.Y(n_11197)
);

A2O1A1Ixp33_ASAP7_75t_L g11198 ( 
.A1(n_10339),
.A2(n_1024),
.B(n_1022),
.C(n_1023),
.Y(n_11198)
);

AOI21xp5_ASAP7_75t_L g11199 ( 
.A1(n_9964),
.A2(n_1022),
.B(n_1025),
.Y(n_11199)
);

CKINVDCx8_ASAP7_75t_R g11200 ( 
.A(n_10330),
.Y(n_11200)
);

NOR2xp33_ASAP7_75t_L g11201 ( 
.A(n_10311),
.B(n_1025),
.Y(n_11201)
);

AOI21xp5_ASAP7_75t_L g11202 ( 
.A1(n_10154),
.A2(n_1026),
.B(n_1027),
.Y(n_11202)
);

AOI21xp5_ASAP7_75t_L g11203 ( 
.A1(n_10157),
.A2(n_1026),
.B(n_1027),
.Y(n_11203)
);

A2O1A1Ixp33_ASAP7_75t_L g11204 ( 
.A1(n_9916),
.A2(n_1030),
.B(n_1028),
.C(n_1029),
.Y(n_11204)
);

AND2x4_ASAP7_75t_L g11205 ( 
.A(n_9980),
.B(n_1030),
.Y(n_11205)
);

A2O1A1Ixp33_ASAP7_75t_L g11206 ( 
.A1(n_9918),
.A2(n_1033),
.B(n_1031),
.C(n_1032),
.Y(n_11206)
);

INVx2_ASAP7_75t_L g11207 ( 
.A(n_10216),
.Y(n_11207)
);

NOR3xp33_ASAP7_75t_SL g11208 ( 
.A(n_10256),
.B(n_1032),
.C(n_1033),
.Y(n_11208)
);

NOR3xp33_ASAP7_75t_SL g11209 ( 
.A(n_10115),
.B(n_1034),
.C(n_1035),
.Y(n_11209)
);

O2A1O1Ixp33_ASAP7_75t_L g11210 ( 
.A1(n_10297),
.A2(n_10304),
.B(n_9938),
.C(n_9944),
.Y(n_11210)
);

AOI21xp5_ASAP7_75t_L g11211 ( 
.A1(n_10159),
.A2(n_1036),
.B(n_1037),
.Y(n_11211)
);

HB1xp67_ASAP7_75t_L g11212 ( 
.A(n_10271),
.Y(n_11212)
);

NOR2xp33_ASAP7_75t_L g11213 ( 
.A(n_10321),
.B(n_10316),
.Y(n_11213)
);

NAND2xp5_ASAP7_75t_L g11214 ( 
.A(n_9919),
.B(n_1036),
.Y(n_11214)
);

OAI22xp5_ASAP7_75t_L g11215 ( 
.A1(n_10252),
.A2(n_1039),
.B1(n_1037),
.B2(n_1038),
.Y(n_11215)
);

OR2x2_ASAP7_75t_L g11216 ( 
.A(n_10165),
.B(n_1038),
.Y(n_11216)
);

NOR3xp33_ASAP7_75t_L g11217 ( 
.A(n_10292),
.B(n_1039),
.C(n_1040),
.Y(n_11217)
);

AOI21xp5_ASAP7_75t_L g11218 ( 
.A1(n_10170),
.A2(n_1040),
.B(n_1042),
.Y(n_11218)
);

INVx1_ASAP7_75t_L g11219 ( 
.A(n_10186),
.Y(n_11219)
);

NOR2xp67_ASAP7_75t_L g11220 ( 
.A(n_9986),
.B(n_1042),
.Y(n_11220)
);

NAND2xp5_ASAP7_75t_L g11221 ( 
.A(n_10268),
.B(n_1043),
.Y(n_11221)
);

AOI21xp5_ASAP7_75t_L g11222 ( 
.A1(n_9885),
.A2(n_1043),
.B(n_1044),
.Y(n_11222)
);

INVx1_ASAP7_75t_L g11223 ( 
.A(n_10458),
.Y(n_11223)
);

INVx1_ASAP7_75t_L g11224 ( 
.A(n_10458),
.Y(n_11224)
);

AND2x4_ASAP7_75t_L g11225 ( 
.A(n_9848),
.B(n_1044),
.Y(n_11225)
);

O2A1O1Ixp33_ASAP7_75t_L g11226 ( 
.A1(n_10534),
.A2(n_1047),
.B(n_1045),
.C(n_1046),
.Y(n_11226)
);

AOI21xp5_ASAP7_75t_L g11227 ( 
.A1(n_9885),
.A2(n_1046),
.B(n_1047),
.Y(n_11227)
);

NAND2xp5_ASAP7_75t_SL g11228 ( 
.A(n_9888),
.B(n_1048),
.Y(n_11228)
);

AOI21xp5_ASAP7_75t_L g11229 ( 
.A1(n_9885),
.A2(n_1048),
.B(n_1049),
.Y(n_11229)
);

INVx1_ASAP7_75t_L g11230 ( 
.A(n_10458),
.Y(n_11230)
);

INVx2_ASAP7_75t_L g11231 ( 
.A(n_10088),
.Y(n_11231)
);

OAI22xp5_ASAP7_75t_L g11232 ( 
.A1(n_9837),
.A2(n_1052),
.B1(n_1050),
.B2(n_1051),
.Y(n_11232)
);

INVx1_ASAP7_75t_L g11233 ( 
.A(n_10458),
.Y(n_11233)
);

A2O1A1Ixp33_ASAP7_75t_L g11234 ( 
.A1(n_9837),
.A2(n_1053),
.B(n_1050),
.C(n_1052),
.Y(n_11234)
);

AOI21xp5_ASAP7_75t_L g11235 ( 
.A1(n_9885),
.A2(n_1053),
.B(n_1054),
.Y(n_11235)
);

OAI22x1_ASAP7_75t_L g11236 ( 
.A1(n_9837),
.A2(n_1056),
.B1(n_1054),
.B2(n_1055),
.Y(n_11236)
);

CKINVDCx5p33_ASAP7_75t_R g11237 ( 
.A(n_10345),
.Y(n_11237)
);

INVx1_ASAP7_75t_L g11238 ( 
.A(n_10458),
.Y(n_11238)
);

NAND2xp5_ASAP7_75t_L g11239 ( 
.A(n_10458),
.B(n_1055),
.Y(n_11239)
);

AOI22xp5_ASAP7_75t_L g11240 ( 
.A1(n_9837),
.A2(n_1059),
.B1(n_1057),
.B2(n_1058),
.Y(n_11240)
);

AOI21xp33_ASAP7_75t_L g11241 ( 
.A1(n_9837),
.A2(n_1057),
.B(n_1058),
.Y(n_11241)
);

BUFx6f_ASAP7_75t_L g11242 ( 
.A(n_10451),
.Y(n_11242)
);

NOR2xp33_ASAP7_75t_L g11243 ( 
.A(n_9837),
.B(n_1059),
.Y(n_11243)
);

NAND2xp5_ASAP7_75t_SL g11244 ( 
.A(n_9888),
.B(n_1060),
.Y(n_11244)
);

NAND2xp5_ASAP7_75t_L g11245 ( 
.A(n_10458),
.B(n_1060),
.Y(n_11245)
);

NAND2xp5_ASAP7_75t_L g11246 ( 
.A(n_10458),
.B(n_1061),
.Y(n_11246)
);

INVx1_ASAP7_75t_L g11247 ( 
.A(n_10458),
.Y(n_11247)
);

NOR3xp33_ASAP7_75t_L g11248 ( 
.A(n_9909),
.B(n_1061),
.C(n_1062),
.Y(n_11248)
);

NAND2xp5_ASAP7_75t_L g11249 ( 
.A(n_10458),
.B(n_1062),
.Y(n_11249)
);

INVx1_ASAP7_75t_SL g11250 ( 
.A(n_10106),
.Y(n_11250)
);

A2O1A1Ixp33_ASAP7_75t_L g11251 ( 
.A1(n_9837),
.A2(n_1065),
.B(n_1063),
.C(n_1064),
.Y(n_11251)
);

INVx1_ASAP7_75t_SL g11252 ( 
.A(n_10106),
.Y(n_11252)
);

AOI21xp5_ASAP7_75t_L g11253 ( 
.A1(n_9885),
.A2(n_1063),
.B(n_1064),
.Y(n_11253)
);

INVx1_ASAP7_75t_L g11254 ( 
.A(n_10458),
.Y(n_11254)
);

OAI22xp5_ASAP7_75t_L g11255 ( 
.A1(n_9837),
.A2(n_1067),
.B1(n_1065),
.B2(n_1066),
.Y(n_11255)
);

A2O1A1Ixp33_ASAP7_75t_L g11256 ( 
.A1(n_9837),
.A2(n_1069),
.B(n_1066),
.C(n_1068),
.Y(n_11256)
);

AOI22xp5_ASAP7_75t_L g11257 ( 
.A1(n_9837),
.A2(n_1070),
.B1(n_1068),
.B2(n_1069),
.Y(n_11257)
);

INVx1_ASAP7_75t_L g11258 ( 
.A(n_10458),
.Y(n_11258)
);

INVx1_ASAP7_75t_SL g11259 ( 
.A(n_10106),
.Y(n_11259)
);

INVx2_ASAP7_75t_L g11260 ( 
.A(n_10088),
.Y(n_11260)
);

INVxp67_ASAP7_75t_SL g11261 ( 
.A(n_10458),
.Y(n_11261)
);

NAND2xp5_ASAP7_75t_L g11262 ( 
.A(n_10458),
.B(n_1070),
.Y(n_11262)
);

BUFx6f_ASAP7_75t_L g11263 ( 
.A(n_10838),
.Y(n_11263)
);

NAND2xp5_ASAP7_75t_L g11264 ( 
.A(n_10737),
.B(n_1071),
.Y(n_11264)
);

AOI21xp5_ASAP7_75t_L g11265 ( 
.A1(n_10542),
.A2(n_1071),
.B(n_1072),
.Y(n_11265)
);

OAI21x1_ASAP7_75t_L g11266 ( 
.A1(n_10582),
.A2(n_1072),
.B(n_1073),
.Y(n_11266)
);

NAND2xp5_ASAP7_75t_L g11267 ( 
.A(n_10560),
.B(n_1073),
.Y(n_11267)
);

OAI21x1_ASAP7_75t_L g11268 ( 
.A1(n_10590),
.A2(n_1074),
.B(n_1075),
.Y(n_11268)
);

AOI211x1_ASAP7_75t_L g11269 ( 
.A1(n_10572),
.A2(n_1077),
.B(n_1074),
.C(n_1076),
.Y(n_11269)
);

OAI21x1_ASAP7_75t_L g11270 ( 
.A1(n_10773),
.A2(n_1076),
.B(n_1077),
.Y(n_11270)
);

OAI21xp5_ASAP7_75t_L g11271 ( 
.A1(n_10979),
.A2(n_11022),
.B(n_11210),
.Y(n_11271)
);

OAI21x1_ASAP7_75t_L g11272 ( 
.A1(n_10735),
.A2(n_1078),
.B(n_1079),
.Y(n_11272)
);

OAI21x1_ASAP7_75t_L g11273 ( 
.A1(n_11043),
.A2(n_1078),
.B(n_1079),
.Y(n_11273)
);

NAND2xp5_ASAP7_75t_L g11274 ( 
.A(n_10575),
.B(n_1080),
.Y(n_11274)
);

NOR2x1_ASAP7_75t_L g11275 ( 
.A(n_10917),
.B(n_1080),
.Y(n_11275)
);

NAND2xp5_ASAP7_75t_L g11276 ( 
.A(n_11261),
.B(n_1081),
.Y(n_11276)
);

NAND2x1_ASAP7_75t_L g11277 ( 
.A(n_11223),
.B(n_1081),
.Y(n_11277)
);

OAI21x1_ASAP7_75t_L g11278 ( 
.A1(n_10791),
.A2(n_1082),
.B(n_1083),
.Y(n_11278)
);

OAI21x1_ASAP7_75t_L g11279 ( 
.A1(n_11161),
.A2(n_1082),
.B(n_1083),
.Y(n_11279)
);

OAI21xp5_ASAP7_75t_L g11280 ( 
.A1(n_10732),
.A2(n_10704),
.B(n_10847),
.Y(n_11280)
);

NAND2x1_ASAP7_75t_L g11281 ( 
.A(n_11224),
.B(n_1084),
.Y(n_11281)
);

BUFx5_ASAP7_75t_L g11282 ( 
.A(n_11058),
.Y(n_11282)
);

OA22x2_ASAP7_75t_L g11283 ( 
.A1(n_10541),
.A2(n_1087),
.B1(n_1084),
.B2(n_1086),
.Y(n_11283)
);

NAND2xp5_ASAP7_75t_SL g11284 ( 
.A(n_10567),
.B(n_11126),
.Y(n_11284)
);

OAI21x1_ASAP7_75t_L g11285 ( 
.A1(n_11162),
.A2(n_1087),
.B(n_1088),
.Y(n_11285)
);

INVx2_ASAP7_75t_L g11286 ( 
.A(n_10599),
.Y(n_11286)
);

AND2x2_ASAP7_75t_L g11287 ( 
.A(n_10571),
.B(n_1089),
.Y(n_11287)
);

AND2x2_ASAP7_75t_L g11288 ( 
.A(n_10570),
.B(n_1089),
.Y(n_11288)
);

AOI21x1_ASAP7_75t_L g11289 ( 
.A1(n_10608),
.A2(n_1090),
.B(n_1091),
.Y(n_11289)
);

NAND2xp5_ASAP7_75t_L g11290 ( 
.A(n_11230),
.B(n_1090),
.Y(n_11290)
);

NOR2x1_ASAP7_75t_SL g11291 ( 
.A(n_11126),
.B(n_10567),
.Y(n_11291)
);

INVxp67_ASAP7_75t_SL g11292 ( 
.A(n_10828),
.Y(n_11292)
);

AND2x4_ASAP7_75t_L g11293 ( 
.A(n_10584),
.B(n_1091),
.Y(n_11293)
);

OAI21xp5_ASAP7_75t_L g11294 ( 
.A1(n_10717),
.A2(n_1092),
.B(n_1093),
.Y(n_11294)
);

OAI21xp5_ASAP7_75t_L g11295 ( 
.A1(n_10710),
.A2(n_1092),
.B(n_1093),
.Y(n_11295)
);

CKINVDCx8_ASAP7_75t_R g11296 ( 
.A(n_10908),
.Y(n_11296)
);

OAI22xp5_ASAP7_75t_L g11297 ( 
.A1(n_10875),
.A2(n_1099),
.B1(n_1097),
.B2(n_1098),
.Y(n_11297)
);

A2O1A1Ixp33_ASAP7_75t_SL g11298 ( 
.A1(n_11243),
.A2(n_1100),
.B(n_1097),
.C(n_1099),
.Y(n_11298)
);

NAND2xp33_ASAP7_75t_SL g11299 ( 
.A(n_11068),
.B(n_1101),
.Y(n_11299)
);

BUFx12f_ASAP7_75t_L g11300 ( 
.A(n_10546),
.Y(n_11300)
);

AND2x4_ASAP7_75t_L g11301 ( 
.A(n_10592),
.B(n_1101),
.Y(n_11301)
);

AND2x2_ASAP7_75t_L g11302 ( 
.A(n_10615),
.B(n_1102),
.Y(n_11302)
);

INVx5_ASAP7_75t_L g11303 ( 
.A(n_10597),
.Y(n_11303)
);

OAI21x1_ASAP7_75t_L g11304 ( 
.A1(n_11189),
.A2(n_11197),
.B(n_11219),
.Y(n_11304)
);

INVx1_ASAP7_75t_L g11305 ( 
.A(n_10612),
.Y(n_11305)
);

OAI21x1_ASAP7_75t_L g11306 ( 
.A1(n_11046),
.A2(n_1103),
.B(n_1104),
.Y(n_11306)
);

AND2x2_ASAP7_75t_L g11307 ( 
.A(n_10654),
.B(n_1103),
.Y(n_11307)
);

CKINVDCx8_ASAP7_75t_R g11308 ( 
.A(n_11237),
.Y(n_11308)
);

NOR2x1_ASAP7_75t_SL g11309 ( 
.A(n_11126),
.B(n_1106),
.Y(n_11309)
);

INVx6_ASAP7_75t_L g11310 ( 
.A(n_10832),
.Y(n_11310)
);

BUFx10_ASAP7_75t_L g11311 ( 
.A(n_10838),
.Y(n_11311)
);

BUFx6f_ASAP7_75t_L g11312 ( 
.A(n_10867),
.Y(n_11312)
);

AOI21xp5_ASAP7_75t_L g11313 ( 
.A1(n_10861),
.A2(n_1106),
.B(n_1107),
.Y(n_11313)
);

OAI21xp5_ASAP7_75t_L g11314 ( 
.A1(n_11222),
.A2(n_1107),
.B(n_1108),
.Y(n_11314)
);

NAND2xp5_ASAP7_75t_L g11315 ( 
.A(n_11233),
.B(n_1109),
.Y(n_11315)
);

BUFx2_ASAP7_75t_L g11316 ( 
.A(n_10581),
.Y(n_11316)
);

NAND2xp5_ASAP7_75t_L g11317 ( 
.A(n_11238),
.B(n_1109),
.Y(n_11317)
);

OAI22xp5_ASAP7_75t_L g11318 ( 
.A1(n_10969),
.A2(n_1112),
.B1(n_1110),
.B2(n_1111),
.Y(n_11318)
);

NAND2xp5_ASAP7_75t_L g11319 ( 
.A(n_11247),
.B(n_11254),
.Y(n_11319)
);

NAND2xp5_ASAP7_75t_L g11320 ( 
.A(n_11258),
.B(n_1110),
.Y(n_11320)
);

BUFx6f_ASAP7_75t_L g11321 ( 
.A(n_10867),
.Y(n_11321)
);

INVx1_ASAP7_75t_L g11322 ( 
.A(n_10545),
.Y(n_11322)
);

CKINVDCx11_ASAP7_75t_R g11323 ( 
.A(n_10672),
.Y(n_11323)
);

NOR2xp33_ASAP7_75t_L g11324 ( 
.A(n_10905),
.B(n_1111),
.Y(n_11324)
);

OAI21x1_ASAP7_75t_L g11325 ( 
.A1(n_11077),
.A2(n_1112),
.B(n_1113),
.Y(n_11325)
);

BUFx2_ASAP7_75t_L g11326 ( 
.A(n_10893),
.Y(n_11326)
);

INVx3_ASAP7_75t_L g11327 ( 
.A(n_10544),
.Y(n_11327)
);

OAI21x1_ASAP7_75t_L g11328 ( 
.A1(n_11034),
.A2(n_1113),
.B(n_1114),
.Y(n_11328)
);

AO21x2_ASAP7_75t_L g11329 ( 
.A1(n_11045),
.A2(n_11117),
.B(n_11104),
.Y(n_11329)
);

NAND2xp5_ASAP7_75t_L g11330 ( 
.A(n_10885),
.B(n_1114),
.Y(n_11330)
);

AOI21x1_ASAP7_75t_L g11331 ( 
.A1(n_10751),
.A2(n_10862),
.B(n_11017),
.Y(n_11331)
);

BUFx3_ASAP7_75t_L g11332 ( 
.A(n_11052),
.Y(n_11332)
);

OAI21x1_ASAP7_75t_L g11333 ( 
.A1(n_10715),
.A2(n_1115),
.B(n_1117),
.Y(n_11333)
);

OAI21x1_ASAP7_75t_L g11334 ( 
.A1(n_11039),
.A2(n_1115),
.B(n_1117),
.Y(n_11334)
);

INVx4_ASAP7_75t_L g11335 ( 
.A(n_10814),
.Y(n_11335)
);

INVx1_ASAP7_75t_L g11336 ( 
.A(n_10548),
.Y(n_11336)
);

NAND2xp5_ASAP7_75t_L g11337 ( 
.A(n_10902),
.B(n_1118),
.Y(n_11337)
);

BUFx6f_ASAP7_75t_L g11338 ( 
.A(n_10958),
.Y(n_11338)
);

NAND2xp5_ASAP7_75t_L g11339 ( 
.A(n_10906),
.B(n_1118),
.Y(n_11339)
);

OAI21x1_ASAP7_75t_L g11340 ( 
.A1(n_11127),
.A2(n_1119),
.B(n_1120),
.Y(n_11340)
);

INVxp67_ASAP7_75t_SL g11341 ( 
.A(n_10634),
.Y(n_11341)
);

INVxp67_ASAP7_75t_L g11342 ( 
.A(n_10937),
.Y(n_11342)
);

OAI21xp33_ASAP7_75t_L g11343 ( 
.A1(n_11248),
.A2(n_1120),
.B(n_1121),
.Y(n_11343)
);

BUFx2_ASAP7_75t_L g11344 ( 
.A(n_10898),
.Y(n_11344)
);

INVx1_ASAP7_75t_SL g11345 ( 
.A(n_10743),
.Y(n_11345)
);

BUFx6f_ASAP7_75t_L g11346 ( 
.A(n_10958),
.Y(n_11346)
);

BUFx2_ASAP7_75t_L g11347 ( 
.A(n_10539),
.Y(n_11347)
);

NAND2xp5_ASAP7_75t_SL g11348 ( 
.A(n_10567),
.B(n_1122),
.Y(n_11348)
);

AO31x2_ASAP7_75t_L g11349 ( 
.A1(n_10929),
.A2(n_1124),
.A3(n_1122),
.B(n_1123),
.Y(n_11349)
);

BUFx4_ASAP7_75t_SL g11350 ( 
.A(n_10719),
.Y(n_11350)
);

OAI21x1_ASAP7_75t_L g11351 ( 
.A1(n_10757),
.A2(n_1123),
.B(n_1124),
.Y(n_11351)
);

AOI21xp5_ASAP7_75t_L g11352 ( 
.A1(n_10806),
.A2(n_1125),
.B(n_1126),
.Y(n_11352)
);

AOI21xp5_ASAP7_75t_L g11353 ( 
.A1(n_10756),
.A2(n_1125),
.B(n_1126),
.Y(n_11353)
);

INVx1_ASAP7_75t_L g11354 ( 
.A(n_10587),
.Y(n_11354)
);

INVx1_ASAP7_75t_L g11355 ( 
.A(n_10588),
.Y(n_11355)
);

INVx1_ASAP7_75t_L g11356 ( 
.A(n_10611),
.Y(n_11356)
);

NAND2x1_ASAP7_75t_L g11357 ( 
.A(n_10766),
.B(n_1127),
.Y(n_11357)
);

INVx3_ASAP7_75t_L g11358 ( 
.A(n_10630),
.Y(n_11358)
);

OAI21x1_ASAP7_75t_L g11359 ( 
.A1(n_11054),
.A2(n_1127),
.B(n_1128),
.Y(n_11359)
);

OAI21x1_ASAP7_75t_L g11360 ( 
.A1(n_11227),
.A2(n_1128),
.B(n_1129),
.Y(n_11360)
);

OA22x2_ASAP7_75t_L g11361 ( 
.A1(n_11236),
.A2(n_1131),
.B1(n_1129),
.B2(n_1130),
.Y(n_11361)
);

AO31x2_ASAP7_75t_L g11362 ( 
.A1(n_10752),
.A2(n_10996),
.A3(n_10980),
.B(n_10783),
.Y(n_11362)
);

AOI21xp5_ASAP7_75t_L g11363 ( 
.A1(n_10685),
.A2(n_1130),
.B(n_1131),
.Y(n_11363)
);

AOI21xp5_ASAP7_75t_L g11364 ( 
.A1(n_10970),
.A2(n_1132),
.B(n_1133),
.Y(n_11364)
);

OAI21x1_ASAP7_75t_L g11365 ( 
.A1(n_11229),
.A2(n_1133),
.B(n_1134),
.Y(n_11365)
);

INVx3_ASAP7_75t_L g11366 ( 
.A(n_11051),
.Y(n_11366)
);

NAND2xp5_ASAP7_75t_L g11367 ( 
.A(n_10892),
.B(n_1134),
.Y(n_11367)
);

AOI22xp5_ASAP7_75t_L g11368 ( 
.A1(n_10865),
.A2(n_1137),
.B1(n_1135),
.B2(n_1136),
.Y(n_11368)
);

AND2x4_ASAP7_75t_L g11369 ( 
.A(n_11260),
.B(n_1135),
.Y(n_11369)
);

OAI21xp5_ASAP7_75t_L g11370 ( 
.A1(n_11235),
.A2(n_1136),
.B(n_1137),
.Y(n_11370)
);

OAI21x1_ASAP7_75t_L g11371 ( 
.A1(n_11253),
.A2(n_1139),
.B(n_1140),
.Y(n_11371)
);

AOI21xp5_ASAP7_75t_L g11372 ( 
.A1(n_11228),
.A2(n_1139),
.B(n_1140),
.Y(n_11372)
);

NAND2x1p5_ASAP7_75t_L g11373 ( 
.A(n_10868),
.B(n_1141),
.Y(n_11373)
);

NAND2xp5_ASAP7_75t_L g11374 ( 
.A(n_10933),
.B(n_1141),
.Y(n_11374)
);

OAI21xp5_ASAP7_75t_L g11375 ( 
.A1(n_10763),
.A2(n_1142),
.B(n_1143),
.Y(n_11375)
);

NAND2x1p5_ASAP7_75t_L g11376 ( 
.A(n_10868),
.B(n_1142),
.Y(n_11376)
);

AOI21xp5_ASAP7_75t_L g11377 ( 
.A1(n_11244),
.A2(n_1143),
.B(n_1144),
.Y(n_11377)
);

AOI21xp5_ASAP7_75t_L g11378 ( 
.A1(n_10754),
.A2(n_1145),
.B(n_1146),
.Y(n_11378)
);

OAI21x1_ASAP7_75t_L g11379 ( 
.A1(n_10936),
.A2(n_1146),
.B(n_1147),
.Y(n_11379)
);

INVx2_ASAP7_75t_L g11380 ( 
.A(n_10625),
.Y(n_11380)
);

NAND2xp5_ASAP7_75t_L g11381 ( 
.A(n_10938),
.B(n_10951),
.Y(n_11381)
);

AO31x2_ASAP7_75t_L g11382 ( 
.A1(n_10923),
.A2(n_1150),
.A3(n_1148),
.B(n_1149),
.Y(n_11382)
);

AOI21xp5_ASAP7_75t_L g11383 ( 
.A1(n_11114),
.A2(n_1148),
.B(n_1149),
.Y(n_11383)
);

BUFx2_ASAP7_75t_L g11384 ( 
.A(n_10667),
.Y(n_11384)
);

NAND2xp5_ASAP7_75t_SL g11385 ( 
.A(n_11187),
.B(n_1150),
.Y(n_11385)
);

NAND2xp5_ASAP7_75t_SL g11386 ( 
.A(n_11187),
.B(n_1152),
.Y(n_11386)
);

OAI21x1_ASAP7_75t_L g11387 ( 
.A1(n_10574),
.A2(n_1152),
.B(n_1153),
.Y(n_11387)
);

AOI21xp5_ASAP7_75t_L g11388 ( 
.A1(n_11057),
.A2(n_1153),
.B(n_1154),
.Y(n_11388)
);

OAI21x1_ASAP7_75t_L g11389 ( 
.A1(n_10871),
.A2(n_1154),
.B(n_1155),
.Y(n_11389)
);

AO22x2_ASAP7_75t_L g11390 ( 
.A1(n_10965),
.A2(n_1157),
.B1(n_1155),
.B2(n_1156),
.Y(n_11390)
);

NAND2xp5_ASAP7_75t_L g11391 ( 
.A(n_10913),
.B(n_1156),
.Y(n_11391)
);

BUFx6f_ASAP7_75t_L g11392 ( 
.A(n_11052),
.Y(n_11392)
);

OR2x2_ASAP7_75t_L g11393 ( 
.A(n_10815),
.B(n_1158),
.Y(n_11393)
);

AOI21xp5_ASAP7_75t_L g11394 ( 
.A1(n_10921),
.A2(n_1159),
.B(n_1160),
.Y(n_11394)
);

AND2x2_ASAP7_75t_L g11395 ( 
.A(n_10662),
.B(n_1159),
.Y(n_11395)
);

OAI21x1_ASAP7_75t_L g11396 ( 
.A1(n_10684),
.A2(n_1160),
.B(n_1161),
.Y(n_11396)
);

OAI21x1_ASAP7_75t_L g11397 ( 
.A1(n_10972),
.A2(n_1161),
.B(n_1162),
.Y(n_11397)
);

NAND2xp5_ASAP7_75t_SL g11398 ( 
.A(n_10640),
.B(n_1162),
.Y(n_11398)
);

AOI21x1_ASAP7_75t_L g11399 ( 
.A1(n_10941),
.A2(n_1163),
.B(n_1164),
.Y(n_11399)
);

OAI21xp5_ASAP7_75t_L g11400 ( 
.A1(n_10798),
.A2(n_1163),
.B(n_1164),
.Y(n_11400)
);

AOI21xp5_ASAP7_75t_L g11401 ( 
.A1(n_10727),
.A2(n_1165),
.B(n_1166),
.Y(n_11401)
);

AND2x2_ASAP7_75t_L g11402 ( 
.A(n_11138),
.B(n_1165),
.Y(n_11402)
);

INVx1_ASAP7_75t_L g11403 ( 
.A(n_10623),
.Y(n_11403)
);

AO31x2_ASAP7_75t_L g11404 ( 
.A1(n_10940),
.A2(n_1169),
.A3(n_1167),
.B(n_1168),
.Y(n_11404)
);

INVx1_ASAP7_75t_L g11405 ( 
.A(n_10686),
.Y(n_11405)
);

AND2x2_ASAP7_75t_L g11406 ( 
.A(n_10768),
.B(n_1168),
.Y(n_11406)
);

OAI21x1_ASAP7_75t_L g11407 ( 
.A1(n_10811),
.A2(n_1169),
.B(n_1170),
.Y(n_11407)
);

OAI21x1_ASAP7_75t_L g11408 ( 
.A1(n_10605),
.A2(n_10679),
.B(n_10551),
.Y(n_11408)
);

NAND2xp5_ASAP7_75t_L g11409 ( 
.A(n_10914),
.B(n_1170),
.Y(n_11409)
);

AND2x4_ASAP7_75t_L g11410 ( 
.A(n_10554),
.B(n_1171),
.Y(n_11410)
);

AOI21xp5_ASAP7_75t_L g11411 ( 
.A1(n_11085),
.A2(n_1171),
.B(n_1172),
.Y(n_11411)
);

AOI21xp5_ASAP7_75t_L g11412 ( 
.A1(n_10628),
.A2(n_1172),
.B(n_1173),
.Y(n_11412)
);

NAND2xp5_ASAP7_75t_L g11413 ( 
.A(n_10924),
.B(n_1174),
.Y(n_11413)
);

NAND2xp5_ASAP7_75t_L g11414 ( 
.A(n_10956),
.B(n_1175),
.Y(n_11414)
);

INVx2_ASAP7_75t_L g11415 ( 
.A(n_10642),
.Y(n_11415)
);

AOI21xp5_ASAP7_75t_L g11416 ( 
.A1(n_10977),
.A2(n_1175),
.B(n_1176),
.Y(n_11416)
);

OAI21x1_ASAP7_75t_L g11417 ( 
.A1(n_10650),
.A2(n_10656),
.B(n_10652),
.Y(n_11417)
);

NAND2x1_ASAP7_75t_L g11418 ( 
.A(n_10767),
.B(n_1176),
.Y(n_11418)
);

AO31x2_ASAP7_75t_L g11419 ( 
.A1(n_10950),
.A2(n_1179),
.A3(n_1177),
.B(n_1178),
.Y(n_11419)
);

AOI21xp5_ASAP7_75t_L g11420 ( 
.A1(n_11226),
.A2(n_1177),
.B(n_1178),
.Y(n_11420)
);

NAND2xp5_ASAP7_75t_L g11421 ( 
.A(n_10821),
.B(n_1179),
.Y(n_11421)
);

BUFx6f_ASAP7_75t_L g11422 ( 
.A(n_11056),
.Y(n_11422)
);

HB1xp67_ASAP7_75t_L g11423 ( 
.A(n_10653),
.Y(n_11423)
);

INVx3_ASAP7_75t_L g11424 ( 
.A(n_11050),
.Y(n_11424)
);

AOI21xp5_ASAP7_75t_L g11425 ( 
.A1(n_11147),
.A2(n_1180),
.B(n_1181),
.Y(n_11425)
);

OAI22xp5_ASAP7_75t_L g11426 ( 
.A1(n_10987),
.A2(n_1182),
.B1(n_1180),
.B2(n_1181),
.Y(n_11426)
);

NAND2xp5_ASAP7_75t_L g11427 ( 
.A(n_10841),
.B(n_1183),
.Y(n_11427)
);

NOR2x1_ASAP7_75t_SL g11428 ( 
.A(n_10661),
.B(n_1183),
.Y(n_11428)
);

OAI22xp5_ASAP7_75t_L g11429 ( 
.A1(n_11004),
.A2(n_1186),
.B1(n_1184),
.B2(n_1185),
.Y(n_11429)
);

AND2x2_ASAP7_75t_L g11430 ( 
.A(n_11186),
.B(n_1184),
.Y(n_11430)
);

INVx2_ASAP7_75t_L g11431 ( 
.A(n_10666),
.Y(n_11431)
);

NAND2xp5_ASAP7_75t_L g11432 ( 
.A(n_10851),
.B(n_1185),
.Y(n_11432)
);

OAI21x1_ASAP7_75t_L g11433 ( 
.A1(n_10673),
.A2(n_10674),
.B(n_10787),
.Y(n_11433)
);

NAND2xp5_ASAP7_75t_L g11434 ( 
.A(n_10859),
.B(n_1187),
.Y(n_11434)
);

INVx1_ASAP7_75t_L g11435 ( 
.A(n_10688),
.Y(n_11435)
);

OAI22xp5_ASAP7_75t_L g11436 ( 
.A1(n_10796),
.A2(n_1190),
.B1(n_1188),
.B2(n_1189),
.Y(n_11436)
);

AND2x2_ASAP7_75t_L g11437 ( 
.A(n_11186),
.B(n_1188),
.Y(n_11437)
);

NAND2xp5_ASAP7_75t_L g11438 ( 
.A(n_10863),
.B(n_1190),
.Y(n_11438)
);

A2O1A1Ixp33_ASAP7_75t_L g11439 ( 
.A1(n_10675),
.A2(n_1193),
.B(n_1191),
.C(n_1192),
.Y(n_11439)
);

OAI21x1_ASAP7_75t_L g11440 ( 
.A1(n_10795),
.A2(n_1191),
.B(n_1192),
.Y(n_11440)
);

INVxp67_ASAP7_75t_L g11441 ( 
.A(n_11103),
.Y(n_11441)
);

OAI21x1_ASAP7_75t_L g11442 ( 
.A1(n_10803),
.A2(n_1193),
.B(n_1194),
.Y(n_11442)
);

NOR2x1_ASAP7_75t_L g11443 ( 
.A(n_11160),
.B(n_1194),
.Y(n_11443)
);

INVx2_ASAP7_75t_L g11444 ( 
.A(n_10681),
.Y(n_11444)
);

BUFx10_ASAP7_75t_L g11445 ( 
.A(n_10695),
.Y(n_11445)
);

NAND2xp5_ASAP7_75t_L g11446 ( 
.A(n_10873),
.B(n_1195),
.Y(n_11446)
);

AOI21xp5_ASAP7_75t_L g11447 ( 
.A1(n_11196),
.A2(n_1195),
.B(n_1196),
.Y(n_11447)
);

NOR2xp67_ASAP7_75t_SL g11448 ( 
.A(n_10746),
.B(n_10591),
.Y(n_11448)
);

INVx2_ASAP7_75t_L g11449 ( 
.A(n_10682),
.Y(n_11449)
);

OAI21x1_ASAP7_75t_L g11450 ( 
.A1(n_10812),
.A2(n_1196),
.B(n_1197),
.Y(n_11450)
);

INVx1_ASAP7_75t_L g11451 ( 
.A(n_10690),
.Y(n_11451)
);

INVxp67_ASAP7_75t_L g11452 ( 
.A(n_11105),
.Y(n_11452)
);

OAI22xp5_ASAP7_75t_L g11453 ( 
.A1(n_10822),
.A2(n_1199),
.B1(n_1197),
.B2(n_1198),
.Y(n_11453)
);

AOI21xp5_ASAP7_75t_L g11454 ( 
.A1(n_11144),
.A2(n_1198),
.B(n_1200),
.Y(n_11454)
);

CKINVDCx5p33_ASAP7_75t_R g11455 ( 
.A(n_10601),
.Y(n_11455)
);

OAI21x1_ASAP7_75t_L g11456 ( 
.A1(n_10843),
.A2(n_1200),
.B(n_1201),
.Y(n_11456)
);

OAI21xp33_ASAP7_75t_L g11457 ( 
.A1(n_11030),
.A2(n_1201),
.B(n_1202),
.Y(n_11457)
);

NAND2xp5_ASAP7_75t_L g11458 ( 
.A(n_10696),
.B(n_1202),
.Y(n_11458)
);

AOI21xp5_ASAP7_75t_L g11459 ( 
.A1(n_10556),
.A2(n_1203),
.B(n_1204),
.Y(n_11459)
);

INVx1_ASAP7_75t_L g11460 ( 
.A(n_10698),
.Y(n_11460)
);

A2O1A1Ixp33_ASAP7_75t_L g11461 ( 
.A1(n_10552),
.A2(n_1206),
.B(n_1204),
.C(n_1205),
.Y(n_11461)
);

OAI21x1_ASAP7_75t_SL g11462 ( 
.A1(n_10741),
.A2(n_1205),
.B(n_1206),
.Y(n_11462)
);

INVx3_ASAP7_75t_L g11463 ( 
.A(n_11050),
.Y(n_11463)
);

BUFx2_ASAP7_75t_L g11464 ( 
.A(n_10949),
.Y(n_11464)
);

OAI21x1_ASAP7_75t_L g11465 ( 
.A1(n_10846),
.A2(n_1207),
.B(n_1208),
.Y(n_11465)
);

AOI21xp5_ASAP7_75t_L g11466 ( 
.A1(n_10576),
.A2(n_1208),
.B(n_1209),
.Y(n_11466)
);

AOI211x1_ASAP7_75t_L g11467 ( 
.A1(n_10895),
.A2(n_1211),
.B(n_1209),
.C(n_1210),
.Y(n_11467)
);

NAND3xp33_ASAP7_75t_L g11468 ( 
.A(n_10724),
.B(n_1210),
.C(n_1211),
.Y(n_11468)
);

OAI21x1_ASAP7_75t_L g11469 ( 
.A1(n_10858),
.A2(n_1212),
.B(n_1213),
.Y(n_11469)
);

A2O1A1Ixp33_ASAP7_75t_L g11470 ( 
.A1(n_10621),
.A2(n_10669),
.B(n_10633),
.C(n_10769),
.Y(n_11470)
);

INVx2_ASAP7_75t_L g11471 ( 
.A(n_10722),
.Y(n_11471)
);

AOI221x1_ASAP7_75t_L g11472 ( 
.A1(n_11035),
.A2(n_1215),
.B1(n_1213),
.B2(n_1214),
.C(n_1216),
.Y(n_11472)
);

INVx1_ASAP7_75t_L g11473 ( 
.A(n_10712),
.Y(n_11473)
);

NAND2xp5_ASAP7_75t_L g11474 ( 
.A(n_10729),
.B(n_1214),
.Y(n_11474)
);

NAND2xp5_ASAP7_75t_L g11475 ( 
.A(n_10731),
.B(n_1215),
.Y(n_11475)
);

BUFx6f_ASAP7_75t_L g11476 ( 
.A(n_11056),
.Y(n_11476)
);

INVxp67_ASAP7_75t_SL g11477 ( 
.A(n_10561),
.Y(n_11477)
);

OAI21x1_ASAP7_75t_L g11478 ( 
.A1(n_10872),
.A2(n_1216),
.B(n_1217),
.Y(n_11478)
);

NAND2xp5_ASAP7_75t_SL g11479 ( 
.A(n_11010),
.B(n_1218),
.Y(n_11479)
);

NAND2xp5_ASAP7_75t_L g11480 ( 
.A(n_10733),
.B(n_10744),
.Y(n_11480)
);

OAI21x1_ASAP7_75t_L g11481 ( 
.A1(n_10878),
.A2(n_1218),
.B(n_1219),
.Y(n_11481)
);

OA21x2_ASAP7_75t_L g11482 ( 
.A1(n_10835),
.A2(n_1219),
.B(n_1220),
.Y(n_11482)
);

AND2x4_ASAP7_75t_L g11483 ( 
.A(n_11231),
.B(n_10747),
.Y(n_11483)
);

NAND2x1_ASAP7_75t_L g11484 ( 
.A(n_10786),
.B(n_1220),
.Y(n_11484)
);

NAND2xp5_ASAP7_75t_SL g11485 ( 
.A(n_10975),
.B(n_1221),
.Y(n_11485)
);

AND2x2_ASAP7_75t_L g11486 ( 
.A(n_10749),
.B(n_1221),
.Y(n_11486)
);

AOI21xp5_ASAP7_75t_L g11487 ( 
.A1(n_10609),
.A2(n_1222),
.B(n_1223),
.Y(n_11487)
);

INVx3_ASAP7_75t_L g11488 ( 
.A(n_10901),
.Y(n_11488)
);

INVx1_ASAP7_75t_SL g11489 ( 
.A(n_11250),
.Y(n_11489)
);

AOI22xp33_ASAP7_75t_L g11490 ( 
.A1(n_11053),
.A2(n_1225),
.B1(n_1222),
.B2(n_1224),
.Y(n_11490)
);

AND2x2_ASAP7_75t_L g11491 ( 
.A(n_10755),
.B(n_1224),
.Y(n_11491)
);

OAI22xp5_ASAP7_75t_L g11492 ( 
.A1(n_10891),
.A2(n_1228),
.B1(n_1225),
.B2(n_1226),
.Y(n_11492)
);

AOI21xp5_ASAP7_75t_L g11493 ( 
.A1(n_11059),
.A2(n_1226),
.B(n_1228),
.Y(n_11493)
);

AOI21xp5_ASAP7_75t_SL g11494 ( 
.A1(n_10547),
.A2(n_1229),
.B(n_1230),
.Y(n_11494)
);

INVx1_ASAP7_75t_L g11495 ( 
.A(n_10718),
.Y(n_11495)
);

AO31x2_ASAP7_75t_L g11496 ( 
.A1(n_10802),
.A2(n_1231),
.A3(n_1229),
.B(n_1230),
.Y(n_11496)
);

INVx2_ASAP7_75t_L g11497 ( 
.A(n_10758),
.Y(n_11497)
);

A2O1A1Ixp33_ASAP7_75t_L g11498 ( 
.A1(n_10998),
.A2(n_11009),
.B(n_10880),
.C(n_10907),
.Y(n_11498)
);

NAND2xp5_ASAP7_75t_L g11499 ( 
.A(n_10761),
.B(n_1231),
.Y(n_11499)
);

AO31x2_ASAP7_75t_L g11500 ( 
.A1(n_10807),
.A2(n_1234),
.A3(n_1232),
.B(n_1233),
.Y(n_11500)
);

NOR2xp33_ASAP7_75t_L g11501 ( 
.A(n_10986),
.B(n_1232),
.Y(n_11501)
);

BUFx3_ASAP7_75t_L g11502 ( 
.A(n_10909),
.Y(n_11502)
);

OAI21xp5_ASAP7_75t_L g11503 ( 
.A1(n_10882),
.A2(n_1233),
.B(n_1235),
.Y(n_11503)
);

INVx1_ASAP7_75t_L g11504 ( 
.A(n_10748),
.Y(n_11504)
);

AO31x2_ASAP7_75t_L g11505 ( 
.A1(n_10850),
.A2(n_1237),
.A3(n_1235),
.B(n_1236),
.Y(n_11505)
);

HB1xp67_ASAP7_75t_L g11506 ( 
.A(n_10764),
.Y(n_11506)
);

OAI21x1_ASAP7_75t_L g11507 ( 
.A1(n_10884),
.A2(n_1236),
.B(n_1237),
.Y(n_11507)
);

AOI21xp5_ASAP7_75t_L g11508 ( 
.A1(n_11076),
.A2(n_1238),
.B(n_1240),
.Y(n_11508)
);

AND2x2_ASAP7_75t_L g11509 ( 
.A(n_11252),
.B(n_1238),
.Y(n_11509)
);

AOI21x1_ASAP7_75t_L g11510 ( 
.A1(n_10713),
.A2(n_1240),
.B(n_1241),
.Y(n_11510)
);

OAI21x1_ASAP7_75t_SL g11511 ( 
.A1(n_11020),
.A2(n_1241),
.B(n_1242),
.Y(n_11511)
);

AO21x1_ASAP7_75t_L g11512 ( 
.A1(n_11042),
.A2(n_10853),
.B(n_10974),
.Y(n_11512)
);

INVx2_ASAP7_75t_L g11513 ( 
.A(n_10765),
.Y(n_11513)
);

BUFx2_ASAP7_75t_L g11514 ( 
.A(n_10725),
.Y(n_11514)
);

OAI21x1_ASAP7_75t_L g11515 ( 
.A1(n_10889),
.A2(n_10896),
.B(n_10894),
.Y(n_11515)
);

AND2x2_ASAP7_75t_L g11516 ( 
.A(n_11259),
.B(n_1242),
.Y(n_11516)
);

AO31x2_ASAP7_75t_L g11517 ( 
.A1(n_10879),
.A2(n_1245),
.A3(n_1243),
.B(n_1244),
.Y(n_11517)
);

OAI21xp5_ASAP7_75t_L g11518 ( 
.A1(n_10899),
.A2(n_10920),
.B(n_10904),
.Y(n_11518)
);

NAND2xp5_ASAP7_75t_L g11519 ( 
.A(n_11028),
.B(n_1243),
.Y(n_11519)
);

AOI22xp5_ASAP7_75t_L g11520 ( 
.A1(n_11217),
.A2(n_1247),
.B1(n_1244),
.B2(n_1246),
.Y(n_11520)
);

AOI21xp5_ASAP7_75t_L g11521 ( 
.A1(n_10852),
.A2(n_1246),
.B(n_1247),
.Y(n_11521)
);

OA21x2_ASAP7_75t_L g11522 ( 
.A1(n_10990),
.A2(n_1248),
.B(n_1249),
.Y(n_11522)
);

OAI21x1_ASAP7_75t_L g11523 ( 
.A1(n_10947),
.A2(n_1248),
.B(n_1249),
.Y(n_11523)
);

A2O1A1Ixp33_ASAP7_75t_L g11524 ( 
.A1(n_10911),
.A2(n_1252),
.B(n_1250),
.C(n_1251),
.Y(n_11524)
);

AOI21x1_ASAP7_75t_L g11525 ( 
.A1(n_10626),
.A2(n_1250),
.B(n_1251),
.Y(n_11525)
);

OAI21x1_ASAP7_75t_L g11526 ( 
.A1(n_10953),
.A2(n_1252),
.B(n_1253),
.Y(n_11526)
);

NAND2xp5_ASAP7_75t_L g11527 ( 
.A(n_11031),
.B(n_1253),
.Y(n_11527)
);

INVx8_ASAP7_75t_L g11528 ( 
.A(n_10948),
.Y(n_11528)
);

OAI21xp5_ASAP7_75t_L g11529 ( 
.A1(n_10959),
.A2(n_1254),
.B(n_1255),
.Y(n_11529)
);

AND2x2_ASAP7_75t_L g11530 ( 
.A(n_11079),
.B(n_1255),
.Y(n_11530)
);

NAND2xp33_ASAP7_75t_L g11531 ( 
.A(n_11023),
.B(n_1256),
.Y(n_11531)
);

INVx1_ASAP7_75t_L g11532 ( 
.A(n_10789),
.Y(n_11532)
);

BUFx6f_ASAP7_75t_L g11533 ( 
.A(n_10901),
.Y(n_11533)
);

NAND2xp5_ASAP7_75t_L g11534 ( 
.A(n_11036),
.B(n_1256),
.Y(n_11534)
);

BUFx6f_ASAP7_75t_L g11535 ( 
.A(n_11049),
.Y(n_11535)
);

NOR2xp33_ASAP7_75t_SL g11536 ( 
.A(n_10631),
.B(n_10837),
.Y(n_11536)
);

NAND2xp5_ASAP7_75t_L g11537 ( 
.A(n_10854),
.B(n_1257),
.Y(n_11537)
);

AOI21xp33_ASAP7_75t_L g11538 ( 
.A1(n_11213),
.A2(n_1257),
.B(n_1258),
.Y(n_11538)
);

NAND2xp5_ASAP7_75t_L g11539 ( 
.A(n_10943),
.B(n_1258),
.Y(n_11539)
);

OAI21xp5_ASAP7_75t_L g11540 ( 
.A1(n_11002),
.A2(n_1259),
.B(n_1260),
.Y(n_11540)
);

INVx4_ASAP7_75t_L g11541 ( 
.A(n_11024),
.Y(n_11541)
);

AOI21xp5_ASAP7_75t_L g11542 ( 
.A1(n_10935),
.A2(n_1259),
.B(n_1260),
.Y(n_11542)
);

OAI21x1_ASAP7_75t_L g11543 ( 
.A1(n_11007),
.A2(n_1261),
.B(n_1262),
.Y(n_11543)
);

NAND2xp5_ASAP7_75t_L g11544 ( 
.A(n_10808),
.B(n_1261),
.Y(n_11544)
);

NAND2xp5_ASAP7_75t_L g11545 ( 
.A(n_11148),
.B(n_1263),
.Y(n_11545)
);

NAND2xp5_ASAP7_75t_L g11546 ( 
.A(n_11164),
.B(n_1263),
.Y(n_11546)
);

NAND2xp5_ASAP7_75t_L g11547 ( 
.A(n_11165),
.B(n_10978),
.Y(n_11547)
);

OAI22x1_ASAP7_75t_L g11548 ( 
.A1(n_11152),
.A2(n_11178),
.B1(n_10706),
.B2(n_11088),
.Y(n_11548)
);

INVx1_ASAP7_75t_L g11549 ( 
.A(n_10543),
.Y(n_11549)
);

OAI21x1_ASAP7_75t_L g11550 ( 
.A1(n_11012),
.A2(n_1264),
.B(n_1265),
.Y(n_11550)
);

OAI22xp5_ASAP7_75t_L g11551 ( 
.A1(n_10569),
.A2(n_1266),
.B1(n_1264),
.B2(n_1265),
.Y(n_11551)
);

AOI21x1_ASAP7_75t_L g11552 ( 
.A1(n_10651),
.A2(n_1267),
.B(n_1268),
.Y(n_11552)
);

AOI22xp5_ASAP7_75t_L g11553 ( 
.A1(n_10957),
.A2(n_1269),
.B1(n_1267),
.B2(n_1268),
.Y(n_11553)
);

OAI21x1_ASAP7_75t_L g11554 ( 
.A1(n_11033),
.A2(n_1269),
.B(n_1270),
.Y(n_11554)
);

O2A1O1Ixp5_ASAP7_75t_L g11555 ( 
.A1(n_10645),
.A2(n_1272),
.B(n_1270),
.C(n_1271),
.Y(n_11555)
);

NAND2xp5_ASAP7_75t_L g11556 ( 
.A(n_11156),
.B(n_1271),
.Y(n_11556)
);

BUFx6f_ASAP7_75t_L g11557 ( 
.A(n_11049),
.Y(n_11557)
);

INVx1_ASAP7_75t_L g11558 ( 
.A(n_11239),
.Y(n_11558)
);

OAI21xp5_ASAP7_75t_L g11559 ( 
.A1(n_11202),
.A2(n_1273),
.B(n_1274),
.Y(n_11559)
);

INVx4_ASAP7_75t_L g11560 ( 
.A(n_11055),
.Y(n_11560)
);

OAI22xp5_ASAP7_75t_L g11561 ( 
.A1(n_10583),
.A2(n_1275),
.B1(n_1273),
.B2(n_1274),
.Y(n_11561)
);

NAND2xp5_ASAP7_75t_SL g11562 ( 
.A(n_11212),
.B(n_1277),
.Y(n_11562)
);

NAND2xp5_ASAP7_75t_L g11563 ( 
.A(n_11155),
.B(n_1277),
.Y(n_11563)
);

NAND2xp5_ASAP7_75t_L g11564 ( 
.A(n_10716),
.B(n_1278),
.Y(n_11564)
);

AOI21xp5_ASAP7_75t_L g11565 ( 
.A1(n_11188),
.A2(n_1278),
.B(n_1279),
.Y(n_11565)
);

OAI21x1_ASAP7_75t_L g11566 ( 
.A1(n_11203),
.A2(n_1279),
.B(n_1280),
.Y(n_11566)
);

OA21x2_ASAP7_75t_L g11567 ( 
.A1(n_10845),
.A2(n_1281),
.B(n_1282),
.Y(n_11567)
);

A2O1A1Ixp33_ASAP7_75t_L g11568 ( 
.A1(n_11102),
.A2(n_1283),
.B(n_1281),
.C(n_1282),
.Y(n_11568)
);

AOI21x1_ASAP7_75t_L g11569 ( 
.A1(n_10657),
.A2(n_1283),
.B(n_1284),
.Y(n_11569)
);

AOI21xp5_ASAP7_75t_L g11570 ( 
.A1(n_10856),
.A2(n_11000),
.B(n_11145),
.Y(n_11570)
);

NAND2xp5_ASAP7_75t_L g11571 ( 
.A(n_11245),
.B(n_1284),
.Y(n_11571)
);

NAND2xp5_ASAP7_75t_L g11572 ( 
.A(n_11246),
.B(n_1285),
.Y(n_11572)
);

OAI22x1_ASAP7_75t_L g11573 ( 
.A1(n_10855),
.A2(n_1287),
.B1(n_1285),
.B2(n_1286),
.Y(n_11573)
);

OAI21x1_ASAP7_75t_L g11574 ( 
.A1(n_11211),
.A2(n_11151),
.B(n_11139),
.Y(n_11574)
);

A2O1A1Ixp33_ASAP7_75t_L g11575 ( 
.A1(n_11108),
.A2(n_1288),
.B(n_1286),
.C(n_1287),
.Y(n_11575)
);

AOI22xp33_ASAP7_75t_L g11576 ( 
.A1(n_10784),
.A2(n_1291),
.B1(n_1289),
.B2(n_1290),
.Y(n_11576)
);

OAI21x1_ASAP7_75t_L g11577 ( 
.A1(n_11153),
.A2(n_1289),
.B(n_1291),
.Y(n_11577)
);

INVxp67_ASAP7_75t_SL g11578 ( 
.A(n_10593),
.Y(n_11578)
);

INVx1_ASAP7_75t_L g11579 ( 
.A(n_11249),
.Y(n_11579)
);

INVx3_ASAP7_75t_L g11580 ( 
.A(n_10916),
.Y(n_11580)
);

AOI21xp5_ASAP7_75t_L g11581 ( 
.A1(n_11157),
.A2(n_1292),
.B(n_1293),
.Y(n_11581)
);

NAND2x1p5_ASAP7_75t_L g11582 ( 
.A(n_10868),
.B(n_1293),
.Y(n_11582)
);

NAND2xp5_ASAP7_75t_L g11583 ( 
.A(n_11262),
.B(n_1294),
.Y(n_11583)
);

CKINVDCx5p33_ASAP7_75t_R g11584 ( 
.A(n_10602),
.Y(n_11584)
);

AOI21xp5_ASAP7_75t_L g11585 ( 
.A1(n_10774),
.A2(n_1294),
.B(n_1295),
.Y(n_11585)
);

AO31x2_ASAP7_75t_L g11586 ( 
.A1(n_10655),
.A2(n_1297),
.A3(n_1295),
.B(n_1296),
.Y(n_11586)
);

OAI21xp5_ASAP7_75t_L g11587 ( 
.A1(n_11037),
.A2(n_11074),
.B(n_11071),
.Y(n_11587)
);

AOI21xp5_ASAP7_75t_L g11588 ( 
.A1(n_10691),
.A2(n_1296),
.B(n_1297),
.Y(n_11588)
);

NAND2xp5_ASAP7_75t_L g11589 ( 
.A(n_10557),
.B(n_1298),
.Y(n_11589)
);

INVx1_ASAP7_75t_L g11590 ( 
.A(n_10643),
.Y(n_11590)
);

OAI21x1_ASAP7_75t_L g11591 ( 
.A1(n_11171),
.A2(n_1298),
.B(n_1299),
.Y(n_11591)
);

NAND2xp5_ASAP7_75t_L g11592 ( 
.A(n_10598),
.B(n_1299),
.Y(n_11592)
);

NAND2xp5_ASAP7_75t_L g11593 ( 
.A(n_10607),
.B(n_1300),
.Y(n_11593)
);

AOI21xp5_ASAP7_75t_SL g11594 ( 
.A1(n_10585),
.A2(n_1300),
.B(n_1302),
.Y(n_11594)
);

OAI21x1_ASAP7_75t_L g11595 ( 
.A1(n_11174),
.A2(n_1302),
.B(n_1303),
.Y(n_11595)
);

OAI21xp33_ASAP7_75t_L g11596 ( 
.A1(n_11080),
.A2(n_1303),
.B(n_1304),
.Y(n_11596)
);

AOI21xp5_ASAP7_75t_L g11597 ( 
.A1(n_11122),
.A2(n_1304),
.B(n_1305),
.Y(n_11597)
);

NAND2xp5_ASAP7_75t_L g11598 ( 
.A(n_10564),
.B(n_1306),
.Y(n_11598)
);

OAI21x1_ASAP7_75t_L g11599 ( 
.A1(n_11218),
.A2(n_1306),
.B(n_1307),
.Y(n_11599)
);

INVx1_ASAP7_75t_L g11600 ( 
.A(n_10705),
.Y(n_11600)
);

OAI21xp5_ASAP7_75t_L g11601 ( 
.A1(n_11086),
.A2(n_1308),
.B(n_1310),
.Y(n_11601)
);

NAND2xp5_ASAP7_75t_SL g11602 ( 
.A(n_10984),
.B(n_11140),
.Y(n_11602)
);

OAI21x1_ASAP7_75t_L g11603 ( 
.A1(n_11192),
.A2(n_1308),
.B(n_1311),
.Y(n_11603)
);

NAND2x1_ASAP7_75t_L g11604 ( 
.A(n_10820),
.B(n_1311),
.Y(n_11604)
);

AOI21xp5_ASAP7_75t_L g11605 ( 
.A1(n_10994),
.A2(n_1312),
.B(n_1314),
.Y(n_11605)
);

NAND2xp5_ASAP7_75t_L g11606 ( 
.A(n_10550),
.B(n_1312),
.Y(n_11606)
);

NAND2xp5_ASAP7_75t_L g11607 ( 
.A(n_10586),
.B(n_10562),
.Y(n_11607)
);

NAND2xp5_ASAP7_75t_L g11608 ( 
.A(n_11180),
.B(n_1314),
.Y(n_11608)
);

INVx1_ASAP7_75t_L g11609 ( 
.A(n_10714),
.Y(n_11609)
);

AO31x2_ASAP7_75t_L g11610 ( 
.A1(n_10993),
.A2(n_1317),
.A3(n_1315),
.B(n_1316),
.Y(n_11610)
);

OAI21x1_ASAP7_75t_L g11611 ( 
.A1(n_11193),
.A2(n_1315),
.B(n_1316),
.Y(n_11611)
);

OAI21x1_ASAP7_75t_L g11612 ( 
.A1(n_11194),
.A2(n_1317),
.B(n_1318),
.Y(n_11612)
);

INVx1_ASAP7_75t_L g11613 ( 
.A(n_10659),
.Y(n_11613)
);

NAND2xp5_ASAP7_75t_L g11614 ( 
.A(n_11183),
.B(n_1318),
.Y(n_11614)
);

OAI21x1_ASAP7_75t_L g11615 ( 
.A1(n_11199),
.A2(n_1319),
.B(n_1320),
.Y(n_11615)
);

OAI21xp5_ASAP7_75t_L g11616 ( 
.A1(n_11090),
.A2(n_1319),
.B(n_1320),
.Y(n_11616)
);

OAI22x1_ASAP7_75t_L g11617 ( 
.A1(n_10860),
.A2(n_1323),
.B1(n_1321),
.B2(n_1322),
.Y(n_11617)
);

INVx3_ASAP7_75t_L g11618 ( 
.A(n_11040),
.Y(n_11618)
);

OAI21x1_ASAP7_75t_L g11619 ( 
.A1(n_11092),
.A2(n_1321),
.B(n_1324),
.Y(n_11619)
);

INVx2_ASAP7_75t_L g11620 ( 
.A(n_10797),
.Y(n_11620)
);

OAI21x1_ASAP7_75t_L g11621 ( 
.A1(n_11097),
.A2(n_1325),
.B(n_1326),
.Y(n_11621)
);

OAI21x1_ASAP7_75t_L g11622 ( 
.A1(n_11099),
.A2(n_1325),
.B(n_1326),
.Y(n_11622)
);

OAI21x1_ASAP7_75t_SL g11623 ( 
.A1(n_10638),
.A2(n_1327),
.B(n_1328),
.Y(n_11623)
);

AND2x2_ASAP7_75t_L g11624 ( 
.A(n_11183),
.B(n_1327),
.Y(n_11624)
);

NAND2xp5_ASAP7_75t_L g11625 ( 
.A(n_10864),
.B(n_1328),
.Y(n_11625)
);

NAND3x1_ASAP7_75t_L g11626 ( 
.A(n_11131),
.B(n_1329),
.C(n_1330),
.Y(n_11626)
);

OAI21x1_ASAP7_75t_L g11627 ( 
.A1(n_11107),
.A2(n_1329),
.B(n_1330),
.Y(n_11627)
);

AOI21x1_ASAP7_75t_SL g11628 ( 
.A1(n_11119),
.A2(n_1331),
.B(n_1332),
.Y(n_11628)
);

NAND2xp5_ASAP7_75t_L g11629 ( 
.A(n_10934),
.B(n_1331),
.Y(n_11629)
);

HB1xp67_ASAP7_75t_L g11630 ( 
.A(n_10734),
.Y(n_11630)
);

AOI21xp5_ASAP7_75t_L g11631 ( 
.A1(n_10994),
.A2(n_1332),
.B(n_1333),
.Y(n_11631)
);

O2A1O1Ixp5_ASAP7_75t_L g11632 ( 
.A1(n_10870),
.A2(n_11241),
.B(n_10721),
.C(n_10579),
.Y(n_11632)
);

OAI21x1_ASAP7_75t_L g11633 ( 
.A1(n_11115),
.A2(n_1334),
.B(n_1335),
.Y(n_11633)
);

NAND2xp5_ASAP7_75t_L g11634 ( 
.A(n_10955),
.B(n_1334),
.Y(n_11634)
);

NAND2xp5_ASAP7_75t_L g11635 ( 
.A(n_10960),
.B(n_1336),
.Y(n_11635)
);

NOR2xp33_ASAP7_75t_L g11636 ( 
.A(n_10594),
.B(n_1336),
.Y(n_11636)
);

AOI21xp5_ASAP7_75t_L g11637 ( 
.A1(n_10603),
.A2(n_1337),
.B(n_1338),
.Y(n_11637)
);

AND2x2_ASAP7_75t_L g11638 ( 
.A(n_11109),
.B(n_1337),
.Y(n_11638)
);

AO31x2_ASAP7_75t_L g11639 ( 
.A1(n_10995),
.A2(n_1342),
.A3(n_1339),
.B(n_1340),
.Y(n_11639)
);

NAND2xp5_ASAP7_75t_L g11640 ( 
.A(n_10966),
.B(n_1339),
.Y(n_11640)
);

AO21x1_ASAP7_75t_L g11641 ( 
.A1(n_10720),
.A2(n_1342),
.B(n_1343),
.Y(n_11641)
);

INVx1_ASAP7_75t_L g11642 ( 
.A(n_10671),
.Y(n_11642)
);

OAI21xp5_ASAP7_75t_L g11643 ( 
.A1(n_11128),
.A2(n_1344),
.B(n_1345),
.Y(n_11643)
);

AND2x2_ASAP7_75t_L g11644 ( 
.A(n_10664),
.B(n_1344),
.Y(n_11644)
);

AO31x2_ASAP7_75t_L g11645 ( 
.A1(n_11006),
.A2(n_1348),
.A3(n_1346),
.B(n_1347),
.Y(n_11645)
);

NAND2xp5_ASAP7_75t_SL g11646 ( 
.A(n_10730),
.B(n_1347),
.Y(n_11646)
);

INVx1_ASAP7_75t_L g11647 ( 
.A(n_10678),
.Y(n_11647)
);

AO31x2_ASAP7_75t_L g11648 ( 
.A1(n_10604),
.A2(n_1351),
.A3(n_1349),
.B(n_1350),
.Y(n_11648)
);

INVx2_ASAP7_75t_L g11649 ( 
.A(n_10805),
.Y(n_11649)
);

OAI21x1_ASAP7_75t_L g11650 ( 
.A1(n_11135),
.A2(n_1349),
.B(n_1350),
.Y(n_11650)
);

NAND2xp5_ASAP7_75t_SL g11651 ( 
.A(n_11070),
.B(n_1351),
.Y(n_11651)
);

NAND2xp5_ASAP7_75t_L g11652 ( 
.A(n_10973),
.B(n_1352),
.Y(n_11652)
);

NAND2xp5_ASAP7_75t_L g11653 ( 
.A(n_10779),
.B(n_10961),
.Y(n_11653)
);

OA22x2_ASAP7_75t_L g11654 ( 
.A1(n_11011),
.A2(n_1354),
.B1(n_1352),
.B2(n_1353),
.Y(n_11654)
);

NAND2xp5_ASAP7_75t_L g11655 ( 
.A(n_10627),
.B(n_1353),
.Y(n_11655)
);

AOI21xp5_ASAP7_75t_L g11656 ( 
.A1(n_10610),
.A2(n_1354),
.B(n_1355),
.Y(n_11656)
);

NOR2x1_ASAP7_75t_L g11657 ( 
.A(n_10613),
.B(n_1355),
.Y(n_11657)
);

NAND2xp5_ASAP7_75t_L g11658 ( 
.A(n_11047),
.B(n_1357),
.Y(n_11658)
);

BUFx6f_ASAP7_75t_L g11659 ( 
.A(n_10776),
.Y(n_11659)
);

NAND2xp5_ASAP7_75t_L g11660 ( 
.A(n_10813),
.B(n_1358),
.Y(n_11660)
);

OAI21xp5_ASAP7_75t_L g11661 ( 
.A1(n_11064),
.A2(n_11094),
.B(n_11078),
.Y(n_11661)
);

NAND2xp5_ASAP7_75t_L g11662 ( 
.A(n_10702),
.B(n_10833),
.Y(n_11662)
);

OAI21x1_ASAP7_75t_L g11663 ( 
.A1(n_10707),
.A2(n_11163),
.B(n_10566),
.Y(n_11663)
);

AOI21xp5_ASAP7_75t_L g11664 ( 
.A1(n_10622),
.A2(n_1358),
.B(n_1359),
.Y(n_11664)
);

OAI22x1_ASAP7_75t_L g11665 ( 
.A1(n_11027),
.A2(n_1362),
.B1(n_1360),
.B2(n_1361),
.Y(n_11665)
);

AOI21x1_ASAP7_75t_L g11666 ( 
.A1(n_10701),
.A2(n_1360),
.B(n_1361),
.Y(n_11666)
);

NAND2x1p5_ASAP7_75t_L g11667 ( 
.A(n_10788),
.B(n_10819),
.Y(n_11667)
);

OAI22x1_ASAP7_75t_L g11668 ( 
.A1(n_11015),
.A2(n_1364),
.B1(n_1362),
.B2(n_1363),
.Y(n_11668)
);

OAI21x1_ASAP7_75t_L g11669 ( 
.A1(n_11214),
.A2(n_10693),
.B(n_10689),
.Y(n_11669)
);

OAI21x1_ASAP7_75t_L g11670 ( 
.A1(n_10694),
.A2(n_1364),
.B(n_1365),
.Y(n_11670)
);

NAND2xp5_ASAP7_75t_L g11671 ( 
.A(n_10839),
.B(n_1365),
.Y(n_11671)
);

NAND2xp5_ASAP7_75t_L g11672 ( 
.A(n_10842),
.B(n_10849),
.Y(n_11672)
);

OAI21x1_ASAP7_75t_L g11673 ( 
.A1(n_10711),
.A2(n_10742),
.B(n_10736),
.Y(n_11673)
);

INVx1_ASAP7_75t_L g11674 ( 
.A(n_10780),
.Y(n_11674)
);

INVx2_ASAP7_75t_L g11675 ( 
.A(n_10781),
.Y(n_11675)
);

OAI21x1_ASAP7_75t_L g11676 ( 
.A1(n_10968),
.A2(n_1366),
.B(n_1367),
.Y(n_11676)
);

OAI21x1_ASAP7_75t_L g11677 ( 
.A1(n_10999),
.A2(n_1366),
.B(n_1367),
.Y(n_11677)
);

NAND2xp5_ASAP7_75t_L g11678 ( 
.A(n_10877),
.B(n_10883),
.Y(n_11678)
);

OAI22xp5_ASAP7_75t_L g11679 ( 
.A1(n_10687),
.A2(n_1370),
.B1(n_1368),
.B2(n_1369),
.Y(n_11679)
);

AO31x2_ASAP7_75t_L g11680 ( 
.A1(n_11204),
.A2(n_1370),
.A3(n_1368),
.B(n_1369),
.Y(n_11680)
);

NAND2xp5_ASAP7_75t_L g11681 ( 
.A(n_10888),
.B(n_1372),
.Y(n_11681)
);

NOR2xp33_ASAP7_75t_L g11682 ( 
.A(n_10649),
.B(n_1372),
.Y(n_11682)
);

OAI21xp5_ASAP7_75t_L g11683 ( 
.A1(n_11206),
.A2(n_1373),
.B(n_1374),
.Y(n_11683)
);

NAND2xp5_ASAP7_75t_L g11684 ( 
.A(n_10890),
.B(n_1373),
.Y(n_11684)
);

INVx3_ASAP7_75t_L g11685 ( 
.A(n_10648),
.Y(n_11685)
);

INVx2_ASAP7_75t_L g11686 ( 
.A(n_10670),
.Y(n_11686)
);

OAI21x1_ASAP7_75t_L g11687 ( 
.A1(n_11216),
.A2(n_1374),
.B(n_1375),
.Y(n_11687)
);

OAI21xp5_ASAP7_75t_L g11688 ( 
.A1(n_10915),
.A2(n_1376),
.B(n_1377),
.Y(n_11688)
);

INVx2_ASAP7_75t_L g11689 ( 
.A(n_10709),
.Y(n_11689)
);

BUFx6f_ASAP7_75t_L g11690 ( 
.A(n_10776),
.Y(n_11690)
);

O2A1O1Ixp33_ASAP7_75t_SL g11691 ( 
.A1(n_11234),
.A2(n_1380),
.B(n_1378),
.C(n_1379),
.Y(n_11691)
);

INVx1_ASAP7_75t_L g11692 ( 
.A(n_10629),
.Y(n_11692)
);

OA21x2_ASAP7_75t_L g11693 ( 
.A1(n_10723),
.A2(n_1378),
.B(n_1380),
.Y(n_11693)
);

OAI21x1_ASAP7_75t_L g11694 ( 
.A1(n_10639),
.A2(n_1382),
.B(n_1383),
.Y(n_11694)
);

NAND2xp5_ASAP7_75t_L g11695 ( 
.A(n_10897),
.B(n_1382),
.Y(n_11695)
);

INVx1_ASAP7_75t_L g11696 ( 
.A(n_10740),
.Y(n_11696)
);

NAND2xp5_ASAP7_75t_L g11697 ( 
.A(n_10903),
.B(n_1383),
.Y(n_11697)
);

OR2x2_ASAP7_75t_L g11698 ( 
.A(n_10614),
.B(n_1384),
.Y(n_11698)
);

NAND2xp5_ASAP7_75t_SL g11699 ( 
.A(n_11095),
.B(n_1385),
.Y(n_11699)
);

AOI22xp5_ASAP7_75t_L g11700 ( 
.A1(n_10782),
.A2(n_1387),
.B1(n_1385),
.B2(n_1386),
.Y(n_11700)
);

AND3x4_ASAP7_75t_L g11701 ( 
.A(n_11166),
.B(n_1386),
.C(n_1387),
.Y(n_11701)
);

OAI21x1_ASAP7_75t_L g11702 ( 
.A1(n_10942),
.A2(n_1388),
.B(n_1389),
.Y(n_11702)
);

OAI21xp5_ASAP7_75t_L g11703 ( 
.A1(n_11201),
.A2(n_1388),
.B(n_1389),
.Y(n_11703)
);

AOI21xp5_ASAP7_75t_L g11704 ( 
.A1(n_11170),
.A2(n_1390),
.B(n_1391),
.Y(n_11704)
);

AND2x4_ASAP7_75t_L g11705 ( 
.A(n_10793),
.B(n_1390),
.Y(n_11705)
);

OAI21x1_ASAP7_75t_L g11706 ( 
.A1(n_11220),
.A2(n_1391),
.B(n_1392),
.Y(n_11706)
);

OAI21x1_ASAP7_75t_L g11707 ( 
.A1(n_11149),
.A2(n_1392),
.B(n_1393),
.Y(n_11707)
);

INVx2_ASAP7_75t_L g11708 ( 
.A(n_10848),
.Y(n_11708)
);

BUFx2_ASAP7_75t_L g11709 ( 
.A(n_10636),
.Y(n_11709)
);

OR2x2_ASAP7_75t_L g11710 ( 
.A(n_10616),
.B(n_1393),
.Y(n_11710)
);

AND2x4_ASAP7_75t_L g11711 ( 
.A(n_10982),
.B(n_1394),
.Y(n_11711)
);

NAND2xp5_ASAP7_75t_L g11712 ( 
.A(n_10912),
.B(n_1394),
.Y(n_11712)
);

NAND2xp5_ASAP7_75t_L g11713 ( 
.A(n_10926),
.B(n_1395),
.Y(n_11713)
);

AOI21xp5_ASAP7_75t_L g11714 ( 
.A1(n_11170),
.A2(n_1395),
.B(n_1396),
.Y(n_11714)
);

OAI21x1_ASAP7_75t_L g11715 ( 
.A1(n_10809),
.A2(n_1397),
.B(n_1398),
.Y(n_11715)
);

AO21x1_ASAP7_75t_L g11716 ( 
.A1(n_11008),
.A2(n_1398),
.B(n_1399),
.Y(n_11716)
);

NAND2xp5_ASAP7_75t_SL g11717 ( 
.A(n_11205),
.B(n_10931),
.Y(n_11717)
);

AOI22xp5_ASAP7_75t_L g11718 ( 
.A1(n_11137),
.A2(n_1401),
.B1(n_1399),
.B2(n_1400),
.Y(n_11718)
);

NAND2xp5_ASAP7_75t_SL g11719 ( 
.A(n_11208),
.B(n_1400),
.Y(n_11719)
);

INVx1_ASAP7_75t_SL g11720 ( 
.A(n_10857),
.Y(n_11720)
);

NAND2x1_ASAP7_75t_L g11721 ( 
.A(n_10820),
.B(n_1401),
.Y(n_11721)
);

NAND2xp5_ASAP7_75t_L g11722 ( 
.A(n_10928),
.B(n_1402),
.Y(n_11722)
);

NAND2xp5_ASAP7_75t_L g11723 ( 
.A(n_10944),
.B(n_1402),
.Y(n_11723)
);

NAND2xp5_ASAP7_75t_L g11724 ( 
.A(n_10946),
.B(n_1403),
.Y(n_11724)
);

AOI21xp5_ASAP7_75t_L g11725 ( 
.A1(n_10635),
.A2(n_1404),
.B(n_1405),
.Y(n_11725)
);

OAI21x1_ASAP7_75t_L g11726 ( 
.A1(n_10810),
.A2(n_1404),
.B(n_1405),
.Y(n_11726)
);

NAND2xp5_ASAP7_75t_L g11727 ( 
.A(n_10952),
.B(n_1406),
.Y(n_11727)
);

OAI21x1_ASAP7_75t_L g11728 ( 
.A1(n_11207),
.A2(n_1406),
.B(n_1407),
.Y(n_11728)
);

INVx1_ASAP7_75t_L g11729 ( 
.A(n_10676),
.Y(n_11729)
);

INVx1_ASAP7_75t_SL g11730 ( 
.A(n_11134),
.Y(n_11730)
);

OAI21x1_ASAP7_75t_L g11731 ( 
.A1(n_10989),
.A2(n_10992),
.B(n_10991),
.Y(n_11731)
);

OAI21x1_ASAP7_75t_L g11732 ( 
.A1(n_10997),
.A2(n_1407),
.B(n_1408),
.Y(n_11732)
);

NAND2xp5_ASAP7_75t_L g11733 ( 
.A(n_10618),
.B(n_1409),
.Y(n_11733)
);

CKINVDCx12_ASAP7_75t_R g11734 ( 
.A(n_10589),
.Y(n_11734)
);

NOR2x1_ASAP7_75t_L g11735 ( 
.A(n_10981),
.B(n_1410),
.Y(n_11735)
);

A2O1A1Ixp33_ASAP7_75t_L g11736 ( 
.A1(n_10800),
.A2(n_1413),
.B(n_1411),
.C(n_1412),
.Y(n_11736)
);

O2A1O1Ixp5_ASAP7_75t_L g11737 ( 
.A1(n_10624),
.A2(n_1414),
.B(n_1411),
.C(n_1413),
.Y(n_11737)
);

OAI21x1_ASAP7_75t_SL g11738 ( 
.A1(n_10646),
.A2(n_1414),
.B(n_1415),
.Y(n_11738)
);

OAI21x1_ASAP7_75t_L g11739 ( 
.A1(n_11005),
.A2(n_1415),
.B(n_1416),
.Y(n_11739)
);

AND2x2_ASAP7_75t_L g11740 ( 
.A(n_11061),
.B(n_1416),
.Y(n_11740)
);

INVx3_ASAP7_75t_L g11741 ( 
.A(n_10559),
.Y(n_11741)
);

OAI21x1_ASAP7_75t_L g11742 ( 
.A1(n_11013),
.A2(n_1418),
.B(n_1419),
.Y(n_11742)
);

AOI21xp5_ASAP7_75t_L g11743 ( 
.A1(n_11111),
.A2(n_1419),
.B(n_1421),
.Y(n_11743)
);

OAI21xp5_ASAP7_75t_L g11744 ( 
.A1(n_11251),
.A2(n_1421),
.B(n_1422),
.Y(n_11744)
);

NAND2xp5_ASAP7_75t_L g11745 ( 
.A(n_11195),
.B(n_1422),
.Y(n_11745)
);

NAND2xp5_ASAP7_75t_L g11746 ( 
.A(n_10925),
.B(n_1423),
.Y(n_11746)
);

AOI21xp5_ASAP7_75t_L g11747 ( 
.A1(n_10699),
.A2(n_1423),
.B(n_1424),
.Y(n_11747)
);

NAND2xp5_ASAP7_75t_L g11748 ( 
.A(n_10927),
.B(n_1424),
.Y(n_11748)
);

OAI21x1_ASAP7_75t_L g11749 ( 
.A1(n_11032),
.A2(n_1425),
.B(n_1426),
.Y(n_11749)
);

A2O1A1Ixp33_ASAP7_75t_L g11750 ( 
.A1(n_10804),
.A2(n_1428),
.B(n_1426),
.C(n_1427),
.Y(n_11750)
);

AO21x2_ASAP7_75t_L g11751 ( 
.A1(n_11120),
.A2(n_1427),
.B(n_1428),
.Y(n_11751)
);

OAI21x1_ASAP7_75t_L g11752 ( 
.A1(n_10869),
.A2(n_1429),
.B(n_1430),
.Y(n_11752)
);

OAI21x1_ASAP7_75t_L g11753 ( 
.A1(n_10840),
.A2(n_1429),
.B(n_1430),
.Y(n_11753)
);

NAND2x1_ASAP7_75t_L g11754 ( 
.A(n_10680),
.B(n_1431),
.Y(n_11754)
);

OA21x2_ASAP7_75t_L g11755 ( 
.A1(n_10876),
.A2(n_1431),
.B(n_1432),
.Y(n_11755)
);

NAND2xp5_ASAP7_75t_L g11756 ( 
.A(n_10954),
.B(n_1432),
.Y(n_11756)
);

AOI21xp5_ASAP7_75t_L g11757 ( 
.A1(n_10918),
.A2(n_1433),
.B(n_1434),
.Y(n_11757)
);

NAND2xp5_ASAP7_75t_L g11758 ( 
.A(n_11069),
.B(n_11096),
.Y(n_11758)
);

OAI21x1_ASAP7_75t_L g11759 ( 
.A1(n_11016),
.A2(n_1433),
.B(n_1434),
.Y(n_11759)
);

A2O1A1Ixp33_ASAP7_75t_L g11760 ( 
.A1(n_10824),
.A2(n_10826),
.B(n_10829),
.C(n_10825),
.Y(n_11760)
);

AND2x4_ASAP7_75t_L g11761 ( 
.A(n_11048),
.B(n_1435),
.Y(n_11761)
);

NAND2xp5_ASAP7_75t_L g11762 ( 
.A(n_11101),
.B(n_1435),
.Y(n_11762)
);

OAI21x1_ASAP7_75t_L g11763 ( 
.A1(n_11019),
.A2(n_10700),
.B(n_11100),
.Y(n_11763)
);

NAND2xp5_ASAP7_75t_L g11764 ( 
.A(n_11106),
.B(n_1436),
.Y(n_11764)
);

NAND2xp5_ASAP7_75t_L g11765 ( 
.A(n_10558),
.B(n_1436),
.Y(n_11765)
);

INVxp67_ASAP7_75t_SL g11766 ( 
.A(n_10658),
.Y(n_11766)
);

AOI21xp5_ASAP7_75t_SL g11767 ( 
.A1(n_11256),
.A2(n_1438),
.B(n_1439),
.Y(n_11767)
);

INVx1_ASAP7_75t_L g11768 ( 
.A(n_10680),
.Y(n_11768)
);

OAI22xp5_ASAP7_75t_L g11769 ( 
.A1(n_10771),
.A2(n_1440),
.B1(n_1438),
.B2(n_1439),
.Y(n_11769)
);

AOI21xp5_ASAP7_75t_L g11770 ( 
.A1(n_11121),
.A2(n_1441),
.B(n_1442),
.Y(n_11770)
);

NAND2xp5_ASAP7_75t_L g11771 ( 
.A(n_11018),
.B(n_11084),
.Y(n_11771)
);

INVx3_ASAP7_75t_L g11772 ( 
.A(n_10559),
.Y(n_11772)
);

OAI21x1_ASAP7_75t_L g11773 ( 
.A1(n_11065),
.A2(n_1442),
.B(n_1443),
.Y(n_11773)
);

OAI21x1_ASAP7_75t_SL g11774 ( 
.A1(n_10647),
.A2(n_1443),
.B(n_1444),
.Y(n_11774)
);

NAND2xp5_ASAP7_75t_L g11775 ( 
.A(n_11136),
.B(n_1445),
.Y(n_11775)
);

OAI22xp5_ASAP7_75t_L g11776 ( 
.A1(n_10578),
.A2(n_1447),
.B1(n_1445),
.B2(n_1446),
.Y(n_11776)
);

BUFx8_ASAP7_75t_L g11777 ( 
.A(n_10619),
.Y(n_11777)
);

NAND2xp5_ASAP7_75t_SL g11778 ( 
.A(n_11060),
.B(n_1446),
.Y(n_11778)
);

OAI22xp5_ASAP7_75t_L g11779 ( 
.A1(n_10775),
.A2(n_1449),
.B1(n_1447),
.B2(n_1448),
.Y(n_11779)
);

OAI22xp5_ASAP7_75t_L g11780 ( 
.A1(n_10778),
.A2(n_1450),
.B1(n_1448),
.B2(n_1449),
.Y(n_11780)
);

NAND2xp5_ASAP7_75t_L g11781 ( 
.A(n_11158),
.B(n_1450),
.Y(n_11781)
);

AOI21xp5_ASAP7_75t_L g11782 ( 
.A1(n_11124),
.A2(n_1451),
.B(n_1452),
.Y(n_11782)
);

AND2x2_ASAP7_75t_L g11783 ( 
.A(n_11091),
.B(n_10573),
.Y(n_11783)
);

OAI22xp5_ASAP7_75t_L g11784 ( 
.A1(n_11240),
.A2(n_11257),
.B1(n_10985),
.B2(n_11190),
.Y(n_11784)
);

NAND2xp5_ASAP7_75t_L g11785 ( 
.A(n_11179),
.B(n_1451),
.Y(n_11785)
);

OA22x2_ASAP7_75t_L g11786 ( 
.A1(n_10589),
.A2(n_1454),
.B1(n_1452),
.B2(n_1453),
.Y(n_11786)
);

OAI21x1_ASAP7_75t_L g11787 ( 
.A1(n_11067),
.A2(n_1454),
.B(n_1455),
.Y(n_11787)
);

AOI21x1_ASAP7_75t_L g11788 ( 
.A1(n_10600),
.A2(n_1455),
.B(n_1456),
.Y(n_11788)
);

OAI21x1_ASAP7_75t_L g11789 ( 
.A1(n_10738),
.A2(n_1456),
.B(n_1457),
.Y(n_11789)
);

AOI221xp5_ASAP7_75t_L g11790 ( 
.A1(n_10563),
.A2(n_1460),
.B1(n_1458),
.B2(n_1459),
.C(n_1461),
.Y(n_11790)
);

INVx2_ASAP7_75t_L g11791 ( 
.A(n_10540),
.Y(n_11791)
);

AOI21xp5_ASAP7_75t_L g11792 ( 
.A1(n_11177),
.A2(n_1458),
.B(n_1460),
.Y(n_11792)
);

OAI21xp5_ASAP7_75t_L g11793 ( 
.A1(n_11198),
.A2(n_11150),
.B(n_11232),
.Y(n_11793)
);

OAI22xp5_ASAP7_75t_L g11794 ( 
.A1(n_11081),
.A2(n_1463),
.B1(n_1461),
.B2(n_1462),
.Y(n_11794)
);

NAND2xp5_ASAP7_75t_L g11795 ( 
.A(n_11021),
.B(n_11029),
.Y(n_11795)
);

OA21x2_ASAP7_75t_L g11796 ( 
.A1(n_11130),
.A2(n_1462),
.B(n_1463),
.Y(n_11796)
);

INVx2_ASAP7_75t_L g11797 ( 
.A(n_11225),
.Y(n_11797)
);

OAI21x1_ASAP7_75t_L g11798 ( 
.A1(n_10549),
.A2(n_1464),
.B(n_1465),
.Y(n_11798)
);

OAI22x1_ASAP7_75t_L g11799 ( 
.A1(n_10988),
.A2(n_1466),
.B1(n_1464),
.B2(n_1465),
.Y(n_11799)
);

BUFx2_ASAP7_75t_L g11800 ( 
.A(n_10565),
.Y(n_11800)
);

OAI22xp5_ASAP7_75t_L g11801 ( 
.A1(n_10983),
.A2(n_1468),
.B1(n_1466),
.B2(n_1467),
.Y(n_11801)
);

NAND2xp33_ASAP7_75t_L g11802 ( 
.A(n_10881),
.B(n_1467),
.Y(n_11802)
);

OR2x2_ASAP7_75t_L g11803 ( 
.A(n_10816),
.B(n_1468),
.Y(n_11803)
);

OAI21xp5_ASAP7_75t_L g11804 ( 
.A1(n_11255),
.A2(n_11026),
.B(n_10794),
.Y(n_11804)
);

NOR2xp33_ASAP7_75t_L g11805 ( 
.A(n_11182),
.B(n_1469),
.Y(n_11805)
);

OAI22xp5_ASAP7_75t_L g11806 ( 
.A1(n_11209),
.A2(n_1472),
.B1(n_1470),
.B2(n_1471),
.Y(n_11806)
);

OAI21x1_ASAP7_75t_L g11807 ( 
.A1(n_10555),
.A2(n_1470),
.B(n_1471),
.Y(n_11807)
);

NAND2xp5_ASAP7_75t_L g11808 ( 
.A(n_11185),
.B(n_1472),
.Y(n_11808)
);

AOI21xp5_ASAP7_75t_L g11809 ( 
.A1(n_11044),
.A2(n_1473),
.B(n_1474),
.Y(n_11809)
);

CKINVDCx8_ASAP7_75t_R g11810 ( 
.A(n_10799),
.Y(n_11810)
);

NAND2xp5_ASAP7_75t_L g11811 ( 
.A(n_11176),
.B(n_11184),
.Y(n_11811)
);

INVx1_ASAP7_75t_SL g11812 ( 
.A(n_11083),
.Y(n_11812)
);

OR2x2_ASAP7_75t_L g11813 ( 
.A(n_10823),
.B(n_1473),
.Y(n_11813)
);

NAND2xp5_ASAP7_75t_L g11814 ( 
.A(n_11062),
.B(n_1474),
.Y(n_11814)
);

AOI21xp33_ASAP7_75t_L g11815 ( 
.A1(n_10770),
.A2(n_1475),
.B(n_1476),
.Y(n_11815)
);

OAI21x1_ASAP7_75t_L g11816 ( 
.A1(n_11132),
.A2(n_1475),
.B(n_1476),
.Y(n_11816)
);

AO31x2_ASAP7_75t_L g11817 ( 
.A1(n_10777),
.A2(n_1479),
.A3(n_1477),
.B(n_1478),
.Y(n_11817)
);

INVx2_ASAP7_75t_L g11818 ( 
.A(n_10945),
.Y(n_11818)
);

BUFx12f_ASAP7_75t_L g11819 ( 
.A(n_10886),
.Y(n_11819)
);

NAND2xp5_ASAP7_75t_L g11820 ( 
.A(n_11066),
.B(n_1477),
.Y(n_11820)
);

INVx1_ASAP7_75t_L g11821 ( 
.A(n_11110),
.Y(n_11821)
);

NOR2xp33_ASAP7_75t_L g11822 ( 
.A(n_10760),
.B(n_1478),
.Y(n_11822)
);

OAI21x1_ASAP7_75t_L g11823 ( 
.A1(n_11098),
.A2(n_1479),
.B(n_1480),
.Y(n_11823)
);

OAI21x1_ASAP7_75t_L g11824 ( 
.A1(n_11221),
.A2(n_1480),
.B(n_1481),
.Y(n_11824)
);

INVx1_ASAP7_75t_L g11825 ( 
.A(n_11110),
.Y(n_11825)
);

NAND2xp5_ASAP7_75t_L g11826 ( 
.A(n_11073),
.B(n_1481),
.Y(n_11826)
);

AOI211x1_ASAP7_75t_L g11827 ( 
.A1(n_10919),
.A2(n_1484),
.B(n_1482),
.C(n_1483),
.Y(n_11827)
);

INVx2_ASAP7_75t_L g11828 ( 
.A(n_10568),
.Y(n_11828)
);

AND2x2_ASAP7_75t_L g11829 ( 
.A(n_10617),
.B(n_1482),
.Y(n_11829)
);

INVx1_ASAP7_75t_L g11830 ( 
.A(n_11082),
.Y(n_11830)
);

OAI22x1_ASAP7_75t_L g11831 ( 
.A1(n_10644),
.A2(n_1486),
.B1(n_1483),
.B2(n_1484),
.Y(n_11831)
);

INVx1_ASAP7_75t_SL g11832 ( 
.A(n_10818),
.Y(n_11832)
);

BUFx3_ASAP7_75t_L g11833 ( 
.A(n_10799),
.Y(n_11833)
);

NOR2x1_ASAP7_75t_SL g11834 ( 
.A(n_10568),
.B(n_1486),
.Y(n_11834)
);

OAI21x1_ASAP7_75t_L g11835 ( 
.A1(n_11089),
.A2(n_1487),
.B(n_1488),
.Y(n_11835)
);

OAI21x1_ASAP7_75t_SL g11836 ( 
.A1(n_10606),
.A2(n_1488),
.B(n_1489),
.Y(n_11836)
);

CKINVDCx5p33_ASAP7_75t_R g11837 ( 
.A(n_10790),
.Y(n_11837)
);

OAI21x1_ASAP7_75t_L g11838 ( 
.A1(n_11093),
.A2(n_1490),
.B(n_1491),
.Y(n_11838)
);

NAND2xp5_ASAP7_75t_L g11839 ( 
.A(n_10962),
.B(n_1490),
.Y(n_11839)
);

NAND2x1p5_ASAP7_75t_L g11840 ( 
.A(n_10939),
.B(n_1492),
.Y(n_11840)
);

NAND2xp5_ASAP7_75t_L g11841 ( 
.A(n_10964),
.B(n_1493),
.Y(n_11841)
);

OAI21x1_ASAP7_75t_L g11842 ( 
.A1(n_11167),
.A2(n_1494),
.B(n_1495),
.Y(n_11842)
);

INVx4_ASAP7_75t_L g11843 ( 
.A(n_10580),
.Y(n_11843)
);

INVx1_ASAP7_75t_L g11844 ( 
.A(n_10830),
.Y(n_11844)
);

BUFx8_ASAP7_75t_L g11845 ( 
.A(n_10817),
.Y(n_11845)
);

AOI21xp5_ASAP7_75t_L g11846 ( 
.A1(n_11191),
.A2(n_1494),
.B(n_1496),
.Y(n_11846)
);

NAND2xp5_ASAP7_75t_L g11847 ( 
.A(n_11141),
.B(n_1496),
.Y(n_11847)
);

NAND2xp5_ASAP7_75t_SL g11848 ( 
.A(n_11060),
.B(n_1497),
.Y(n_11848)
);

OAI21xp5_ASAP7_75t_L g11849 ( 
.A1(n_10844),
.A2(n_1498),
.B(n_1499),
.Y(n_11849)
);

BUFx6f_ASAP7_75t_L g11850 ( 
.A(n_10817),
.Y(n_11850)
);

NAND2xp5_ASAP7_75t_L g11851 ( 
.A(n_11123),
.B(n_1498),
.Y(n_11851)
);

INVx4_ASAP7_75t_L g11852 ( 
.A(n_10580),
.Y(n_11852)
);

AO21x1_ASAP7_75t_L g11853 ( 
.A1(n_10692),
.A2(n_1499),
.B(n_1500),
.Y(n_11853)
);

NAND2xp5_ASAP7_75t_L g11854 ( 
.A(n_11129),
.B(n_11142),
.Y(n_11854)
);

INVx5_ASAP7_75t_L g11855 ( 
.A(n_10881),
.Y(n_11855)
);

NAND2xp5_ASAP7_75t_L g11856 ( 
.A(n_11169),
.B(n_1500),
.Y(n_11856)
);

AOI21xp5_ASAP7_75t_L g11857 ( 
.A1(n_11075),
.A2(n_1501),
.B(n_1502),
.Y(n_11857)
);

AOI21xp5_ASAP7_75t_L g11858 ( 
.A1(n_10665),
.A2(n_1501),
.B(n_1502),
.Y(n_11858)
);

OAI21x1_ASAP7_75t_L g11859 ( 
.A1(n_10831),
.A2(n_11001),
.B(n_11215),
.Y(n_11859)
);

AND2x4_ASAP7_75t_L g11860 ( 
.A(n_11464),
.B(n_10553),
.Y(n_11860)
);

OAI21x1_ASAP7_75t_L g11861 ( 
.A1(n_11304),
.A2(n_11173),
.B(n_11172),
.Y(n_11861)
);

OR2x6_ASAP7_75t_L g11862 ( 
.A(n_11528),
.B(n_11087),
.Y(n_11862)
);

OAI21x1_ASAP7_75t_L g11863 ( 
.A1(n_11271),
.A2(n_11175),
.B(n_11154),
.Y(n_11863)
);

AND2x2_ASAP7_75t_L g11864 ( 
.A(n_11326),
.B(n_10637),
.Y(n_11864)
);

OAI21x1_ASAP7_75t_L g11865 ( 
.A1(n_11396),
.A2(n_11146),
.B(n_11041),
.Y(n_11865)
);

BUFx6f_ASAP7_75t_L g11866 ( 
.A(n_11323),
.Y(n_11866)
);

AOI22xp33_ASAP7_75t_L g11867 ( 
.A1(n_11815),
.A2(n_10910),
.B1(n_10971),
.B2(n_10967),
.Y(n_11867)
);

INVx3_ASAP7_75t_L g11868 ( 
.A(n_11332),
.Y(n_11868)
);

INVx1_ASAP7_75t_L g11869 ( 
.A(n_11506),
.Y(n_11869)
);

INVxp67_ASAP7_75t_SL g11870 ( 
.A(n_11292),
.Y(n_11870)
);

INVx1_ASAP7_75t_L g11871 ( 
.A(n_11322),
.Y(n_11871)
);

AO21x2_ASAP7_75t_L g11872 ( 
.A1(n_11291),
.A2(n_11159),
.B(n_10596),
.Y(n_11872)
);

BUFx2_ASAP7_75t_L g11873 ( 
.A(n_11344),
.Y(n_11873)
);

BUFx6f_ASAP7_75t_L g11874 ( 
.A(n_11392),
.Y(n_11874)
);

AO21x2_ASAP7_75t_L g11875 ( 
.A1(n_11284),
.A2(n_10874),
.B(n_10728),
.Y(n_11875)
);

OAI21x1_ASAP7_75t_L g11876 ( 
.A1(n_11268),
.A2(n_11025),
.B(n_10745),
.Y(n_11876)
);

BUFx2_ASAP7_75t_SL g11877 ( 
.A(n_11303),
.Y(n_11877)
);

INVxp67_ASAP7_75t_SL g11878 ( 
.A(n_11341),
.Y(n_11878)
);

OR2x6_ASAP7_75t_L g11879 ( 
.A(n_11528),
.B(n_11087),
.Y(n_11879)
);

BUFx6f_ASAP7_75t_L g11880 ( 
.A(n_11392),
.Y(n_11880)
);

INVx1_ASAP7_75t_L g11881 ( 
.A(n_11336),
.Y(n_11881)
);

OAI21x1_ASAP7_75t_L g11882 ( 
.A1(n_11266),
.A2(n_10726),
.B(n_10663),
.Y(n_11882)
);

NAND2x1p5_ASAP7_75t_L g11883 ( 
.A(n_11855),
.B(n_10792),
.Y(n_11883)
);

NAND2xp5_ASAP7_75t_SL g11884 ( 
.A(n_11855),
.B(n_10632),
.Y(n_11884)
);

OAI21x1_ASAP7_75t_L g11885 ( 
.A1(n_11574),
.A2(n_11696),
.B(n_11515),
.Y(n_11885)
);

BUFx2_ASAP7_75t_L g11886 ( 
.A(n_11347),
.Y(n_11886)
);

INVx1_ASAP7_75t_L g11887 ( 
.A(n_11354),
.Y(n_11887)
);

INVx1_ASAP7_75t_L g11888 ( 
.A(n_11355),
.Y(n_11888)
);

AOI21xp33_ASAP7_75t_L g11889 ( 
.A1(n_11280),
.A2(n_11118),
.B(n_10930),
.Y(n_11889)
);

INVx2_ASAP7_75t_L g11890 ( 
.A(n_11513),
.Y(n_11890)
);

INVx1_ASAP7_75t_L g11891 ( 
.A(n_11356),
.Y(n_11891)
);

OAI21x1_ASAP7_75t_L g11892 ( 
.A1(n_11270),
.A2(n_11408),
.B(n_11669),
.Y(n_11892)
);

INVx1_ASAP7_75t_SL g11893 ( 
.A(n_11730),
.Y(n_11893)
);

INVx1_ASAP7_75t_L g11894 ( 
.A(n_11403),
.Y(n_11894)
);

INVx2_ASAP7_75t_L g11895 ( 
.A(n_11405),
.Y(n_11895)
);

INVx2_ASAP7_75t_L g11896 ( 
.A(n_11435),
.Y(n_11896)
);

INVx1_ASAP7_75t_SL g11897 ( 
.A(n_11345),
.Y(n_11897)
);

BUFx3_ASAP7_75t_L g11898 ( 
.A(n_11300),
.Y(n_11898)
);

INVx3_ASAP7_75t_L g11899 ( 
.A(n_11366),
.Y(n_11899)
);

BUFx3_ASAP7_75t_L g11900 ( 
.A(n_11845),
.Y(n_11900)
);

BUFx6f_ASAP7_75t_L g11901 ( 
.A(n_11422),
.Y(n_11901)
);

INVx8_ASAP7_75t_L g11902 ( 
.A(n_11303),
.Y(n_11902)
);

OA21x2_ASAP7_75t_L g11903 ( 
.A1(n_11673),
.A2(n_10641),
.B(n_10750),
.Y(n_11903)
);

INVx2_ASAP7_75t_L g11904 ( 
.A(n_11451),
.Y(n_11904)
);

OAI21x1_ASAP7_75t_L g11905 ( 
.A1(n_11433),
.A2(n_11113),
.B(n_11038),
.Y(n_11905)
);

AND2x4_ASAP7_75t_L g11906 ( 
.A(n_11514),
.B(n_10577),
.Y(n_11906)
);

AO21x2_ASAP7_75t_L g11907 ( 
.A1(n_11329),
.A2(n_10772),
.B(n_10759),
.Y(n_11907)
);

INVx1_ASAP7_75t_SL g11908 ( 
.A(n_11832),
.Y(n_11908)
);

BUFx12f_ASAP7_75t_L g11909 ( 
.A(n_11311),
.Y(n_11909)
);

INVx2_ASAP7_75t_L g11910 ( 
.A(n_11460),
.Y(n_11910)
);

AND2x4_ASAP7_75t_L g11911 ( 
.A(n_11384),
.B(n_10632),
.Y(n_11911)
);

NAND2xp5_ASAP7_75t_L g11912 ( 
.A(n_11342),
.B(n_11316),
.Y(n_11912)
);

INVx1_ASAP7_75t_L g11913 ( 
.A(n_11473),
.Y(n_11913)
);

INVx1_ASAP7_75t_L g11914 ( 
.A(n_11495),
.Y(n_11914)
);

BUFx2_ASAP7_75t_L g11915 ( 
.A(n_11667),
.Y(n_11915)
);

INVx2_ASAP7_75t_L g11916 ( 
.A(n_11504),
.Y(n_11916)
);

INVx2_ASAP7_75t_L g11917 ( 
.A(n_11305),
.Y(n_11917)
);

CKINVDCx10_ASAP7_75t_R g11918 ( 
.A(n_11350),
.Y(n_11918)
);

NAND2x1p5_ASAP7_75t_L g11919 ( 
.A(n_11489),
.B(n_10801),
.Y(n_11919)
);

INVx1_ASAP7_75t_L g11920 ( 
.A(n_11423),
.Y(n_11920)
);

OAI21x1_ASAP7_75t_L g11921 ( 
.A1(n_11417),
.A2(n_11116),
.B(n_10836),
.Y(n_11921)
);

OAI21x1_ASAP7_75t_L g11922 ( 
.A1(n_11331),
.A2(n_10785),
.B(n_11003),
.Y(n_11922)
);

NAND2x1p5_ASAP7_75t_L g11923 ( 
.A(n_11448),
.B(n_10827),
.Y(n_11923)
);

INVx2_ASAP7_75t_L g11924 ( 
.A(n_11286),
.Y(n_11924)
);

BUFx4f_ASAP7_75t_SL g11925 ( 
.A(n_11819),
.Y(n_11925)
);

BUFx2_ASAP7_75t_L g11926 ( 
.A(n_11768),
.Y(n_11926)
);

INVx1_ASAP7_75t_L g11927 ( 
.A(n_11477),
.Y(n_11927)
);

NOR2xp33_ASAP7_75t_L g11928 ( 
.A(n_11653),
.B(n_11393),
.Y(n_11928)
);

INVx1_ASAP7_75t_L g11929 ( 
.A(n_11380),
.Y(n_11929)
);

INVx6_ASAP7_75t_L g11930 ( 
.A(n_11445),
.Y(n_11930)
);

INVx3_ASAP7_75t_SL g11931 ( 
.A(n_11837),
.Y(n_11931)
);

AO21x1_ASAP7_75t_L g11932 ( 
.A1(n_11802),
.A2(n_10887),
.B(n_10866),
.Y(n_11932)
);

INVx8_ASAP7_75t_L g11933 ( 
.A(n_11263),
.Y(n_11933)
);

OAI21x1_ASAP7_75t_SL g11934 ( 
.A1(n_11309),
.A2(n_10753),
.B(n_10703),
.Y(n_11934)
);

OAI21x1_ASAP7_75t_L g11935 ( 
.A1(n_11265),
.A2(n_10762),
.B(n_10739),
.Y(n_11935)
);

BUFx8_ASAP7_75t_L g11936 ( 
.A(n_11263),
.Y(n_11936)
);

INVx1_ASAP7_75t_L g11937 ( 
.A(n_11415),
.Y(n_11937)
);

BUFx3_ASAP7_75t_L g11938 ( 
.A(n_11296),
.Y(n_11938)
);

INVx3_ASAP7_75t_L g11939 ( 
.A(n_11358),
.Y(n_11939)
);

BUFx6f_ASAP7_75t_L g11940 ( 
.A(n_11422),
.Y(n_11940)
);

OAI21xp5_ASAP7_75t_L g11941 ( 
.A1(n_11394),
.A2(n_10881),
.B(n_10595),
.Y(n_11941)
);

INVx2_ASAP7_75t_L g11942 ( 
.A(n_11431),
.Y(n_11942)
);

BUFx2_ASAP7_75t_L g11943 ( 
.A(n_11441),
.Y(n_11943)
);

INVx1_ASAP7_75t_L g11944 ( 
.A(n_11444),
.Y(n_11944)
);

INVx1_ASAP7_75t_SL g11945 ( 
.A(n_11502),
.Y(n_11945)
);

INVx1_ASAP7_75t_L g11946 ( 
.A(n_11449),
.Y(n_11946)
);

INVx8_ASAP7_75t_L g11947 ( 
.A(n_11312),
.Y(n_11947)
);

BUFx12f_ASAP7_75t_L g11948 ( 
.A(n_11777),
.Y(n_11948)
);

OAI21x1_ASAP7_75t_L g11949 ( 
.A1(n_11587),
.A2(n_10683),
.B(n_10668),
.Y(n_11949)
);

NAND2x1p5_ASAP7_75t_L g11950 ( 
.A(n_11327),
.B(n_10660),
.Y(n_11950)
);

AO21x2_ASAP7_75t_L g11951 ( 
.A1(n_11264),
.A2(n_10620),
.B(n_11168),
.Y(n_11951)
);

NAND2x1p5_ASAP7_75t_L g11952 ( 
.A(n_11709),
.B(n_10660),
.Y(n_11952)
);

INVx1_ASAP7_75t_L g11953 ( 
.A(n_11471),
.Y(n_11953)
);

NAND2x1p5_ASAP7_75t_L g11954 ( 
.A(n_11580),
.B(n_10677),
.Y(n_11954)
);

BUFx6f_ASAP7_75t_L g11955 ( 
.A(n_11476),
.Y(n_11955)
);

OAI21x1_ASAP7_75t_L g11956 ( 
.A1(n_11518),
.A2(n_10976),
.B(n_10963),
.Y(n_11956)
);

INVx2_ASAP7_75t_SL g11957 ( 
.A(n_11618),
.Y(n_11957)
);

BUFx6f_ASAP7_75t_L g11958 ( 
.A(n_11476),
.Y(n_11958)
);

OAI21x1_ASAP7_75t_L g11959 ( 
.A1(n_11272),
.A2(n_11133),
.B(n_11112),
.Y(n_11959)
);

INVx2_ASAP7_75t_L g11960 ( 
.A(n_11497),
.Y(n_11960)
);

INVx2_ASAP7_75t_SL g11961 ( 
.A(n_11424),
.Y(n_11961)
);

INVx1_ASAP7_75t_L g11962 ( 
.A(n_11480),
.Y(n_11962)
);

INVx4_ASAP7_75t_L g11963 ( 
.A(n_11455),
.Y(n_11963)
);

INVx3_ASAP7_75t_L g11964 ( 
.A(n_11685),
.Y(n_11964)
);

HB1xp67_ASAP7_75t_L g11965 ( 
.A(n_11483),
.Y(n_11965)
);

INVx1_ASAP7_75t_SL g11966 ( 
.A(n_11812),
.Y(n_11966)
);

AOI22x1_ASAP7_75t_L g11967 ( 
.A1(n_11704),
.A2(n_11014),
.B1(n_10708),
.B2(n_11063),
.Y(n_11967)
);

OAI21x1_ASAP7_75t_L g11968 ( 
.A1(n_11663),
.A2(n_11143),
.B(n_10922),
.Y(n_11968)
);

OAI21xp5_ASAP7_75t_L g11969 ( 
.A1(n_11401),
.A2(n_10932),
.B(n_10900),
.Y(n_11969)
);

INVx2_ASAP7_75t_L g11970 ( 
.A(n_11282),
.Y(n_11970)
);

BUFx6f_ASAP7_75t_L g11971 ( 
.A(n_11533),
.Y(n_11971)
);

INVxp67_ASAP7_75t_SL g11972 ( 
.A(n_11452),
.Y(n_11972)
);

NOR2xp33_ASAP7_75t_L g11973 ( 
.A(n_11335),
.B(n_10677),
.Y(n_11973)
);

INVx1_ASAP7_75t_L g11974 ( 
.A(n_11532),
.Y(n_11974)
);

AO21x2_ASAP7_75t_L g11975 ( 
.A1(n_11714),
.A2(n_10834),
.B(n_11072),
.Y(n_11975)
);

INVx8_ASAP7_75t_L g11976 ( 
.A(n_11312),
.Y(n_11976)
);

INVx1_ASAP7_75t_SL g11977 ( 
.A(n_11584),
.Y(n_11977)
);

AO21x2_ASAP7_75t_L g11978 ( 
.A1(n_11276),
.A2(n_10830),
.B(n_11181),
.Y(n_11978)
);

BUFx2_ASAP7_75t_L g11979 ( 
.A(n_11630),
.Y(n_11979)
);

INVx3_ASAP7_75t_SL g11980 ( 
.A(n_11541),
.Y(n_11980)
);

INVx2_ASAP7_75t_SL g11981 ( 
.A(n_11463),
.Y(n_11981)
);

AND2x2_ASAP7_75t_L g11982 ( 
.A(n_11600),
.B(n_10697),
.Y(n_11982)
);

AO21x2_ASAP7_75t_L g11983 ( 
.A1(n_11290),
.A2(n_11125),
.B(n_10697),
.Y(n_11983)
);

CKINVDCx11_ASAP7_75t_R g11984 ( 
.A(n_11308),
.Y(n_11984)
);

AO21x2_ASAP7_75t_L g11985 ( 
.A1(n_11315),
.A2(n_11200),
.B(n_11242),
.Y(n_11985)
);

AOI22x1_ASAP7_75t_L g11986 ( 
.A1(n_11573),
.A2(n_11242),
.B1(n_1505),
.B2(n_1503),
.Y(n_11986)
);

AO21x2_ASAP7_75t_L g11987 ( 
.A1(n_11317),
.A2(n_1503),
.B(n_1504),
.Y(n_11987)
);

INVx4_ASAP7_75t_L g11988 ( 
.A(n_11560),
.Y(n_11988)
);

CKINVDCx5p33_ASAP7_75t_R g11989 ( 
.A(n_11810),
.Y(n_11989)
);

INVx1_ASAP7_75t_L g11990 ( 
.A(n_11319),
.Y(n_11990)
);

INVx3_ASAP7_75t_L g11991 ( 
.A(n_11533),
.Y(n_11991)
);

INVx1_ASAP7_75t_SL g11992 ( 
.A(n_11720),
.Y(n_11992)
);

OAI21x1_ASAP7_75t_L g11993 ( 
.A1(n_11279),
.A2(n_11285),
.B(n_11278),
.Y(n_11993)
);

INVx1_ASAP7_75t_L g11994 ( 
.A(n_11282),
.Y(n_11994)
);

INVx3_ASAP7_75t_L g11995 ( 
.A(n_11535),
.Y(n_11995)
);

INVx2_ASAP7_75t_L g11996 ( 
.A(n_11282),
.Y(n_11996)
);

AO21x2_ASAP7_75t_L g11997 ( 
.A1(n_11320),
.A2(n_1504),
.B(n_1505),
.Y(n_11997)
);

OR3x4_ASAP7_75t_SL g11998 ( 
.A(n_11766),
.B(n_1506),
.C(n_1507),
.Y(n_11998)
);

BUFx6f_ASAP7_75t_L g11999 ( 
.A(n_11535),
.Y(n_11999)
);

OAI21x1_ASAP7_75t_L g12000 ( 
.A1(n_11397),
.A2(n_1507),
.B(n_1508),
.Y(n_12000)
);

INVx1_ASAP7_75t_L g12001 ( 
.A(n_11282),
.Y(n_12001)
);

INVx1_ASAP7_75t_L g12002 ( 
.A(n_11381),
.Y(n_12002)
);

INVx4_ASAP7_75t_L g12003 ( 
.A(n_11321),
.Y(n_12003)
);

BUFx3_ASAP7_75t_L g12004 ( 
.A(n_11310),
.Y(n_12004)
);

NAND2xp5_ASAP7_75t_L g12005 ( 
.A(n_11549),
.B(n_1508),
.Y(n_12005)
);

AO21x1_ASAP7_75t_L g12006 ( 
.A1(n_11822),
.A2(n_1509),
.B(n_1510),
.Y(n_12006)
);

CKINVDCx5p33_ASAP7_75t_R g12007 ( 
.A(n_11321),
.Y(n_12007)
);

INVx4_ASAP7_75t_L g12008 ( 
.A(n_11338),
.Y(n_12008)
);

OAI21xp5_ASAP7_75t_L g12009 ( 
.A1(n_11416),
.A2(n_1509),
.B(n_1510),
.Y(n_12009)
);

OAI21x1_ASAP7_75t_L g12010 ( 
.A1(n_11399),
.A2(n_11389),
.B(n_11334),
.Y(n_12010)
);

OAI21xp5_ASAP7_75t_L g12011 ( 
.A1(n_11493),
.A2(n_1511),
.B(n_1512),
.Y(n_12011)
);

AOI21x1_ASAP7_75t_L g12012 ( 
.A1(n_11699),
.A2(n_1511),
.B(n_1512),
.Y(n_12012)
);

INVx4_ASAP7_75t_L g12013 ( 
.A(n_11338),
.Y(n_12013)
);

INVx2_ASAP7_75t_L g12014 ( 
.A(n_11620),
.Y(n_12014)
);

INVx3_ASAP7_75t_L g12015 ( 
.A(n_11557),
.Y(n_12015)
);

BUFx3_ASAP7_75t_L g12016 ( 
.A(n_11833),
.Y(n_12016)
);

INVx2_ASAP7_75t_L g12017 ( 
.A(n_11649),
.Y(n_12017)
);

BUFx6f_ASAP7_75t_SL g12018 ( 
.A(n_11711),
.Y(n_12018)
);

NAND3xp33_ASAP7_75t_SL g12019 ( 
.A(n_11512),
.B(n_1513),
.C(n_1514),
.Y(n_12019)
);

INVx3_ASAP7_75t_L g12020 ( 
.A(n_11557),
.Y(n_12020)
);

OA21x2_ASAP7_75t_L g12021 ( 
.A1(n_11844),
.A2(n_1514),
.B(n_1515),
.Y(n_12021)
);

INVx4_ASAP7_75t_L g12022 ( 
.A(n_11346),
.Y(n_12022)
);

OAI21x1_ASAP7_75t_L g12023 ( 
.A1(n_11351),
.A2(n_1515),
.B(n_1517),
.Y(n_12023)
);

INVx4_ASAP7_75t_L g12024 ( 
.A(n_11346),
.Y(n_12024)
);

OAI21x1_ASAP7_75t_L g12025 ( 
.A1(n_11340),
.A2(n_1517),
.B(n_1518),
.Y(n_12025)
);

AO21x2_ASAP7_75t_L g12026 ( 
.A1(n_11267),
.A2(n_1518),
.B(n_1519),
.Y(n_12026)
);

OA21x2_ASAP7_75t_L g12027 ( 
.A1(n_11821),
.A2(n_1519),
.B(n_1520),
.Y(n_12027)
);

CKINVDCx16_ASAP7_75t_R g12028 ( 
.A(n_11536),
.Y(n_12028)
);

INVx5_ASAP7_75t_L g12029 ( 
.A(n_11659),
.Y(n_12029)
);

AND2x4_ASAP7_75t_L g12030 ( 
.A(n_11609),
.B(n_1521),
.Y(n_12030)
);

INVx3_ASAP7_75t_L g12031 ( 
.A(n_11843),
.Y(n_12031)
);

INVx3_ASAP7_75t_SL g12032 ( 
.A(n_11293),
.Y(n_12032)
);

OAI21x1_ASAP7_75t_SL g12033 ( 
.A1(n_11716),
.A2(n_11641),
.B(n_11853),
.Y(n_12033)
);

AOI22xp33_ASAP7_75t_L g12034 ( 
.A1(n_11793),
.A2(n_1523),
.B1(n_1521),
.B2(n_1522),
.Y(n_12034)
);

CKINVDCx5p33_ASAP7_75t_R g12035 ( 
.A(n_11659),
.Y(n_12035)
);

INVx1_ASAP7_75t_L g12036 ( 
.A(n_11613),
.Y(n_12036)
);

INVx1_ASAP7_75t_L g12037 ( 
.A(n_11642),
.Y(n_12037)
);

OAI21xp5_ASAP7_75t_L g12038 ( 
.A1(n_11508),
.A2(n_1522),
.B(n_1523),
.Y(n_12038)
);

BUFx3_ASAP7_75t_L g12039 ( 
.A(n_11690),
.Y(n_12039)
);

INVx4_ASAP7_75t_L g12040 ( 
.A(n_11690),
.Y(n_12040)
);

BUFx8_ASAP7_75t_L g12041 ( 
.A(n_11740),
.Y(n_12041)
);

NAND2xp5_ASAP7_75t_L g12042 ( 
.A(n_11558),
.B(n_1524),
.Y(n_12042)
);

INVx1_ASAP7_75t_SL g12043 ( 
.A(n_11800),
.Y(n_12043)
);

NAND2x1p5_ASAP7_75t_L g12044 ( 
.A(n_11275),
.B(n_1525),
.Y(n_12044)
);

BUFx6f_ASAP7_75t_L g12045 ( 
.A(n_11850),
.Y(n_12045)
);

NAND2x1p5_ASAP7_75t_L g12046 ( 
.A(n_11604),
.B(n_1526),
.Y(n_12046)
);

INVx3_ASAP7_75t_SL g12047 ( 
.A(n_11301),
.Y(n_12047)
);

OAI21x1_ASAP7_75t_L g12048 ( 
.A1(n_11359),
.A2(n_1527),
.B(n_1528),
.Y(n_12048)
);

INVx1_ASAP7_75t_L g12049 ( 
.A(n_11647),
.Y(n_12049)
);

BUFx3_ASAP7_75t_L g12050 ( 
.A(n_11850),
.Y(n_12050)
);

INVx1_ASAP7_75t_L g12051 ( 
.A(n_11674),
.Y(n_12051)
);

BUFx6f_ASAP7_75t_L g12052 ( 
.A(n_11741),
.Y(n_12052)
);

AND2x4_ASAP7_75t_L g12053 ( 
.A(n_11686),
.B(n_11689),
.Y(n_12053)
);

INVx2_ASAP7_75t_SL g12054 ( 
.A(n_11708),
.Y(n_12054)
);

INVx1_ASAP7_75t_L g12055 ( 
.A(n_11579),
.Y(n_12055)
);

INVx2_ASAP7_75t_L g12056 ( 
.A(n_11675),
.Y(n_12056)
);

OAI21x1_ASAP7_75t_L g12057 ( 
.A1(n_11325),
.A2(n_1527),
.B(n_1529),
.Y(n_12057)
);

NAND2x1p5_ASAP7_75t_L g12058 ( 
.A(n_11721),
.B(n_1529),
.Y(n_12058)
);

INVx8_ASAP7_75t_L g12059 ( 
.A(n_11705),
.Y(n_12059)
);

BUFx12f_ASAP7_75t_L g12060 ( 
.A(n_11840),
.Y(n_12060)
);

INVx2_ASAP7_75t_L g12061 ( 
.A(n_11590),
.Y(n_12061)
);

NAND2x1p5_ASAP7_75t_L g12062 ( 
.A(n_11754),
.B(n_1530),
.Y(n_12062)
);

INVx6_ASAP7_75t_L g12063 ( 
.A(n_11852),
.Y(n_12063)
);

AND2x4_ASAP7_75t_L g12064 ( 
.A(n_11828),
.B(n_1530),
.Y(n_12064)
);

OAI21x1_ASAP7_75t_L g12065 ( 
.A1(n_11379),
.A2(n_1531),
.B(n_1532),
.Y(n_12065)
);

INVx1_ASAP7_75t_L g12066 ( 
.A(n_11547),
.Y(n_12066)
);

AO21x2_ASAP7_75t_L g12067 ( 
.A1(n_11458),
.A2(n_1531),
.B(n_1532),
.Y(n_12067)
);

INVx2_ASAP7_75t_L g12068 ( 
.A(n_11692),
.Y(n_12068)
);

OAI21xp5_ASAP7_75t_L g12069 ( 
.A1(n_11352),
.A2(n_1533),
.B(n_1534),
.Y(n_12069)
);

INVx1_ASAP7_75t_L g12070 ( 
.A(n_11474),
.Y(n_12070)
);

NOR2x1_ASAP7_75t_R g12071 ( 
.A(n_11651),
.B(n_1533),
.Y(n_12071)
);

INVx1_ASAP7_75t_L g12072 ( 
.A(n_11475),
.Y(n_12072)
);

OAI21x1_ASAP7_75t_L g12073 ( 
.A1(n_11407),
.A2(n_1534),
.B(n_1535),
.Y(n_12073)
);

INVx2_ASAP7_75t_L g12074 ( 
.A(n_11729),
.Y(n_12074)
);

OAI21x1_ASAP7_75t_L g12075 ( 
.A1(n_11333),
.A2(n_1536),
.B(n_1537),
.Y(n_12075)
);

INVx1_ASAP7_75t_L g12076 ( 
.A(n_11499),
.Y(n_12076)
);

AOI22x1_ASAP7_75t_L g12077 ( 
.A1(n_11617),
.A2(n_11799),
.B1(n_11353),
.B2(n_11665),
.Y(n_12077)
);

OAI21xp5_ASAP7_75t_L g12078 ( 
.A1(n_11487),
.A2(n_1536),
.B(n_1537),
.Y(n_12078)
);

INVx4_ASAP7_75t_L g12079 ( 
.A(n_11772),
.Y(n_12079)
);

INVx2_ASAP7_75t_SL g12080 ( 
.A(n_11488),
.Y(n_12080)
);

INVx1_ASAP7_75t_L g12081 ( 
.A(n_11522),
.Y(n_12081)
);

INVx1_ASAP7_75t_L g12082 ( 
.A(n_11825),
.Y(n_12082)
);

OAI21x1_ASAP7_75t_L g12083 ( 
.A1(n_11273),
.A2(n_1538),
.B(n_1539),
.Y(n_12083)
);

BUFx3_ASAP7_75t_L g12084 ( 
.A(n_11783),
.Y(n_12084)
);

INVx8_ASAP7_75t_L g12085 ( 
.A(n_11761),
.Y(n_12085)
);

INVx1_ASAP7_75t_L g12086 ( 
.A(n_11486),
.Y(n_12086)
);

OA21x2_ASAP7_75t_L g12087 ( 
.A1(n_11731),
.A2(n_1538),
.B(n_1539),
.Y(n_12087)
);

BUFx2_ASAP7_75t_R g12088 ( 
.A(n_11602),
.Y(n_12088)
);

INVx1_ASAP7_75t_L g12089 ( 
.A(n_11491),
.Y(n_12089)
);

NAND2xp5_ASAP7_75t_L g12090 ( 
.A(n_11830),
.B(n_1540),
.Y(n_12090)
);

CKINVDCx5p33_ASAP7_75t_R g12091 ( 
.A(n_11734),
.Y(n_12091)
);

CKINVDCx16_ASAP7_75t_R g12092 ( 
.A(n_11299),
.Y(n_12092)
);

BUFx3_ASAP7_75t_L g12093 ( 
.A(n_11791),
.Y(n_12093)
);

AND2x2_ASAP7_75t_L g12094 ( 
.A(n_11797),
.B(n_1540),
.Y(n_12094)
);

NAND2xp5_ASAP7_75t_L g12095 ( 
.A(n_11607),
.B(n_1541),
.Y(n_12095)
);

OR2x2_ASAP7_75t_L g12096 ( 
.A(n_11274),
.B(n_1542),
.Y(n_12096)
);

BUFx2_ASAP7_75t_SL g12097 ( 
.A(n_11430),
.Y(n_12097)
);

OAI21x1_ASAP7_75t_L g12098 ( 
.A1(n_11306),
.A2(n_1542),
.B(n_1544),
.Y(n_12098)
);

NOR2xp33_ASAP7_75t_L g12099 ( 
.A(n_11672),
.B(n_1544),
.Y(n_12099)
);

INVx1_ASAP7_75t_L g12100 ( 
.A(n_11544),
.Y(n_12100)
);

INVx2_ASAP7_75t_L g12101 ( 
.A(n_11818),
.Y(n_12101)
);

BUFx12f_ASAP7_75t_L g12102 ( 
.A(n_11437),
.Y(n_12102)
);

HB1xp67_ASAP7_75t_L g12103 ( 
.A(n_11578),
.Y(n_12103)
);

BUFx3_ASAP7_75t_L g12104 ( 
.A(n_11624),
.Y(n_12104)
);

INVx1_ASAP7_75t_L g12105 ( 
.A(n_11482),
.Y(n_12105)
);

BUFx8_ASAP7_75t_L g12106 ( 
.A(n_11644),
.Y(n_12106)
);

NOR2xp33_ASAP7_75t_L g12107 ( 
.A(n_11678),
.B(n_1545),
.Y(n_12107)
);

OAI21x1_ASAP7_75t_L g12108 ( 
.A1(n_11328),
.A2(n_1545),
.B(n_1546),
.Y(n_12108)
);

BUFx12f_ASAP7_75t_L g12109 ( 
.A(n_11509),
.Y(n_12109)
);

AND2x2_ASAP7_75t_L g12110 ( 
.A(n_11287),
.B(n_1547),
.Y(n_12110)
);

INVx2_ASAP7_75t_L g12111 ( 
.A(n_11302),
.Y(n_12111)
);

INVx1_ASAP7_75t_L g12112 ( 
.A(n_11330),
.Y(n_12112)
);

AOI21x1_ASAP7_75t_L g12113 ( 
.A1(n_11562),
.A2(n_1547),
.B(n_1548),
.Y(n_12113)
);

INVx2_ASAP7_75t_L g12114 ( 
.A(n_11337),
.Y(n_12114)
);

AND2x4_ASAP7_75t_L g12115 ( 
.A(n_11369),
.B(n_1548),
.Y(n_12115)
);

AO21x2_ASAP7_75t_L g12116 ( 
.A1(n_11339),
.A2(n_11479),
.B(n_11375),
.Y(n_12116)
);

NOR2xp33_ASAP7_75t_L g12117 ( 
.A(n_11662),
.B(n_1549),
.Y(n_12117)
);

AO21x2_ASAP7_75t_L g12118 ( 
.A1(n_11462),
.A2(n_1549),
.B(n_1550),
.Y(n_12118)
);

OAI21x1_ASAP7_75t_L g12119 ( 
.A1(n_11360),
.A2(n_1551),
.B(n_1552),
.Y(n_12119)
);

HB1xp67_ASAP7_75t_L g12120 ( 
.A(n_11796),
.Y(n_12120)
);

CKINVDCx6p67_ASAP7_75t_R g12121 ( 
.A(n_11548),
.Y(n_12121)
);

INVxp67_ASAP7_75t_SL g12122 ( 
.A(n_11391),
.Y(n_12122)
);

OAI21x1_ASAP7_75t_L g12123 ( 
.A1(n_11365),
.A2(n_1551),
.B(n_1552),
.Y(n_12123)
);

INVx1_ASAP7_75t_L g12124 ( 
.A(n_11409),
.Y(n_12124)
);

AOI22x1_ASAP7_75t_L g12125 ( 
.A1(n_11363),
.A2(n_1555),
.B1(n_1553),
.B2(n_1554),
.Y(n_12125)
);

INVx2_ASAP7_75t_L g12126 ( 
.A(n_11614),
.Y(n_12126)
);

INVx1_ASAP7_75t_L g12127 ( 
.A(n_11413),
.Y(n_12127)
);

OAI21x1_ASAP7_75t_L g12128 ( 
.A1(n_11371),
.A2(n_1553),
.B(n_1555),
.Y(n_12128)
);

INVx1_ASAP7_75t_L g12129 ( 
.A(n_11414),
.Y(n_12129)
);

INVx1_ASAP7_75t_L g12130 ( 
.A(n_11421),
.Y(n_12130)
);

BUFx2_ASAP7_75t_L g12131 ( 
.A(n_11288),
.Y(n_12131)
);

OAI21xp5_ASAP7_75t_L g12132 ( 
.A1(n_11378),
.A2(n_1556),
.B(n_1557),
.Y(n_12132)
);

OAI21x1_ASAP7_75t_L g12133 ( 
.A1(n_11702),
.A2(n_1556),
.B(n_1558),
.Y(n_12133)
);

OAI21x1_ASAP7_75t_L g12134 ( 
.A1(n_11687),
.A2(n_1558),
.B(n_1559),
.Y(n_12134)
);

BUFx3_ASAP7_75t_L g12135 ( 
.A(n_11395),
.Y(n_12135)
);

OAI21x1_ASAP7_75t_L g12136 ( 
.A1(n_11566),
.A2(n_1559),
.B(n_1560),
.Y(n_12136)
);

INVx1_ASAP7_75t_L g12137 ( 
.A(n_11427),
.Y(n_12137)
);

AO21x2_ASAP7_75t_L g12138 ( 
.A1(n_11447),
.A2(n_1561),
.B(n_1562),
.Y(n_12138)
);

OAI21x1_ASAP7_75t_L g12139 ( 
.A1(n_11440),
.A2(n_1562),
.B(n_1563),
.Y(n_12139)
);

INVx2_ASAP7_75t_SL g12140 ( 
.A(n_11307),
.Y(n_12140)
);

INVx1_ASAP7_75t_L g12141 ( 
.A(n_11432),
.Y(n_12141)
);

AO21x2_ASAP7_75t_L g12142 ( 
.A1(n_11295),
.A2(n_11538),
.B(n_11374),
.Y(n_12142)
);

BUFx3_ASAP7_75t_L g12143 ( 
.A(n_11516),
.Y(n_12143)
);

INVx2_ASAP7_75t_L g12144 ( 
.A(n_11410),
.Y(n_12144)
);

OAI21x1_ASAP7_75t_L g12145 ( 
.A1(n_11442),
.A2(n_1563),
.B(n_1564),
.Y(n_12145)
);

INVx1_ASAP7_75t_L g12146 ( 
.A(n_11434),
.Y(n_12146)
);

HB1xp67_ASAP7_75t_L g12147 ( 
.A(n_11563),
.Y(n_12147)
);

HB1xp67_ASAP7_75t_L g12148 ( 
.A(n_11438),
.Y(n_12148)
);

BUFx12f_ASAP7_75t_L g12149 ( 
.A(n_11803),
.Y(n_12149)
);

INVx1_ASAP7_75t_SL g12150 ( 
.A(n_11402),
.Y(n_12150)
);

CKINVDCx20_ASAP7_75t_R g12151 ( 
.A(n_11811),
.Y(n_12151)
);

NAND2xp5_ASAP7_75t_L g12152 ( 
.A(n_11795),
.B(n_1564),
.Y(n_12152)
);

CKINVDCx20_ASAP7_75t_R g12153 ( 
.A(n_11854),
.Y(n_12153)
);

INVx3_ASAP7_75t_L g12154 ( 
.A(n_11698),
.Y(n_12154)
);

INVx1_ASAP7_75t_SL g12155 ( 
.A(n_11530),
.Y(n_12155)
);

OAI21x1_ASAP7_75t_L g12156 ( 
.A1(n_11450),
.A2(n_1565),
.B(n_1566),
.Y(n_12156)
);

INVx1_ASAP7_75t_L g12157 ( 
.A(n_11446),
.Y(n_12157)
);

AOI22x1_ASAP7_75t_L g12158 ( 
.A1(n_11668),
.A2(n_1567),
.B1(n_1565),
.B2(n_1566),
.Y(n_12158)
);

INVx2_ASAP7_75t_L g12159 ( 
.A(n_11277),
.Y(n_12159)
);

OAI21xp5_ASAP7_75t_L g12160 ( 
.A1(n_11498),
.A2(n_1567),
.B(n_1568),
.Y(n_12160)
);

BUFx6f_ASAP7_75t_L g12161 ( 
.A(n_11701),
.Y(n_12161)
);

OAI21x1_ASAP7_75t_L g12162 ( 
.A1(n_11456),
.A2(n_1569),
.B(n_1570),
.Y(n_12162)
);

INVx3_ASAP7_75t_L g12163 ( 
.A(n_11710),
.Y(n_12163)
);

OAI21xp5_ASAP7_75t_L g12164 ( 
.A1(n_11570),
.A2(n_1572),
.B(n_1573),
.Y(n_12164)
);

AO21x1_ASAP7_75t_SL g12165 ( 
.A1(n_11661),
.A2(n_1572),
.B(n_1573),
.Y(n_12165)
);

HB1xp67_ASAP7_75t_L g12166 ( 
.A(n_11519),
.Y(n_12166)
);

INVx3_ASAP7_75t_L g12167 ( 
.A(n_11281),
.Y(n_12167)
);

OAI21x1_ASAP7_75t_L g12168 ( 
.A1(n_11465),
.A2(n_1574),
.B(n_1575),
.Y(n_12168)
);

CKINVDCx5p33_ASAP7_75t_R g12169 ( 
.A(n_11682),
.Y(n_12169)
);

OR2x2_ASAP7_75t_L g12170 ( 
.A(n_11771),
.B(n_1574),
.Y(n_12170)
);

OAI21x1_ASAP7_75t_L g12171 ( 
.A1(n_11469),
.A2(n_1575),
.B(n_1576),
.Y(n_12171)
);

HB1xp67_ASAP7_75t_L g12172 ( 
.A(n_11527),
.Y(n_12172)
);

OAI21x1_ASAP7_75t_L g12173 ( 
.A1(n_11478),
.A2(n_1576),
.B(n_1577),
.Y(n_12173)
);

BUFx3_ASAP7_75t_L g12174 ( 
.A(n_11406),
.Y(n_12174)
);

INVx4_ASAP7_75t_L g12175 ( 
.A(n_11373),
.Y(n_12175)
);

INVx2_ASAP7_75t_L g12176 ( 
.A(n_11367),
.Y(n_12176)
);

CKINVDCx20_ASAP7_75t_R g12177 ( 
.A(n_11717),
.Y(n_12177)
);

BUFx6f_ASAP7_75t_L g12178 ( 
.A(n_11376),
.Y(n_12178)
);

INVx2_ASAP7_75t_L g12179 ( 
.A(n_11537),
.Y(n_12179)
);

INVx1_ASAP7_75t_L g12180 ( 
.A(n_11534),
.Y(n_12180)
);

INVx1_ASAP7_75t_SL g12181 ( 
.A(n_11813),
.Y(n_12181)
);

AO21x2_ASAP7_75t_L g12182 ( 
.A1(n_11294),
.A2(n_1577),
.B(n_1578),
.Y(n_12182)
);

INVx2_ASAP7_75t_SL g12183 ( 
.A(n_11556),
.Y(n_12183)
);

INVx3_ASAP7_75t_L g12184 ( 
.A(n_11357),
.Y(n_12184)
);

INVx1_ASAP7_75t_L g12185 ( 
.A(n_11545),
.Y(n_12185)
);

INVx1_ASAP7_75t_L g12186 ( 
.A(n_11546),
.Y(n_12186)
);

BUFx3_ASAP7_75t_L g12187 ( 
.A(n_11638),
.Y(n_12187)
);

BUFx2_ASAP7_75t_L g12188 ( 
.A(n_11763),
.Y(n_12188)
);

INVx2_ASAP7_75t_L g12189 ( 
.A(n_11418),
.Y(n_12189)
);

INVx1_ASAP7_75t_L g12190 ( 
.A(n_11349),
.Y(n_12190)
);

AND2x2_ASAP7_75t_L g12191 ( 
.A(n_11829),
.B(n_1578),
.Y(n_12191)
);

AND2x2_ASAP7_75t_L g12192 ( 
.A(n_11657),
.B(n_11324),
.Y(n_12192)
);

INVx2_ASAP7_75t_L g12193 ( 
.A(n_11484),
.Y(n_12193)
);

INVx2_ASAP7_75t_SL g12194 ( 
.A(n_11608),
.Y(n_12194)
);

AO21x2_ASAP7_75t_L g12195 ( 
.A1(n_11703),
.A2(n_11398),
.B(n_11348),
.Y(n_12195)
);

NAND2xp5_ASAP7_75t_L g12196 ( 
.A(n_11539),
.B(n_1579),
.Y(n_12196)
);

BUFx2_ASAP7_75t_L g12197 ( 
.A(n_11582),
.Y(n_12197)
);

BUFx8_ASAP7_75t_L g12198 ( 
.A(n_11428),
.Y(n_12198)
);

AND2x2_ASAP7_75t_L g12199 ( 
.A(n_11501),
.B(n_1580),
.Y(n_12199)
);

OAI21x1_ASAP7_75t_L g12200 ( 
.A1(n_11481),
.A2(n_1580),
.B(n_1582),
.Y(n_12200)
);

INVx1_ASAP7_75t_L g12201 ( 
.A(n_11349),
.Y(n_12201)
);

BUFx12f_ASAP7_75t_L g12202 ( 
.A(n_11735),
.Y(n_12202)
);

AND2x4_ASAP7_75t_L g12203 ( 
.A(n_11670),
.B(n_1582),
.Y(n_12203)
);

INVx1_ASAP7_75t_L g12204 ( 
.A(n_11586),
.Y(n_12204)
);

AOI22x1_ASAP7_75t_L g12205 ( 
.A1(n_11313),
.A2(n_1585),
.B1(n_1583),
.B2(n_1584),
.Y(n_12205)
);

OA21x2_ASAP7_75t_L g12206 ( 
.A1(n_11472),
.A2(n_1583),
.B(n_1585),
.Y(n_12206)
);

OR2x6_ASAP7_75t_L g12207 ( 
.A(n_11605),
.B(n_1586),
.Y(n_12207)
);

BUFx3_ASAP7_75t_L g12208 ( 
.A(n_11658),
.Y(n_12208)
);

OAI21x1_ASAP7_75t_L g12209 ( 
.A1(n_11507),
.A2(n_1586),
.B(n_1587),
.Y(n_12209)
);

INVx2_ASAP7_75t_L g12210 ( 
.A(n_11715),
.Y(n_12210)
);

CKINVDCx11_ASAP7_75t_R g12211 ( 
.A(n_11784),
.Y(n_12211)
);

OAI21x1_ASAP7_75t_L g12212 ( 
.A1(n_11523),
.A2(n_1588),
.B(n_1589),
.Y(n_12212)
);

OAI21x1_ASAP7_75t_L g12213 ( 
.A1(n_11526),
.A2(n_1588),
.B(n_1590),
.Y(n_12213)
);

INVx2_ASAP7_75t_L g12214 ( 
.A(n_11726),
.Y(n_12214)
);

NOR2xp67_ASAP7_75t_SL g12215 ( 
.A(n_11594),
.B(n_1590),
.Y(n_12215)
);

AO21x2_ASAP7_75t_L g12216 ( 
.A1(n_11314),
.A2(n_1591),
.B(n_1592),
.Y(n_12216)
);

OA21x2_ASAP7_75t_L g12217 ( 
.A1(n_11732),
.A2(n_11742),
.B(n_11739),
.Y(n_12217)
);

INVx1_ASAP7_75t_SL g12218 ( 
.A(n_11758),
.Y(n_12218)
);

AOI22x1_ASAP7_75t_L g12219 ( 
.A1(n_11364),
.A2(n_1593),
.B1(n_1591),
.B2(n_1592),
.Y(n_12219)
);

INVx1_ASAP7_75t_L g12220 ( 
.A(n_11586),
.Y(n_12220)
);

INVx1_ASAP7_75t_L g12221 ( 
.A(n_11835),
.Y(n_12221)
);

AO21x2_ASAP7_75t_L g12222 ( 
.A1(n_11370),
.A2(n_11743),
.B(n_11400),
.Y(n_12222)
);

AO21x2_ASAP7_75t_L g12223 ( 
.A1(n_11485),
.A2(n_1594),
.B(n_1595),
.Y(n_12223)
);

AO21x2_ASAP7_75t_L g12224 ( 
.A1(n_11559),
.A2(n_1594),
.B(n_1595),
.Y(n_12224)
);

INVx1_ASAP7_75t_L g12225 ( 
.A(n_11838),
.Y(n_12225)
);

OAI21x1_ASAP7_75t_L g12226 ( 
.A1(n_11543),
.A2(n_1596),
.B(n_1597),
.Y(n_12226)
);

OAI21x1_ASAP7_75t_L g12227 ( 
.A1(n_11550),
.A2(n_1596),
.B(n_1597),
.Y(n_12227)
);

OAI21x1_ASAP7_75t_L g12228 ( 
.A1(n_11554),
.A2(n_1598),
.B(n_1599),
.Y(n_12228)
);

INVx3_ASAP7_75t_L g12229 ( 
.A(n_11759),
.Y(n_12229)
);

INVx2_ASAP7_75t_L g12230 ( 
.A(n_11749),
.Y(n_12230)
);

OAI21x1_ASAP7_75t_L g12231 ( 
.A1(n_11577),
.A2(n_1599),
.B(n_1600),
.Y(n_12231)
);

BUFx8_ASAP7_75t_L g12232 ( 
.A(n_11834),
.Y(n_12232)
);

INVx4_ASAP7_75t_L g12233 ( 
.A(n_11786),
.Y(n_12233)
);

NAND2xp5_ASAP7_75t_SL g12234 ( 
.A(n_11804),
.B(n_1600),
.Y(n_12234)
);

INVx5_ASAP7_75t_L g12235 ( 
.A(n_11443),
.Y(n_12235)
);

AND2x4_ASAP7_75t_L g12236 ( 
.A(n_11824),
.B(n_1602),
.Y(n_12236)
);

OAI21x1_ASAP7_75t_L g12237 ( 
.A1(n_11591),
.A2(n_1602),
.B(n_1603),
.Y(n_12237)
);

BUFx8_ASAP7_75t_L g12238 ( 
.A(n_11831),
.Y(n_12238)
);

OAI21x1_ASAP7_75t_L g12239 ( 
.A1(n_11595),
.A2(n_1603),
.B(n_1604),
.Y(n_12239)
);

INVx1_ASAP7_75t_SL g12240 ( 
.A(n_11589),
.Y(n_12240)
);

INVx3_ASAP7_75t_L g12241 ( 
.A(n_11755),
.Y(n_12241)
);

BUFx2_ASAP7_75t_SL g12242 ( 
.A(n_11385),
.Y(n_12242)
);

AO21x2_ASAP7_75t_L g12243 ( 
.A1(n_11503),
.A2(n_1604),
.B(n_1605),
.Y(n_12243)
);

INVx2_ASAP7_75t_SL g12244 ( 
.A(n_11571),
.Y(n_12244)
);

BUFx6f_ASAP7_75t_L g12245 ( 
.A(n_11386),
.Y(n_12245)
);

INVx4_ASAP7_75t_L g12246 ( 
.A(n_11654),
.Y(n_12246)
);

OAI21xp5_ASAP7_75t_L g12247 ( 
.A1(n_11632),
.A2(n_1605),
.B(n_1606),
.Y(n_12247)
);

CKINVDCx5p33_ASAP7_75t_R g12248 ( 
.A(n_11764),
.Y(n_12248)
);

OAI21xp5_ASAP7_75t_L g12249 ( 
.A1(n_11470),
.A2(n_1606),
.B(n_1607),
.Y(n_12249)
);

NAND2xp5_ASAP7_75t_L g12250 ( 
.A(n_11564),
.B(n_1607),
.Y(n_12250)
);

BUFx2_ASAP7_75t_L g12251 ( 
.A(n_11572),
.Y(n_12251)
);

AO21x2_ASAP7_75t_L g12252 ( 
.A1(n_11529),
.A2(n_1608),
.B(n_1609),
.Y(n_12252)
);

BUFx3_ASAP7_75t_L g12253 ( 
.A(n_11847),
.Y(n_12253)
);

OAI21x1_ASAP7_75t_L g12254 ( 
.A1(n_11603),
.A2(n_1608),
.B(n_1609),
.Y(n_12254)
);

INVx1_ASAP7_75t_L g12255 ( 
.A(n_11390),
.Y(n_12255)
);

OAI21x1_ASAP7_75t_L g12256 ( 
.A1(n_11611),
.A2(n_1610),
.B(n_1611),
.Y(n_12256)
);

BUFx6f_ASAP7_75t_L g12257 ( 
.A(n_11583),
.Y(n_12257)
);

NAND2xp5_ASAP7_75t_L g12258 ( 
.A(n_11660),
.B(n_1610),
.Y(n_12258)
);

BUFx12f_ASAP7_75t_L g12259 ( 
.A(n_11805),
.Y(n_12259)
);

OAI21x1_ASAP7_75t_L g12260 ( 
.A1(n_11612),
.A2(n_11619),
.B(n_11615),
.Y(n_12260)
);

OAI21x1_ASAP7_75t_L g12261 ( 
.A1(n_11621),
.A2(n_1611),
.B(n_1612),
.Y(n_12261)
);

AOI21x1_ASAP7_75t_L g12262 ( 
.A1(n_11289),
.A2(n_1612),
.B(n_1613),
.Y(n_12262)
);

INVx1_ASAP7_75t_L g12263 ( 
.A(n_11693),
.Y(n_12263)
);

OR2x2_ASAP7_75t_L g12264 ( 
.A(n_11598),
.B(n_1613),
.Y(n_12264)
);

NAND2x1p5_ASAP7_75t_L g12265 ( 
.A(n_11789),
.B(n_1614),
.Y(n_12265)
);

INVx2_ASAP7_75t_L g12266 ( 
.A(n_11707),
.Y(n_12266)
);

BUFx3_ASAP7_75t_L g12267 ( 
.A(n_11765),
.Y(n_12267)
);

INVx1_ASAP7_75t_L g12268 ( 
.A(n_11728),
.Y(n_12268)
);

BUFx2_ASAP7_75t_L g12269 ( 
.A(n_11859),
.Y(n_12269)
);

BUFx3_ASAP7_75t_L g12270 ( 
.A(n_11839),
.Y(n_12270)
);

INVx2_ASAP7_75t_L g12271 ( 
.A(n_11706),
.Y(n_12271)
);

NAND2xp5_ASAP7_75t_L g12272 ( 
.A(n_11606),
.B(n_1614),
.Y(n_12272)
);

OAI21x1_ASAP7_75t_L g12273 ( 
.A1(n_11622),
.A2(n_1615),
.B(n_1616),
.Y(n_12273)
);

CKINVDCx5p33_ASAP7_75t_R g12274 ( 
.A(n_11841),
.Y(n_12274)
);

INVxp67_ASAP7_75t_SL g12275 ( 
.A(n_11599),
.Y(n_12275)
);

INVx2_ASAP7_75t_L g12276 ( 
.A(n_11525),
.Y(n_12276)
);

OAI21x1_ASAP7_75t_L g12277 ( 
.A1(n_11627),
.A2(n_1615),
.B(n_1616),
.Y(n_12277)
);

INVxp67_ASAP7_75t_SL g12278 ( 
.A(n_11633),
.Y(n_12278)
);

INVx2_ASAP7_75t_L g12279 ( 
.A(n_11552),
.Y(n_12279)
);

INVx2_ASAP7_75t_L g12280 ( 
.A(n_11569),
.Y(n_12280)
);

NAND2x1p5_ASAP7_75t_L g12281 ( 
.A(n_11778),
.B(n_1617),
.Y(n_12281)
);

BUFx3_ASAP7_75t_L g12282 ( 
.A(n_11851),
.Y(n_12282)
);

INVx2_ASAP7_75t_L g12283 ( 
.A(n_11666),
.Y(n_12283)
);

BUFx3_ASAP7_75t_L g12284 ( 
.A(n_11856),
.Y(n_12284)
);

BUFx10_ASAP7_75t_L g12285 ( 
.A(n_11636),
.Y(n_12285)
);

OAI21x1_ASAP7_75t_L g12286 ( 
.A1(n_11650),
.A2(n_1617),
.B(n_1618),
.Y(n_12286)
);

CKINVDCx6p67_ASAP7_75t_R g12287 ( 
.A(n_11848),
.Y(n_12287)
);

NAND2x1p5_ASAP7_75t_L g12288 ( 
.A(n_11816),
.B(n_1618),
.Y(n_12288)
);

NAND2x1p5_ASAP7_75t_L g12289 ( 
.A(n_11567),
.B(n_1619),
.Y(n_12289)
);

INVx1_ASAP7_75t_L g12290 ( 
.A(n_11871),
.Y(n_12290)
);

INVx1_ASAP7_75t_L g12291 ( 
.A(n_11881),
.Y(n_12291)
);

INVx2_ASAP7_75t_L g12292 ( 
.A(n_11926),
.Y(n_12292)
);

AO21x2_ASAP7_75t_L g12293 ( 
.A1(n_12081),
.A2(n_12105),
.B(n_12019),
.Y(n_12293)
);

CKINVDCx20_ASAP7_75t_R g12294 ( 
.A(n_11984),
.Y(n_12294)
);

OAI21xp5_ASAP7_75t_L g12295 ( 
.A1(n_12249),
.A2(n_11597),
.B(n_11425),
.Y(n_12295)
);

OAI21x1_ASAP7_75t_L g12296 ( 
.A1(n_11885),
.A2(n_11628),
.B(n_11387),
.Y(n_12296)
);

INVx1_ASAP7_75t_L g12297 ( 
.A(n_11887),
.Y(n_12297)
);

OAI221xp5_ASAP7_75t_L g12298 ( 
.A1(n_12160),
.A2(n_12247),
.B1(n_12164),
.B2(n_12038),
.C(n_12011),
.Y(n_12298)
);

BUFx3_ASAP7_75t_L g12299 ( 
.A(n_11948),
.Y(n_12299)
);

OAI22xp5_ASAP7_75t_L g12300 ( 
.A1(n_12235),
.A2(n_11368),
.B1(n_11490),
.B2(n_11700),
.Y(n_12300)
);

INVxp67_ASAP7_75t_SL g12301 ( 
.A(n_12103),
.Y(n_12301)
);

AO21x2_ASAP7_75t_L g12302 ( 
.A1(n_12120),
.A2(n_11688),
.B(n_11757),
.Y(n_12302)
);

NAND2xp5_ASAP7_75t_L g12303 ( 
.A(n_11878),
.B(n_11733),
.Y(n_12303)
);

AND2x2_ASAP7_75t_L g12304 ( 
.A(n_11873),
.B(n_11593),
.Y(n_12304)
);

CKINVDCx5p33_ASAP7_75t_R g12305 ( 
.A(n_11918),
.Y(n_12305)
);

OAI21x1_ASAP7_75t_L g12306 ( 
.A1(n_11892),
.A2(n_11588),
.B(n_11752),
.Y(n_12306)
);

OAI21x1_ASAP7_75t_L g12307 ( 
.A1(n_11970),
.A2(n_11626),
.B(n_11753),
.Y(n_12307)
);

AOI22xp5_ASAP7_75t_L g12308 ( 
.A1(n_12215),
.A2(n_11343),
.B1(n_11531),
.B2(n_11794),
.Y(n_12308)
);

NAND2xp5_ASAP7_75t_L g12309 ( 
.A(n_12122),
.B(n_11671),
.Y(n_12309)
);

INVx2_ASAP7_75t_L g12310 ( 
.A(n_12159),
.Y(n_12310)
);

AO21x2_ASAP7_75t_L g12311 ( 
.A1(n_12263),
.A2(n_11511),
.B(n_11540),
.Y(n_12311)
);

OR2x6_ASAP7_75t_L g12312 ( 
.A(n_11877),
.B(n_11494),
.Y(n_12312)
);

OAI21xp5_ASAP7_75t_L g12313 ( 
.A1(n_11889),
.A2(n_11468),
.B(n_11521),
.Y(n_12313)
);

OAI21x1_ASAP7_75t_L g12314 ( 
.A1(n_11996),
.A2(n_11631),
.B(n_11773),
.Y(n_12314)
);

OA21x2_ASAP7_75t_L g12315 ( 
.A1(n_12269),
.A2(n_11555),
.B(n_11681),
.Y(n_12315)
);

OA21x2_ASAP7_75t_L g12316 ( 
.A1(n_12188),
.A2(n_11695),
.B(n_11684),
.Y(n_12316)
);

NAND2xp5_ASAP7_75t_SL g12317 ( 
.A(n_12028),
.B(n_11592),
.Y(n_12317)
);

OAI21x1_ASAP7_75t_L g12318 ( 
.A1(n_11994),
.A2(n_12001),
.B(n_12241),
.Y(n_12318)
);

OAI21x1_ASAP7_75t_L g12319 ( 
.A1(n_12229),
.A2(n_11787),
.B(n_11676),
.Y(n_12319)
);

INVx3_ASAP7_75t_SL g12320 ( 
.A(n_11902),
.Y(n_12320)
);

AND2x2_ASAP7_75t_L g12321 ( 
.A(n_11886),
.B(n_11697),
.Y(n_12321)
);

AOI222xp33_ASAP7_75t_L g12322 ( 
.A1(n_12078),
.A2(n_11596),
.B1(n_11683),
.B2(n_11492),
.C1(n_11744),
.C2(n_11616),
.Y(n_12322)
);

AND2x2_ASAP7_75t_L g12323 ( 
.A(n_11979),
.B(n_11712),
.Y(n_12323)
);

INVx1_ASAP7_75t_L g12324 ( 
.A(n_11888),
.Y(n_12324)
);

BUFx2_ASAP7_75t_L g12325 ( 
.A(n_11919),
.Y(n_12325)
);

OAI22xp5_ASAP7_75t_L g12326 ( 
.A1(n_12235),
.A2(n_11524),
.B1(n_11553),
.B2(n_11439),
.Y(n_12326)
);

OAI22xp5_ASAP7_75t_L g12327 ( 
.A1(n_12233),
.A2(n_11461),
.B1(n_11467),
.B2(n_11568),
.Y(n_12327)
);

OAI22xp5_ASAP7_75t_L g12328 ( 
.A1(n_12177),
.A2(n_11575),
.B1(n_11718),
.B2(n_11520),
.Y(n_12328)
);

INVx2_ASAP7_75t_L g12329 ( 
.A(n_11895),
.Y(n_12329)
);

OAI21x1_ASAP7_75t_L g12330 ( 
.A1(n_12266),
.A2(n_11677),
.B(n_11823),
.Y(n_12330)
);

AOI21xp5_ASAP7_75t_L g12331 ( 
.A1(n_12222),
.A2(n_11767),
.B(n_11643),
.Y(n_12331)
);

INVx2_ASAP7_75t_L g12332 ( 
.A(n_11896),
.Y(n_12332)
);

OAI21x1_ASAP7_75t_L g12333 ( 
.A1(n_11993),
.A2(n_11842),
.B(n_11510),
.Y(n_12333)
);

NAND2x1p5_ASAP7_75t_L g12334 ( 
.A(n_11915),
.B(n_11646),
.Y(n_12334)
);

OAI21xp5_ASAP7_75t_L g12335 ( 
.A1(n_11949),
.A2(n_11542),
.B(n_11420),
.Y(n_12335)
);

OAI21x1_ASAP7_75t_L g12336 ( 
.A1(n_12204),
.A2(n_12220),
.B(n_12010),
.Y(n_12336)
);

A2O1A1Ixp33_ASAP7_75t_L g12337 ( 
.A1(n_11941),
.A2(n_12009),
.B(n_12234),
.C(n_11725),
.Y(n_12337)
);

NAND2xp5_ASAP7_75t_L g12338 ( 
.A(n_12066),
.B(n_11713),
.Y(n_12338)
);

OAI21xp5_ASAP7_75t_L g12339 ( 
.A1(n_11863),
.A2(n_11809),
.B(n_11601),
.Y(n_12339)
);

INVx3_ASAP7_75t_L g12340 ( 
.A(n_12079),
.Y(n_12340)
);

INVx2_ASAP7_75t_L g12341 ( 
.A(n_11904),
.Y(n_12341)
);

NOR2xp67_ASAP7_75t_L g12342 ( 
.A(n_12202),
.B(n_11722),
.Y(n_12342)
);

NAND2xp5_ASAP7_75t_L g12343 ( 
.A(n_12124),
.B(n_11723),
.Y(n_12343)
);

OAI21x1_ASAP7_75t_L g12344 ( 
.A1(n_12271),
.A2(n_11861),
.B(n_12190),
.Y(n_12344)
);

INVx1_ASAP7_75t_L g12345 ( 
.A(n_11891),
.Y(n_12345)
);

OAI21x1_ASAP7_75t_L g12346 ( 
.A1(n_12201),
.A2(n_11565),
.B(n_11377),
.Y(n_12346)
);

OAI21xp5_ASAP7_75t_L g12347 ( 
.A1(n_12069),
.A2(n_11585),
.B(n_11637),
.Y(n_12347)
);

INVx1_ASAP7_75t_L g12348 ( 
.A(n_11894),
.Y(n_12348)
);

OAI21x1_ASAP7_75t_L g12349 ( 
.A1(n_12210),
.A2(n_11372),
.B(n_11454),
.Y(n_12349)
);

AO21x2_ASAP7_75t_L g12350 ( 
.A1(n_12033),
.A2(n_11747),
.B(n_11298),
.Y(n_12350)
);

HB1xp67_ASAP7_75t_L g12351 ( 
.A(n_12230),
.Y(n_12351)
);

INVx1_ASAP7_75t_L g12352 ( 
.A(n_11913),
.Y(n_12352)
);

OAI21x1_ASAP7_75t_L g12353 ( 
.A1(n_12214),
.A2(n_11748),
.B(n_11746),
.Y(n_12353)
);

OAI21x1_ASAP7_75t_L g12354 ( 
.A1(n_11968),
.A2(n_11756),
.B(n_11798),
.Y(n_12354)
);

INVx3_ASAP7_75t_L g12355 ( 
.A(n_12003),
.Y(n_12355)
);

INVx1_ASAP7_75t_L g12356 ( 
.A(n_11914),
.Y(n_12356)
);

OAI21x1_ASAP7_75t_L g12357 ( 
.A1(n_12268),
.A2(n_11807),
.B(n_11388),
.Y(n_12357)
);

BUFx12f_ASAP7_75t_L g12358 ( 
.A(n_11866),
.Y(n_12358)
);

BUFx3_ASAP7_75t_L g12359 ( 
.A(n_11866),
.Y(n_12359)
);

OAI21x1_ASAP7_75t_L g12360 ( 
.A1(n_12260),
.A2(n_11383),
.B(n_11857),
.Y(n_12360)
);

AO31x2_ASAP7_75t_L g12361 ( 
.A1(n_12006),
.A2(n_11806),
.A3(n_11318),
.B(n_11561),
.Y(n_12361)
);

INVx2_ASAP7_75t_SL g12362 ( 
.A(n_11930),
.Y(n_12362)
);

NOR2x1_ASAP7_75t_SL g12363 ( 
.A(n_11875),
.B(n_11751),
.Y(n_12363)
);

NAND2x1p5_ASAP7_75t_L g12364 ( 
.A(n_11884),
.B(n_11719),
.Y(n_12364)
);

AOI22xp33_ASAP7_75t_L g12365 ( 
.A1(n_12211),
.A2(n_11849),
.B1(n_11297),
.B2(n_11457),
.Y(n_12365)
);

OAI21x1_ASAP7_75t_L g12366 ( 
.A1(n_12221),
.A2(n_11581),
.B(n_11411),
.Y(n_12366)
);

INVx1_ASAP7_75t_SL g12367 ( 
.A(n_12088),
.Y(n_12367)
);

OAI21x1_ASAP7_75t_SL g12368 ( 
.A1(n_11932),
.A2(n_11466),
.B(n_11459),
.Y(n_12368)
);

NAND2xp5_ASAP7_75t_L g12369 ( 
.A(n_12127),
.B(n_11724),
.Y(n_12369)
);

OR2x2_ASAP7_75t_L g12370 ( 
.A(n_11912),
.B(n_11745),
.Y(n_12370)
);

NOR2xp67_ASAP7_75t_L g12371 ( 
.A(n_11988),
.B(n_11727),
.Y(n_12371)
);

OR2x2_ASAP7_75t_L g12372 ( 
.A(n_11920),
.B(n_11655),
.Y(n_12372)
);

CKINVDCx5p33_ASAP7_75t_R g12373 ( 
.A(n_11938),
.Y(n_12373)
);

AOI21xp5_ASAP7_75t_L g12374 ( 
.A1(n_12132),
.A2(n_11907),
.B(n_11664),
.Y(n_12374)
);

INVx2_ASAP7_75t_L g12375 ( 
.A(n_11910),
.Y(n_12375)
);

INVx2_ASAP7_75t_L g12376 ( 
.A(n_11916),
.Y(n_12376)
);

NAND2xp5_ASAP7_75t_L g12377 ( 
.A(n_12129),
.B(n_12130),
.Y(n_12377)
);

INVx1_ASAP7_75t_L g12378 ( 
.A(n_11869),
.Y(n_12378)
);

OA21x2_ASAP7_75t_L g12379 ( 
.A1(n_12082),
.A2(n_11820),
.B(n_11814),
.Y(n_12379)
);

NAND2xp33_ASAP7_75t_SL g12380 ( 
.A(n_12246),
.B(n_11625),
.Y(n_12380)
);

OAI21x1_ASAP7_75t_L g12381 ( 
.A1(n_12225),
.A2(n_11412),
.B(n_11361),
.Y(n_12381)
);

INVx2_ASAP7_75t_L g12382 ( 
.A(n_12189),
.Y(n_12382)
);

NAND2xp5_ASAP7_75t_L g12383 ( 
.A(n_12137),
.B(n_11826),
.Y(n_12383)
);

INVx1_ASAP7_75t_L g12384 ( 
.A(n_11974),
.Y(n_12384)
);

OAI21x1_ASAP7_75t_L g12385 ( 
.A1(n_11882),
.A2(n_11694),
.B(n_11788),
.Y(n_12385)
);

INVx1_ASAP7_75t_L g12386 ( 
.A(n_12036),
.Y(n_12386)
);

INVx2_ASAP7_75t_SL g12387 ( 
.A(n_12063),
.Y(n_12387)
);

AOI21xp5_ASAP7_75t_L g12388 ( 
.A1(n_12206),
.A2(n_11656),
.B(n_11770),
.Y(n_12388)
);

OAI21x1_ASAP7_75t_L g12389 ( 
.A1(n_12276),
.A2(n_12280),
.B(n_12279),
.Y(n_12389)
);

INVx1_ASAP7_75t_L g12390 ( 
.A(n_12037),
.Y(n_12390)
);

OAI21x1_ASAP7_75t_L g12391 ( 
.A1(n_12283),
.A2(n_11792),
.B(n_11782),
.Y(n_12391)
);

OAI21xp5_ASAP7_75t_L g12392 ( 
.A1(n_12275),
.A2(n_11634),
.B(n_11629),
.Y(n_12392)
);

INVx2_ASAP7_75t_L g12393 ( 
.A(n_12193),
.Y(n_12393)
);

A2O1A1Ixp33_ASAP7_75t_L g12394 ( 
.A1(n_12161),
.A2(n_11760),
.B(n_11750),
.C(n_11736),
.Y(n_12394)
);

AND2x2_ASAP7_75t_L g12395 ( 
.A(n_12043),
.B(n_11762),
.Y(n_12395)
);

OAI22xp33_ASAP7_75t_L g12396 ( 
.A1(n_12092),
.A2(n_11283),
.B1(n_11679),
.B2(n_11551),
.Y(n_12396)
);

OAI21x1_ASAP7_75t_L g12397 ( 
.A1(n_12278),
.A2(n_11956),
.B(n_11921),
.Y(n_12397)
);

INVx2_ASAP7_75t_L g12398 ( 
.A(n_11927),
.Y(n_12398)
);

NAND2x1p5_ASAP7_75t_L g12399 ( 
.A(n_11992),
.B(n_11846),
.Y(n_12399)
);

OAI21x1_ASAP7_75t_L g12400 ( 
.A1(n_11959),
.A2(n_12068),
.B(n_12061),
.Y(n_12400)
);

AND2x2_ASAP7_75t_L g12401 ( 
.A(n_11965),
.B(n_11775),
.Y(n_12401)
);

HB1xp67_ASAP7_75t_L g12402 ( 
.A(n_11870),
.Y(n_12402)
);

AND2x2_ASAP7_75t_L g12403 ( 
.A(n_11943),
.B(n_11781),
.Y(n_12403)
);

AOI22xp5_ASAP7_75t_L g12404 ( 
.A1(n_11978),
.A2(n_11429),
.B1(n_11426),
.B2(n_11779),
.Y(n_12404)
);

INVxp67_ASAP7_75t_L g12405 ( 
.A(n_11903),
.Y(n_12405)
);

INVx2_ASAP7_75t_L g12406 ( 
.A(n_11890),
.Y(n_12406)
);

OAI21x1_ASAP7_75t_L g12407 ( 
.A1(n_11899),
.A2(n_11738),
.B(n_11623),
.Y(n_12407)
);

INVx1_ASAP7_75t_L g12408 ( 
.A(n_12049),
.Y(n_12408)
);

OAI21x1_ASAP7_75t_L g12409 ( 
.A1(n_12051),
.A2(n_11774),
.B(n_11737),
.Y(n_12409)
);

OAI21xp5_ASAP7_75t_L g12410 ( 
.A1(n_12117),
.A2(n_11640),
.B(n_11635),
.Y(n_12410)
);

OAI21x1_ASAP7_75t_L g12411 ( 
.A1(n_11876),
.A2(n_11652),
.B(n_11785),
.Y(n_12411)
);

INVx1_ASAP7_75t_L g12412 ( 
.A(n_11962),
.Y(n_12412)
);

OAI21x1_ASAP7_75t_L g12413 ( 
.A1(n_12055),
.A2(n_12167),
.B(n_11952),
.Y(n_12413)
);

NAND2xp5_ASAP7_75t_L g12414 ( 
.A(n_12141),
.B(n_11808),
.Y(n_12414)
);

INVx1_ASAP7_75t_L g12415 ( 
.A(n_11917),
.Y(n_12415)
);

NOR2xp33_ASAP7_75t_L g12416 ( 
.A(n_11980),
.B(n_11436),
.Y(n_12416)
);

INVx1_ASAP7_75t_L g12417 ( 
.A(n_11929),
.Y(n_12417)
);

OAI21x1_ASAP7_75t_L g12418 ( 
.A1(n_11964),
.A2(n_11836),
.B(n_11858),
.Y(n_12418)
);

OAI21xp5_ASAP7_75t_L g12419 ( 
.A1(n_12099),
.A2(n_11453),
.B(n_11790),
.Y(n_12419)
);

NOR3xp33_ASAP7_75t_L g12420 ( 
.A(n_11905),
.B(n_11801),
.C(n_11780),
.Y(n_12420)
);

OAI21x1_ASAP7_75t_L g12421 ( 
.A1(n_11950),
.A2(n_11576),
.B(n_11769),
.Y(n_12421)
);

OR2x2_ASAP7_75t_L g12422 ( 
.A(n_12154),
.B(n_11680),
.Y(n_12422)
);

HB1xp67_ASAP7_75t_L g12423 ( 
.A(n_12217),
.Y(n_12423)
);

OAI21x1_ASAP7_75t_SL g12424 ( 
.A1(n_12255),
.A2(n_11776),
.B(n_11362),
.Y(n_12424)
);

INVx2_ASAP7_75t_SL g12425 ( 
.A(n_11936),
.Y(n_12425)
);

INVx1_ASAP7_75t_L g12426 ( 
.A(n_11937),
.Y(n_12426)
);

BUFx2_ASAP7_75t_L g12427 ( 
.A(n_11883),
.Y(n_12427)
);

NAND2xp5_ASAP7_75t_L g12428 ( 
.A(n_12146),
.B(n_11362),
.Y(n_12428)
);

OA21x2_ASAP7_75t_L g12429 ( 
.A1(n_12002),
.A2(n_11680),
.B(n_11404),
.Y(n_12429)
);

AOI22xp33_ASAP7_75t_L g12430 ( 
.A1(n_12077),
.A2(n_11827),
.B1(n_11691),
.B2(n_11639),
.Y(n_12430)
);

OAI21x1_ASAP7_75t_L g12431 ( 
.A1(n_11939),
.A2(n_12179),
.B(n_12176),
.Y(n_12431)
);

AND2x2_ASAP7_75t_L g12432 ( 
.A(n_12084),
.B(n_11382),
.Y(n_12432)
);

OA21x2_ASAP7_75t_L g12433 ( 
.A1(n_11944),
.A2(n_11404),
.B(n_11382),
.Y(n_12433)
);

OAI21x1_ASAP7_75t_L g12434 ( 
.A1(n_11935),
.A2(n_11496),
.B(n_11419),
.Y(n_12434)
);

OAI21x1_ASAP7_75t_L g12435 ( 
.A1(n_12056),
.A2(n_11496),
.B(n_11419),
.Y(n_12435)
);

OAI21x1_ASAP7_75t_L g12436 ( 
.A1(n_12114),
.A2(n_11505),
.B(n_11500),
.Y(n_12436)
);

INVx1_ASAP7_75t_L g12437 ( 
.A(n_11946),
.Y(n_12437)
);

AOI21xp5_ASAP7_75t_L g12438 ( 
.A1(n_12142),
.A2(n_11639),
.B(n_11610),
.Y(n_12438)
);

OAI21x1_ASAP7_75t_SL g12439 ( 
.A1(n_12021),
.A2(n_11269),
.B(n_11817),
.Y(n_12439)
);

OAI21x1_ASAP7_75t_L g12440 ( 
.A1(n_11924),
.A2(n_11505),
.B(n_11500),
.Y(n_12440)
);

INVx2_ASAP7_75t_L g12441 ( 
.A(n_11942),
.Y(n_12441)
);

BUFx6f_ASAP7_75t_L g12442 ( 
.A(n_11900),
.Y(n_12442)
);

OAI21x1_ASAP7_75t_L g12443 ( 
.A1(n_11960),
.A2(n_11517),
.B(n_11645),
.Y(n_12443)
);

AO21x1_ASAP7_75t_L g12444 ( 
.A1(n_12192),
.A2(n_11817),
.B(n_11517),
.Y(n_12444)
);

NAND2xp5_ASAP7_75t_L g12445 ( 
.A(n_12157),
.B(n_11648),
.Y(n_12445)
);

AND2x4_ASAP7_75t_L g12446 ( 
.A(n_12053),
.B(n_11648),
.Y(n_12446)
);

INVx1_ASAP7_75t_L g12447 ( 
.A(n_11953),
.Y(n_12447)
);

OAI21x1_ASAP7_75t_SL g12448 ( 
.A1(n_12027),
.A2(n_11610),
.B(n_11645),
.Y(n_12448)
);

AND2x4_ASAP7_75t_L g12449 ( 
.A(n_11957),
.B(n_1620),
.Y(n_12449)
);

OAI21xp5_ASAP7_75t_SL g12450 ( 
.A1(n_11867),
.A2(n_1620),
.B(n_1621),
.Y(n_12450)
);

OAI21x1_ASAP7_75t_L g12451 ( 
.A1(n_11954),
.A2(n_1621),
.B(n_1622),
.Y(n_12451)
);

AND2x2_ASAP7_75t_L g12452 ( 
.A(n_11864),
.B(n_1622),
.Y(n_12452)
);

INVx1_ASAP7_75t_L g12453 ( 
.A(n_12074),
.Y(n_12453)
);

OAI21x1_ASAP7_75t_L g12454 ( 
.A1(n_12070),
.A2(n_1623),
.B(n_1624),
.Y(n_12454)
);

INVx2_ASAP7_75t_L g12455 ( 
.A(n_12014),
.Y(n_12455)
);

OAI21x1_ASAP7_75t_L g12456 ( 
.A1(n_12072),
.A2(n_1623),
.B(n_1624),
.Y(n_12456)
);

OAI21x1_ASAP7_75t_L g12457 ( 
.A1(n_12076),
.A2(n_1625),
.B(n_1626),
.Y(n_12457)
);

CKINVDCx5p33_ASAP7_75t_R g12458 ( 
.A(n_11989),
.Y(n_12458)
);

AO32x2_ASAP7_75t_L g12459 ( 
.A1(n_12183),
.A2(n_1627),
.A3(n_1625),
.B1(n_1626),
.B2(n_1628),
.Y(n_12459)
);

OAI21x1_ASAP7_75t_L g12460 ( 
.A1(n_12180),
.A2(n_12186),
.B(n_12185),
.Y(n_12460)
);

OA21x2_ASAP7_75t_L g12461 ( 
.A1(n_11990),
.A2(n_1627),
.B(n_1629),
.Y(n_12461)
);

INVx1_ASAP7_75t_L g12462 ( 
.A(n_12100),
.Y(n_12462)
);

INVx1_ASAP7_75t_L g12463 ( 
.A(n_12148),
.Y(n_12463)
);

OR2x2_ASAP7_75t_L g12464 ( 
.A(n_12163),
.B(n_1629),
.Y(n_12464)
);

INVx2_ASAP7_75t_L g12465 ( 
.A(n_12017),
.Y(n_12465)
);

OA21x2_ASAP7_75t_L g12466 ( 
.A1(n_11928),
.A2(n_12091),
.B(n_12112),
.Y(n_12466)
);

CKINVDCx16_ASAP7_75t_R g12467 ( 
.A(n_11998),
.Y(n_12467)
);

OAI21x1_ASAP7_75t_SL g12468 ( 
.A1(n_12012),
.A2(n_1630),
.B(n_1631),
.Y(n_12468)
);

OAI21x1_ASAP7_75t_L g12469 ( 
.A1(n_12184),
.A2(n_1631),
.B(n_1632),
.Y(n_12469)
);

OAI21x1_ASAP7_75t_L g12470 ( 
.A1(n_12133),
.A2(n_1633),
.B(n_1634),
.Y(n_12470)
);

AOI22xp33_ASAP7_75t_L g12471 ( 
.A1(n_12116),
.A2(n_1635),
.B1(n_1633),
.B2(n_1634),
.Y(n_12471)
);

INVx2_ASAP7_75t_L g12472 ( 
.A(n_12054),
.Y(n_12472)
);

INVx1_ASAP7_75t_L g12473 ( 
.A(n_12166),
.Y(n_12473)
);

CKINVDCx20_ASAP7_75t_R g12474 ( 
.A(n_11925),
.Y(n_12474)
);

OAI21x1_ASAP7_75t_L g12475 ( 
.A1(n_12126),
.A2(n_1635),
.B(n_1636),
.Y(n_12475)
);

OAI21x1_ASAP7_75t_L g12476 ( 
.A1(n_12073),
.A2(n_1637),
.B(n_1638),
.Y(n_12476)
);

OAI22xp5_ASAP7_75t_SL g12477 ( 
.A1(n_12161),
.A2(n_1639),
.B1(n_1637),
.B2(n_1638),
.Y(n_12477)
);

AO21x2_ASAP7_75t_L g12478 ( 
.A1(n_12005),
.A2(n_1639),
.B(n_1640),
.Y(n_12478)
);

AND2x2_ASAP7_75t_L g12479 ( 
.A(n_12093),
.B(n_1640),
.Y(n_12479)
);

OAI21xp5_ASAP7_75t_L g12480 ( 
.A1(n_12107),
.A2(n_1641),
.B(n_1642),
.Y(n_12480)
);

NAND2xp5_ASAP7_75t_L g12481 ( 
.A(n_12172),
.B(n_1641),
.Y(n_12481)
);

INVx1_ASAP7_75t_L g12482 ( 
.A(n_12086),
.Y(n_12482)
);

OA21x2_ASAP7_75t_L g12483 ( 
.A1(n_11972),
.A2(n_1642),
.B(n_1643),
.Y(n_12483)
);

INVx2_ASAP7_75t_L g12484 ( 
.A(n_12101),
.Y(n_12484)
);

INVx1_ASAP7_75t_L g12485 ( 
.A(n_12089),
.Y(n_12485)
);

NAND2xp5_ASAP7_75t_L g12486 ( 
.A(n_12147),
.B(n_1643),
.Y(n_12486)
);

INVx1_ASAP7_75t_L g12487 ( 
.A(n_12087),
.Y(n_12487)
);

OAI21x1_ASAP7_75t_L g12488 ( 
.A1(n_12134),
.A2(n_1644),
.B(n_1645),
.Y(n_12488)
);

AOI22xp33_ASAP7_75t_L g12489 ( 
.A1(n_12125),
.A2(n_1647),
.B1(n_1644),
.B2(n_1646),
.Y(n_12489)
);

BUFx6f_ASAP7_75t_L g12490 ( 
.A(n_11909),
.Y(n_12490)
);

BUFx6f_ASAP7_75t_L g12491 ( 
.A(n_11898),
.Y(n_12491)
);

OAI21xp5_ASAP7_75t_L g12492 ( 
.A1(n_11922),
.A2(n_1646),
.B(n_1648),
.Y(n_12492)
);

NAND2xp5_ASAP7_75t_L g12493 ( 
.A(n_12218),
.B(n_1648),
.Y(n_12493)
);

NOR2xp33_ASAP7_75t_L g12494 ( 
.A(n_11931),
.B(n_1649),
.Y(n_12494)
);

INVx3_ASAP7_75t_L g12495 ( 
.A(n_12008),
.Y(n_12495)
);

AO21x2_ASAP7_75t_L g12496 ( 
.A1(n_12042),
.A2(n_1650),
.B(n_1651),
.Y(n_12496)
);

AO31x2_ASAP7_75t_L g12497 ( 
.A1(n_12251),
.A2(n_1652),
.A3(n_1650),
.B(n_1651),
.Y(n_12497)
);

OAI21x1_ASAP7_75t_L g12498 ( 
.A1(n_12065),
.A2(n_1652),
.B(n_1653),
.Y(n_12498)
);

INVx2_ASAP7_75t_L g12499 ( 
.A(n_11985),
.Y(n_12499)
);

BUFx8_ASAP7_75t_L g12500 ( 
.A(n_12018),
.Y(n_12500)
);

BUFx2_ASAP7_75t_SL g12501 ( 
.A(n_11963),
.Y(n_12501)
);

O2A1O1Ixp5_ASAP7_75t_L g12502 ( 
.A1(n_12175),
.A2(n_11969),
.B(n_12203),
.C(n_12236),
.Y(n_12502)
);

NAND2xp5_ASAP7_75t_L g12503 ( 
.A(n_12194),
.B(n_1653),
.Y(n_12503)
);

BUFx12f_ASAP7_75t_L g12504 ( 
.A(n_12232),
.Y(n_12504)
);

AO31x2_ASAP7_75t_L g12505 ( 
.A1(n_12197),
.A2(n_1656),
.A3(n_1654),
.B(n_1655),
.Y(n_12505)
);

INVx1_ASAP7_75t_L g12506 ( 
.A(n_12111),
.Y(n_12506)
);

OR2x6_ASAP7_75t_L g12507 ( 
.A(n_11923),
.B(n_1654),
.Y(n_12507)
);

NAND2x1p5_ASAP7_75t_L g12508 ( 
.A(n_11897),
.B(n_1655),
.Y(n_12508)
);

AOI22xp33_ASAP7_75t_L g12509 ( 
.A1(n_12195),
.A2(n_1660),
.B1(n_1658),
.B2(n_1659),
.Y(n_12509)
);

OAI21xp5_ASAP7_75t_L g12510 ( 
.A1(n_11865),
.A2(n_1658),
.B(n_1659),
.Y(n_12510)
);

OAI22xp33_ASAP7_75t_L g12511 ( 
.A1(n_12121),
.A2(n_1662),
.B1(n_1660),
.B2(n_1661),
.Y(n_12511)
);

OAI21x1_ASAP7_75t_L g12512 ( 
.A1(n_12023),
.A2(n_1661),
.B(n_1663),
.Y(n_12512)
);

NOR2xp33_ASAP7_75t_L g12513 ( 
.A(n_12004),
.B(n_1664),
.Y(n_12513)
);

AO31x2_ASAP7_75t_L g12514 ( 
.A1(n_12040),
.A2(n_1666),
.A3(n_1664),
.B(n_1665),
.Y(n_12514)
);

AOI22xp33_ASAP7_75t_L g12515 ( 
.A1(n_12238),
.A2(n_1668),
.B1(n_1666),
.B2(n_1667),
.Y(n_12515)
);

OAI21x1_ASAP7_75t_L g12516 ( 
.A1(n_12025),
.A2(n_1667),
.B(n_1669),
.Y(n_12516)
);

OAI21xp5_ASAP7_75t_L g12517 ( 
.A1(n_12044),
.A2(n_1669),
.B(n_1670),
.Y(n_12517)
);

INVx2_ASAP7_75t_L g12518 ( 
.A(n_12104),
.Y(n_12518)
);

NOR2xp33_ASAP7_75t_L g12519 ( 
.A(n_12240),
.B(n_1670),
.Y(n_12519)
);

AND2x4_ASAP7_75t_L g12520 ( 
.A(n_11911),
.B(n_12031),
.Y(n_12520)
);

INVx1_ASAP7_75t_L g12521 ( 
.A(n_12181),
.Y(n_12521)
);

BUFx2_ASAP7_75t_SL g12522 ( 
.A(n_12029),
.Y(n_12522)
);

A2O1A1Ixp33_ASAP7_75t_L g12523 ( 
.A1(n_12242),
.A2(n_1673),
.B(n_1671),
.C(n_1672),
.Y(n_12523)
);

OAI21x1_ASAP7_75t_L g12524 ( 
.A1(n_12048),
.A2(n_1671),
.B(n_1672),
.Y(n_12524)
);

OAI21x1_ASAP7_75t_L g12525 ( 
.A1(n_12108),
.A2(n_1674),
.B(n_1675),
.Y(n_12525)
);

NOR2xp67_ASAP7_75t_L g12526 ( 
.A(n_12029),
.B(n_12013),
.Y(n_12526)
);

OAI21x1_ASAP7_75t_L g12527 ( 
.A1(n_12289),
.A2(n_1675),
.B(n_1676),
.Y(n_12527)
);

OA21x2_ASAP7_75t_L g12528 ( 
.A1(n_12131),
.A2(n_1676),
.B(n_1677),
.Y(n_12528)
);

INVx2_ASAP7_75t_SL g12529 ( 
.A(n_12059),
.Y(n_12529)
);

BUFx8_ASAP7_75t_L g12530 ( 
.A(n_12110),
.Y(n_12530)
);

INVx2_ASAP7_75t_L g12531 ( 
.A(n_11982),
.Y(n_12531)
);

OR2x6_ASAP7_75t_L g12532 ( 
.A(n_12097),
.B(n_1677),
.Y(n_12532)
);

INVx1_ASAP7_75t_L g12533 ( 
.A(n_12144),
.Y(n_12533)
);

OA21x2_ASAP7_75t_L g12534 ( 
.A1(n_12090),
.A2(n_1678),
.B(n_1679),
.Y(n_12534)
);

AOI22xp33_ASAP7_75t_L g12535 ( 
.A1(n_12182),
.A2(n_1680),
.B1(n_1678),
.B2(n_1679),
.Y(n_12535)
);

O2A1O1Ixp33_ASAP7_75t_SL g12536 ( 
.A1(n_11893),
.A2(n_1683),
.B(n_1681),
.C(n_1682),
.Y(n_12536)
);

AOI21xp5_ASAP7_75t_L g12537 ( 
.A1(n_12138),
.A2(n_12224),
.B(n_12216),
.Y(n_12537)
);

AO31x2_ASAP7_75t_L g12538 ( 
.A1(n_12022),
.A2(n_1684),
.A3(n_1681),
.B(n_1682),
.Y(n_12538)
);

INVx2_ASAP7_75t_L g12539 ( 
.A(n_12257),
.Y(n_12539)
);

NAND2xp5_ASAP7_75t_L g12540 ( 
.A(n_12244),
.B(n_1684),
.Y(n_12540)
);

OAI21x1_ASAP7_75t_L g12541 ( 
.A1(n_12075),
.A2(n_1686),
.B(n_1687),
.Y(n_12541)
);

OAI21x1_ASAP7_75t_L g12542 ( 
.A1(n_12000),
.A2(n_1686),
.B(n_1688),
.Y(n_12542)
);

BUFx3_ASAP7_75t_L g12543 ( 
.A(n_12016),
.Y(n_12543)
);

AOI22xp33_ASAP7_75t_L g12544 ( 
.A1(n_12219),
.A2(n_12243),
.B1(n_12252),
.B2(n_12205),
.Y(n_12544)
);

OAI21x1_ASAP7_75t_SL g12545 ( 
.A1(n_12080),
.A2(n_1689),
.B(n_1690),
.Y(n_12545)
);

BUFx12f_ASAP7_75t_L g12546 ( 
.A(n_12264),
.Y(n_12546)
);

NAND2xp5_ASAP7_75t_L g12547 ( 
.A(n_12150),
.B(n_1689),
.Y(n_12547)
);

OAI21x1_ASAP7_75t_L g12548 ( 
.A1(n_12057),
.A2(n_12098),
.B(n_12083),
.Y(n_12548)
);

OR2x2_ASAP7_75t_L g12549 ( 
.A(n_12155),
.B(n_1691),
.Y(n_12549)
);

BUFx3_ASAP7_75t_L g12550 ( 
.A(n_11933),
.Y(n_12550)
);

NAND2xp33_ASAP7_75t_SL g12551 ( 
.A(n_11872),
.B(n_12178),
.Y(n_12551)
);

INVx1_ASAP7_75t_L g12552 ( 
.A(n_11906),
.Y(n_12552)
);

AOI21xp5_ASAP7_75t_L g12553 ( 
.A1(n_12207),
.A2(n_1691),
.B(n_1692),
.Y(n_12553)
);

OAI21x1_ASAP7_75t_L g12554 ( 
.A1(n_12262),
.A2(n_1693),
.B(n_1694),
.Y(n_12554)
);

OAI21x1_ASAP7_75t_L g12555 ( 
.A1(n_12119),
.A2(n_1693),
.B(n_1695),
.Y(n_12555)
);

OAI21x1_ASAP7_75t_L g12556 ( 
.A1(n_12123),
.A2(n_1695),
.B(n_1696),
.Y(n_12556)
);

BUFx6f_ASAP7_75t_SL g12557 ( 
.A(n_11862),
.Y(n_12557)
);

INVx1_ASAP7_75t_L g12558 ( 
.A(n_12140),
.Y(n_12558)
);

NAND2xp5_ASAP7_75t_L g12559 ( 
.A(n_12270),
.B(n_1696),
.Y(n_12559)
);

INVx1_ASAP7_75t_L g12560 ( 
.A(n_11860),
.Y(n_12560)
);

NAND2xp5_ASAP7_75t_L g12561 ( 
.A(n_12282),
.B(n_1697),
.Y(n_12561)
);

OAI21x1_ASAP7_75t_L g12562 ( 
.A1(n_12128),
.A2(n_1697),
.B(n_1698),
.Y(n_12562)
);

OAI21x1_ASAP7_75t_L g12563 ( 
.A1(n_12136),
.A2(n_1698),
.B(n_1699),
.Y(n_12563)
);

INVx2_ASAP7_75t_SL g12564 ( 
.A(n_11947),
.Y(n_12564)
);

INVx2_ASAP7_75t_L g12565 ( 
.A(n_12257),
.Y(n_12565)
);

NAND2xp5_ASAP7_75t_L g12566 ( 
.A(n_12284),
.B(n_1699),
.Y(n_12566)
);

HB1xp67_ASAP7_75t_L g12567 ( 
.A(n_12143),
.Y(n_12567)
);

AOI22xp5_ASAP7_75t_L g12568 ( 
.A1(n_11983),
.A2(n_11975),
.B1(n_12287),
.B2(n_12034),
.Y(n_12568)
);

BUFx3_ASAP7_75t_L g12569 ( 
.A(n_11976),
.Y(n_12569)
);

INVx1_ASAP7_75t_L g12570 ( 
.A(n_12170),
.Y(n_12570)
);

INVx2_ASAP7_75t_SL g12571 ( 
.A(n_12007),
.Y(n_12571)
);

BUFx2_ASAP7_75t_L g12572 ( 
.A(n_12135),
.Y(n_12572)
);

INVx1_ASAP7_75t_L g12573 ( 
.A(n_12067),
.Y(n_12573)
);

AND2x4_ASAP7_75t_L g12574 ( 
.A(n_11961),
.B(n_1700),
.Y(n_12574)
);

BUFx2_ASAP7_75t_L g12575 ( 
.A(n_12041),
.Y(n_12575)
);

INVx1_ASAP7_75t_L g12576 ( 
.A(n_12026),
.Y(n_12576)
);

AND2x4_ASAP7_75t_L g12577 ( 
.A(n_11981),
.B(n_1700),
.Y(n_12577)
);

OAI21x1_ASAP7_75t_L g12578 ( 
.A1(n_12139),
.A2(n_1701),
.B(n_1702),
.Y(n_12578)
);

OAI21x1_ASAP7_75t_SL g12579 ( 
.A1(n_11934),
.A2(n_1701),
.B(n_1702),
.Y(n_12579)
);

BUFx2_ASAP7_75t_L g12580 ( 
.A(n_12109),
.Y(n_12580)
);

AOI21xp33_ASAP7_75t_L g12581 ( 
.A1(n_12071),
.A2(n_11967),
.B(n_12169),
.Y(n_12581)
);

INVx1_ASAP7_75t_L g12582 ( 
.A(n_11987),
.Y(n_12582)
);

NAND2xp5_ASAP7_75t_L g12583 ( 
.A(n_12253),
.B(n_1703),
.Y(n_12583)
);

CKINVDCx6p67_ASAP7_75t_R g12584 ( 
.A(n_12060),
.Y(n_12584)
);

NOR2xp33_ASAP7_75t_L g12585 ( 
.A(n_11966),
.B(n_1704),
.Y(n_12585)
);

BUFx6f_ASAP7_75t_L g12586 ( 
.A(n_11874),
.Y(n_12586)
);

AO31x2_ASAP7_75t_L g12587 ( 
.A1(n_12024),
.A2(n_1706),
.A3(n_1704),
.B(n_1705),
.Y(n_12587)
);

OAI21xp5_ASAP7_75t_L g12588 ( 
.A1(n_12196),
.A2(n_1705),
.B(n_1707),
.Y(n_12588)
);

AOI22x1_ASAP7_75t_L g12589 ( 
.A1(n_12178),
.A2(n_12058),
.B1(n_12062),
.B2(n_12046),
.Y(n_12589)
);

OAI21x1_ASAP7_75t_L g12590 ( 
.A1(n_12145),
.A2(n_1707),
.B(n_1708),
.Y(n_12590)
);

INVx1_ASAP7_75t_L g12591 ( 
.A(n_11997),
.Y(n_12591)
);

NAND2xp5_ASAP7_75t_L g12592 ( 
.A(n_12208),
.B(n_12153),
.Y(n_12592)
);

INVx2_ASAP7_75t_SL g12593 ( 
.A(n_11879),
.Y(n_12593)
);

BUFx2_ASAP7_75t_L g12594 ( 
.A(n_12149),
.Y(n_12594)
);

INVx2_ASAP7_75t_L g12595 ( 
.A(n_12174),
.Y(n_12595)
);

NAND2xp5_ASAP7_75t_SL g12596 ( 
.A(n_11908),
.B(n_1708),
.Y(n_12596)
);

CKINVDCx5p33_ASAP7_75t_R g12597 ( 
.A(n_11977),
.Y(n_12597)
);

INVx1_ASAP7_75t_L g12598 ( 
.A(n_11868),
.Y(n_12598)
);

AO22x2_ASAP7_75t_L g12599 ( 
.A1(n_11945),
.A2(n_1711),
.B1(n_1709),
.B2(n_1710),
.Y(n_12599)
);

OAI21x1_ASAP7_75t_L g12600 ( 
.A1(n_12156),
.A2(n_1709),
.B(n_1710),
.Y(n_12600)
);

INVx1_ASAP7_75t_L g12601 ( 
.A(n_12094),
.Y(n_12601)
);

OAI21x1_ASAP7_75t_L g12602 ( 
.A1(n_12162),
.A2(n_1711),
.B(n_1712),
.Y(n_12602)
);

INVx1_ASAP7_75t_L g12603 ( 
.A(n_12187),
.Y(n_12603)
);

OAI211xp5_ASAP7_75t_SL g12604 ( 
.A1(n_12095),
.A2(n_1715),
.B(n_1713),
.C(n_1714),
.Y(n_12604)
);

AO21x1_ASAP7_75t_L g12605 ( 
.A1(n_12152),
.A2(n_1713),
.B(n_1714),
.Y(n_12605)
);

INVx1_ASAP7_75t_L g12606 ( 
.A(n_12096),
.Y(n_12606)
);

CKINVDCx5p33_ASAP7_75t_R g12607 ( 
.A(n_12035),
.Y(n_12607)
);

HB1xp67_ASAP7_75t_L g12608 ( 
.A(n_11951),
.Y(n_12608)
);

O2A1O1Ixp5_ASAP7_75t_L g12609 ( 
.A1(n_12113),
.A2(n_1717),
.B(n_1715),
.C(n_1716),
.Y(n_12609)
);

CKINVDCx6p67_ASAP7_75t_R g12610 ( 
.A(n_12032),
.Y(n_12610)
);

AOI21xp5_ASAP7_75t_L g12611 ( 
.A1(n_12118),
.A2(n_12223),
.B(n_12272),
.Y(n_12611)
);

INVx2_ASAP7_75t_L g12612 ( 
.A(n_12052),
.Y(n_12612)
);

OAI21x1_ASAP7_75t_SL g12613 ( 
.A1(n_11986),
.A2(n_1716),
.B(n_1717),
.Y(n_12613)
);

AND2x4_ASAP7_75t_L g12614 ( 
.A(n_11991),
.B(n_1718),
.Y(n_12614)
);

AOI21xp5_ASAP7_75t_L g12615 ( 
.A1(n_12258),
.A2(n_1718),
.B(n_1719),
.Y(n_12615)
);

INVxp67_ASAP7_75t_SL g12616 ( 
.A(n_12245),
.Y(n_12616)
);

CKINVDCx5p33_ASAP7_75t_R g12617 ( 
.A(n_12102),
.Y(n_12617)
);

OAI22xp33_ASAP7_75t_L g12618 ( 
.A1(n_12245),
.A2(n_1722),
.B1(n_1719),
.B2(n_1721),
.Y(n_12618)
);

NOR2xp67_ASAP7_75t_L g12619 ( 
.A(n_12259),
.B(n_1721),
.Y(n_12619)
);

NOR2x1_ASAP7_75t_SL g12620 ( 
.A(n_12165),
.B(n_1722),
.Y(n_12620)
);

NAND3xp33_ASAP7_75t_L g12621 ( 
.A(n_12158),
.B(n_12198),
.C(n_12250),
.Y(n_12621)
);

OAI21x1_ASAP7_75t_L g12622 ( 
.A1(n_12168),
.A2(n_1723),
.B(n_1724),
.Y(n_12622)
);

INVx1_ASAP7_75t_L g12623 ( 
.A(n_12030),
.Y(n_12623)
);

NOR2x1_ASAP7_75t_L g12624 ( 
.A(n_12267),
.B(n_1723),
.Y(n_12624)
);

AO21x2_ASAP7_75t_L g12625 ( 
.A1(n_12171),
.A2(n_1724),
.B(n_1725),
.Y(n_12625)
);

OA21x2_ASAP7_75t_L g12626 ( 
.A1(n_11973),
.A2(n_1725),
.B(n_1726),
.Y(n_12626)
);

AND2x4_ASAP7_75t_L g12627 ( 
.A(n_11995),
.B(n_1727),
.Y(n_12627)
);

CKINVDCx5p33_ASAP7_75t_R g12628 ( 
.A(n_11874),
.Y(n_12628)
);

AND2x4_ASAP7_75t_L g12629 ( 
.A(n_12015),
.B(n_1728),
.Y(n_12629)
);

BUFx3_ASAP7_75t_L g12630 ( 
.A(n_12047),
.Y(n_12630)
);

INVx2_ASAP7_75t_L g12631 ( 
.A(n_12052),
.Y(n_12631)
);

OAI21x1_ASAP7_75t_L g12632 ( 
.A1(n_12173),
.A2(n_1728),
.B(n_1729),
.Y(n_12632)
);

HB1xp67_ASAP7_75t_L g12633 ( 
.A(n_12200),
.Y(n_12633)
);

NOR2xp33_ASAP7_75t_L g12634 ( 
.A(n_12285),
.B(n_1729),
.Y(n_12634)
);

NAND3xp33_ASAP7_75t_SL g12635 ( 
.A(n_12248),
.B(n_1730),
.C(n_1731),
.Y(n_12635)
);

AO31x2_ASAP7_75t_L g12636 ( 
.A1(n_12039),
.A2(n_1732),
.A3(n_1730),
.B(n_1731),
.Y(n_12636)
);

OAI21x1_ASAP7_75t_L g12637 ( 
.A1(n_12209),
.A2(n_1733),
.B(n_1734),
.Y(n_12637)
);

AOI21x1_ASAP7_75t_L g12638 ( 
.A1(n_12199),
.A2(n_1733),
.B(n_1734),
.Y(n_12638)
);

OAI22xp5_ASAP7_75t_L g12639 ( 
.A1(n_12288),
.A2(n_1737),
.B1(n_1735),
.B2(n_1736),
.Y(n_12639)
);

AOI22xp33_ASAP7_75t_L g12640 ( 
.A1(n_12274),
.A2(n_1739),
.B1(n_1737),
.B2(n_1738),
.Y(n_12640)
);

INVx1_ASAP7_75t_L g12641 ( 
.A(n_12212),
.Y(n_12641)
);

INVx2_ASAP7_75t_L g12642 ( 
.A(n_12050),
.Y(n_12642)
);

INVx1_ASAP7_75t_L g12643 ( 
.A(n_12213),
.Y(n_12643)
);

AND2x2_ASAP7_75t_L g12644 ( 
.A(n_12020),
.B(n_1739),
.Y(n_12644)
);

NAND2x1p5_ASAP7_75t_L g12645 ( 
.A(n_11880),
.B(n_1741),
.Y(n_12645)
);

NAND2xp5_ASAP7_75t_L g12646 ( 
.A(n_12151),
.B(n_1741),
.Y(n_12646)
);

INVx2_ASAP7_75t_L g12647 ( 
.A(n_11880),
.Y(n_12647)
);

INVx3_ASAP7_75t_L g12648 ( 
.A(n_11901),
.Y(n_12648)
);

INVx3_ASAP7_75t_L g12649 ( 
.A(n_11901),
.Y(n_12649)
);

AO31x2_ASAP7_75t_L g12650 ( 
.A1(n_12226),
.A2(n_1745),
.A3(n_1742),
.B(n_1743),
.Y(n_12650)
);

INVx1_ASAP7_75t_L g12651 ( 
.A(n_12227),
.Y(n_12651)
);

AO31x2_ASAP7_75t_L g12652 ( 
.A1(n_12228),
.A2(n_1746),
.A3(n_1743),
.B(n_1745),
.Y(n_12652)
);

INVx1_ASAP7_75t_L g12653 ( 
.A(n_12231),
.Y(n_12653)
);

INVx1_ASAP7_75t_L g12654 ( 
.A(n_12237),
.Y(n_12654)
);

OAI21xp5_ASAP7_75t_L g12655 ( 
.A1(n_12239),
.A2(n_1746),
.B(n_1747),
.Y(n_12655)
);

INVx2_ASAP7_75t_L g12656 ( 
.A(n_11940),
.Y(n_12656)
);

AOI221xp5_ASAP7_75t_L g12657 ( 
.A1(n_12281),
.A2(n_1749),
.B1(n_1747),
.B2(n_1748),
.C(n_1750),
.Y(n_12657)
);

OAI21x1_ASAP7_75t_L g12658 ( 
.A1(n_12254),
.A2(n_1748),
.B(n_1750),
.Y(n_12658)
);

OAI21x1_ASAP7_75t_L g12659 ( 
.A1(n_12256),
.A2(n_1751),
.B(n_1752),
.Y(n_12659)
);

OAI22xp5_ASAP7_75t_L g12660 ( 
.A1(n_12265),
.A2(n_1753),
.B1(n_1751),
.B2(n_1752),
.Y(n_12660)
);

AND2x2_ASAP7_75t_L g12661 ( 
.A(n_11940),
.B(n_1753),
.Y(n_12661)
);

OAI21x1_ASAP7_75t_L g12662 ( 
.A1(n_12261),
.A2(n_1754),
.B(n_1755),
.Y(n_12662)
);

AND2x4_ASAP7_75t_L g12663 ( 
.A(n_12630),
.B(n_11955),
.Y(n_12663)
);

OAI21x1_ASAP7_75t_L g12664 ( 
.A1(n_12318),
.A2(n_12277),
.B(n_12273),
.Y(n_12664)
);

INVxp33_ASAP7_75t_L g12665 ( 
.A(n_12490),
.Y(n_12665)
);

OA21x2_ASAP7_75t_L g12666 ( 
.A1(n_12405),
.A2(n_12286),
.B(n_12191),
.Y(n_12666)
);

INVx1_ASAP7_75t_L g12667 ( 
.A(n_12384),
.Y(n_12667)
);

NAND2xp5_ASAP7_75t_L g12668 ( 
.A(n_12611),
.B(n_12064),
.Y(n_12668)
);

A2O1A1Ixp33_ASAP7_75t_L g12669 ( 
.A1(n_12331),
.A2(n_12115),
.B(n_12085),
.C(n_11958),
.Y(n_12669)
);

OAI21xp5_ASAP7_75t_L g12670 ( 
.A1(n_12374),
.A2(n_12106),
.B(n_11958),
.Y(n_12670)
);

INVx1_ASAP7_75t_SL g12671 ( 
.A(n_12522),
.Y(n_12671)
);

AOI21xp5_ASAP7_75t_L g12672 ( 
.A1(n_12298),
.A2(n_11971),
.B(n_11955),
.Y(n_12672)
);

INVx1_ASAP7_75t_L g12673 ( 
.A(n_12290),
.Y(n_12673)
);

INVx2_ASAP7_75t_SL g12674 ( 
.A(n_12500),
.Y(n_12674)
);

OAI21xp5_ASAP7_75t_L g12675 ( 
.A1(n_12337),
.A2(n_11999),
.B(n_11971),
.Y(n_12675)
);

INVx1_ASAP7_75t_L g12676 ( 
.A(n_12291),
.Y(n_12676)
);

AND2x2_ASAP7_75t_L g12677 ( 
.A(n_12427),
.B(n_11999),
.Y(n_12677)
);

OR2x6_ASAP7_75t_L g12678 ( 
.A(n_12532),
.B(n_12045),
.Y(n_12678)
);

OAI21xp5_ASAP7_75t_L g12679 ( 
.A1(n_12537),
.A2(n_12502),
.B(n_12568),
.Y(n_12679)
);

OA21x2_ASAP7_75t_L g12680 ( 
.A1(n_12413),
.A2(n_12045),
.B(n_1754),
.Y(n_12680)
);

NAND2xp5_ASAP7_75t_L g12681 ( 
.A(n_12379),
.B(n_1755),
.Y(n_12681)
);

OAI21x1_ASAP7_75t_L g12682 ( 
.A1(n_12336),
.A2(n_12400),
.B(n_12344),
.Y(n_12682)
);

INVx1_ASAP7_75t_L g12683 ( 
.A(n_12297),
.Y(n_12683)
);

INVx1_ASAP7_75t_L g12684 ( 
.A(n_12324),
.Y(n_12684)
);

INVx1_ASAP7_75t_L g12685 ( 
.A(n_12345),
.Y(n_12685)
);

INVx1_ASAP7_75t_L g12686 ( 
.A(n_12348),
.Y(n_12686)
);

OAI21x1_ASAP7_75t_L g12687 ( 
.A1(n_12397),
.A2(n_1756),
.B(n_1757),
.Y(n_12687)
);

OAI22xp33_ASAP7_75t_L g12688 ( 
.A1(n_12467),
.A2(n_1758),
.B1(n_1756),
.B2(n_1757),
.Y(n_12688)
);

AOI21xp5_ASAP7_75t_L g12689 ( 
.A1(n_12335),
.A2(n_12339),
.B(n_12295),
.Y(n_12689)
);

A2O1A1Ixp33_ASAP7_75t_L g12690 ( 
.A1(n_12394),
.A2(n_1760),
.B(n_1758),
.C(n_1759),
.Y(n_12690)
);

INVx2_ASAP7_75t_SL g12691 ( 
.A(n_12442),
.Y(n_12691)
);

OA21x2_ASAP7_75t_L g12692 ( 
.A1(n_12460),
.A2(n_1759),
.B(n_1761),
.Y(n_12692)
);

AO21x2_ASAP7_75t_L g12693 ( 
.A1(n_12608),
.A2(n_12423),
.B(n_12582),
.Y(n_12693)
);

INVx1_ASAP7_75t_SL g12694 ( 
.A(n_12367),
.Y(n_12694)
);

NAND2xp5_ASAP7_75t_L g12695 ( 
.A(n_12316),
.B(n_1761),
.Y(n_12695)
);

HB1xp67_ASAP7_75t_L g12696 ( 
.A(n_12402),
.Y(n_12696)
);

CKINVDCx5p33_ASAP7_75t_R g12697 ( 
.A(n_12305),
.Y(n_12697)
);

BUFx12f_ASAP7_75t_L g12698 ( 
.A(n_12358),
.Y(n_12698)
);

INVx1_ASAP7_75t_L g12699 ( 
.A(n_12352),
.Y(n_12699)
);

BUFx2_ASAP7_75t_L g12700 ( 
.A(n_12610),
.Y(n_12700)
);

NAND2x1p5_ASAP7_75t_L g12701 ( 
.A(n_12572),
.B(n_1762),
.Y(n_12701)
);

NAND2xp5_ASAP7_75t_L g12702 ( 
.A(n_12428),
.B(n_1762),
.Y(n_12702)
);

INVx2_ASAP7_75t_L g12703 ( 
.A(n_12431),
.Y(n_12703)
);

AOI21xp5_ASAP7_75t_L g12704 ( 
.A1(n_12313),
.A2(n_1763),
.B(n_1764),
.Y(n_12704)
);

HB1xp67_ASAP7_75t_L g12705 ( 
.A(n_12633),
.Y(n_12705)
);

NAND2xp5_ASAP7_75t_L g12706 ( 
.A(n_12463),
.B(n_1763),
.Y(n_12706)
);

AOI21xp5_ASAP7_75t_L g12707 ( 
.A1(n_12347),
.A2(n_1764),
.B(n_1765),
.Y(n_12707)
);

AO21x2_ASAP7_75t_L g12708 ( 
.A1(n_12591),
.A2(n_1765),
.B(n_1766),
.Y(n_12708)
);

NAND2xp5_ASAP7_75t_L g12709 ( 
.A(n_12473),
.B(n_1766),
.Y(n_12709)
);

OAI21x1_ASAP7_75t_L g12710 ( 
.A1(n_12389),
.A2(n_1767),
.B(n_1768),
.Y(n_12710)
);

OR2x2_ASAP7_75t_L g12711 ( 
.A(n_12422),
.B(n_1767),
.Y(n_12711)
);

AO21x2_ASAP7_75t_L g12712 ( 
.A1(n_12576),
.A2(n_1768),
.B(n_1769),
.Y(n_12712)
);

AOI21xp5_ASAP7_75t_L g12713 ( 
.A1(n_12388),
.A2(n_1769),
.B(n_1770),
.Y(n_12713)
);

OA21x2_ASAP7_75t_L g12714 ( 
.A1(n_12411),
.A2(n_1770),
.B(n_1771),
.Y(n_12714)
);

INVx3_ASAP7_75t_L g12715 ( 
.A(n_12442),
.Y(n_12715)
);

OAI21xp33_ASAP7_75t_L g12716 ( 
.A1(n_12404),
.A2(n_12450),
.B(n_12544),
.Y(n_12716)
);

AND2x2_ASAP7_75t_L g12717 ( 
.A(n_12325),
.B(n_1771),
.Y(n_12717)
);

AOI21xp5_ASAP7_75t_L g12718 ( 
.A1(n_12368),
.A2(n_1772),
.B(n_1773),
.Y(n_12718)
);

NAND2xp5_ASAP7_75t_SL g12719 ( 
.A(n_12551),
.B(n_12380),
.Y(n_12719)
);

OAI21xp5_ASAP7_75t_L g12720 ( 
.A1(n_12438),
.A2(n_1773),
.B(n_1774),
.Y(n_12720)
);

OAI21x1_ASAP7_75t_L g12721 ( 
.A1(n_12436),
.A2(n_1775),
.B(n_1776),
.Y(n_12721)
);

INVx2_ASAP7_75t_L g12722 ( 
.A(n_12382),
.Y(n_12722)
);

INVx2_ASAP7_75t_L g12723 ( 
.A(n_12393),
.Y(n_12723)
);

OA21x2_ASAP7_75t_L g12724 ( 
.A1(n_12499),
.A2(n_1775),
.B(n_1776),
.Y(n_12724)
);

NAND2xp5_ASAP7_75t_L g12725 ( 
.A(n_12573),
.B(n_1777),
.Y(n_12725)
);

INVx1_ASAP7_75t_L g12726 ( 
.A(n_12356),
.Y(n_12726)
);

NAND2xp5_ASAP7_75t_L g12727 ( 
.A(n_12462),
.B(n_1777),
.Y(n_12727)
);

AOI21xp5_ASAP7_75t_L g12728 ( 
.A1(n_12350),
.A2(n_1778),
.B(n_1779),
.Y(n_12728)
);

INVx2_ASAP7_75t_L g12729 ( 
.A(n_12310),
.Y(n_12729)
);

NAND2xp5_ASAP7_75t_L g12730 ( 
.A(n_12570),
.B(n_1778),
.Y(n_12730)
);

OAI21x1_ASAP7_75t_L g12731 ( 
.A1(n_12435),
.A2(n_1779),
.B(n_1780),
.Y(n_12731)
);

INVx2_ASAP7_75t_L g12732 ( 
.A(n_12455),
.Y(n_12732)
);

OA21x2_ASAP7_75t_L g12733 ( 
.A1(n_12301),
.A2(n_1781),
.B(n_1782),
.Y(n_12733)
);

INVx2_ASAP7_75t_L g12734 ( 
.A(n_12465),
.Y(n_12734)
);

AO21x2_ASAP7_75t_L g12735 ( 
.A1(n_12363),
.A2(n_1781),
.B(n_1782),
.Y(n_12735)
);

OAI21x1_ASAP7_75t_L g12736 ( 
.A1(n_12440),
.A2(n_1783),
.B(n_1784),
.Y(n_12736)
);

NAND2xp5_ASAP7_75t_L g12737 ( 
.A(n_12392),
.B(n_1783),
.Y(n_12737)
);

INVx2_ASAP7_75t_L g12738 ( 
.A(n_12484),
.Y(n_12738)
);

OR2x6_ASAP7_75t_L g12739 ( 
.A(n_12532),
.B(n_1785),
.Y(n_12739)
);

AOI21xp5_ASAP7_75t_L g12740 ( 
.A1(n_12326),
.A2(n_1785),
.B(n_1786),
.Y(n_12740)
);

OA21x2_ASAP7_75t_L g12741 ( 
.A1(n_12487),
.A2(n_1786),
.B(n_1787),
.Y(n_12741)
);

AOI22x1_ASAP7_75t_L g12742 ( 
.A1(n_12424),
.A2(n_1789),
.B1(n_1787),
.B2(n_1788),
.Y(n_12742)
);

NAND2xp5_ASAP7_75t_L g12743 ( 
.A(n_12606),
.B(n_12444),
.Y(n_12743)
);

INVx2_ASAP7_75t_L g12744 ( 
.A(n_12441),
.Y(n_12744)
);

AND2x4_ASAP7_75t_L g12745 ( 
.A(n_12526),
.B(n_1788),
.Y(n_12745)
);

AO31x2_ASAP7_75t_L g12746 ( 
.A1(n_12605),
.A2(n_1791),
.A3(n_1789),
.B(n_1790),
.Y(n_12746)
);

BUFx3_ASAP7_75t_L g12747 ( 
.A(n_12299),
.Y(n_12747)
);

OAI21x1_ASAP7_75t_SL g12748 ( 
.A1(n_12579),
.A2(n_1790),
.B(n_1791),
.Y(n_12748)
);

BUFx12f_ASAP7_75t_L g12749 ( 
.A(n_12504),
.Y(n_12749)
);

INVx1_ASAP7_75t_L g12750 ( 
.A(n_12386),
.Y(n_12750)
);

INVx1_ASAP7_75t_L g12751 ( 
.A(n_12390),
.Y(n_12751)
);

OR2x2_ASAP7_75t_L g12752 ( 
.A(n_12445),
.B(n_1792),
.Y(n_12752)
);

INVx1_ASAP7_75t_L g12753 ( 
.A(n_12408),
.Y(n_12753)
);

AOI221xp5_ASAP7_75t_L g12754 ( 
.A1(n_12396),
.A2(n_1795),
.B1(n_1793),
.B2(n_1794),
.C(n_1796),
.Y(n_12754)
);

NAND2xp5_ASAP7_75t_L g12755 ( 
.A(n_12323),
.B(n_1796),
.Y(n_12755)
);

NAND2xp5_ASAP7_75t_L g12756 ( 
.A(n_12353),
.B(n_1797),
.Y(n_12756)
);

BUFx8_ASAP7_75t_L g12757 ( 
.A(n_12490),
.Y(n_12757)
);

CKINVDCx5p33_ASAP7_75t_R g12758 ( 
.A(n_12458),
.Y(n_12758)
);

INVx3_ASAP7_75t_L g12759 ( 
.A(n_12491),
.Y(n_12759)
);

INVx1_ASAP7_75t_L g12760 ( 
.A(n_12412),
.Y(n_12760)
);

OA21x2_ASAP7_75t_L g12761 ( 
.A1(n_12292),
.A2(n_1797),
.B(n_1798),
.Y(n_12761)
);

OA21x2_ASAP7_75t_L g12762 ( 
.A1(n_12317),
.A2(n_1798),
.B(n_1799),
.Y(n_12762)
);

HB1xp67_ASAP7_75t_L g12763 ( 
.A(n_12433),
.Y(n_12763)
);

INVx1_ASAP7_75t_L g12764 ( 
.A(n_12417),
.Y(n_12764)
);

INVx2_ASAP7_75t_SL g12765 ( 
.A(n_12359),
.Y(n_12765)
);

OAI21x1_ASAP7_75t_L g12766 ( 
.A1(n_12443),
.A2(n_1799),
.B(n_1801),
.Y(n_12766)
);

CKINVDCx14_ASAP7_75t_R g12767 ( 
.A(n_12294),
.Y(n_12767)
);

AOI21xp5_ASAP7_75t_L g12768 ( 
.A1(n_12302),
.A2(n_1801),
.B(n_1802),
.Y(n_12768)
);

OAI21x1_ASAP7_75t_SL g12769 ( 
.A1(n_12466),
.A2(n_1802),
.B(n_1803),
.Y(n_12769)
);

INVx1_ASAP7_75t_L g12770 ( 
.A(n_12426),
.Y(n_12770)
);

BUFx5_ASAP7_75t_L g12771 ( 
.A(n_12550),
.Y(n_12771)
);

INVx1_ASAP7_75t_L g12772 ( 
.A(n_12437),
.Y(n_12772)
);

NAND2xp5_ASAP7_75t_L g12773 ( 
.A(n_12401),
.B(n_1803),
.Y(n_12773)
);

BUFx3_ASAP7_75t_L g12774 ( 
.A(n_12474),
.Y(n_12774)
);

INVx1_ASAP7_75t_L g12775 ( 
.A(n_12447),
.Y(n_12775)
);

OAI21x1_ASAP7_75t_L g12776 ( 
.A1(n_12434),
.A2(n_1804),
.B(n_1805),
.Y(n_12776)
);

INVx2_ASAP7_75t_L g12777 ( 
.A(n_12406),
.Y(n_12777)
);

NAND2xp5_ASAP7_75t_L g12778 ( 
.A(n_12377),
.B(n_1806),
.Y(n_12778)
);

OA21x2_ASAP7_75t_L g12779 ( 
.A1(n_12616),
.A2(n_1806),
.B(n_1807),
.Y(n_12779)
);

INVx2_ASAP7_75t_L g12780 ( 
.A(n_12329),
.Y(n_12780)
);

AOI21xp5_ASAP7_75t_L g12781 ( 
.A1(n_12327),
.A2(n_1807),
.B(n_1809),
.Y(n_12781)
);

NAND2xp5_ASAP7_75t_L g12782 ( 
.A(n_12432),
.B(n_1809),
.Y(n_12782)
);

INVx3_ASAP7_75t_L g12783 ( 
.A(n_12491),
.Y(n_12783)
);

OAI21x1_ASAP7_75t_L g12784 ( 
.A1(n_12354),
.A2(n_1810),
.B(n_1811),
.Y(n_12784)
);

INVx1_ASAP7_75t_L g12785 ( 
.A(n_12378),
.Y(n_12785)
);

INVx1_ASAP7_75t_L g12786 ( 
.A(n_12482),
.Y(n_12786)
);

INVx2_ASAP7_75t_L g12787 ( 
.A(n_12332),
.Y(n_12787)
);

OAI21x1_ASAP7_75t_L g12788 ( 
.A1(n_12333),
.A2(n_1810),
.B(n_1811),
.Y(n_12788)
);

AOI21xp5_ASAP7_75t_L g12789 ( 
.A1(n_12419),
.A2(n_1813),
.B(n_1814),
.Y(n_12789)
);

NAND2xp5_ASAP7_75t_L g12790 ( 
.A(n_12641),
.B(n_1813),
.Y(n_12790)
);

INVx2_ASAP7_75t_L g12791 ( 
.A(n_12341),
.Y(n_12791)
);

INVx1_ASAP7_75t_L g12792 ( 
.A(n_12485),
.Y(n_12792)
);

INVx1_ASAP7_75t_L g12793 ( 
.A(n_12375),
.Y(n_12793)
);

INVx1_ASAP7_75t_L g12794 ( 
.A(n_12376),
.Y(n_12794)
);

OAI21xp5_ASAP7_75t_L g12795 ( 
.A1(n_12510),
.A2(n_12360),
.B(n_12492),
.Y(n_12795)
);

OAI21x1_ASAP7_75t_L g12796 ( 
.A1(n_12330),
.A2(n_1814),
.B(n_1815),
.Y(n_12796)
);

NOR2xp33_ASAP7_75t_L g12797 ( 
.A(n_12320),
.B(n_12584),
.Y(n_12797)
);

INVx2_ASAP7_75t_L g12798 ( 
.A(n_12446),
.Y(n_12798)
);

AOI21x1_ASAP7_75t_L g12799 ( 
.A1(n_12594),
.A2(n_1816),
.B(n_1817),
.Y(n_12799)
);

INVx1_ASAP7_75t_L g12800 ( 
.A(n_12398),
.Y(n_12800)
);

OAI21x1_ASAP7_75t_L g12801 ( 
.A1(n_12319),
.A2(n_1817),
.B(n_1818),
.Y(n_12801)
);

A2O1A1Ixp33_ASAP7_75t_L g12802 ( 
.A1(n_12420),
.A2(n_1820),
.B(n_1818),
.C(n_1819),
.Y(n_12802)
);

NOR2xp33_ASAP7_75t_L g12803 ( 
.A(n_12557),
.B(n_1820),
.Y(n_12803)
);

AOI21xp5_ASAP7_75t_L g12804 ( 
.A1(n_12312),
.A2(n_12328),
.B(n_12300),
.Y(n_12804)
);

CKINVDCx20_ASAP7_75t_R g12805 ( 
.A(n_12607),
.Y(n_12805)
);

OR2x6_ASAP7_75t_L g12806 ( 
.A(n_12507),
.B(n_1821),
.Y(n_12806)
);

AOI21xp5_ASAP7_75t_L g12807 ( 
.A1(n_12312),
.A2(n_1821),
.B(n_1822),
.Y(n_12807)
);

INVx1_ASAP7_75t_L g12808 ( 
.A(n_12415),
.Y(n_12808)
);

INVx2_ASAP7_75t_L g12809 ( 
.A(n_12472),
.Y(n_12809)
);

OR2x6_ASAP7_75t_L g12810 ( 
.A(n_12507),
.B(n_1822),
.Y(n_12810)
);

OA21x2_ASAP7_75t_L g12811 ( 
.A1(n_12351),
.A2(n_1823),
.B(n_1824),
.Y(n_12811)
);

AOI21xp5_ASAP7_75t_L g12812 ( 
.A1(n_12480),
.A2(n_12523),
.B(n_12604),
.Y(n_12812)
);

INVx2_ASAP7_75t_L g12813 ( 
.A(n_12539),
.Y(n_12813)
);

AND2x4_ASAP7_75t_L g12814 ( 
.A(n_12593),
.B(n_1823),
.Y(n_12814)
);

NAND2xp5_ASAP7_75t_L g12815 ( 
.A(n_12643),
.B(n_1824),
.Y(n_12815)
);

OAI21x1_ASAP7_75t_L g12816 ( 
.A1(n_12651),
.A2(n_1825),
.B(n_1826),
.Y(n_12816)
);

HB1xp67_ASAP7_75t_L g12817 ( 
.A(n_12653),
.Y(n_12817)
);

NAND2xp5_ASAP7_75t_SL g12818 ( 
.A(n_12362),
.B(n_1825),
.Y(n_12818)
);

AOI21xp5_ASAP7_75t_L g12819 ( 
.A1(n_12322),
.A2(n_1826),
.B(n_1827),
.Y(n_12819)
);

INVx1_ASAP7_75t_L g12820 ( 
.A(n_12453),
.Y(n_12820)
);

OAI21x1_ASAP7_75t_L g12821 ( 
.A1(n_12654),
.A2(n_1828),
.B(n_1829),
.Y(n_12821)
);

AND2x2_ASAP7_75t_L g12822 ( 
.A(n_12340),
.B(n_1828),
.Y(n_12822)
);

AND2x4_ASAP7_75t_L g12823 ( 
.A(n_12355),
.B(n_1829),
.Y(n_12823)
);

INVx1_ASAP7_75t_L g12824 ( 
.A(n_12506),
.Y(n_12824)
);

OA21x2_ASAP7_75t_L g12825 ( 
.A1(n_12307),
.A2(n_12592),
.B(n_12381),
.Y(n_12825)
);

INVx1_ASAP7_75t_L g12826 ( 
.A(n_12429),
.Y(n_12826)
);

INVx2_ASAP7_75t_L g12827 ( 
.A(n_12565),
.Y(n_12827)
);

INVx2_ASAP7_75t_L g12828 ( 
.A(n_12531),
.Y(n_12828)
);

AOI21x1_ASAP7_75t_L g12829 ( 
.A1(n_12580),
.A2(n_1830),
.B(n_1831),
.Y(n_12829)
);

AND2x2_ASAP7_75t_L g12830 ( 
.A(n_12321),
.B(n_1830),
.Y(n_12830)
);

NOR2x1_ASAP7_75t_R g12831 ( 
.A(n_12575),
.B(n_1831),
.Y(n_12831)
);

AO31x2_ASAP7_75t_L g12832 ( 
.A1(n_12647),
.A2(n_1835),
.A3(n_1832),
.B(n_1834),
.Y(n_12832)
);

INVx3_ASAP7_75t_L g12833 ( 
.A(n_12520),
.Y(n_12833)
);

OA21x2_ASAP7_75t_L g12834 ( 
.A1(n_12598),
.A2(n_1832),
.B(n_1834),
.Y(n_12834)
);

HB1xp67_ASAP7_75t_L g12835 ( 
.A(n_12293),
.Y(n_12835)
);

INVxp33_ASAP7_75t_L g12836 ( 
.A(n_12416),
.Y(n_12836)
);

AO31x2_ASAP7_75t_L g12837 ( 
.A1(n_12656),
.A2(n_12519),
.A3(n_12486),
.B(n_12481),
.Y(n_12837)
);

NAND2xp5_ASAP7_75t_L g12838 ( 
.A(n_12309),
.B(n_1837),
.Y(n_12838)
);

AOI21xp5_ASAP7_75t_L g12839 ( 
.A1(n_12511),
.A2(n_1837),
.B(n_1838),
.Y(n_12839)
);

INVx1_ASAP7_75t_L g12840 ( 
.A(n_12521),
.Y(n_12840)
);

AOI22xp33_ASAP7_75t_L g12841 ( 
.A1(n_12311),
.A2(n_1840),
.B1(n_1838),
.B2(n_1839),
.Y(n_12841)
);

NAND2xp5_ASAP7_75t_L g12842 ( 
.A(n_12403),
.B(n_1839),
.Y(n_12842)
);

OAI21xp5_ASAP7_75t_L g12843 ( 
.A1(n_12621),
.A2(n_1840),
.B(n_1841),
.Y(n_12843)
);

BUFx6f_ASAP7_75t_L g12844 ( 
.A(n_12425),
.Y(n_12844)
);

AOI21xp5_ASAP7_75t_L g12845 ( 
.A1(n_12588),
.A2(n_1841),
.B(n_1842),
.Y(n_12845)
);

INVx1_ASAP7_75t_L g12846 ( 
.A(n_12461),
.Y(n_12846)
);

NAND2xp5_ASAP7_75t_L g12847 ( 
.A(n_12338),
.B(n_1842),
.Y(n_12847)
);

INVx1_ASAP7_75t_L g12848 ( 
.A(n_12372),
.Y(n_12848)
);

OAI21xp5_ASAP7_75t_L g12849 ( 
.A1(n_12346),
.A2(n_1843),
.B(n_1844),
.Y(n_12849)
);

AOI22xp33_ASAP7_75t_L g12850 ( 
.A1(n_12365),
.A2(n_1845),
.B1(n_1843),
.B2(n_1844),
.Y(n_12850)
);

OA21x2_ASAP7_75t_L g12851 ( 
.A1(n_12303),
.A2(n_1845),
.B(n_1846),
.Y(n_12851)
);

INVx1_ASAP7_75t_L g12852 ( 
.A(n_12409),
.Y(n_12852)
);

INVx1_ASAP7_75t_L g12853 ( 
.A(n_12533),
.Y(n_12853)
);

INVx2_ASAP7_75t_L g12854 ( 
.A(n_12364),
.Y(n_12854)
);

HB1xp67_ASAP7_75t_L g12855 ( 
.A(n_12315),
.Y(n_12855)
);

OR2x2_ASAP7_75t_L g12856 ( 
.A(n_12370),
.B(n_12343),
.Y(n_12856)
);

AOI21xp5_ASAP7_75t_L g12857 ( 
.A1(n_12615),
.A2(n_12553),
.B(n_12391),
.Y(n_12857)
);

INVx2_ASAP7_75t_L g12858 ( 
.A(n_12642),
.Y(n_12858)
);

AND2x4_ASAP7_75t_L g12859 ( 
.A(n_12495),
.B(n_1846),
.Y(n_12859)
);

AND2x2_ASAP7_75t_L g12860 ( 
.A(n_12304),
.B(n_1847),
.Y(n_12860)
);

AND2x2_ASAP7_75t_L g12861 ( 
.A(n_12567),
.B(n_1848),
.Y(n_12861)
);

OAI21x1_ASAP7_75t_L g12862 ( 
.A1(n_12314),
.A2(n_1848),
.B(n_1849),
.Y(n_12862)
);

NAND2xp5_ASAP7_75t_L g12863 ( 
.A(n_12395),
.B(n_1849),
.Y(n_12863)
);

BUFx3_ASAP7_75t_L g12864 ( 
.A(n_12543),
.Y(n_12864)
);

AND2x2_ASAP7_75t_L g12865 ( 
.A(n_12612),
.B(n_1850),
.Y(n_12865)
);

INVx1_ASAP7_75t_L g12866 ( 
.A(n_12448),
.Y(n_12866)
);

INVx2_ASAP7_75t_L g12867 ( 
.A(n_12407),
.Y(n_12867)
);

INVx2_ASAP7_75t_L g12868 ( 
.A(n_12518),
.Y(n_12868)
);

OAI22xp5_ASAP7_75t_L g12869 ( 
.A1(n_12430),
.A2(n_1852),
.B1(n_1850),
.B2(n_1851),
.Y(n_12869)
);

AOI21xp5_ASAP7_75t_L g12870 ( 
.A1(n_12517),
.A2(n_1851),
.B(n_1852),
.Y(n_12870)
);

OAI21x1_ASAP7_75t_L g12871 ( 
.A1(n_12357),
.A2(n_1854),
.B(n_1855),
.Y(n_12871)
);

A2O1A1Ixp33_ASAP7_75t_L g12872 ( 
.A1(n_12308),
.A2(n_1856),
.B(n_1854),
.C(n_1855),
.Y(n_12872)
);

NAND2xp5_ASAP7_75t_L g12873 ( 
.A(n_12369),
.B(n_1857),
.Y(n_12873)
);

AOI21xp5_ASAP7_75t_L g12874 ( 
.A1(n_12471),
.A2(n_12536),
.B(n_12655),
.Y(n_12874)
);

OAI21x1_ASAP7_75t_SL g12875 ( 
.A1(n_12620),
.A2(n_1857),
.B(n_1858),
.Y(n_12875)
);

NOR2xp33_ASAP7_75t_L g12876 ( 
.A(n_12501),
.B(n_1858),
.Y(n_12876)
);

INVx1_ASAP7_75t_L g12877 ( 
.A(n_12548),
.Y(n_12877)
);

INVx8_ASAP7_75t_L g12878 ( 
.A(n_12661),
.Y(n_12878)
);

OAI21xp5_ASAP7_75t_L g12879 ( 
.A1(n_12366),
.A2(n_1859),
.B(n_1860),
.Y(n_12879)
);

NAND2xp5_ASAP7_75t_L g12880 ( 
.A(n_12383),
.B(n_1859),
.Y(n_12880)
);

AOI21x1_ASAP7_75t_L g12881 ( 
.A1(n_12342),
.A2(n_12528),
.B(n_12619),
.Y(n_12881)
);

HB1xp67_ASAP7_75t_L g12882 ( 
.A(n_12483),
.Y(n_12882)
);

AOI21xp5_ASAP7_75t_L g12883 ( 
.A1(n_12596),
.A2(n_1860),
.B(n_1861),
.Y(n_12883)
);

AND2x2_ASAP7_75t_L g12884 ( 
.A(n_12631),
.B(n_1861),
.Y(n_12884)
);

HB1xp67_ASAP7_75t_L g12885 ( 
.A(n_12626),
.Y(n_12885)
);

CKINVDCx5p33_ASAP7_75t_R g12886 ( 
.A(n_12597),
.Y(n_12886)
);

INVx2_ASAP7_75t_L g12887 ( 
.A(n_12552),
.Y(n_12887)
);

NAND2xp5_ASAP7_75t_L g12888 ( 
.A(n_12414),
.B(n_1862),
.Y(n_12888)
);

AOI21xp5_ASAP7_75t_L g12889 ( 
.A1(n_12581),
.A2(n_12635),
.B(n_12509),
.Y(n_12889)
);

INVx2_ASAP7_75t_L g12890 ( 
.A(n_12560),
.Y(n_12890)
);

AND2x2_ASAP7_75t_L g12891 ( 
.A(n_12595),
.B(n_1863),
.Y(n_12891)
);

OAI21xp5_ASAP7_75t_L g12892 ( 
.A1(n_12349),
.A2(n_1864),
.B(n_1865),
.Y(n_12892)
);

OA21x2_ASAP7_75t_L g12893 ( 
.A1(n_12385),
.A2(n_12371),
.B(n_12603),
.Y(n_12893)
);

AND2x2_ASAP7_75t_L g12894 ( 
.A(n_12558),
.B(n_12623),
.Y(n_12894)
);

INVx1_ASAP7_75t_L g12895 ( 
.A(n_12601),
.Y(n_12895)
);

OAI21x1_ASAP7_75t_L g12896 ( 
.A1(n_12296),
.A2(n_1864),
.B(n_1865),
.Y(n_12896)
);

OA21x2_ASAP7_75t_L g12897 ( 
.A1(n_12410),
.A2(n_1866),
.B(n_1867),
.Y(n_12897)
);

BUFx3_ASAP7_75t_L g12898 ( 
.A(n_12569),
.Y(n_12898)
);

INVx3_ASAP7_75t_L g12899 ( 
.A(n_12586),
.Y(n_12899)
);

INVx1_ASAP7_75t_L g12900 ( 
.A(n_12439),
.Y(n_12900)
);

INVx1_ASAP7_75t_L g12901 ( 
.A(n_12464),
.Y(n_12901)
);

INVx1_ASAP7_75t_L g12902 ( 
.A(n_12497),
.Y(n_12902)
);

AOI21x1_ASAP7_75t_L g12903 ( 
.A1(n_12624),
.A2(n_12493),
.B(n_12559),
.Y(n_12903)
);

NAND2xp5_ASAP7_75t_L g12904 ( 
.A(n_12534),
.B(n_1866),
.Y(n_12904)
);

OA21x2_ASAP7_75t_L g12905 ( 
.A1(n_12306),
.A2(n_1867),
.B(n_1869),
.Y(n_12905)
);

NAND2xp5_ASAP7_75t_L g12906 ( 
.A(n_12478),
.B(n_12496),
.Y(n_12906)
);

AND2x2_ASAP7_75t_L g12907 ( 
.A(n_12334),
.B(n_12648),
.Y(n_12907)
);

AOI22xp33_ASAP7_75t_L g12908 ( 
.A1(n_12589),
.A2(n_1871),
.B1(n_1869),
.B2(n_1870),
.Y(n_12908)
);

AOI21x1_ASAP7_75t_L g12909 ( 
.A1(n_12561),
.A2(n_1870),
.B(n_1871),
.Y(n_12909)
);

INVx1_ASAP7_75t_L g12910 ( 
.A(n_12497),
.Y(n_12910)
);

NAND2xp5_ASAP7_75t_L g12911 ( 
.A(n_12503),
.B(n_1872),
.Y(n_12911)
);

INVx1_ASAP7_75t_L g12912 ( 
.A(n_12549),
.Y(n_12912)
);

NAND2xp5_ASAP7_75t_L g12913 ( 
.A(n_12540),
.B(n_1872),
.Y(n_12913)
);

INVx1_ASAP7_75t_L g12914 ( 
.A(n_12505),
.Y(n_12914)
);

NAND2x1p5_ASAP7_75t_L g12915 ( 
.A(n_12387),
.B(n_1873),
.Y(n_12915)
);

CKINVDCx5p33_ASAP7_75t_R g12916 ( 
.A(n_12373),
.Y(n_12916)
);

BUFx2_ASAP7_75t_R g12917 ( 
.A(n_12617),
.Y(n_12917)
);

INVx2_ASAP7_75t_L g12918 ( 
.A(n_12649),
.Y(n_12918)
);

AOI22xp33_ASAP7_75t_L g12919 ( 
.A1(n_12399),
.A2(n_1875),
.B1(n_1873),
.B2(n_1874),
.Y(n_12919)
);

HB1xp67_ASAP7_75t_L g12920 ( 
.A(n_12505),
.Y(n_12920)
);

INVx2_ASAP7_75t_L g12921 ( 
.A(n_12586),
.Y(n_12921)
);

INVx1_ASAP7_75t_L g12922 ( 
.A(n_12547),
.Y(n_12922)
);

INVx1_ASAP7_75t_L g12923 ( 
.A(n_12650),
.Y(n_12923)
);

AO21x2_ASAP7_75t_L g12924 ( 
.A1(n_12566),
.A2(n_1874),
.B(n_1875),
.Y(n_12924)
);

INVx1_ASAP7_75t_SL g12925 ( 
.A(n_12546),
.Y(n_12925)
);

OAI21x1_ASAP7_75t_L g12926 ( 
.A1(n_12418),
.A2(n_1876),
.B(n_1877),
.Y(n_12926)
);

BUFx3_ASAP7_75t_L g12927 ( 
.A(n_12628),
.Y(n_12927)
);

AND2x2_ASAP7_75t_L g12928 ( 
.A(n_12529),
.B(n_12452),
.Y(n_12928)
);

AO31x2_ASAP7_75t_L g12929 ( 
.A1(n_12494),
.A2(n_1878),
.A3(n_1876),
.B(n_1877),
.Y(n_12929)
);

NAND2xp5_ASAP7_75t_L g12930 ( 
.A(n_12583),
.B(n_1879),
.Y(n_12930)
);

INVx2_ASAP7_75t_L g12931 ( 
.A(n_12469),
.Y(n_12931)
);

AOI21xp5_ASAP7_75t_L g12932 ( 
.A1(n_12657),
.A2(n_1879),
.B(n_1880),
.Y(n_12932)
);

AO31x2_ASAP7_75t_L g12933 ( 
.A1(n_12634),
.A2(n_1882),
.A3(n_1880),
.B(n_1881),
.Y(n_12933)
);

INVx1_ASAP7_75t_L g12934 ( 
.A(n_12650),
.Y(n_12934)
);

AO21x2_ASAP7_75t_L g12935 ( 
.A1(n_12646),
.A2(n_1881),
.B(n_1882),
.Y(n_12935)
);

NOR2x1_ASAP7_75t_R g12936 ( 
.A(n_12614),
.B(n_1883),
.Y(n_12936)
);

INVx1_ASAP7_75t_L g12937 ( 
.A(n_12652),
.Y(n_12937)
);

AOI21x1_ASAP7_75t_L g12938 ( 
.A1(n_12638),
.A2(n_1883),
.B(n_1884),
.Y(n_12938)
);

INVx1_ASAP7_75t_L g12939 ( 
.A(n_12652),
.Y(n_12939)
);

INVx1_ASAP7_75t_L g12940 ( 
.A(n_12459),
.Y(n_12940)
);

AOI21xp5_ASAP7_75t_L g12941 ( 
.A1(n_12609),
.A2(n_1884),
.B(n_1885),
.Y(n_12941)
);

BUFx6f_ASAP7_75t_L g12942 ( 
.A(n_12627),
.Y(n_12942)
);

AOI21xp5_ASAP7_75t_L g12943 ( 
.A1(n_12535),
.A2(n_1885),
.B(n_1886),
.Y(n_12943)
);

A2O1A1Ixp33_ASAP7_75t_L g12944 ( 
.A1(n_12515),
.A2(n_1888),
.B(n_1886),
.C(n_1887),
.Y(n_12944)
);

INVx2_ASAP7_75t_L g12945 ( 
.A(n_12644),
.Y(n_12945)
);

INVx3_ASAP7_75t_L g12946 ( 
.A(n_12571),
.Y(n_12946)
);

CKINVDCx6p67_ASAP7_75t_R g12947 ( 
.A(n_12479),
.Y(n_12947)
);

NOR2xp33_ASAP7_75t_L g12948 ( 
.A(n_12564),
.B(n_1888),
.Y(n_12948)
);

NOR2x1_ASAP7_75t_SL g12949 ( 
.A(n_12625),
.B(n_1889),
.Y(n_12949)
);

AOI21x1_ASAP7_75t_L g12950 ( 
.A1(n_12599),
.A2(n_1890),
.B(n_1891),
.Y(n_12950)
);

CKINVDCx11_ASAP7_75t_R g12951 ( 
.A(n_12629),
.Y(n_12951)
);

BUFx2_ASAP7_75t_SL g12952 ( 
.A(n_12574),
.Y(n_12952)
);

OAI21x1_ASAP7_75t_L g12953 ( 
.A1(n_12508),
.A2(n_1890),
.B(n_1891),
.Y(n_12953)
);

NAND2xp5_ASAP7_75t_L g12954 ( 
.A(n_12361),
.B(n_1892),
.Y(n_12954)
);

AND2x4_ASAP7_75t_L g12955 ( 
.A(n_12449),
.B(n_1892),
.Y(n_12955)
);

INVx2_ASAP7_75t_L g12956 ( 
.A(n_12454),
.Y(n_12956)
);

AO31x2_ASAP7_75t_L g12957 ( 
.A1(n_12585),
.A2(n_1896),
.A3(n_1894),
.B(n_1895),
.Y(n_12957)
);

AND2x2_ASAP7_75t_L g12958 ( 
.A(n_12421),
.B(n_1894),
.Y(n_12958)
);

INVx1_ASAP7_75t_L g12959 ( 
.A(n_12459),
.Y(n_12959)
);

INVx1_ASAP7_75t_L g12960 ( 
.A(n_12554),
.Y(n_12960)
);

AOI21xp33_ASAP7_75t_SL g12961 ( 
.A1(n_12477),
.A2(n_1896),
.B(n_1897),
.Y(n_12961)
);

NAND3xp33_ASAP7_75t_L g12962 ( 
.A(n_12489),
.B(n_1897),
.C(n_1898),
.Y(n_12962)
);

OAI21x1_ASAP7_75t_L g12963 ( 
.A1(n_12456),
.A2(n_1898),
.B(n_1899),
.Y(n_12963)
);

OR2x2_ASAP7_75t_L g12964 ( 
.A(n_12361),
.B(n_1899),
.Y(n_12964)
);

INVx1_ASAP7_75t_L g12965 ( 
.A(n_12457),
.Y(n_12965)
);

AO31x2_ASAP7_75t_L g12966 ( 
.A1(n_12639),
.A2(n_1902),
.A3(n_1900),
.B(n_1901),
.Y(n_12966)
);

OAI21xp5_ASAP7_75t_L g12967 ( 
.A1(n_12470),
.A2(n_1900),
.B(n_1902),
.Y(n_12967)
);

OAI21x1_ASAP7_75t_L g12968 ( 
.A1(n_12475),
.A2(n_1903),
.B(n_1904),
.Y(n_12968)
);

NAND2xp5_ASAP7_75t_L g12969 ( 
.A(n_12577),
.B(n_1903),
.Y(n_12969)
);

HB1xp67_ASAP7_75t_L g12970 ( 
.A(n_12514),
.Y(n_12970)
);

INVx2_ASAP7_75t_L g12971 ( 
.A(n_12451),
.Y(n_12971)
);

INVx2_ASAP7_75t_L g12972 ( 
.A(n_12545),
.Y(n_12972)
);

AO31x2_ASAP7_75t_L g12973 ( 
.A1(n_12660),
.A2(n_1906),
.A3(n_1904),
.B(n_1905),
.Y(n_12973)
);

AOI22xp33_ASAP7_75t_L g12974 ( 
.A1(n_12613),
.A2(n_1908),
.B1(n_1905),
.B2(n_1906),
.Y(n_12974)
);

INVx1_ASAP7_75t_L g12975 ( 
.A(n_12636),
.Y(n_12975)
);

NAND2xp5_ASAP7_75t_L g12976 ( 
.A(n_12514),
.B(n_1908),
.Y(n_12976)
);

OA21x2_ASAP7_75t_L g12977 ( 
.A1(n_12476),
.A2(n_1909),
.B(n_1910),
.Y(n_12977)
);

AND2x4_ASAP7_75t_L g12978 ( 
.A(n_12527),
.B(n_12488),
.Y(n_12978)
);

NAND2xp5_ASAP7_75t_L g12979 ( 
.A(n_12538),
.B(n_1909),
.Y(n_12979)
);

INVx1_ASAP7_75t_L g12980 ( 
.A(n_12636),
.Y(n_12980)
);

AO21x2_ASAP7_75t_L g12981 ( 
.A1(n_12468),
.A2(n_1910),
.B(n_1911),
.Y(n_12981)
);

AOI222xp33_ASAP7_75t_L g12982 ( 
.A1(n_12640),
.A2(n_1915),
.B1(n_1917),
.B2(n_1912),
.C1(n_1914),
.C2(n_1916),
.Y(n_12982)
);

INVx1_ASAP7_75t_L g12983 ( 
.A(n_12538),
.Y(n_12983)
);

AND2x2_ASAP7_75t_L g12984 ( 
.A(n_12513),
.B(n_1912),
.Y(n_12984)
);

OA21x2_ASAP7_75t_L g12985 ( 
.A1(n_12498),
.A2(n_1915),
.B(n_1917),
.Y(n_12985)
);

INVx2_ASAP7_75t_L g12986 ( 
.A(n_12516),
.Y(n_12986)
);

INVx2_ASAP7_75t_L g12987 ( 
.A(n_12524),
.Y(n_12987)
);

INVx1_ASAP7_75t_L g12988 ( 
.A(n_12587),
.Y(n_12988)
);

OAI21x1_ASAP7_75t_L g12989 ( 
.A1(n_12512),
.A2(n_1918),
.B(n_1919),
.Y(n_12989)
);

NAND2xp5_ASAP7_75t_L g12990 ( 
.A(n_12587),
.B(n_1920),
.Y(n_12990)
);

HB1xp67_ASAP7_75t_L g12991 ( 
.A(n_12525),
.Y(n_12991)
);

INVx2_ASAP7_75t_L g12992 ( 
.A(n_12542),
.Y(n_12992)
);

AND2x2_ASAP7_75t_L g12993 ( 
.A(n_12555),
.B(n_1922),
.Y(n_12993)
);

A2O1A1Ixp33_ASAP7_75t_L g12994 ( 
.A1(n_12556),
.A2(n_1925),
.B(n_1923),
.C(n_1924),
.Y(n_12994)
);

AOI21xp5_ASAP7_75t_L g12995 ( 
.A1(n_12618),
.A2(n_1924),
.B(n_1925),
.Y(n_12995)
);

OAI21x1_ASAP7_75t_L g12996 ( 
.A1(n_12541),
.A2(n_1926),
.B(n_1927),
.Y(n_12996)
);

OA21x2_ASAP7_75t_L g12997 ( 
.A1(n_12562),
.A2(n_1926),
.B(n_1927),
.Y(n_12997)
);

INVx2_ASAP7_75t_L g12998 ( 
.A(n_12563),
.Y(n_12998)
);

A2O1A1Ixp33_ASAP7_75t_L g12999 ( 
.A1(n_12578),
.A2(n_1930),
.B(n_1928),
.C(n_1929),
.Y(n_12999)
);

NAND2xp5_ASAP7_75t_L g13000 ( 
.A(n_12590),
.B(n_1928),
.Y(n_13000)
);

OAI21xp5_ASAP7_75t_L g13001 ( 
.A1(n_12600),
.A2(n_1929),
.B(n_1931),
.Y(n_13001)
);

AND2x4_ASAP7_75t_L g13002 ( 
.A(n_12602),
.B(n_1931),
.Y(n_13002)
);

AOI21xp5_ASAP7_75t_L g13003 ( 
.A1(n_12622),
.A2(n_1932),
.B(n_1933),
.Y(n_13003)
);

INVx1_ASAP7_75t_SL g13004 ( 
.A(n_12645),
.Y(n_13004)
);

INVx1_ASAP7_75t_L g13005 ( 
.A(n_12632),
.Y(n_13005)
);

INVx2_ASAP7_75t_L g13006 ( 
.A(n_12637),
.Y(n_13006)
);

OA21x2_ASAP7_75t_L g13007 ( 
.A1(n_12658),
.A2(n_1933),
.B(n_1934),
.Y(n_13007)
);

OAI21xp5_ASAP7_75t_L g13008 ( 
.A1(n_12659),
.A2(n_1934),
.B(n_1935),
.Y(n_13008)
);

BUFx2_ASAP7_75t_L g13009 ( 
.A(n_12530),
.Y(n_13009)
);

AND2x4_ASAP7_75t_L g13010 ( 
.A(n_12662),
.B(n_1935),
.Y(n_13010)
);

AOI21x1_ASAP7_75t_L g13011 ( 
.A1(n_12526),
.A2(n_1936),
.B(n_1937),
.Y(n_13011)
);

AO21x2_ASAP7_75t_L g13012 ( 
.A1(n_12608),
.A2(n_1936),
.B(n_1938),
.Y(n_13012)
);

NAND2xp5_ASAP7_75t_L g13013 ( 
.A(n_12611),
.B(n_1938),
.Y(n_13013)
);

AO31x2_ASAP7_75t_L g13014 ( 
.A1(n_12363),
.A2(n_1941),
.A3(n_1939),
.B(n_1940),
.Y(n_13014)
);

OR2x2_ASAP7_75t_L g13015 ( 
.A(n_12856),
.B(n_1939),
.Y(n_13015)
);

AOI21x1_ASAP7_75t_L g13016 ( 
.A1(n_12719),
.A2(n_1941),
.B(n_1942),
.Y(n_13016)
);

INVx1_ASAP7_75t_L g13017 ( 
.A(n_12667),
.Y(n_13017)
);

HB1xp67_ASAP7_75t_L g13018 ( 
.A(n_13014),
.Y(n_13018)
);

OR2x2_ASAP7_75t_L g13019 ( 
.A(n_12848),
.B(n_1943),
.Y(n_13019)
);

HB1xp67_ASAP7_75t_L g13020 ( 
.A(n_13014),
.Y(n_13020)
);

INVx1_ASAP7_75t_L g13021 ( 
.A(n_12673),
.Y(n_13021)
);

AND2x2_ASAP7_75t_L g13022 ( 
.A(n_12671),
.B(n_1943),
.Y(n_13022)
);

OAI21x1_ASAP7_75t_L g13023 ( 
.A1(n_12682),
.A2(n_1944),
.B(n_1945),
.Y(n_13023)
);

INVx1_ASAP7_75t_L g13024 ( 
.A(n_12676),
.Y(n_13024)
);

AND2x2_ASAP7_75t_L g13025 ( 
.A(n_12700),
.B(n_1944),
.Y(n_13025)
);

INVx1_ASAP7_75t_L g13026 ( 
.A(n_12683),
.Y(n_13026)
);

INVx2_ASAP7_75t_L g13027 ( 
.A(n_12771),
.Y(n_13027)
);

NAND2xp5_ASAP7_75t_L g13028 ( 
.A(n_12851),
.B(n_12965),
.Y(n_13028)
);

OAI21x1_ASAP7_75t_L g13029 ( 
.A1(n_12881),
.A2(n_1945),
.B(n_1946),
.Y(n_13029)
);

HB1xp67_ASAP7_75t_L g13030 ( 
.A(n_12696),
.Y(n_13030)
);

INVx1_ASAP7_75t_L g13031 ( 
.A(n_12684),
.Y(n_13031)
);

AOI22xp33_ASAP7_75t_L g13032 ( 
.A1(n_12716),
.A2(n_1948),
.B1(n_1946),
.B2(n_1947),
.Y(n_13032)
);

INVx2_ASAP7_75t_L g13033 ( 
.A(n_12771),
.Y(n_13033)
);

INVx2_ASAP7_75t_L g13034 ( 
.A(n_12771),
.Y(n_13034)
);

OA21x2_ASAP7_75t_L g13035 ( 
.A1(n_12679),
.A2(n_1947),
.B(n_1948),
.Y(n_13035)
);

INVxp67_ASAP7_75t_SL g13036 ( 
.A(n_12855),
.Y(n_13036)
);

INVx1_ASAP7_75t_L g13037 ( 
.A(n_12685),
.Y(n_13037)
);

INVx1_ASAP7_75t_L g13038 ( 
.A(n_12686),
.Y(n_13038)
);

INVx2_ASAP7_75t_L g13039 ( 
.A(n_12844),
.Y(n_13039)
);

BUFx2_ASAP7_75t_L g13040 ( 
.A(n_12749),
.Y(n_13040)
);

INVx1_ASAP7_75t_L g13041 ( 
.A(n_12699),
.Y(n_13041)
);

AOI21x1_ASAP7_75t_L g13042 ( 
.A1(n_12835),
.A2(n_1949),
.B(n_1951),
.Y(n_13042)
);

BUFx6f_ASAP7_75t_L g13043 ( 
.A(n_12698),
.Y(n_13043)
);

INVx1_ASAP7_75t_L g13044 ( 
.A(n_12726),
.Y(n_13044)
);

HB1xp67_ASAP7_75t_L g13045 ( 
.A(n_12735),
.Y(n_13045)
);

INVx2_ASAP7_75t_L g13046 ( 
.A(n_12844),
.Y(n_13046)
);

AND2x2_ASAP7_75t_L g13047 ( 
.A(n_12833),
.B(n_1949),
.Y(n_13047)
);

INVx5_ASAP7_75t_L g13048 ( 
.A(n_12674),
.Y(n_13048)
);

INVx2_ASAP7_75t_L g13049 ( 
.A(n_12765),
.Y(n_13049)
);

INVx2_ASAP7_75t_L g13050 ( 
.A(n_12907),
.Y(n_13050)
);

INVx2_ASAP7_75t_SL g13051 ( 
.A(n_12757),
.Y(n_13051)
);

INVx2_ASAP7_75t_L g13052 ( 
.A(n_12677),
.Y(n_13052)
);

INVx1_ASAP7_75t_L g13053 ( 
.A(n_12750),
.Y(n_13053)
);

INVx1_ASAP7_75t_L g13054 ( 
.A(n_12751),
.Y(n_13054)
);

INVx2_ASAP7_75t_L g13055 ( 
.A(n_12747),
.Y(n_13055)
);

HB1xp67_ASAP7_75t_L g13056 ( 
.A(n_12705),
.Y(n_13056)
);

HB1xp67_ASAP7_75t_L g13057 ( 
.A(n_12905),
.Y(n_13057)
);

INVx1_ASAP7_75t_L g13058 ( 
.A(n_12753),
.Y(n_13058)
);

INVx1_ASAP7_75t_L g13059 ( 
.A(n_12764),
.Y(n_13059)
);

INVx2_ASAP7_75t_L g13060 ( 
.A(n_12759),
.Y(n_13060)
);

HB1xp67_ASAP7_75t_L g13061 ( 
.A(n_12885),
.Y(n_13061)
);

INVx2_ASAP7_75t_L g13062 ( 
.A(n_12783),
.Y(n_13062)
);

INVx2_ASAP7_75t_SL g13063 ( 
.A(n_12878),
.Y(n_13063)
);

NAND2xp5_ASAP7_75t_L g13064 ( 
.A(n_12940),
.B(n_12959),
.Y(n_13064)
);

INVx2_ASAP7_75t_L g13065 ( 
.A(n_12918),
.Y(n_13065)
);

AND2x2_ASAP7_75t_L g13066 ( 
.A(n_12854),
.B(n_1951),
.Y(n_13066)
);

HB1xp67_ASAP7_75t_L g13067 ( 
.A(n_12692),
.Y(n_13067)
);

INVx2_ASAP7_75t_L g13068 ( 
.A(n_12715),
.Y(n_13068)
);

OAI21x1_ASAP7_75t_L g13069 ( 
.A1(n_12826),
.A2(n_12798),
.B(n_12866),
.Y(n_13069)
);

AO21x2_ASAP7_75t_L g13070 ( 
.A1(n_12882),
.A2(n_1952),
.B(n_1953),
.Y(n_13070)
);

NAND2xp5_ASAP7_75t_L g13071 ( 
.A(n_13013),
.B(n_1952),
.Y(n_13071)
);

INVx2_ASAP7_75t_L g13072 ( 
.A(n_12680),
.Y(n_13072)
);

BUFx6f_ASAP7_75t_L g13073 ( 
.A(n_12774),
.Y(n_13073)
);

NOR2xp33_ASAP7_75t_L g13074 ( 
.A(n_12665),
.B(n_1953),
.Y(n_13074)
);

HB1xp67_ASAP7_75t_L g13075 ( 
.A(n_12991),
.Y(n_13075)
);

OAI22xp5_ASAP7_75t_L g13076 ( 
.A1(n_12689),
.A2(n_1956),
.B1(n_1954),
.B2(n_1955),
.Y(n_13076)
);

OAI21x1_ASAP7_75t_L g13077 ( 
.A1(n_12703),
.A2(n_1954),
.B(n_1955),
.Y(n_13077)
);

AO21x1_ASAP7_75t_L g13078 ( 
.A1(n_12768),
.A2(n_1956),
.B(n_1957),
.Y(n_13078)
);

INVx1_ASAP7_75t_L g13079 ( 
.A(n_12770),
.Y(n_13079)
);

OR2x2_ASAP7_75t_L g13080 ( 
.A(n_12711),
.B(n_1958),
.Y(n_13080)
);

INVx1_ASAP7_75t_L g13081 ( 
.A(n_12772),
.Y(n_13081)
);

INVx1_ASAP7_75t_L g13082 ( 
.A(n_12775),
.Y(n_13082)
);

INVx2_ASAP7_75t_L g13083 ( 
.A(n_12899),
.Y(n_13083)
);

OAI21x1_ASAP7_75t_L g13084 ( 
.A1(n_12867),
.A2(n_1959),
.B(n_1960),
.Y(n_13084)
);

AOI22xp33_ASAP7_75t_L g13085 ( 
.A1(n_12754),
.A2(n_1961),
.B1(n_1959),
.B2(n_1960),
.Y(n_13085)
);

INVx1_ASAP7_75t_L g13086 ( 
.A(n_12786),
.Y(n_13086)
);

INVx2_ASAP7_75t_SL g13087 ( 
.A(n_12878),
.Y(n_13087)
);

OAI21x1_ASAP7_75t_SL g13088 ( 
.A1(n_12769),
.A2(n_1961),
.B(n_1962),
.Y(n_13088)
);

AND2x2_ASAP7_75t_L g13089 ( 
.A(n_12813),
.B(n_1963),
.Y(n_13089)
);

INVx1_ASAP7_75t_L g13090 ( 
.A(n_12792),
.Y(n_13090)
);

INVxp67_ASAP7_75t_L g13091 ( 
.A(n_12831),
.Y(n_13091)
);

INVx2_ASAP7_75t_L g13092 ( 
.A(n_12946),
.Y(n_13092)
);

AO21x2_ASAP7_75t_L g13093 ( 
.A1(n_12693),
.A2(n_1963),
.B(n_1964),
.Y(n_13093)
);

OAI21x1_ASAP7_75t_L g13094 ( 
.A1(n_12893),
.A2(n_1964),
.B(n_1965),
.Y(n_13094)
);

INVx3_ASAP7_75t_L g13095 ( 
.A(n_12864),
.Y(n_13095)
);

OR2x2_ASAP7_75t_L g13096 ( 
.A(n_12906),
.B(n_1966),
.Y(n_13096)
);

INVx1_ASAP7_75t_L g13097 ( 
.A(n_12760),
.Y(n_13097)
);

INVx2_ASAP7_75t_L g13098 ( 
.A(n_12691),
.Y(n_13098)
);

AND2x2_ASAP7_75t_L g13099 ( 
.A(n_12827),
.B(n_1966),
.Y(n_13099)
);

NAND2xp5_ASAP7_75t_L g13100 ( 
.A(n_12970),
.B(n_1967),
.Y(n_13100)
);

INVx1_ASAP7_75t_L g13101 ( 
.A(n_12785),
.Y(n_13101)
);

AO21x2_ASAP7_75t_L g13102 ( 
.A1(n_12763),
.A2(n_1967),
.B(n_1968),
.Y(n_13102)
);

NAND2xp5_ASAP7_75t_L g13103 ( 
.A(n_12920),
.B(n_1968),
.Y(n_13103)
);

INVx1_ASAP7_75t_L g13104 ( 
.A(n_12808),
.Y(n_13104)
);

OAI21x1_ASAP7_75t_L g13105 ( 
.A1(n_12743),
.A2(n_1969),
.B(n_1970),
.Y(n_13105)
);

BUFx2_ASAP7_75t_L g13106 ( 
.A(n_12678),
.Y(n_13106)
);

INVx2_ASAP7_75t_L g13107 ( 
.A(n_12921),
.Y(n_13107)
);

INVx4_ASAP7_75t_L g13108 ( 
.A(n_12697),
.Y(n_13108)
);

INVx1_ASAP7_75t_L g13109 ( 
.A(n_12820),
.Y(n_13109)
);

OR2x6_ASAP7_75t_L g13110 ( 
.A(n_12678),
.B(n_12806),
.Y(n_13110)
);

NAND2x1_ASAP7_75t_L g13111 ( 
.A(n_12825),
.B(n_12846),
.Y(n_13111)
);

INVx2_ASAP7_75t_L g13112 ( 
.A(n_12926),
.Y(n_13112)
);

NAND2xp5_ASAP7_75t_L g13113 ( 
.A(n_12914),
.B(n_1969),
.Y(n_13113)
);

BUFx3_ASAP7_75t_L g13114 ( 
.A(n_13009),
.Y(n_13114)
);

INVx2_ASAP7_75t_L g13115 ( 
.A(n_12925),
.Y(n_13115)
);

INVx2_ASAP7_75t_L g13116 ( 
.A(n_12858),
.Y(n_13116)
);

INVx2_ASAP7_75t_L g13117 ( 
.A(n_12664),
.Y(n_13117)
);

INVxp67_ASAP7_75t_L g13118 ( 
.A(n_12779),
.Y(n_13118)
);

INVx2_ASAP7_75t_L g13119 ( 
.A(n_12745),
.Y(n_13119)
);

AND2x2_ASAP7_75t_L g13120 ( 
.A(n_12694),
.B(n_1971),
.Y(n_13120)
);

OR2x2_ASAP7_75t_L g13121 ( 
.A(n_12752),
.B(n_12828),
.Y(n_13121)
);

INVx1_ASAP7_75t_L g13122 ( 
.A(n_12895),
.Y(n_13122)
);

OAI21x1_ASAP7_75t_L g13123 ( 
.A1(n_12852),
.A2(n_1972),
.B(n_1973),
.Y(n_13123)
);

INVx1_ASAP7_75t_L g13124 ( 
.A(n_12824),
.Y(n_13124)
);

INVx1_ASAP7_75t_L g13125 ( 
.A(n_12901),
.Y(n_13125)
);

INVx3_ASAP7_75t_L g13126 ( 
.A(n_12898),
.Y(n_13126)
);

HB1xp67_ASAP7_75t_L g13127 ( 
.A(n_12714),
.Y(n_13127)
);

INVx1_ASAP7_75t_L g13128 ( 
.A(n_12853),
.Y(n_13128)
);

INVx2_ASAP7_75t_L g13129 ( 
.A(n_12945),
.Y(n_13129)
);

AOI21x1_ASAP7_75t_L g13130 ( 
.A1(n_12681),
.A2(n_12695),
.B(n_12950),
.Y(n_13130)
);

INVx2_ASAP7_75t_SL g13131 ( 
.A(n_12927),
.Y(n_13131)
);

INVx1_ASAP7_75t_L g13132 ( 
.A(n_12912),
.Y(n_13132)
);

INVx1_ASAP7_75t_L g13133 ( 
.A(n_12793),
.Y(n_13133)
);

NAND2xp5_ASAP7_75t_L g13134 ( 
.A(n_12983),
.B(n_1972),
.Y(n_13134)
);

INVx1_ASAP7_75t_L g13135 ( 
.A(n_12794),
.Y(n_13135)
);

INVx1_ASAP7_75t_L g13136 ( 
.A(n_12800),
.Y(n_13136)
);

NAND2xp5_ASAP7_75t_L g13137 ( 
.A(n_12988),
.B(n_1973),
.Y(n_13137)
);

HB1xp67_ASAP7_75t_L g13138 ( 
.A(n_12811),
.Y(n_13138)
);

INVx1_ASAP7_75t_L g13139 ( 
.A(n_12840),
.Y(n_13139)
);

OAI222xp33_ASAP7_75t_L g13140 ( 
.A1(n_12804),
.A2(n_1976),
.B1(n_1978),
.B2(n_1974),
.C1(n_1975),
.C2(n_1977),
.Y(n_13140)
);

AND2x2_ASAP7_75t_L g13141 ( 
.A(n_12868),
.B(n_1974),
.Y(n_13141)
);

INVx1_ASAP7_75t_L g13142 ( 
.A(n_12923),
.Y(n_13142)
);

AOI22xp5_ASAP7_75t_L g13143 ( 
.A1(n_12819),
.A2(n_1978),
.B1(n_1975),
.B2(n_1977),
.Y(n_13143)
);

BUFx3_ASAP7_75t_L g13144 ( 
.A(n_12805),
.Y(n_13144)
);

INVx1_ASAP7_75t_L g13145 ( 
.A(n_12934),
.Y(n_13145)
);

INVx1_ASAP7_75t_L g13146 ( 
.A(n_12937),
.Y(n_13146)
);

AND2x2_ASAP7_75t_L g13147 ( 
.A(n_12894),
.B(n_1979),
.Y(n_13147)
);

INVx4_ASAP7_75t_SL g13148 ( 
.A(n_12929),
.Y(n_13148)
);

INVx1_ASAP7_75t_L g13149 ( 
.A(n_12939),
.Y(n_13149)
);

AND2x4_ASAP7_75t_L g13150 ( 
.A(n_12663),
.B(n_1979),
.Y(n_13150)
);

OAI22xp5_ASAP7_75t_L g13151 ( 
.A1(n_12841),
.A2(n_1982),
.B1(n_1980),
.B2(n_1981),
.Y(n_13151)
);

INVx1_ASAP7_75t_L g13152 ( 
.A(n_12741),
.Y(n_13152)
);

INVx1_ASAP7_75t_L g13153 ( 
.A(n_12780),
.Y(n_13153)
);

INVx1_ASAP7_75t_L g13154 ( 
.A(n_12787),
.Y(n_13154)
);

OA21x2_ASAP7_75t_L g13155 ( 
.A1(n_12900),
.A2(n_12668),
.B(n_12670),
.Y(n_13155)
);

INVx1_ASAP7_75t_L g13156 ( 
.A(n_12791),
.Y(n_13156)
);

INVx2_ASAP7_75t_L g13157 ( 
.A(n_12722),
.Y(n_13157)
);

INVx2_ASAP7_75t_L g13158 ( 
.A(n_12723),
.Y(n_13158)
);

OR2x2_ASAP7_75t_L g13159 ( 
.A(n_12837),
.B(n_1981),
.Y(n_13159)
);

INVx1_ASAP7_75t_L g13160 ( 
.A(n_12732),
.Y(n_13160)
);

BUFx5_ASAP7_75t_L g13161 ( 
.A(n_12822),
.Y(n_13161)
);

INVx1_ASAP7_75t_L g13162 ( 
.A(n_12734),
.Y(n_13162)
);

INVx2_ASAP7_75t_L g13163 ( 
.A(n_12729),
.Y(n_13163)
);

NAND2xp5_ASAP7_75t_L g13164 ( 
.A(n_12975),
.B(n_1983),
.Y(n_13164)
);

INVx2_ASAP7_75t_L g13165 ( 
.A(n_12931),
.Y(n_13165)
);

INVx1_ASAP7_75t_L g13166 ( 
.A(n_12738),
.Y(n_13166)
);

INVx1_ASAP7_75t_L g13167 ( 
.A(n_12744),
.Y(n_13167)
);

AND2x2_ASAP7_75t_L g13168 ( 
.A(n_12887),
.B(n_1984),
.Y(n_13168)
);

INVx1_ASAP7_75t_L g13169 ( 
.A(n_12777),
.Y(n_13169)
);

INVx1_ASAP7_75t_L g13170 ( 
.A(n_12902),
.Y(n_13170)
);

INVx1_ASAP7_75t_L g13171 ( 
.A(n_12910),
.Y(n_13171)
);

INVx1_ASAP7_75t_L g13172 ( 
.A(n_12817),
.Y(n_13172)
);

INVx1_ASAP7_75t_L g13173 ( 
.A(n_12960),
.Y(n_13173)
);

INVx1_ASAP7_75t_L g13174 ( 
.A(n_12980),
.Y(n_13174)
);

AO31x2_ASAP7_75t_L g13175 ( 
.A1(n_12954),
.A2(n_1986),
.A3(n_1984),
.B(n_1985),
.Y(n_13175)
);

INVx1_ASAP7_75t_L g13176 ( 
.A(n_12733),
.Y(n_13176)
);

BUFx6f_ASAP7_75t_L g13177 ( 
.A(n_12814),
.Y(n_13177)
);

INVx1_ASAP7_75t_L g13178 ( 
.A(n_12724),
.Y(n_13178)
);

INVx1_ASAP7_75t_L g13179 ( 
.A(n_12922),
.Y(n_13179)
);

INVx2_ASAP7_75t_L g13180 ( 
.A(n_12809),
.Y(n_13180)
);

INVx2_ASAP7_75t_L g13181 ( 
.A(n_12978),
.Y(n_13181)
);

HB1xp67_ASAP7_75t_L g13182 ( 
.A(n_12666),
.Y(n_13182)
);

INVx2_ASAP7_75t_L g13183 ( 
.A(n_12890),
.Y(n_13183)
);

CKINVDCx8_ASAP7_75t_R g13184 ( 
.A(n_12806),
.Y(n_13184)
);

INVx1_ASAP7_75t_L g13185 ( 
.A(n_12834),
.Y(n_13185)
);

AND2x2_ASAP7_75t_L g13186 ( 
.A(n_12837),
.B(n_1985),
.Y(n_13186)
);

CKINVDCx5p33_ASAP7_75t_R g13187 ( 
.A(n_12767),
.Y(n_13187)
);

INVx1_ASAP7_75t_L g13188 ( 
.A(n_12731),
.Y(n_13188)
);

OAI21x1_ASAP7_75t_L g13189 ( 
.A1(n_12877),
.A2(n_1987),
.B(n_1989),
.Y(n_13189)
);

NAND3x1_ASAP7_75t_L g13190 ( 
.A(n_12903),
.B(n_1987),
.C(n_1990),
.Y(n_13190)
);

INVx1_ASAP7_75t_L g13191 ( 
.A(n_12736),
.Y(n_13191)
);

AOI21xp5_ASAP7_75t_L g13192 ( 
.A1(n_12857),
.A2(n_1990),
.B(n_1991),
.Y(n_13192)
);

INVx1_ASAP7_75t_L g13193 ( 
.A(n_12766),
.Y(n_13193)
);

INVx1_ASAP7_75t_L g13194 ( 
.A(n_12721),
.Y(n_13194)
);

INVx3_ASAP7_75t_L g13195 ( 
.A(n_12942),
.Y(n_13195)
);

AND2x2_ASAP7_75t_L g13196 ( 
.A(n_12971),
.B(n_12947),
.Y(n_13196)
);

INVx1_ASAP7_75t_L g13197 ( 
.A(n_13012),
.Y(n_13197)
);

INVx1_ASAP7_75t_L g13198 ( 
.A(n_12776),
.Y(n_13198)
);

INVx1_ASAP7_75t_L g13199 ( 
.A(n_12725),
.Y(n_13199)
);

BUFx3_ASAP7_75t_L g13200 ( 
.A(n_12951),
.Y(n_13200)
);

INVx2_ASAP7_75t_L g13201 ( 
.A(n_12942),
.Y(n_13201)
);

INVx1_ASAP7_75t_L g13202 ( 
.A(n_12708),
.Y(n_13202)
);

OA21x2_ASAP7_75t_L g13203 ( 
.A1(n_12672),
.A2(n_1991),
.B(n_1992),
.Y(n_13203)
);

INVx1_ASAP7_75t_SL g13204 ( 
.A(n_12917),
.Y(n_13204)
);

INVx1_ASAP7_75t_L g13205 ( 
.A(n_12712),
.Y(n_13205)
);

INVx2_ASAP7_75t_SL g13206 ( 
.A(n_12928),
.Y(n_13206)
);

AND2x2_ASAP7_75t_L g13207 ( 
.A(n_12669),
.B(n_12972),
.Y(n_13207)
);

AOI22xp33_ASAP7_75t_L g13208 ( 
.A1(n_12795),
.A2(n_12836),
.B1(n_12812),
.B2(n_12704),
.Y(n_13208)
);

AND2x2_ASAP7_75t_L g13209 ( 
.A(n_12956),
.B(n_1993),
.Y(n_13209)
);

INVx1_ASAP7_75t_L g13210 ( 
.A(n_12977),
.Y(n_13210)
);

INVx2_ASAP7_75t_L g13211 ( 
.A(n_12862),
.Y(n_13211)
);

BUFx2_ASAP7_75t_L g13212 ( 
.A(n_12739),
.Y(n_13212)
);

INVx2_ASAP7_75t_L g13213 ( 
.A(n_12801),
.Y(n_13213)
);

NAND2xp5_ASAP7_75t_L g13214 ( 
.A(n_12958),
.B(n_1993),
.Y(n_13214)
);

INVx2_ASAP7_75t_L g13215 ( 
.A(n_12871),
.Y(n_13215)
);

INVxp67_ASAP7_75t_L g13216 ( 
.A(n_12949),
.Y(n_13216)
);

INVx1_ASAP7_75t_L g13217 ( 
.A(n_12985),
.Y(n_13217)
);

INVx2_ASAP7_75t_L g13218 ( 
.A(n_12784),
.Y(n_13218)
);

INVx1_ASAP7_75t_L g13219 ( 
.A(n_12997),
.Y(n_13219)
);

INVx1_ASAP7_75t_L g13220 ( 
.A(n_13007),
.Y(n_13220)
);

NAND2x1_ASAP7_75t_L g13221 ( 
.A(n_12986),
.B(n_1994),
.Y(n_13221)
);

INVxp67_ASAP7_75t_L g13222 ( 
.A(n_12762),
.Y(n_13222)
);

INVx3_ASAP7_75t_L g13223 ( 
.A(n_12823),
.Y(n_13223)
);

INVx1_ASAP7_75t_L g13224 ( 
.A(n_13005),
.Y(n_13224)
);

BUFx2_ASAP7_75t_L g13225 ( 
.A(n_12739),
.Y(n_13225)
);

INVx1_ASAP7_75t_SL g13226 ( 
.A(n_12952),
.Y(n_13226)
);

BUFx2_ASAP7_75t_L g13227 ( 
.A(n_12675),
.Y(n_13227)
);

INVx2_ASAP7_75t_L g13228 ( 
.A(n_12687),
.Y(n_13228)
);

OA21x2_ASAP7_75t_L g13229 ( 
.A1(n_12782),
.A2(n_1994),
.B(n_1995),
.Y(n_13229)
);

NOR2xp33_ASAP7_75t_L g13230 ( 
.A(n_12797),
.B(n_12964),
.Y(n_13230)
);

OAI21x1_ASAP7_75t_L g13231 ( 
.A1(n_12987),
.A2(n_1995),
.B(n_1996),
.Y(n_13231)
);

OAI21x1_ASAP7_75t_L g13232 ( 
.A1(n_12992),
.A2(n_1996),
.B(n_1997),
.Y(n_13232)
);

INVx2_ASAP7_75t_L g13233 ( 
.A(n_12710),
.Y(n_13233)
);

BUFx3_ASAP7_75t_L g13234 ( 
.A(n_12886),
.Y(n_13234)
);

INVx1_ASAP7_75t_L g13235 ( 
.A(n_12938),
.Y(n_13235)
);

AND2x2_ASAP7_75t_L g13236 ( 
.A(n_12830),
.B(n_1997),
.Y(n_13236)
);

INVx3_ASAP7_75t_L g13237 ( 
.A(n_12859),
.Y(n_13237)
);

CKINVDCx5p33_ASAP7_75t_R g13238 ( 
.A(n_12758),
.Y(n_13238)
);

AND2x4_ASAP7_75t_L g13239 ( 
.A(n_13004),
.B(n_1998),
.Y(n_13239)
);

INVx1_ASAP7_75t_L g13240 ( 
.A(n_12788),
.Y(n_13240)
);

INVx1_ASAP7_75t_L g13241 ( 
.A(n_12727),
.Y(n_13241)
);

INVx1_ASAP7_75t_L g13242 ( 
.A(n_12896),
.Y(n_13242)
);

INVx1_ASAP7_75t_L g13243 ( 
.A(n_12998),
.Y(n_13243)
);

INVx1_ASAP7_75t_SL g13244 ( 
.A(n_12701),
.Y(n_13244)
);

NAND2xp5_ASAP7_75t_L g13245 ( 
.A(n_12889),
.B(n_12924),
.Y(n_13245)
);

INVx1_ASAP7_75t_L g13246 ( 
.A(n_13006),
.Y(n_13246)
);

INVx3_ASAP7_75t_L g13247 ( 
.A(n_12916),
.Y(n_13247)
);

INVx3_ASAP7_75t_L g13248 ( 
.A(n_12810),
.Y(n_13248)
);

OA21x2_ASAP7_75t_L g13249 ( 
.A1(n_12702),
.A2(n_1998),
.B(n_1999),
.Y(n_13249)
);

OAI21x1_ASAP7_75t_L g13250 ( 
.A1(n_13011),
.A2(n_1999),
.B(n_2000),
.Y(n_13250)
);

INVx2_ASAP7_75t_SL g13251 ( 
.A(n_12861),
.Y(n_13251)
);

INVx1_ASAP7_75t_L g13252 ( 
.A(n_12904),
.Y(n_13252)
);

INVx1_ASAP7_75t_L g13253 ( 
.A(n_12761),
.Y(n_13253)
);

OAI21x1_ASAP7_75t_L g13254 ( 
.A1(n_12796),
.A2(n_2000),
.B(n_2001),
.Y(n_13254)
);

INVx1_ASAP7_75t_L g13255 ( 
.A(n_12976),
.Y(n_13255)
);

INVx2_ASAP7_75t_L g13256 ( 
.A(n_12875),
.Y(n_13256)
);

INVx2_ASAP7_75t_L g13257 ( 
.A(n_12865),
.Y(n_13257)
);

INVx2_ASAP7_75t_L g13258 ( 
.A(n_12884),
.Y(n_13258)
);

INVx2_ASAP7_75t_L g13259 ( 
.A(n_12816),
.Y(n_13259)
);

HB1xp67_ASAP7_75t_L g13260 ( 
.A(n_12897),
.Y(n_13260)
);

INVx1_ASAP7_75t_L g13261 ( 
.A(n_12979),
.Y(n_13261)
);

INVx2_ASAP7_75t_L g13262 ( 
.A(n_12821),
.Y(n_13262)
);

INVx3_ASAP7_75t_L g13263 ( 
.A(n_12810),
.Y(n_13263)
);

HB1xp67_ASAP7_75t_L g13264 ( 
.A(n_13002),
.Y(n_13264)
);

INVx1_ASAP7_75t_L g13265 ( 
.A(n_12990),
.Y(n_13265)
);

HB1xp67_ASAP7_75t_L g13266 ( 
.A(n_13010),
.Y(n_13266)
);

INVx2_ASAP7_75t_L g13267 ( 
.A(n_12891),
.Y(n_13267)
);

OAI21x1_ASAP7_75t_L g13268 ( 
.A1(n_12756),
.A2(n_2001),
.B(n_2002),
.Y(n_13268)
);

INVx2_ASAP7_75t_L g13269 ( 
.A(n_12915),
.Y(n_13269)
);

INVx1_ASAP7_75t_L g13270 ( 
.A(n_12706),
.Y(n_13270)
);

INVx1_ASAP7_75t_L g13271 ( 
.A(n_12709),
.Y(n_13271)
);

INVx1_ASAP7_75t_L g13272 ( 
.A(n_12790),
.Y(n_13272)
);

INVx2_ASAP7_75t_SL g13273 ( 
.A(n_12717),
.Y(n_13273)
);

INVx1_ASAP7_75t_SL g13274 ( 
.A(n_12860),
.Y(n_13274)
);

AND2x2_ASAP7_75t_L g13275 ( 
.A(n_12892),
.B(n_2002),
.Y(n_13275)
);

AND2x2_ASAP7_75t_L g13276 ( 
.A(n_12879),
.B(n_2003),
.Y(n_13276)
);

INVx2_ASAP7_75t_L g13277 ( 
.A(n_12742),
.Y(n_13277)
);

OA21x2_ASAP7_75t_L g13278 ( 
.A1(n_12815),
.A2(n_12728),
.B(n_12730),
.Y(n_13278)
);

INVx2_ASAP7_75t_SL g13279 ( 
.A(n_12955),
.Y(n_13279)
);

INVx2_ASAP7_75t_L g13280 ( 
.A(n_12748),
.Y(n_13280)
);

INVx1_ASAP7_75t_L g13281 ( 
.A(n_12832),
.Y(n_13281)
);

INVx1_ASAP7_75t_L g13282 ( 
.A(n_12832),
.Y(n_13282)
);

INVx6_ASAP7_75t_L g13283 ( 
.A(n_12984),
.Y(n_13283)
);

INVx2_ASAP7_75t_L g13284 ( 
.A(n_12909),
.Y(n_13284)
);

INVx1_ASAP7_75t_L g13285 ( 
.A(n_13000),
.Y(n_13285)
);

HB1xp67_ASAP7_75t_L g13286 ( 
.A(n_12935),
.Y(n_13286)
);

INVxp67_ASAP7_75t_L g13287 ( 
.A(n_12936),
.Y(n_13287)
);

AO31x2_ASAP7_75t_L g13288 ( 
.A1(n_12737),
.A2(n_2005),
.A3(n_2003),
.B(n_2004),
.Y(n_13288)
);

AO21x2_ASAP7_75t_L g13289 ( 
.A1(n_12688),
.A2(n_2004),
.B(n_2005),
.Y(n_13289)
);

AND2x2_ASAP7_75t_L g13290 ( 
.A(n_12849),
.B(n_2006),
.Y(n_13290)
);

INVx1_ASAP7_75t_L g13291 ( 
.A(n_12746),
.Y(n_13291)
);

AND2x2_ASAP7_75t_L g13292 ( 
.A(n_12773),
.B(n_2006),
.Y(n_13292)
);

OAI21x1_ASAP7_75t_L g13293 ( 
.A1(n_12829),
.A2(n_2007),
.B(n_2008),
.Y(n_13293)
);

INVx3_ASAP7_75t_L g13294 ( 
.A(n_12799),
.Y(n_13294)
);

OAI21xp33_ASAP7_75t_SL g13295 ( 
.A1(n_12720),
.A2(n_2008),
.B(n_2009),
.Y(n_13295)
);

INVx1_ASAP7_75t_L g13296 ( 
.A(n_12746),
.Y(n_13296)
);

AO31x2_ASAP7_75t_L g13297 ( 
.A1(n_12718),
.A2(n_2011),
.A3(n_2009),
.B(n_2010),
.Y(n_13297)
);

AND2x4_ASAP7_75t_L g13298 ( 
.A(n_12807),
.B(n_2012),
.Y(n_13298)
);

OAI21x1_ASAP7_75t_L g13299 ( 
.A1(n_12778),
.A2(n_2012),
.B(n_2013),
.Y(n_13299)
);

OR2x6_ASAP7_75t_L g13300 ( 
.A(n_12781),
.B(n_2013),
.Y(n_13300)
);

INVx1_ASAP7_75t_L g13301 ( 
.A(n_12989),
.Y(n_13301)
);

NOR2xp33_ASAP7_75t_L g13302 ( 
.A(n_12803),
.B(n_2014),
.Y(n_13302)
);

INVx1_ASAP7_75t_L g13303 ( 
.A(n_12996),
.Y(n_13303)
);

AOI22xp33_ASAP7_75t_L g13304 ( 
.A1(n_12707),
.A2(n_2016),
.B1(n_2014),
.B2(n_2015),
.Y(n_13304)
);

HB1xp67_ASAP7_75t_L g13305 ( 
.A(n_12981),
.Y(n_13305)
);

AND2x2_ASAP7_75t_L g13306 ( 
.A(n_12842),
.B(n_2016),
.Y(n_13306)
);

INVx2_ASAP7_75t_L g13307 ( 
.A(n_12993),
.Y(n_13307)
);

INVx3_ASAP7_75t_L g13308 ( 
.A(n_12953),
.Y(n_13308)
);

AND2x2_ASAP7_75t_L g13309 ( 
.A(n_12755),
.B(n_2017),
.Y(n_13309)
);

INVx2_ASAP7_75t_L g13310 ( 
.A(n_12963),
.Y(n_13310)
);

INVx2_ASAP7_75t_L g13311 ( 
.A(n_12968),
.Y(n_13311)
);

INVx1_ASAP7_75t_L g13312 ( 
.A(n_12838),
.Y(n_13312)
);

AOI22xp33_ASAP7_75t_L g13313 ( 
.A1(n_12789),
.A2(n_2019),
.B1(n_2017),
.B2(n_2018),
.Y(n_13313)
);

INVx2_ASAP7_75t_L g13314 ( 
.A(n_12929),
.Y(n_13314)
);

INVx2_ASAP7_75t_L g13315 ( 
.A(n_12933),
.Y(n_13315)
);

NAND2xp5_ASAP7_75t_L g13316 ( 
.A(n_12874),
.B(n_2018),
.Y(n_13316)
);

INVx1_ASAP7_75t_L g13317 ( 
.A(n_12847),
.Y(n_13317)
);

INVx1_ASAP7_75t_L g13318 ( 
.A(n_12873),
.Y(n_13318)
);

INVx1_ASAP7_75t_L g13319 ( 
.A(n_12880),
.Y(n_13319)
);

BUFx2_ASAP7_75t_L g13320 ( 
.A(n_12933),
.Y(n_13320)
);

AND2x2_ASAP7_75t_L g13321 ( 
.A(n_12863),
.B(n_2020),
.Y(n_13321)
);

AND2x2_ASAP7_75t_L g13322 ( 
.A(n_12888),
.B(n_12876),
.Y(n_13322)
);

AO21x1_ASAP7_75t_SL g13323 ( 
.A1(n_12908),
.A2(n_2021),
.B(n_2022),
.Y(n_13323)
);

BUFx2_ASAP7_75t_L g13324 ( 
.A(n_12957),
.Y(n_13324)
);

INVx4_ASAP7_75t_L g13325 ( 
.A(n_12948),
.Y(n_13325)
);

INVx1_ASAP7_75t_L g13326 ( 
.A(n_12911),
.Y(n_13326)
);

INVx2_ASAP7_75t_L g13327 ( 
.A(n_12957),
.Y(n_13327)
);

INVx1_ASAP7_75t_L g13328 ( 
.A(n_12913),
.Y(n_13328)
);

INVx1_ASAP7_75t_L g13329 ( 
.A(n_12930),
.Y(n_13329)
);

INVx1_ASAP7_75t_L g13330 ( 
.A(n_12941),
.Y(n_13330)
);

INVx2_ASAP7_75t_SL g13331 ( 
.A(n_12969),
.Y(n_13331)
);

INVx1_ASAP7_75t_L g13332 ( 
.A(n_12966),
.Y(n_13332)
);

INVxp67_ASAP7_75t_L g13333 ( 
.A(n_12818),
.Y(n_13333)
);

CKINVDCx5p33_ASAP7_75t_R g13334 ( 
.A(n_12869),
.Y(n_13334)
);

INVx1_ASAP7_75t_L g13335 ( 
.A(n_12966),
.Y(n_13335)
);

AND2x2_ASAP7_75t_L g13336 ( 
.A(n_12967),
.B(n_2023),
.Y(n_13336)
);

INVx1_ASAP7_75t_L g13337 ( 
.A(n_12973),
.Y(n_13337)
);

INVx3_ASAP7_75t_L g13338 ( 
.A(n_12973),
.Y(n_13338)
);

OAI21x1_ASAP7_75t_L g13339 ( 
.A1(n_13003),
.A2(n_2023),
.B(n_2024),
.Y(n_13339)
);

INVx1_ASAP7_75t_L g13340 ( 
.A(n_13001),
.Y(n_13340)
);

INVx1_ASAP7_75t_L g13341 ( 
.A(n_13008),
.Y(n_13341)
);

INVx1_ASAP7_75t_L g13342 ( 
.A(n_12713),
.Y(n_13342)
);

INVx3_ASAP7_75t_L g13343 ( 
.A(n_12961),
.Y(n_13343)
);

INVx3_ASAP7_75t_L g13344 ( 
.A(n_12843),
.Y(n_13344)
);

INVx3_ASAP7_75t_L g13345 ( 
.A(n_12690),
.Y(n_13345)
);

INVx1_ASAP7_75t_L g13346 ( 
.A(n_12994),
.Y(n_13346)
);

INVx1_ASAP7_75t_L g13347 ( 
.A(n_12999),
.Y(n_13347)
);

NOR2xp33_ASAP7_75t_L g13348 ( 
.A(n_12740),
.B(n_2024),
.Y(n_13348)
);

AO21x2_ASAP7_75t_L g13349 ( 
.A1(n_12802),
.A2(n_2025),
.B(n_2026),
.Y(n_13349)
);

INVx1_ASAP7_75t_L g13350 ( 
.A(n_12872),
.Y(n_13350)
);

OAI21x1_ASAP7_75t_L g13351 ( 
.A1(n_12845),
.A2(n_12870),
.B(n_12839),
.Y(n_13351)
);

AND2x2_ASAP7_75t_L g13352 ( 
.A(n_12850),
.B(n_12919),
.Y(n_13352)
);

INVx1_ASAP7_75t_L g13353 ( 
.A(n_12962),
.Y(n_13353)
);

INVx1_ASAP7_75t_L g13354 ( 
.A(n_12883),
.Y(n_13354)
);

INVx2_ASAP7_75t_L g13355 ( 
.A(n_12974),
.Y(n_13355)
);

INVx1_ASAP7_75t_L g13356 ( 
.A(n_12932),
.Y(n_13356)
);

BUFx3_ASAP7_75t_L g13357 ( 
.A(n_12995),
.Y(n_13357)
);

HB1xp67_ASAP7_75t_L g13358 ( 
.A(n_12943),
.Y(n_13358)
);

OR2x2_ASAP7_75t_L g13359 ( 
.A(n_12944),
.B(n_2026),
.Y(n_13359)
);

INVx1_ASAP7_75t_L g13360 ( 
.A(n_12982),
.Y(n_13360)
);

AOI22xp33_ASAP7_75t_SL g13361 ( 
.A1(n_12689),
.A2(n_2029),
.B1(n_2027),
.B2(n_2028),
.Y(n_13361)
);

INVx1_ASAP7_75t_L g13362 ( 
.A(n_12667),
.Y(n_13362)
);

OAI221xp5_ASAP7_75t_L g13363 ( 
.A1(n_13208),
.A2(n_2031),
.B1(n_2027),
.B2(n_2030),
.C(n_2032),
.Y(n_13363)
);

OAI22xp5_ASAP7_75t_L g13364 ( 
.A1(n_13190),
.A2(n_2032),
.B1(n_2030),
.B2(n_2031),
.Y(n_13364)
);

AND2x4_ASAP7_75t_L g13365 ( 
.A(n_13200),
.B(n_2033),
.Y(n_13365)
);

AOI22xp33_ASAP7_75t_L g13366 ( 
.A1(n_13360),
.A2(n_2035),
.B1(n_2033),
.B2(n_2034),
.Y(n_13366)
);

AOI22xp33_ASAP7_75t_L g13367 ( 
.A1(n_13358),
.A2(n_2036),
.B1(n_2034),
.B2(n_2035),
.Y(n_13367)
);

INVx4_ASAP7_75t_SL g13368 ( 
.A(n_13043),
.Y(n_13368)
);

AOI22xp33_ASAP7_75t_SL g13369 ( 
.A1(n_13227),
.A2(n_2038),
.B1(n_2036),
.B2(n_2037),
.Y(n_13369)
);

HB1xp67_ASAP7_75t_L g13370 ( 
.A(n_13212),
.Y(n_13370)
);

AOI22xp33_ASAP7_75t_L g13371 ( 
.A1(n_13344),
.A2(n_2041),
.B1(n_2038),
.B2(n_2039),
.Y(n_13371)
);

CKINVDCx5p33_ASAP7_75t_R g13372 ( 
.A(n_13187),
.Y(n_13372)
);

OAI22xp33_ASAP7_75t_L g13373 ( 
.A1(n_13111),
.A2(n_2043),
.B1(n_2039),
.B2(n_2041),
.Y(n_13373)
);

INVx1_ASAP7_75t_L g13374 ( 
.A(n_13030),
.Y(n_13374)
);

AOI22xp33_ASAP7_75t_L g13375 ( 
.A1(n_13345),
.A2(n_2045),
.B1(n_2043),
.B2(n_2044),
.Y(n_13375)
);

OAI22xp33_ASAP7_75t_L g13376 ( 
.A1(n_13245),
.A2(n_2047),
.B1(n_2044),
.B2(n_2046),
.Y(n_13376)
);

OAI211xp5_ASAP7_75t_L g13377 ( 
.A1(n_13222),
.A2(n_2048),
.B(n_2046),
.C(n_2047),
.Y(n_13377)
);

NAND2xp5_ASAP7_75t_L g13378 ( 
.A(n_13343),
.B(n_2048),
.Y(n_13378)
);

OAI22xp33_ASAP7_75t_L g13379 ( 
.A1(n_13138),
.A2(n_2051),
.B1(n_2049),
.B2(n_2050),
.Y(n_13379)
);

AND2x4_ASAP7_75t_L g13380 ( 
.A(n_13048),
.B(n_13114),
.Y(n_13380)
);

INVx5_ASAP7_75t_SL g13381 ( 
.A(n_13043),
.Y(n_13381)
);

INVx2_ASAP7_75t_L g13382 ( 
.A(n_13048),
.Y(n_13382)
);

AOI22xp33_ASAP7_75t_SL g13383 ( 
.A1(n_13305),
.A2(n_2052),
.B1(n_2049),
.B2(n_2050),
.Y(n_13383)
);

AOI221xp5_ASAP7_75t_L g13384 ( 
.A1(n_13118),
.A2(n_2054),
.B1(n_2052),
.B2(n_2053),
.C(n_2055),
.Y(n_13384)
);

AOI22xp33_ASAP7_75t_L g13385 ( 
.A1(n_13357),
.A2(n_2055),
.B1(n_2053),
.B2(n_2054),
.Y(n_13385)
);

OAI21xp33_ASAP7_75t_L g13386 ( 
.A1(n_13064),
.A2(n_2056),
.B(n_2057),
.Y(n_13386)
);

AND2x2_ASAP7_75t_L g13387 ( 
.A(n_13226),
.B(n_2057),
.Y(n_13387)
);

INVx2_ASAP7_75t_SL g13388 ( 
.A(n_13051),
.Y(n_13388)
);

OAI22xp33_ASAP7_75t_L g13389 ( 
.A1(n_13260),
.A2(n_2060),
.B1(n_2058),
.B2(n_2059),
.Y(n_13389)
);

OAI21x1_ASAP7_75t_L g13390 ( 
.A1(n_13069),
.A2(n_2058),
.B(n_2059),
.Y(n_13390)
);

AOI22xp33_ASAP7_75t_L g13391 ( 
.A1(n_13356),
.A2(n_13350),
.B1(n_13347),
.B2(n_13346),
.Y(n_13391)
);

INVx1_ASAP7_75t_L g13392 ( 
.A(n_13061),
.Y(n_13392)
);

INVx1_ASAP7_75t_L g13393 ( 
.A(n_13174),
.Y(n_13393)
);

NOR2xp33_ASAP7_75t_R g13394 ( 
.A(n_13184),
.B(n_2060),
.Y(n_13394)
);

INVx1_ASAP7_75t_L g13395 ( 
.A(n_13170),
.Y(n_13395)
);

OAI221xp5_ASAP7_75t_L g13396 ( 
.A1(n_13316),
.A2(n_2063),
.B1(n_2061),
.B2(n_2062),
.C(n_2064),
.Y(n_13396)
);

INVx1_ASAP7_75t_L g13397 ( 
.A(n_13171),
.Y(n_13397)
);

INVx2_ASAP7_75t_L g13398 ( 
.A(n_13126),
.Y(n_13398)
);

OAI222xp33_ASAP7_75t_L g13399 ( 
.A1(n_13324),
.A2(n_2065),
.B1(n_2067),
.B2(n_2061),
.C1(n_2063),
.C2(n_2066),
.Y(n_13399)
);

OAI221xp5_ASAP7_75t_L g13400 ( 
.A1(n_13032),
.A2(n_2068),
.B1(n_2065),
.B2(n_2067),
.C(n_2069),
.Y(n_13400)
);

NOR2xp33_ASAP7_75t_L g13401 ( 
.A(n_13204),
.B(n_2070),
.Y(n_13401)
);

AOI22xp33_ASAP7_75t_SL g13402 ( 
.A1(n_13127),
.A2(n_2072),
.B1(n_2070),
.B2(n_2071),
.Y(n_13402)
);

AOI22xp33_ASAP7_75t_SL g13403 ( 
.A1(n_13320),
.A2(n_2074),
.B1(n_2072),
.B2(n_2073),
.Y(n_13403)
);

INVx1_ASAP7_75t_L g13404 ( 
.A(n_13142),
.Y(n_13404)
);

AOI22xp33_ASAP7_75t_SL g13405 ( 
.A1(n_13067),
.A2(n_2075),
.B1(n_2073),
.B2(n_2074),
.Y(n_13405)
);

INVx3_ASAP7_75t_L g13406 ( 
.A(n_13177),
.Y(n_13406)
);

OAI21xp5_ASAP7_75t_SL g13407 ( 
.A1(n_13340),
.A2(n_2075),
.B(n_2076),
.Y(n_13407)
);

OAI22xp33_ASAP7_75t_L g13408 ( 
.A1(n_13341),
.A2(n_2078),
.B1(n_2076),
.B2(n_2077),
.Y(n_13408)
);

INVx1_ASAP7_75t_L g13409 ( 
.A(n_13145),
.Y(n_13409)
);

NOR2xp33_ASAP7_75t_L g13410 ( 
.A(n_13040),
.B(n_2077),
.Y(n_13410)
);

OAI22xp5_ASAP7_75t_L g13411 ( 
.A1(n_13334),
.A2(n_13202),
.B1(n_13205),
.B2(n_13197),
.Y(n_13411)
);

AOI22xp5_ASAP7_75t_L g13412 ( 
.A1(n_13035),
.A2(n_2081),
.B1(n_2079),
.B2(n_2080),
.Y(n_13412)
);

AOI22xp33_ASAP7_75t_L g13413 ( 
.A1(n_13330),
.A2(n_2081),
.B1(n_2079),
.B2(n_2080),
.Y(n_13413)
);

INVx4_ASAP7_75t_SL g13414 ( 
.A(n_13175),
.Y(n_13414)
);

OA21x2_ASAP7_75t_L g13415 ( 
.A1(n_13036),
.A2(n_2082),
.B(n_2083),
.Y(n_13415)
);

INVx3_ASAP7_75t_L g13416 ( 
.A(n_13177),
.Y(n_13416)
);

AOI22xp33_ASAP7_75t_L g13417 ( 
.A1(n_13353),
.A2(n_2084),
.B1(n_2082),
.B2(n_2083),
.Y(n_13417)
);

INVx2_ASAP7_75t_L g13418 ( 
.A(n_13095),
.Y(n_13418)
);

AO21x2_ASAP7_75t_L g13419 ( 
.A1(n_13186),
.A2(n_2084),
.B(n_2085),
.Y(n_13419)
);

NAND2xp5_ASAP7_75t_L g13420 ( 
.A(n_13225),
.B(n_2085),
.Y(n_13420)
);

AO21x2_ASAP7_75t_L g13421 ( 
.A1(n_13286),
.A2(n_2086),
.B(n_2087),
.Y(n_13421)
);

NAND2xp5_ASAP7_75t_L g13422 ( 
.A(n_13277),
.B(n_2086),
.Y(n_13422)
);

AOI22xp33_ASAP7_75t_L g13423 ( 
.A1(n_13106),
.A2(n_2090),
.B1(n_2088),
.B2(n_2089),
.Y(n_13423)
);

AND2x4_ASAP7_75t_SL g13424 ( 
.A(n_13073),
.B(n_2089),
.Y(n_13424)
);

OAI211xp5_ASAP7_75t_L g13425 ( 
.A1(n_13143),
.A2(n_2092),
.B(n_2090),
.C(n_2091),
.Y(n_13425)
);

NAND2xp5_ASAP7_75t_L g13426 ( 
.A(n_13216),
.B(n_13273),
.Y(n_13426)
);

OAI22xp33_ASAP7_75t_L g13427 ( 
.A1(n_13057),
.A2(n_2095),
.B1(n_2092),
.B2(n_2094),
.Y(n_13427)
);

INVx1_ASAP7_75t_L g13428 ( 
.A(n_13146),
.Y(n_13428)
);

AOI221xp5_ASAP7_75t_SL g13429 ( 
.A1(n_13192),
.A2(n_2096),
.B1(n_2094),
.B2(n_2095),
.C(n_2097),
.Y(n_13429)
);

AND2x2_ASAP7_75t_L g13430 ( 
.A(n_13110),
.B(n_2097),
.Y(n_13430)
);

OAI211xp5_ASAP7_75t_L g13431 ( 
.A1(n_13361),
.A2(n_2100),
.B(n_2098),
.C(n_2099),
.Y(n_13431)
);

AND2x2_ASAP7_75t_L g13432 ( 
.A(n_13110),
.B(n_2098),
.Y(n_13432)
);

OAI211xp5_ASAP7_75t_SL g13433 ( 
.A1(n_13342),
.A2(n_2101),
.B(n_2099),
.C(n_2100),
.Y(n_13433)
);

OAI22xp5_ASAP7_75t_L g13434 ( 
.A1(n_13294),
.A2(n_2103),
.B1(n_2101),
.B2(n_2102),
.Y(n_13434)
);

INVx8_ASAP7_75t_L g13435 ( 
.A(n_13150),
.Y(n_13435)
);

AND2x2_ASAP7_75t_L g13436 ( 
.A(n_13115),
.B(n_2102),
.Y(n_13436)
);

AOI22xp33_ASAP7_75t_L g13437 ( 
.A1(n_13355),
.A2(n_2106),
.B1(n_2104),
.B2(n_2105),
.Y(n_13437)
);

INVx1_ASAP7_75t_L g13438 ( 
.A(n_13149),
.Y(n_13438)
);

OAI21x1_ASAP7_75t_L g13439 ( 
.A1(n_13094),
.A2(n_2104),
.B(n_2105),
.Y(n_13439)
);

AOI21xp33_ASAP7_75t_L g13440 ( 
.A1(n_13230),
.A2(n_2106),
.B(n_2107),
.Y(n_13440)
);

OAI211xp5_ASAP7_75t_L g13441 ( 
.A1(n_13295),
.A2(n_2109),
.B(n_2107),
.C(n_2108),
.Y(n_13441)
);

AND2x2_ASAP7_75t_L g13442 ( 
.A(n_13195),
.B(n_2108),
.Y(n_13442)
);

AOI21x1_ASAP7_75t_L g13443 ( 
.A1(n_13045),
.A2(n_2110),
.B(n_2111),
.Y(n_13443)
);

INVx2_ASAP7_75t_L g13444 ( 
.A(n_13161),
.Y(n_13444)
);

OAI21x1_ASAP7_75t_L g13445 ( 
.A1(n_13028),
.A2(n_2110),
.B(n_2111),
.Y(n_13445)
);

AOI22xp33_ASAP7_75t_L g13446 ( 
.A1(n_13352),
.A2(n_2114),
.B1(n_2112),
.B2(n_2113),
.Y(n_13446)
);

AOI22xp33_ASAP7_75t_L g13447 ( 
.A1(n_13207),
.A2(n_2114),
.B1(n_2112),
.B2(n_2113),
.Y(n_13447)
);

AO21x1_ASAP7_75t_L g13448 ( 
.A1(n_13159),
.A2(n_2115),
.B(n_2116),
.Y(n_13448)
);

INVx1_ASAP7_75t_L g13449 ( 
.A(n_13056),
.Y(n_13449)
);

HB1xp67_ASAP7_75t_L g13450 ( 
.A(n_13264),
.Y(n_13450)
);

AOI22xp33_ASAP7_75t_SL g13451 ( 
.A1(n_13338),
.A2(n_2117),
.B1(n_2115),
.B2(n_2116),
.Y(n_13451)
);

INVx2_ASAP7_75t_SL g13452 ( 
.A(n_13073),
.Y(n_13452)
);

OAI211xp5_ASAP7_75t_SL g13453 ( 
.A1(n_13354),
.A2(n_2119),
.B(n_2117),
.C(n_2118),
.Y(n_13453)
);

AND2x2_ASAP7_75t_L g13454 ( 
.A(n_13039),
.B(n_2118),
.Y(n_13454)
);

AOI22xp33_ASAP7_75t_SL g13455 ( 
.A1(n_13155),
.A2(n_2121),
.B1(n_2119),
.B2(n_2120),
.Y(n_13455)
);

OR2x2_ASAP7_75t_L g13456 ( 
.A(n_13121),
.B(n_2120),
.Y(n_13456)
);

INVxp67_ASAP7_75t_L g13457 ( 
.A(n_13070),
.Y(n_13457)
);

OAI22xp33_ASAP7_75t_L g13458 ( 
.A1(n_13176),
.A2(n_13152),
.B1(n_13185),
.B2(n_13182),
.Y(n_13458)
);

AOI22xp33_ASAP7_75t_L g13459 ( 
.A1(n_13196),
.A2(n_2123),
.B1(n_2121),
.B2(n_2122),
.Y(n_13459)
);

AND2x4_ASAP7_75t_SL g13460 ( 
.A(n_13108),
.B(n_2122),
.Y(n_13460)
);

INVx1_ASAP7_75t_L g13461 ( 
.A(n_13017),
.Y(n_13461)
);

OR2x2_ASAP7_75t_L g13462 ( 
.A(n_13331),
.B(n_2124),
.Y(n_13462)
);

NAND2xp5_ASAP7_75t_L g13463 ( 
.A(n_13251),
.B(n_2124),
.Y(n_13463)
);

AND2x2_ASAP7_75t_L g13464 ( 
.A(n_13046),
.B(n_2125),
.Y(n_13464)
);

OAI221xp5_ASAP7_75t_L g13465 ( 
.A1(n_13313),
.A2(n_2128),
.B1(n_2126),
.B2(n_2127),
.C(n_2129),
.Y(n_13465)
);

NAND2xp5_ASAP7_75t_L g13466 ( 
.A(n_13274),
.B(n_2126),
.Y(n_13466)
);

AND2x2_ASAP7_75t_L g13467 ( 
.A(n_13248),
.B(n_2127),
.Y(n_13467)
);

AOI22xp33_ASAP7_75t_L g13468 ( 
.A1(n_13050),
.A2(n_2131),
.B1(n_2129),
.B2(n_2130),
.Y(n_13468)
);

OAI211xp5_ASAP7_75t_L g13469 ( 
.A1(n_13085),
.A2(n_2132),
.B(n_2130),
.C(n_2131),
.Y(n_13469)
);

OAI221xp5_ASAP7_75t_L g13470 ( 
.A1(n_13304),
.A2(n_2135),
.B1(n_2133),
.B2(n_2134),
.C(n_2136),
.Y(n_13470)
);

AOI221xp5_ASAP7_75t_L g13471 ( 
.A1(n_13140),
.A2(n_2137),
.B1(n_2133),
.B2(n_2134),
.C(n_2138),
.Y(n_13471)
);

OAI22xp5_ASAP7_75t_L g13472 ( 
.A1(n_13333),
.A2(n_2139),
.B1(n_2137),
.B2(n_2138),
.Y(n_13472)
);

AND2x4_ASAP7_75t_SL g13473 ( 
.A(n_13247),
.B(n_2139),
.Y(n_13473)
);

OAI22xp5_ASAP7_75t_L g13474 ( 
.A1(n_13253),
.A2(n_2142),
.B1(n_2140),
.B2(n_2141),
.Y(n_13474)
);

AND2x2_ASAP7_75t_L g13475 ( 
.A(n_13263),
.B(n_2140),
.Y(n_13475)
);

AOI22xp33_ASAP7_75t_L g13476 ( 
.A1(n_13052),
.A2(n_2143),
.B1(n_2141),
.B2(n_2142),
.Y(n_13476)
);

AOI22xp33_ASAP7_75t_L g13477 ( 
.A1(n_13278),
.A2(n_2145),
.B1(n_2143),
.B2(n_2144),
.Y(n_13477)
);

OAI221xp5_ASAP7_75t_L g13478 ( 
.A1(n_13210),
.A2(n_2147),
.B1(n_2144),
.B2(n_2146),
.C(n_2148),
.Y(n_13478)
);

AOI221xp5_ASAP7_75t_L g13479 ( 
.A1(n_13332),
.A2(n_2150),
.B1(n_2148),
.B2(n_2149),
.C(n_2151),
.Y(n_13479)
);

AOI22xp33_ASAP7_75t_SL g13480 ( 
.A1(n_13351),
.A2(n_2151),
.B1(n_2149),
.B2(n_2150),
.Y(n_13480)
);

OAI22xp33_ASAP7_75t_L g13481 ( 
.A1(n_13335),
.A2(n_2154),
.B1(n_2152),
.B2(n_2153),
.Y(n_13481)
);

OAI22xp5_ASAP7_75t_L g13482 ( 
.A1(n_13049),
.A2(n_2154),
.B1(n_2152),
.B2(n_2153),
.Y(n_13482)
);

AOI22xp5_ASAP7_75t_L g13483 ( 
.A1(n_13093),
.A2(n_2157),
.B1(n_2155),
.B2(n_2156),
.Y(n_13483)
);

OAI21x1_ASAP7_75t_L g13484 ( 
.A1(n_13181),
.A2(n_2155),
.B(n_2156),
.Y(n_13484)
);

OAI22xp5_ASAP7_75t_L g13485 ( 
.A1(n_13244),
.A2(n_13092),
.B1(n_13178),
.B2(n_13098),
.Y(n_13485)
);

AOI221xp5_ASAP7_75t_L g13486 ( 
.A1(n_13337),
.A2(n_2159),
.B1(n_2157),
.B2(n_2158),
.C(n_2160),
.Y(n_13486)
);

NAND3xp33_ASAP7_75t_L g13487 ( 
.A(n_13217),
.B(n_2158),
.C(n_2161),
.Y(n_13487)
);

AND2x4_ASAP7_75t_L g13488 ( 
.A(n_13055),
.B(n_2162),
.Y(n_13488)
);

OAI221xp5_ASAP7_75t_L g13489 ( 
.A1(n_13219),
.A2(n_2164),
.B1(n_2162),
.B2(n_2163),
.C(n_2165),
.Y(n_13489)
);

AOI22xp33_ASAP7_75t_L g13490 ( 
.A1(n_13206),
.A2(n_2165),
.B1(n_2163),
.B2(n_2164),
.Y(n_13490)
);

INVx1_ASAP7_75t_L g13491 ( 
.A(n_13021),
.Y(n_13491)
);

INVx1_ASAP7_75t_SL g13492 ( 
.A(n_13144),
.Y(n_13492)
);

AOI22xp33_ASAP7_75t_SL g13493 ( 
.A1(n_13220),
.A2(n_2168),
.B1(n_2166),
.B2(n_2167),
.Y(n_13493)
);

NAND2xp5_ASAP7_75t_L g13494 ( 
.A(n_13256),
.B(n_2166),
.Y(n_13494)
);

INVx2_ASAP7_75t_L g13495 ( 
.A(n_13161),
.Y(n_13495)
);

AOI222xp33_ASAP7_75t_L g13496 ( 
.A1(n_13148),
.A2(n_2170),
.B1(n_2172),
.B2(n_2168),
.C1(n_2169),
.C2(n_2171),
.Y(n_13496)
);

AOI22xp33_ASAP7_75t_L g13497 ( 
.A1(n_13063),
.A2(n_2172),
.B1(n_2169),
.B2(n_2171),
.Y(n_13497)
);

OR2x2_ASAP7_75t_L g13498 ( 
.A(n_13252),
.B(n_2173),
.Y(n_13498)
);

OR2x6_ASAP7_75t_L g13499 ( 
.A(n_13087),
.B(n_2173),
.Y(n_13499)
);

NAND2xp5_ASAP7_75t_SL g13500 ( 
.A(n_13161),
.B(n_2174),
.Y(n_13500)
);

NOR2x1_ASAP7_75t_R g13501 ( 
.A(n_13234),
.B(n_13325),
.Y(n_13501)
);

INVxp67_ASAP7_75t_L g13502 ( 
.A(n_13102),
.Y(n_13502)
);

AOI22xp5_ASAP7_75t_L g13503 ( 
.A1(n_13289),
.A2(n_2177),
.B1(n_2175),
.B2(n_2176),
.Y(n_13503)
);

AND2x2_ASAP7_75t_L g13504 ( 
.A(n_13201),
.B(n_2176),
.Y(n_13504)
);

NAND2xp5_ASAP7_75t_L g13505 ( 
.A(n_13280),
.B(n_2177),
.Y(n_13505)
);

INVx2_ASAP7_75t_L g13506 ( 
.A(n_13131),
.Y(n_13506)
);

AOI22xp33_ASAP7_75t_L g13507 ( 
.A1(n_13255),
.A2(n_2181),
.B1(n_2178),
.B2(n_2180),
.Y(n_13507)
);

O2A1O1Ixp5_ASAP7_75t_L g13508 ( 
.A1(n_13078),
.A2(n_2181),
.B(n_2178),
.C(n_2180),
.Y(n_13508)
);

AOI22xp33_ASAP7_75t_L g13509 ( 
.A1(n_13261),
.A2(n_2184),
.B1(n_2182),
.B2(n_2183),
.Y(n_13509)
);

OAI22xp5_ASAP7_75t_L g13510 ( 
.A1(n_13060),
.A2(n_2184),
.B1(n_2182),
.B2(n_2183),
.Y(n_13510)
);

INVx3_ASAP7_75t_L g13511 ( 
.A(n_13223),
.Y(n_13511)
);

OAI221xp5_ASAP7_75t_L g13512 ( 
.A1(n_13265),
.A2(n_2187),
.B1(n_2185),
.B2(n_2186),
.C(n_2188),
.Y(n_13512)
);

AND2x2_ASAP7_75t_L g13513 ( 
.A(n_13062),
.B(n_2185),
.Y(n_13513)
);

NOR2xp33_ASAP7_75t_L g13514 ( 
.A(n_13091),
.B(n_2188),
.Y(n_13514)
);

AOI21xp5_ASAP7_75t_L g13515 ( 
.A1(n_13221),
.A2(n_2189),
.B(n_2190),
.Y(n_13515)
);

AOI22xp33_ASAP7_75t_SL g13516 ( 
.A1(n_13275),
.A2(n_2191),
.B1(n_2189),
.B2(n_2190),
.Y(n_13516)
);

INVx2_ASAP7_75t_L g13517 ( 
.A(n_13237),
.Y(n_13517)
);

INVx2_ASAP7_75t_L g13518 ( 
.A(n_13119),
.Y(n_13518)
);

AOI22xp5_ASAP7_75t_L g13519 ( 
.A1(n_13349),
.A2(n_2193),
.B1(n_2191),
.B2(n_2192),
.Y(n_13519)
);

OAI21x1_ASAP7_75t_L g13520 ( 
.A1(n_13165),
.A2(n_2192),
.B(n_2193),
.Y(n_13520)
);

OAI221xp5_ASAP7_75t_L g13521 ( 
.A1(n_13359),
.A2(n_2196),
.B1(n_2194),
.B2(n_2195),
.C(n_2197),
.Y(n_13521)
);

AOI22xp5_ASAP7_75t_L g13522 ( 
.A1(n_13076),
.A2(n_2196),
.B1(n_2194),
.B2(n_2195),
.Y(n_13522)
);

NAND3xp33_ASAP7_75t_L g13523 ( 
.A(n_13072),
.B(n_2198),
.C(n_2199),
.Y(n_13523)
);

AOI221xp5_ASAP7_75t_L g13524 ( 
.A1(n_13291),
.A2(n_2201),
.B1(n_2199),
.B2(n_2200),
.C(n_2202),
.Y(n_13524)
);

AOI221xp5_ASAP7_75t_L g13525 ( 
.A1(n_13296),
.A2(n_2203),
.B1(n_2201),
.B2(n_2202),
.C(n_2204),
.Y(n_13525)
);

AND2x2_ASAP7_75t_L g13526 ( 
.A(n_13068),
.B(n_2203),
.Y(n_13526)
);

AOI221xp5_ASAP7_75t_L g13527 ( 
.A1(n_13284),
.A2(n_13088),
.B1(n_13314),
.B2(n_13327),
.C(n_13315),
.Y(n_13527)
);

BUFx2_ASAP7_75t_L g13528 ( 
.A(n_13266),
.Y(n_13528)
);

OAI22xp5_ASAP7_75t_L g13529 ( 
.A1(n_13083),
.A2(n_2206),
.B1(n_2204),
.B2(n_2205),
.Y(n_13529)
);

AOI22xp5_ASAP7_75t_L g13530 ( 
.A1(n_13348),
.A2(n_2207),
.B1(n_2205),
.B2(n_2206),
.Y(n_13530)
);

INVxp67_ASAP7_75t_SL g13531 ( 
.A(n_13287),
.Y(n_13531)
);

OAI221xp5_ASAP7_75t_L g13532 ( 
.A1(n_13235),
.A2(n_2210),
.B1(n_2208),
.B2(n_2209),
.C(n_2211),
.Y(n_13532)
);

OA21x2_ASAP7_75t_L g13533 ( 
.A1(n_13105),
.A2(n_2208),
.B(n_2210),
.Y(n_13533)
);

OAI22xp5_ASAP7_75t_L g13534 ( 
.A1(n_13203),
.A2(n_2213),
.B1(n_2211),
.B2(n_2212),
.Y(n_13534)
);

OR2x2_ASAP7_75t_L g13535 ( 
.A(n_13129),
.B(n_2212),
.Y(n_13535)
);

OAI211xp5_ASAP7_75t_L g13536 ( 
.A1(n_13130),
.A2(n_2215),
.B(n_2213),
.C(n_2214),
.Y(n_13536)
);

AOI221xp5_ASAP7_75t_L g13537 ( 
.A1(n_13075),
.A2(n_13285),
.B1(n_13172),
.B2(n_13125),
.C(n_13018),
.Y(n_13537)
);

OAI211xp5_ASAP7_75t_L g13538 ( 
.A1(n_13016),
.A2(n_2216),
.B(n_2214),
.C(n_2215),
.Y(n_13538)
);

AOI221xp5_ASAP7_75t_L g13539 ( 
.A1(n_13020),
.A2(n_2218),
.B1(n_2216),
.B2(n_2217),
.C(n_2220),
.Y(n_13539)
);

AND2x2_ASAP7_75t_L g13540 ( 
.A(n_13307),
.B(n_2217),
.Y(n_13540)
);

AOI21xp5_ASAP7_75t_L g13541 ( 
.A1(n_13071),
.A2(n_2218),
.B(n_2220),
.Y(n_13541)
);

NAND2xp5_ASAP7_75t_L g13542 ( 
.A(n_13257),
.B(n_2221),
.Y(n_13542)
);

AOI211xp5_ASAP7_75t_SL g13543 ( 
.A1(n_13151),
.A2(n_2223),
.B(n_2221),
.C(n_2222),
.Y(n_13543)
);

AND2x4_ASAP7_75t_L g13544 ( 
.A(n_13279),
.B(n_2222),
.Y(n_13544)
);

AOI21x1_ASAP7_75t_L g13545 ( 
.A1(n_13042),
.A2(n_2223),
.B(n_2224),
.Y(n_13545)
);

INVx1_ASAP7_75t_L g13546 ( 
.A(n_13024),
.Y(n_13546)
);

AND2x4_ASAP7_75t_L g13547 ( 
.A(n_13269),
.B(n_13267),
.Y(n_13547)
);

OAI22xp5_ASAP7_75t_L g13548 ( 
.A1(n_13283),
.A2(n_2227),
.B1(n_2225),
.B2(n_2226),
.Y(n_13548)
);

BUFx2_ASAP7_75t_L g13549 ( 
.A(n_13027),
.Y(n_13549)
);

AOI22xp33_ASAP7_75t_L g13550 ( 
.A1(n_13300),
.A2(n_2228),
.B1(n_2226),
.B2(n_2227),
.Y(n_13550)
);

OAI22xp5_ASAP7_75t_L g13551 ( 
.A1(n_13300),
.A2(n_2231),
.B1(n_2229),
.B2(n_2230),
.Y(n_13551)
);

OAI21xp5_ASAP7_75t_L g13552 ( 
.A1(n_13029),
.A2(n_13023),
.B(n_13096),
.Y(n_13552)
);

INVx2_ASAP7_75t_L g13553 ( 
.A(n_13033),
.Y(n_13553)
);

NAND3xp33_ASAP7_75t_L g13554 ( 
.A(n_13243),
.B(n_2229),
.C(n_2231),
.Y(n_13554)
);

OAI22xp5_ASAP7_75t_L g13555 ( 
.A1(n_13308),
.A2(n_2235),
.B1(n_2233),
.B2(n_2234),
.Y(n_13555)
);

AOI22xp33_ASAP7_75t_L g13556 ( 
.A1(n_13312),
.A2(n_2236),
.B1(n_2233),
.B2(n_2234),
.Y(n_13556)
);

OAI22xp5_ASAP7_75t_L g13557 ( 
.A1(n_13259),
.A2(n_2238),
.B1(n_2236),
.B2(n_2237),
.Y(n_13557)
);

AOI221xp5_ASAP7_75t_L g13558 ( 
.A1(n_13132),
.A2(n_2239),
.B1(n_2237),
.B2(n_2238),
.C(n_2240),
.Y(n_13558)
);

AND2x2_ASAP7_75t_L g13559 ( 
.A(n_13258),
.B(n_2239),
.Y(n_13559)
);

AND2x2_ASAP7_75t_L g13560 ( 
.A(n_13107),
.B(n_2241),
.Y(n_13560)
);

AOI22xp33_ASAP7_75t_L g13561 ( 
.A1(n_13317),
.A2(n_2243),
.B1(n_2241),
.B2(n_2242),
.Y(n_13561)
);

INVx3_ASAP7_75t_L g13562 ( 
.A(n_13034),
.Y(n_13562)
);

OAI211xp5_ASAP7_75t_L g13563 ( 
.A1(n_13103),
.A2(n_2244),
.B(n_2242),
.C(n_2243),
.Y(n_13563)
);

AOI22xp5_ASAP7_75t_L g13564 ( 
.A1(n_13148),
.A2(n_2246),
.B1(n_2244),
.B2(n_2245),
.Y(n_13564)
);

INVx2_ASAP7_75t_L g13565 ( 
.A(n_13065),
.Y(n_13565)
);

OAI22x1_ASAP7_75t_L g13566 ( 
.A1(n_13262),
.A2(n_13271),
.B1(n_13270),
.B2(n_13239),
.Y(n_13566)
);

AOI22xp33_ASAP7_75t_L g13567 ( 
.A1(n_13318),
.A2(n_2247),
.B1(n_2245),
.B2(n_2246),
.Y(n_13567)
);

INVx1_ASAP7_75t_L g13568 ( 
.A(n_13026),
.Y(n_13568)
);

INVx1_ASAP7_75t_L g13569 ( 
.A(n_13031),
.Y(n_13569)
);

NAND2xp5_ASAP7_75t_SL g13570 ( 
.A(n_13322),
.B(n_2247),
.Y(n_13570)
);

OAI21x1_ASAP7_75t_L g13571 ( 
.A1(n_13117),
.A2(n_2249),
.B(n_2250),
.Y(n_13571)
);

OAI22xp5_ASAP7_75t_L g13572 ( 
.A1(n_13218),
.A2(n_2251),
.B1(n_2249),
.B2(n_2250),
.Y(n_13572)
);

AOI221xp5_ASAP7_75t_L g13573 ( 
.A1(n_13100),
.A2(n_2254),
.B1(n_2251),
.B2(n_2252),
.C(n_2255),
.Y(n_13573)
);

BUFx4f_ASAP7_75t_L g13574 ( 
.A(n_13025),
.Y(n_13574)
);

HB1xp67_ASAP7_75t_L g13575 ( 
.A(n_13281),
.Y(n_13575)
);

AOI21xp5_ASAP7_75t_L g13576 ( 
.A1(n_13164),
.A2(n_13113),
.B(n_13134),
.Y(n_13576)
);

OAI22xp33_ASAP7_75t_L g13577 ( 
.A1(n_13213),
.A2(n_2257),
.B1(n_2255),
.B2(n_2256),
.Y(n_13577)
);

OAI211xp5_ASAP7_75t_L g13578 ( 
.A1(n_13336),
.A2(n_13290),
.B(n_13276),
.C(n_13229),
.Y(n_13578)
);

AOI22xp33_ASAP7_75t_SL g13579 ( 
.A1(n_13311),
.A2(n_2259),
.B1(n_2256),
.B2(n_2258),
.Y(n_13579)
);

AOI21xp5_ASAP7_75t_SL g13580 ( 
.A1(n_13298),
.A2(n_2258),
.B(n_2259),
.Y(n_13580)
);

AND2x2_ASAP7_75t_L g13581 ( 
.A(n_13326),
.B(n_2260),
.Y(n_13581)
);

AND2x4_ASAP7_75t_L g13582 ( 
.A(n_13047),
.B(n_2262),
.Y(n_13582)
);

AOI22xp33_ASAP7_75t_L g13583 ( 
.A1(n_13319),
.A2(n_2264),
.B1(n_2262),
.B2(n_2263),
.Y(n_13583)
);

NAND2xp5_ASAP7_75t_L g13584 ( 
.A(n_13249),
.B(n_2263),
.Y(n_13584)
);

AOI22xp33_ASAP7_75t_L g13585 ( 
.A1(n_13329),
.A2(n_2266),
.B1(n_2264),
.B2(n_2265),
.Y(n_13585)
);

AOI22xp33_ASAP7_75t_L g13586 ( 
.A1(n_13328),
.A2(n_2267),
.B1(n_2265),
.B2(n_2266),
.Y(n_13586)
);

AND2x2_ASAP7_75t_L g13587 ( 
.A(n_13241),
.B(n_13272),
.Y(n_13587)
);

OAI22xp5_ASAP7_75t_L g13588 ( 
.A1(n_13188),
.A2(n_2269),
.B1(n_2267),
.B2(n_2268),
.Y(n_13588)
);

AND2x2_ASAP7_75t_L g13589 ( 
.A(n_13022),
.B(n_13199),
.Y(n_13589)
);

AND2x2_ASAP7_75t_L g13590 ( 
.A(n_13233),
.B(n_13116),
.Y(n_13590)
);

OAI21x1_ASAP7_75t_L g13591 ( 
.A1(n_13224),
.A2(n_2268),
.B(n_2269),
.Y(n_13591)
);

INVx1_ASAP7_75t_L g13592 ( 
.A(n_13037),
.Y(n_13592)
);

INVx1_ASAP7_75t_L g13593 ( 
.A(n_13038),
.Y(n_13593)
);

AOI22xp33_ASAP7_75t_L g13594 ( 
.A1(n_13310),
.A2(n_2273),
.B1(n_2270),
.B2(n_2271),
.Y(n_13594)
);

OAI22xp5_ASAP7_75t_L g13595 ( 
.A1(n_13191),
.A2(n_2273),
.B1(n_2270),
.B2(n_2271),
.Y(n_13595)
);

OAI22xp33_ASAP7_75t_L g13596 ( 
.A1(n_13242),
.A2(n_2276),
.B1(n_2274),
.B2(n_2275),
.Y(n_13596)
);

INVx1_ASAP7_75t_L g13597 ( 
.A(n_13041),
.Y(n_13597)
);

AOI22xp5_ASAP7_75t_L g13598 ( 
.A1(n_13211),
.A2(n_2277),
.B1(n_2274),
.B2(n_2275),
.Y(n_13598)
);

AOI21xp5_ASAP7_75t_L g13599 ( 
.A1(n_13137),
.A2(n_2277),
.B(n_2278),
.Y(n_13599)
);

INVx1_ASAP7_75t_L g13600 ( 
.A(n_13044),
.Y(n_13600)
);

OAI22xp33_ASAP7_75t_L g13601 ( 
.A1(n_13228),
.A2(n_2280),
.B1(n_2278),
.B2(n_2279),
.Y(n_13601)
);

INVx1_ASAP7_75t_L g13602 ( 
.A(n_13053),
.Y(n_13602)
);

OA21x2_ASAP7_75t_L g13603 ( 
.A1(n_13282),
.A2(n_2280),
.B(n_2281),
.Y(n_13603)
);

OR2x2_ASAP7_75t_L g13604 ( 
.A(n_13015),
.B(n_2281),
.Y(n_13604)
);

AOI22xp33_ASAP7_75t_SL g13605 ( 
.A1(n_13301),
.A2(n_2284),
.B1(n_2282),
.B2(n_2283),
.Y(n_13605)
);

AOI22xp33_ASAP7_75t_SL g13606 ( 
.A1(n_13303),
.A2(n_2286),
.B1(n_2284),
.B2(n_2285),
.Y(n_13606)
);

OAI22xp5_ASAP7_75t_L g13607 ( 
.A1(n_13193),
.A2(n_2287),
.B1(n_2285),
.B2(n_2286),
.Y(n_13607)
);

AOI222xp33_ASAP7_75t_L g13608 ( 
.A1(n_13302),
.A2(n_2289),
.B1(n_2291),
.B2(n_2287),
.C1(n_2288),
.C2(n_2290),
.Y(n_13608)
);

AO31x2_ASAP7_75t_L g13609 ( 
.A1(n_13173),
.A2(n_2291),
.A3(n_2289),
.B(n_2290),
.Y(n_13609)
);

INVx1_ASAP7_75t_SL g13610 ( 
.A(n_13120),
.Y(n_13610)
);

NAND2xp5_ASAP7_75t_L g13611 ( 
.A(n_13240),
.B(n_2292),
.Y(n_13611)
);

AND2x2_ASAP7_75t_L g13612 ( 
.A(n_13112),
.B(n_2292),
.Y(n_13612)
);

NAND3xp33_ASAP7_75t_L g13613 ( 
.A(n_13246),
.B(n_2293),
.C(n_2294),
.Y(n_13613)
);

OAI22xp33_ASAP7_75t_L g13614 ( 
.A1(n_13194),
.A2(n_2295),
.B1(n_2293),
.B2(n_2294),
.Y(n_13614)
);

INVx2_ASAP7_75t_SL g13615 ( 
.A(n_13238),
.Y(n_13615)
);

AOI22xp33_ASAP7_75t_L g13616 ( 
.A1(n_13215),
.A2(n_13179),
.B1(n_13198),
.B2(n_13180),
.Y(n_13616)
);

INVx1_ASAP7_75t_L g13617 ( 
.A(n_13054),
.Y(n_13617)
);

AND2x2_ASAP7_75t_L g13618 ( 
.A(n_13066),
.B(n_2296),
.Y(n_13618)
);

AOI22xp33_ASAP7_75t_L g13619 ( 
.A1(n_13183),
.A2(n_2299),
.B1(n_2297),
.B2(n_2298),
.Y(n_13619)
);

INVx2_ASAP7_75t_L g13620 ( 
.A(n_13157),
.Y(n_13620)
);

INVx2_ASAP7_75t_SL g13621 ( 
.A(n_13380),
.Y(n_13621)
);

AND2x2_ASAP7_75t_L g13622 ( 
.A(n_13382),
.B(n_13158),
.Y(n_13622)
);

AND2x4_ASAP7_75t_L g13623 ( 
.A(n_13388),
.B(n_13141),
.Y(n_13623)
);

INVx2_ASAP7_75t_L g13624 ( 
.A(n_13528),
.Y(n_13624)
);

INVx1_ASAP7_75t_L g13625 ( 
.A(n_13450),
.Y(n_13625)
);

BUFx3_ASAP7_75t_L g13626 ( 
.A(n_13435),
.Y(n_13626)
);

AND2x2_ASAP7_75t_L g13627 ( 
.A(n_13531),
.B(n_13574),
.Y(n_13627)
);

INVx1_ASAP7_75t_L g13628 ( 
.A(n_13575),
.Y(n_13628)
);

INVx2_ASAP7_75t_L g13629 ( 
.A(n_13406),
.Y(n_13629)
);

CKINVDCx6p67_ASAP7_75t_R g13630 ( 
.A(n_13499),
.Y(n_13630)
);

INVx2_ASAP7_75t_SL g13631 ( 
.A(n_13435),
.Y(n_13631)
);

NAND2xp5_ASAP7_75t_L g13632 ( 
.A(n_13370),
.B(n_13209),
.Y(n_13632)
);

BUFx2_ASAP7_75t_L g13633 ( 
.A(n_13501),
.Y(n_13633)
);

AND2x2_ASAP7_75t_L g13634 ( 
.A(n_13492),
.B(n_13163),
.Y(n_13634)
);

AND2x2_ASAP7_75t_L g13635 ( 
.A(n_13416),
.B(n_13321),
.Y(n_13635)
);

INVx1_ASAP7_75t_L g13636 ( 
.A(n_13374),
.Y(n_13636)
);

INVx2_ASAP7_75t_SL g13637 ( 
.A(n_13368),
.Y(n_13637)
);

INVxp67_ASAP7_75t_L g13638 ( 
.A(n_13419),
.Y(n_13638)
);

INVx2_ASAP7_75t_L g13639 ( 
.A(n_13452),
.Y(n_13639)
);

AND2x2_ASAP7_75t_L g13640 ( 
.A(n_13511),
.B(n_13398),
.Y(n_13640)
);

INVxp67_ASAP7_75t_L g13641 ( 
.A(n_13421),
.Y(n_13641)
);

AND2x2_ASAP7_75t_L g13642 ( 
.A(n_13418),
.B(n_13506),
.Y(n_13642)
);

INVx3_ASAP7_75t_L g13643 ( 
.A(n_13381),
.Y(n_13643)
);

INVx2_ASAP7_75t_L g13644 ( 
.A(n_13372),
.Y(n_13644)
);

AOI22xp33_ASAP7_75t_L g13645 ( 
.A1(n_13391),
.A2(n_13154),
.B1(n_13156),
.B2(n_13153),
.Y(n_13645)
);

INVx2_ASAP7_75t_L g13646 ( 
.A(n_13517),
.Y(n_13646)
);

INVxp33_ASAP7_75t_L g13647 ( 
.A(n_13394),
.Y(n_13647)
);

INVx1_ASAP7_75t_L g13648 ( 
.A(n_13449),
.Y(n_13648)
);

NOR2xp33_ASAP7_75t_L g13649 ( 
.A(n_13381),
.B(n_13019),
.Y(n_13649)
);

INVx3_ASAP7_75t_SL g13650 ( 
.A(n_13368),
.Y(n_13650)
);

NAND2xp5_ASAP7_75t_L g13651 ( 
.A(n_13455),
.B(n_13610),
.Y(n_13651)
);

OR2x2_ASAP7_75t_L g13652 ( 
.A(n_13518),
.B(n_13160),
.Y(n_13652)
);

OR2x2_ASAP7_75t_L g13653 ( 
.A(n_13426),
.B(n_13162),
.Y(n_13653)
);

AND2x2_ASAP7_75t_L g13654 ( 
.A(n_13589),
.B(n_13292),
.Y(n_13654)
);

AND2x2_ASAP7_75t_L g13655 ( 
.A(n_13615),
.B(n_13306),
.Y(n_13655)
);

BUFx6f_ASAP7_75t_L g13656 ( 
.A(n_13365),
.Y(n_13656)
);

AOI22xp33_ASAP7_75t_L g13657 ( 
.A1(n_13411),
.A2(n_13167),
.B1(n_13169),
.B2(n_13166),
.Y(n_13657)
);

AND2x2_ASAP7_75t_L g13658 ( 
.A(n_13547),
.B(n_13309),
.Y(n_13658)
);

INVx2_ASAP7_75t_L g13659 ( 
.A(n_13387),
.Y(n_13659)
);

NAND2xp5_ASAP7_75t_L g13660 ( 
.A(n_13480),
.B(n_13175),
.Y(n_13660)
);

INVx1_ASAP7_75t_L g13661 ( 
.A(n_13392),
.Y(n_13661)
);

AND2x2_ASAP7_75t_L g13662 ( 
.A(n_13430),
.B(n_13147),
.Y(n_13662)
);

AND2x2_ASAP7_75t_L g13663 ( 
.A(n_13432),
.B(n_13236),
.Y(n_13663)
);

NAND2xp5_ASAP7_75t_L g13664 ( 
.A(n_13376),
.B(n_13457),
.Y(n_13664)
);

AND2x2_ASAP7_75t_L g13665 ( 
.A(n_13552),
.B(n_13074),
.Y(n_13665)
);

HB1xp67_ASAP7_75t_L g13666 ( 
.A(n_13414),
.Y(n_13666)
);

NAND2xp5_ASAP7_75t_L g13667 ( 
.A(n_13502),
.B(n_13168),
.Y(n_13667)
);

AND2x2_ASAP7_75t_L g13668 ( 
.A(n_13587),
.B(n_13089),
.Y(n_13668)
);

BUFx2_ASAP7_75t_L g13669 ( 
.A(n_13499),
.Y(n_13669)
);

INVx2_ASAP7_75t_L g13670 ( 
.A(n_13467),
.Y(n_13670)
);

INVx2_ASAP7_75t_L g13671 ( 
.A(n_13475),
.Y(n_13671)
);

INVx1_ASAP7_75t_L g13672 ( 
.A(n_13535),
.Y(n_13672)
);

INVx2_ASAP7_75t_L g13673 ( 
.A(n_13444),
.Y(n_13673)
);

INVx2_ASAP7_75t_L g13674 ( 
.A(n_13495),
.Y(n_13674)
);

INVx3_ASAP7_75t_L g13675 ( 
.A(n_13544),
.Y(n_13675)
);

OR2x2_ASAP7_75t_L g13676 ( 
.A(n_13494),
.B(n_13139),
.Y(n_13676)
);

HB1xp67_ASAP7_75t_L g13677 ( 
.A(n_13414),
.Y(n_13677)
);

INVx2_ASAP7_75t_SL g13678 ( 
.A(n_13460),
.Y(n_13678)
);

INVx2_ASAP7_75t_L g13679 ( 
.A(n_13549),
.Y(n_13679)
);

INVx2_ASAP7_75t_L g13680 ( 
.A(n_13562),
.Y(n_13680)
);

NAND2xp5_ASAP7_75t_L g13681 ( 
.A(n_13407),
.B(n_13288),
.Y(n_13681)
);

AND2x2_ASAP7_75t_L g13682 ( 
.A(n_13590),
.B(n_13099),
.Y(n_13682)
);

OAI21xp5_ASAP7_75t_L g13683 ( 
.A1(n_13508),
.A2(n_13293),
.B(n_13268),
.Y(n_13683)
);

NOR2xp33_ASAP7_75t_L g13684 ( 
.A(n_13578),
.B(n_13214),
.Y(n_13684)
);

AND2x2_ASAP7_75t_L g13685 ( 
.A(n_13485),
.B(n_13133),
.Y(n_13685)
);

INVx3_ASAP7_75t_L g13686 ( 
.A(n_13488),
.Y(n_13686)
);

AND2x2_ASAP7_75t_L g13687 ( 
.A(n_13436),
.B(n_13135),
.Y(n_13687)
);

INVx4_ASAP7_75t_L g13688 ( 
.A(n_13424),
.Y(n_13688)
);

INVx3_ASAP7_75t_L g13689 ( 
.A(n_13582),
.Y(n_13689)
);

BUFx2_ASAP7_75t_L g13690 ( 
.A(n_13415),
.Y(n_13690)
);

AND2x2_ASAP7_75t_L g13691 ( 
.A(n_13566),
.B(n_13136),
.Y(n_13691)
);

INVx1_ASAP7_75t_L g13692 ( 
.A(n_13462),
.Y(n_13692)
);

INVxp67_ASAP7_75t_L g13693 ( 
.A(n_13410),
.Y(n_13693)
);

OR2x2_ASAP7_75t_L g13694 ( 
.A(n_13456),
.B(n_13122),
.Y(n_13694)
);

BUFx2_ASAP7_75t_L g13695 ( 
.A(n_13415),
.Y(n_13695)
);

INVx2_ASAP7_75t_L g13696 ( 
.A(n_13560),
.Y(n_13696)
);

BUFx3_ASAP7_75t_L g13697 ( 
.A(n_13473),
.Y(n_13697)
);

AND2x2_ASAP7_75t_L g13698 ( 
.A(n_13513),
.B(n_13299),
.Y(n_13698)
);

INVx1_ASAP7_75t_L g13699 ( 
.A(n_13393),
.Y(n_13699)
);

INVxp67_ASAP7_75t_L g13700 ( 
.A(n_13500),
.Y(n_13700)
);

HB1xp67_ASAP7_75t_L g13701 ( 
.A(n_13603),
.Y(n_13701)
);

INVx2_ASAP7_75t_L g13702 ( 
.A(n_13526),
.Y(n_13702)
);

AND2x2_ASAP7_75t_L g13703 ( 
.A(n_13565),
.B(n_13104),
.Y(n_13703)
);

AND2x2_ASAP7_75t_L g13704 ( 
.A(n_13553),
.B(n_13109),
.Y(n_13704)
);

AND2x2_ASAP7_75t_L g13705 ( 
.A(n_13618),
.B(n_13124),
.Y(n_13705)
);

INVx1_ASAP7_75t_L g13706 ( 
.A(n_13395),
.Y(n_13706)
);

INVx1_ASAP7_75t_L g13707 ( 
.A(n_13397),
.Y(n_13707)
);

NAND2xp5_ASAP7_75t_L g13708 ( 
.A(n_13477),
.B(n_13288),
.Y(n_13708)
);

AND2x2_ASAP7_75t_L g13709 ( 
.A(n_13442),
.B(n_13128),
.Y(n_13709)
);

INVx1_ASAP7_75t_L g13710 ( 
.A(n_13404),
.Y(n_13710)
);

AO21x2_ASAP7_75t_L g13711 ( 
.A1(n_13458),
.A2(n_13059),
.B(n_13058),
.Y(n_13711)
);

INVx2_ASAP7_75t_SL g13712 ( 
.A(n_13454),
.Y(n_13712)
);

INVx1_ASAP7_75t_L g13713 ( 
.A(n_13409),
.Y(n_13713)
);

INVx2_ASAP7_75t_SL g13714 ( 
.A(n_13464),
.Y(n_13714)
);

AND2x2_ASAP7_75t_L g13715 ( 
.A(n_13581),
.B(n_13079),
.Y(n_13715)
);

INVx2_ASAP7_75t_L g13716 ( 
.A(n_13559),
.Y(n_13716)
);

INVx1_ASAP7_75t_L g13717 ( 
.A(n_13428),
.Y(n_13717)
);

BUFx3_ASAP7_75t_L g13718 ( 
.A(n_13504),
.Y(n_13718)
);

INVx1_ASAP7_75t_L g13719 ( 
.A(n_13438),
.Y(n_13719)
);

OR2x2_ASAP7_75t_L g13720 ( 
.A(n_13420),
.B(n_13080),
.Y(n_13720)
);

HB1xp67_ASAP7_75t_L g13721 ( 
.A(n_13603),
.Y(n_13721)
);

BUFx2_ASAP7_75t_SL g13722 ( 
.A(n_13448),
.Y(n_13722)
);

INVx1_ASAP7_75t_L g13723 ( 
.A(n_13461),
.Y(n_13723)
);

AND2x2_ASAP7_75t_L g13724 ( 
.A(n_13612),
.B(n_13081),
.Y(n_13724)
);

NAND2xp5_ASAP7_75t_L g13725 ( 
.A(n_13599),
.B(n_13082),
.Y(n_13725)
);

AND2x2_ASAP7_75t_L g13726 ( 
.A(n_13540),
.B(n_13086),
.Y(n_13726)
);

AND2x2_ASAP7_75t_L g13727 ( 
.A(n_13620),
.B(n_13090),
.Y(n_13727)
);

INVx1_ASAP7_75t_L g13728 ( 
.A(n_13491),
.Y(n_13728)
);

HB1xp67_ASAP7_75t_L g13729 ( 
.A(n_13390),
.Y(n_13729)
);

OR2x2_ASAP7_75t_L g13730 ( 
.A(n_13505),
.B(n_13097),
.Y(n_13730)
);

INVx2_ASAP7_75t_L g13731 ( 
.A(n_13484),
.Y(n_13731)
);

INVx2_ASAP7_75t_L g13732 ( 
.A(n_13520),
.Y(n_13732)
);

INVx1_ASAP7_75t_L g13733 ( 
.A(n_13546),
.Y(n_13733)
);

INVx1_ASAP7_75t_L g13734 ( 
.A(n_13568),
.Y(n_13734)
);

INVx1_ASAP7_75t_L g13735 ( 
.A(n_13569),
.Y(n_13735)
);

INVx1_ASAP7_75t_L g13736 ( 
.A(n_13592),
.Y(n_13736)
);

INVx1_ASAP7_75t_L g13737 ( 
.A(n_13593),
.Y(n_13737)
);

HB1xp67_ASAP7_75t_L g13738 ( 
.A(n_13443),
.Y(n_13738)
);

AND2x2_ASAP7_75t_L g13739 ( 
.A(n_13445),
.B(n_13101),
.Y(n_13739)
);

INVx1_ASAP7_75t_L g13740 ( 
.A(n_13597),
.Y(n_13740)
);

AND2x2_ASAP7_75t_L g13741 ( 
.A(n_13401),
.B(n_13362),
.Y(n_13741)
);

AO21x2_ASAP7_75t_L g13742 ( 
.A1(n_13373),
.A2(n_13189),
.B(n_13123),
.Y(n_13742)
);

AND2x2_ASAP7_75t_L g13743 ( 
.A(n_13514),
.B(n_13077),
.Y(n_13743)
);

INVx1_ASAP7_75t_L g13744 ( 
.A(n_13600),
.Y(n_13744)
);

INVxp67_ASAP7_75t_SL g13745 ( 
.A(n_13570),
.Y(n_13745)
);

INVxp67_ASAP7_75t_SL g13746 ( 
.A(n_13533),
.Y(n_13746)
);

AND2x2_ASAP7_75t_L g13747 ( 
.A(n_13616),
.B(n_13231),
.Y(n_13747)
);

INVx1_ASAP7_75t_L g13748 ( 
.A(n_13602),
.Y(n_13748)
);

AND2x4_ASAP7_75t_SL g13749 ( 
.A(n_13503),
.B(n_13323),
.Y(n_13749)
);

INVx1_ASAP7_75t_L g13750 ( 
.A(n_13617),
.Y(n_13750)
);

AND2x2_ASAP7_75t_L g13751 ( 
.A(n_13533),
.B(n_13542),
.Y(n_13751)
);

AND2x4_ASAP7_75t_L g13752 ( 
.A(n_13463),
.B(n_13232),
.Y(n_13752)
);

OAI22xp5_ASAP7_75t_L g13753 ( 
.A1(n_13412),
.A2(n_13297),
.B1(n_13339),
.B2(n_13250),
.Y(n_13753)
);

INVx1_ASAP7_75t_L g13754 ( 
.A(n_13498),
.Y(n_13754)
);

INVx2_ASAP7_75t_L g13755 ( 
.A(n_13604),
.Y(n_13755)
);

INVx2_ASAP7_75t_L g13756 ( 
.A(n_13571),
.Y(n_13756)
);

AND2x2_ASAP7_75t_L g13757 ( 
.A(n_13576),
.B(n_13084),
.Y(n_13757)
);

BUFx6f_ASAP7_75t_L g13758 ( 
.A(n_13466),
.Y(n_13758)
);

INVx2_ASAP7_75t_L g13759 ( 
.A(n_13591),
.Y(n_13759)
);

NAND2xp5_ASAP7_75t_L g13760 ( 
.A(n_13541),
.B(n_13297),
.Y(n_13760)
);

AND2x2_ASAP7_75t_L g13761 ( 
.A(n_13611),
.B(n_13254),
.Y(n_13761)
);

OR2x6_ASAP7_75t_L g13762 ( 
.A(n_13580),
.B(n_2297),
.Y(n_13762)
);

AND2x2_ASAP7_75t_L g13763 ( 
.A(n_13422),
.B(n_2298),
.Y(n_13763)
);

INVxp33_ASAP7_75t_SL g13764 ( 
.A(n_13364),
.Y(n_13764)
);

AND2x2_ASAP7_75t_L g13765 ( 
.A(n_13527),
.B(n_2299),
.Y(n_13765)
);

INVx2_ASAP7_75t_L g13766 ( 
.A(n_13439),
.Y(n_13766)
);

INVx1_ASAP7_75t_L g13767 ( 
.A(n_13609),
.Y(n_13767)
);

INVx4_ASAP7_75t_L g13768 ( 
.A(n_13378),
.Y(n_13768)
);

AND2x2_ASAP7_75t_L g13769 ( 
.A(n_13537),
.B(n_2300),
.Y(n_13769)
);

BUFx3_ASAP7_75t_L g13770 ( 
.A(n_13584),
.Y(n_13770)
);

OR2x2_ASAP7_75t_L g13771 ( 
.A(n_13534),
.B(n_2301),
.Y(n_13771)
);

BUFx2_ASAP7_75t_L g13772 ( 
.A(n_13609),
.Y(n_13772)
);

OR2x2_ASAP7_75t_L g13773 ( 
.A(n_13523),
.B(n_2301),
.Y(n_13773)
);

AND2x2_ASAP7_75t_L g13774 ( 
.A(n_13516),
.B(n_2302),
.Y(n_13774)
);

AND2x2_ASAP7_75t_L g13775 ( 
.A(n_13459),
.B(n_2302),
.Y(n_13775)
);

OR2x2_ASAP7_75t_L g13776 ( 
.A(n_13554),
.B(n_2303),
.Y(n_13776)
);

NAND2xp5_ASAP7_75t_L g13777 ( 
.A(n_13536),
.B(n_2303),
.Y(n_13777)
);

AND2x4_ASAP7_75t_L g13778 ( 
.A(n_13487),
.B(n_2304),
.Y(n_13778)
);

HB1xp67_ASAP7_75t_L g13779 ( 
.A(n_13545),
.Y(n_13779)
);

INVx1_ASAP7_75t_L g13780 ( 
.A(n_13613),
.Y(n_13780)
);

INVxp67_ASAP7_75t_SL g13781 ( 
.A(n_13515),
.Y(n_13781)
);

NAND2xp5_ASAP7_75t_L g13782 ( 
.A(n_13389),
.B(n_2304),
.Y(n_13782)
);

INVx1_ASAP7_75t_L g13783 ( 
.A(n_13555),
.Y(n_13783)
);

OR2x2_ASAP7_75t_L g13784 ( 
.A(n_13519),
.B(n_2305),
.Y(n_13784)
);

AND2x4_ASAP7_75t_L g13785 ( 
.A(n_13564),
.B(n_2305),
.Y(n_13785)
);

AND2x2_ASAP7_75t_L g13786 ( 
.A(n_13369),
.B(n_2306),
.Y(n_13786)
);

INVx3_ASAP7_75t_L g13787 ( 
.A(n_13399),
.Y(n_13787)
);

INVxp67_ASAP7_75t_L g13788 ( 
.A(n_13377),
.Y(n_13788)
);

OR2x2_ASAP7_75t_L g13789 ( 
.A(n_13386),
.B(n_2306),
.Y(n_13789)
);

AND2x2_ASAP7_75t_L g13790 ( 
.A(n_13366),
.B(n_2307),
.Y(n_13790)
);

INVx2_ASAP7_75t_L g13791 ( 
.A(n_13483),
.Y(n_13791)
);

BUFx3_ASAP7_75t_L g13792 ( 
.A(n_13521),
.Y(n_13792)
);

OR2x2_ASAP7_75t_L g13793 ( 
.A(n_13557),
.B(n_2308),
.Y(n_13793)
);

BUFx3_ASAP7_75t_L g13794 ( 
.A(n_13530),
.Y(n_13794)
);

NAND2xp5_ASAP7_75t_L g13795 ( 
.A(n_13496),
.B(n_2308),
.Y(n_13795)
);

INVx2_ASAP7_75t_L g13796 ( 
.A(n_13598),
.Y(n_13796)
);

AND2x2_ASAP7_75t_L g13797 ( 
.A(n_13437),
.B(n_2309),
.Y(n_13797)
);

BUFx3_ASAP7_75t_L g13798 ( 
.A(n_13396),
.Y(n_13798)
);

INVx1_ASAP7_75t_L g13799 ( 
.A(n_13474),
.Y(n_13799)
);

OR2x2_ASAP7_75t_L g13800 ( 
.A(n_13434),
.B(n_2310),
.Y(n_13800)
);

AND2x2_ASAP7_75t_L g13801 ( 
.A(n_13367),
.B(n_2310),
.Y(n_13801)
);

NAND2xp5_ASAP7_75t_L g13802 ( 
.A(n_13379),
.B(n_2311),
.Y(n_13802)
);

AND2x4_ASAP7_75t_SL g13803 ( 
.A(n_13550),
.B(n_2312),
.Y(n_13803)
);

INVx1_ASAP7_75t_L g13804 ( 
.A(n_13572),
.Y(n_13804)
);

INVx1_ASAP7_75t_L g13805 ( 
.A(n_13427),
.Y(n_13805)
);

AND2x2_ASAP7_75t_L g13806 ( 
.A(n_13451),
.B(n_13383),
.Y(n_13806)
);

OAI211xp5_ASAP7_75t_L g13807 ( 
.A1(n_13471),
.A2(n_2314),
.B(n_2312),
.C(n_2313),
.Y(n_13807)
);

AND2x2_ASAP7_75t_L g13808 ( 
.A(n_13446),
.B(n_2313),
.Y(n_13808)
);

NAND2xp5_ASAP7_75t_L g13809 ( 
.A(n_13408),
.B(n_2314),
.Y(n_13809)
);

INVxp67_ASAP7_75t_L g13810 ( 
.A(n_13538),
.Y(n_13810)
);

INVx1_ASAP7_75t_L g13811 ( 
.A(n_13588),
.Y(n_13811)
);

AND2x2_ASAP7_75t_L g13812 ( 
.A(n_13579),
.B(n_2315),
.Y(n_13812)
);

INVx2_ASAP7_75t_L g13813 ( 
.A(n_13478),
.Y(n_13813)
);

INVx2_ASAP7_75t_L g13814 ( 
.A(n_13489),
.Y(n_13814)
);

INVx2_ASAP7_75t_SL g13815 ( 
.A(n_13551),
.Y(n_13815)
);

INVx1_ASAP7_75t_L g13816 ( 
.A(n_13595),
.Y(n_13816)
);

INVxp67_ASAP7_75t_L g13817 ( 
.A(n_13441),
.Y(n_13817)
);

INVx1_ASAP7_75t_L g13818 ( 
.A(n_13607),
.Y(n_13818)
);

INVx1_ASAP7_75t_L g13819 ( 
.A(n_13481),
.Y(n_13819)
);

AND2x2_ASAP7_75t_L g13820 ( 
.A(n_13402),
.B(n_2315),
.Y(n_13820)
);

INVx1_ASAP7_75t_L g13821 ( 
.A(n_13596),
.Y(n_13821)
);

INVx2_ASAP7_75t_L g13822 ( 
.A(n_13548),
.Y(n_13822)
);

INVx3_ASAP7_75t_L g13823 ( 
.A(n_13405),
.Y(n_13823)
);

INVx2_ASAP7_75t_L g13824 ( 
.A(n_13650),
.Y(n_13824)
);

NOR2xp33_ASAP7_75t_L g13825 ( 
.A(n_13643),
.B(n_13440),
.Y(n_13825)
);

INVxp67_ASAP7_75t_SL g13826 ( 
.A(n_13697),
.Y(n_13826)
);

INVx1_ASAP7_75t_L g13827 ( 
.A(n_13625),
.Y(n_13827)
);

BUFx12f_ASAP7_75t_L g13828 ( 
.A(n_13637),
.Y(n_13828)
);

INVx2_ASAP7_75t_L g13829 ( 
.A(n_13688),
.Y(n_13829)
);

NAND2xp5_ASAP7_75t_L g13830 ( 
.A(n_13787),
.B(n_13429),
.Y(n_13830)
);

AND2x2_ASAP7_75t_L g13831 ( 
.A(n_13630),
.B(n_13423),
.Y(n_13831)
);

OR2x2_ASAP7_75t_L g13832 ( 
.A(n_13624),
.B(n_13563),
.Y(n_13832)
);

INVx1_ASAP7_75t_L g13833 ( 
.A(n_13701),
.Y(n_13833)
);

NAND2xp5_ASAP7_75t_L g13834 ( 
.A(n_13669),
.B(n_13608),
.Y(n_13834)
);

AND2x2_ASAP7_75t_L g13835 ( 
.A(n_13627),
.B(n_13605),
.Y(n_13835)
);

NAND2xp5_ASAP7_75t_L g13836 ( 
.A(n_13722),
.B(n_13403),
.Y(n_13836)
);

AND2x4_ASAP7_75t_SL g13837 ( 
.A(n_13656),
.B(n_13447),
.Y(n_13837)
);

AND2x2_ASAP7_75t_L g13838 ( 
.A(n_13621),
.B(n_13606),
.Y(n_13838)
);

INVx1_ASAP7_75t_L g13839 ( 
.A(n_13721),
.Y(n_13839)
);

NAND2xp5_ASAP7_75t_L g13840 ( 
.A(n_13675),
.B(n_13806),
.Y(n_13840)
);

AND2x2_ASAP7_75t_L g13841 ( 
.A(n_13647),
.B(n_13543),
.Y(n_13841)
);

INVxp67_ASAP7_75t_SL g13842 ( 
.A(n_13656),
.Y(n_13842)
);

INVx3_ASAP7_75t_L g13843 ( 
.A(n_13626),
.Y(n_13843)
);

OR2x2_ASAP7_75t_L g13844 ( 
.A(n_13651),
.B(n_13659),
.Y(n_13844)
);

INVx1_ASAP7_75t_L g13845 ( 
.A(n_13666),
.Y(n_13845)
);

INVx2_ASAP7_75t_L g13846 ( 
.A(n_13678),
.Y(n_13846)
);

NAND2xp5_ASAP7_75t_L g13847 ( 
.A(n_13823),
.B(n_13614),
.Y(n_13847)
);

NOR2xp33_ASAP7_75t_L g13848 ( 
.A(n_13764),
.B(n_13363),
.Y(n_13848)
);

AND2x2_ASAP7_75t_L g13849 ( 
.A(n_13633),
.B(n_13493),
.Y(n_13849)
);

INVx2_ASAP7_75t_L g13850 ( 
.A(n_13631),
.Y(n_13850)
);

NAND2xp5_ASAP7_75t_SL g13851 ( 
.A(n_13623),
.B(n_13384),
.Y(n_13851)
);

INVxp67_ASAP7_75t_L g13852 ( 
.A(n_13762),
.Y(n_13852)
);

INVx2_ASAP7_75t_L g13853 ( 
.A(n_13686),
.Y(n_13853)
);

HB1xp67_ASAP7_75t_L g13854 ( 
.A(n_13711),
.Y(n_13854)
);

INVx1_ASAP7_75t_L g13855 ( 
.A(n_13677),
.Y(n_13855)
);

INVx1_ASAP7_75t_L g13856 ( 
.A(n_13690),
.Y(n_13856)
);

OR2x6_ASAP7_75t_SL g13857 ( 
.A(n_13720),
.B(n_13472),
.Y(n_13857)
);

INVx1_ASAP7_75t_SL g13858 ( 
.A(n_13762),
.Y(n_13858)
);

INVx2_ASAP7_75t_L g13859 ( 
.A(n_13718),
.Y(n_13859)
);

INVx1_ASAP7_75t_L g13860 ( 
.A(n_13695),
.Y(n_13860)
);

AND2x2_ASAP7_75t_L g13861 ( 
.A(n_13640),
.B(n_13413),
.Y(n_13861)
);

AND2x2_ASAP7_75t_L g13862 ( 
.A(n_13663),
.B(n_13490),
.Y(n_13862)
);

AND2x2_ASAP7_75t_L g13863 ( 
.A(n_13658),
.B(n_13385),
.Y(n_13863)
);

HB1xp67_ASAP7_75t_L g13864 ( 
.A(n_13679),
.Y(n_13864)
);

NOR2xp33_ASAP7_75t_L g13865 ( 
.A(n_13817),
.B(n_13425),
.Y(n_13865)
);

INVx1_ASAP7_75t_L g13866 ( 
.A(n_13628),
.Y(n_13866)
);

HB1xp67_ASAP7_75t_L g13867 ( 
.A(n_13689),
.Y(n_13867)
);

AND2x2_ASAP7_75t_L g13868 ( 
.A(n_13635),
.B(n_13497),
.Y(n_13868)
);

AOI22xp33_ASAP7_75t_L g13869 ( 
.A1(n_13798),
.A2(n_13539),
.B1(n_13486),
.B2(n_13479),
.Y(n_13869)
);

INVx1_ASAP7_75t_L g13870 ( 
.A(n_13694),
.Y(n_13870)
);

INVx1_ASAP7_75t_L g13871 ( 
.A(n_13755),
.Y(n_13871)
);

AOI22xp33_ASAP7_75t_L g13872 ( 
.A1(n_13794),
.A2(n_13433),
.B1(n_13470),
.B2(n_13465),
.Y(n_13872)
);

AND2x2_ASAP7_75t_L g13873 ( 
.A(n_13662),
.B(n_13482),
.Y(n_13873)
);

INVx1_ASAP7_75t_L g13874 ( 
.A(n_13692),
.Y(n_13874)
);

INVxp67_ASAP7_75t_L g13875 ( 
.A(n_13649),
.Y(n_13875)
);

NAND2xp5_ASAP7_75t_L g13876 ( 
.A(n_13810),
.B(n_13573),
.Y(n_13876)
);

INVx1_ASAP7_75t_L g13877 ( 
.A(n_13672),
.Y(n_13877)
);

INVx1_ASAP7_75t_L g13878 ( 
.A(n_13772),
.Y(n_13878)
);

NAND2xp5_ASAP7_75t_L g13879 ( 
.A(n_13788),
.B(n_13577),
.Y(n_13879)
);

AND2x2_ASAP7_75t_L g13880 ( 
.A(n_13642),
.B(n_13510),
.Y(n_13880)
);

AND2x2_ASAP7_75t_L g13881 ( 
.A(n_13654),
.B(n_13529),
.Y(n_13881)
);

NAND2xp5_ASAP7_75t_L g13882 ( 
.A(n_13749),
.B(n_13601),
.Y(n_13882)
);

INVxp67_ASAP7_75t_SL g13883 ( 
.A(n_13641),
.Y(n_13883)
);

AND2x2_ASAP7_75t_L g13884 ( 
.A(n_13639),
.B(n_13468),
.Y(n_13884)
);

AND2x2_ASAP7_75t_L g13885 ( 
.A(n_13655),
.B(n_13594),
.Y(n_13885)
);

INVxp67_ASAP7_75t_SL g13886 ( 
.A(n_13638),
.Y(n_13886)
);

AND2x2_ASAP7_75t_L g13887 ( 
.A(n_13629),
.B(n_13417),
.Y(n_13887)
);

AND2x2_ASAP7_75t_L g13888 ( 
.A(n_13634),
.B(n_13522),
.Y(n_13888)
);

AND2x2_ASAP7_75t_L g13889 ( 
.A(n_13682),
.B(n_13668),
.Y(n_13889)
);

AND2x2_ASAP7_75t_L g13890 ( 
.A(n_13644),
.B(n_13476),
.Y(n_13890)
);

AOI22xp33_ASAP7_75t_L g13891 ( 
.A1(n_13792),
.A2(n_13453),
.B1(n_13525),
.B2(n_13524),
.Y(n_13891)
);

BUFx6f_ASAP7_75t_L g13892 ( 
.A(n_13758),
.Y(n_13892)
);

INVx2_ASAP7_75t_L g13893 ( 
.A(n_13670),
.Y(n_13893)
);

NAND2xp5_ASAP7_75t_L g13894 ( 
.A(n_13745),
.B(n_13558),
.Y(n_13894)
);

INVx2_ASAP7_75t_L g13895 ( 
.A(n_13671),
.Y(n_13895)
);

INVx1_ASAP7_75t_L g13896 ( 
.A(n_13754),
.Y(n_13896)
);

BUFx2_ASAP7_75t_L g13897 ( 
.A(n_13742),
.Y(n_13897)
);

INVx1_ASAP7_75t_L g13898 ( 
.A(n_13705),
.Y(n_13898)
);

OR2x2_ASAP7_75t_L g13899 ( 
.A(n_13805),
.B(n_13532),
.Y(n_13899)
);

AOI22xp33_ASAP7_75t_L g13900 ( 
.A1(n_13791),
.A2(n_13400),
.B1(n_13375),
.B2(n_13371),
.Y(n_13900)
);

NOR2xp67_ASAP7_75t_L g13901 ( 
.A(n_13712),
.B(n_13714),
.Y(n_13901)
);

NAND2xp5_ASAP7_75t_L g13902 ( 
.A(n_13781),
.B(n_13556),
.Y(n_13902)
);

INVx2_ASAP7_75t_L g13903 ( 
.A(n_13622),
.Y(n_13903)
);

AND2x2_ASAP7_75t_L g13904 ( 
.A(n_13741),
.B(n_13561),
.Y(n_13904)
);

INVx1_ASAP7_75t_L g13905 ( 
.A(n_13636),
.Y(n_13905)
);

AND2x2_ASAP7_75t_L g13906 ( 
.A(n_13698),
.B(n_13567),
.Y(n_13906)
);

INVx2_ASAP7_75t_L g13907 ( 
.A(n_13680),
.Y(n_13907)
);

INVx2_ASAP7_75t_L g13908 ( 
.A(n_13702),
.Y(n_13908)
);

OAI22xp5_ASAP7_75t_L g13909 ( 
.A1(n_13660),
.A2(n_13507),
.B1(n_13509),
.B2(n_13583),
.Y(n_13909)
);

INVx1_ASAP7_75t_SL g13910 ( 
.A(n_13757),
.Y(n_13910)
);

AND2x2_ASAP7_75t_L g13911 ( 
.A(n_13743),
.B(n_13700),
.Y(n_13911)
);

INVxp67_ASAP7_75t_SL g13912 ( 
.A(n_13738),
.Y(n_13912)
);

INVxp67_ASAP7_75t_SL g13913 ( 
.A(n_13729),
.Y(n_13913)
);

INVx1_ASAP7_75t_L g13914 ( 
.A(n_13648),
.Y(n_13914)
);

AND2x2_ASAP7_75t_L g13915 ( 
.A(n_13716),
.B(n_13585),
.Y(n_13915)
);

AND2x2_ASAP7_75t_L g13916 ( 
.A(n_13696),
.B(n_13586),
.Y(n_13916)
);

INVx1_ASAP7_75t_L g13917 ( 
.A(n_13661),
.Y(n_13917)
);

HB1xp67_ASAP7_75t_L g13918 ( 
.A(n_13758),
.Y(n_13918)
);

INVx1_ASAP7_75t_L g13919 ( 
.A(n_13715),
.Y(n_13919)
);

AND2x2_ASAP7_75t_L g13920 ( 
.A(n_13646),
.B(n_13619),
.Y(n_13920)
);

OR2x2_ASAP7_75t_L g13921 ( 
.A(n_13632),
.B(n_13512),
.Y(n_13921)
);

AND2x2_ASAP7_75t_L g13922 ( 
.A(n_13687),
.B(n_13431),
.Y(n_13922)
);

NOR2xp33_ASAP7_75t_L g13923 ( 
.A(n_13693),
.B(n_13469),
.Y(n_13923)
);

AND2x2_ASAP7_75t_L g13924 ( 
.A(n_13709),
.B(n_2316),
.Y(n_13924)
);

INVx1_ASAP7_75t_L g13925 ( 
.A(n_13726),
.Y(n_13925)
);

AND2x2_ASAP7_75t_L g13926 ( 
.A(n_13731),
.B(n_13685),
.Y(n_13926)
);

HB1xp67_ASAP7_75t_L g13927 ( 
.A(n_13759),
.Y(n_13927)
);

AND2x2_ASAP7_75t_L g13928 ( 
.A(n_13768),
.B(n_2316),
.Y(n_13928)
);

NAND2xp5_ASAP7_75t_L g13929 ( 
.A(n_13778),
.B(n_13815),
.Y(n_13929)
);

INVx2_ASAP7_75t_L g13930 ( 
.A(n_13724),
.Y(n_13930)
);

NAND2xp5_ASAP7_75t_L g13931 ( 
.A(n_13765),
.B(n_13819),
.Y(n_13931)
);

INVx1_ASAP7_75t_L g13932 ( 
.A(n_13703),
.Y(n_13932)
);

INVx3_ASAP7_75t_L g13933 ( 
.A(n_13652),
.Y(n_13933)
);

INVx5_ASAP7_75t_L g13934 ( 
.A(n_13769),
.Y(n_13934)
);

AND2x2_ASAP7_75t_L g13935 ( 
.A(n_13752),
.B(n_2317),
.Y(n_13935)
);

NAND2xp5_ASAP7_75t_L g13936 ( 
.A(n_13821),
.B(n_13684),
.Y(n_13936)
);

INVx1_ASAP7_75t_L g13937 ( 
.A(n_13727),
.Y(n_13937)
);

INVx1_ASAP7_75t_L g13938 ( 
.A(n_13746),
.Y(n_13938)
);

HB1xp67_ASAP7_75t_L g13939 ( 
.A(n_13756),
.Y(n_13939)
);

INVx2_ASAP7_75t_L g13940 ( 
.A(n_13653),
.Y(n_13940)
);

AOI22xp33_ASAP7_75t_L g13941 ( 
.A1(n_13813),
.A2(n_2319),
.B1(n_2317),
.B2(n_2318),
.Y(n_13941)
);

AND2x2_ASAP7_75t_L g13942 ( 
.A(n_13822),
.B(n_2318),
.Y(n_13942)
);

AND2x2_ASAP7_75t_L g13943 ( 
.A(n_13691),
.B(n_2319),
.Y(n_13943)
);

INVx1_ASAP7_75t_L g13944 ( 
.A(n_13676),
.Y(n_13944)
);

OAI22xp5_ASAP7_75t_L g13945 ( 
.A1(n_13664),
.A2(n_2322),
.B1(n_2320),
.B2(n_2321),
.Y(n_13945)
);

AND2x2_ASAP7_75t_L g13946 ( 
.A(n_13761),
.B(n_2320),
.Y(n_13946)
);

NAND2xp5_ASAP7_75t_L g13947 ( 
.A(n_13785),
.B(n_2321),
.Y(n_13947)
);

INVx2_ASAP7_75t_L g13948 ( 
.A(n_13673),
.Y(n_13948)
);

INVx1_ASAP7_75t_L g13949 ( 
.A(n_13730),
.Y(n_13949)
);

OR2x2_ASAP7_75t_L g13950 ( 
.A(n_13667),
.B(n_13783),
.Y(n_13950)
);

INVx1_ASAP7_75t_L g13951 ( 
.A(n_13767),
.Y(n_13951)
);

INVx2_ASAP7_75t_L g13952 ( 
.A(n_13674),
.Y(n_13952)
);

OR2x2_ASAP7_75t_SL g13953 ( 
.A(n_13779),
.B(n_2322),
.Y(n_13953)
);

INVx3_ASAP7_75t_L g13954 ( 
.A(n_13704),
.Y(n_13954)
);

AND2x4_ASAP7_75t_L g13955 ( 
.A(n_13732),
.B(n_2323),
.Y(n_13955)
);

INVxp67_ASAP7_75t_L g13956 ( 
.A(n_13747),
.Y(n_13956)
);

INVxp67_ASAP7_75t_L g13957 ( 
.A(n_13777),
.Y(n_13957)
);

INVx1_ASAP7_75t_L g13958 ( 
.A(n_13699),
.Y(n_13958)
);

AND2x4_ASAP7_75t_L g13959 ( 
.A(n_13739),
.B(n_2323),
.Y(n_13959)
);

INVx3_ASAP7_75t_L g13960 ( 
.A(n_13766),
.Y(n_13960)
);

AND2x2_ASAP7_75t_L g13961 ( 
.A(n_13770),
.B(n_2324),
.Y(n_13961)
);

OR2x2_ASAP7_75t_L g13962 ( 
.A(n_13811),
.B(n_2324),
.Y(n_13962)
);

AND2x2_ASAP7_75t_L g13963 ( 
.A(n_13665),
.B(n_2325),
.Y(n_13963)
);

AND2x2_ASAP7_75t_L g13964 ( 
.A(n_13804),
.B(n_2326),
.Y(n_13964)
);

AND2x2_ASAP7_75t_L g13965 ( 
.A(n_13780),
.B(n_2326),
.Y(n_13965)
);

INVx2_ASAP7_75t_L g13966 ( 
.A(n_13763),
.Y(n_13966)
);

INVx2_ASAP7_75t_L g13967 ( 
.A(n_13706),
.Y(n_13967)
);

INVx2_ASAP7_75t_L g13968 ( 
.A(n_13707),
.Y(n_13968)
);

OAI222xp33_ASAP7_75t_L g13969 ( 
.A1(n_13760),
.A2(n_2329),
.B1(n_2331),
.B2(n_2327),
.C1(n_2328),
.C2(n_2330),
.Y(n_13969)
);

AOI22xp33_ASAP7_75t_L g13970 ( 
.A1(n_13814),
.A2(n_2330),
.B1(n_2328),
.B2(n_2329),
.Y(n_13970)
);

INVx2_ASAP7_75t_R g13971 ( 
.A(n_13710),
.Y(n_13971)
);

AOI22xp33_ASAP7_75t_L g13972 ( 
.A1(n_13796),
.A2(n_2333),
.B1(n_2331),
.B2(n_2332),
.Y(n_13972)
);

OR2x2_ASAP7_75t_L g13973 ( 
.A(n_13816),
.B(n_2332),
.Y(n_13973)
);

INVx1_ASAP7_75t_L g13974 ( 
.A(n_13713),
.Y(n_13974)
);

NOR2xp33_ASAP7_75t_L g13975 ( 
.A(n_13795),
.B(n_2333),
.Y(n_13975)
);

INVx1_ASAP7_75t_L g13976 ( 
.A(n_13717),
.Y(n_13976)
);

INVx1_ASAP7_75t_L g13977 ( 
.A(n_13719),
.Y(n_13977)
);

OR2x2_ASAP7_75t_L g13978 ( 
.A(n_13818),
.B(n_2334),
.Y(n_13978)
);

AND2x2_ASAP7_75t_L g13979 ( 
.A(n_13799),
.B(n_2335),
.Y(n_13979)
);

INVx2_ASAP7_75t_L g13980 ( 
.A(n_13824),
.Y(n_13980)
);

INVx2_ASAP7_75t_L g13981 ( 
.A(n_13828),
.Y(n_13981)
);

HB1xp67_ASAP7_75t_L g13982 ( 
.A(n_13854),
.Y(n_13982)
);

AND2x2_ASAP7_75t_L g13983 ( 
.A(n_13826),
.B(n_13858),
.Y(n_13983)
);

HB1xp67_ASAP7_75t_L g13984 ( 
.A(n_13901),
.Y(n_13984)
);

INVx3_ASAP7_75t_L g13985 ( 
.A(n_13892),
.Y(n_13985)
);

INVx1_ASAP7_75t_L g13986 ( 
.A(n_13867),
.Y(n_13986)
);

NAND2xp5_ASAP7_75t_L g13987 ( 
.A(n_13842),
.B(n_13751),
.Y(n_13987)
);

INVx1_ASAP7_75t_L g13988 ( 
.A(n_13864),
.Y(n_13988)
);

INVx2_ASAP7_75t_L g13989 ( 
.A(n_13843),
.Y(n_13989)
);

NAND2xp5_ASAP7_75t_L g13990 ( 
.A(n_13852),
.B(n_13681),
.Y(n_13990)
);

NAND2xp5_ASAP7_75t_L g13991 ( 
.A(n_13846),
.B(n_13708),
.Y(n_13991)
);

INVx1_ASAP7_75t_L g13992 ( 
.A(n_13951),
.Y(n_13992)
);

AND2x4_ASAP7_75t_SL g13993 ( 
.A(n_13892),
.B(n_13774),
.Y(n_13993)
);

INVxp67_ASAP7_75t_L g13994 ( 
.A(n_13857),
.Y(n_13994)
);

INVx1_ASAP7_75t_L g13995 ( 
.A(n_13845),
.Y(n_13995)
);

AND2x2_ASAP7_75t_L g13996 ( 
.A(n_13838),
.B(n_13683),
.Y(n_13996)
);

HB1xp67_ASAP7_75t_L g13997 ( 
.A(n_13971),
.Y(n_13997)
);

AND2x2_ASAP7_75t_L g13998 ( 
.A(n_13829),
.B(n_13645),
.Y(n_13998)
);

BUFx2_ASAP7_75t_L g13999 ( 
.A(n_13897),
.Y(n_13999)
);

NAND2xp5_ASAP7_75t_L g14000 ( 
.A(n_13934),
.B(n_13820),
.Y(n_14000)
);

AND2x2_ASAP7_75t_L g14001 ( 
.A(n_13889),
.B(n_13850),
.Y(n_14001)
);

NAND2xp5_ASAP7_75t_L g14002 ( 
.A(n_13934),
.B(n_13812),
.Y(n_14002)
);

INVx1_ASAP7_75t_L g14003 ( 
.A(n_13855),
.Y(n_14003)
);

AND2x2_ASAP7_75t_L g14004 ( 
.A(n_13831),
.B(n_13911),
.Y(n_14004)
);

AND2x2_ASAP7_75t_L g14005 ( 
.A(n_13853),
.B(n_13657),
.Y(n_14005)
);

AND2x2_ASAP7_75t_L g14006 ( 
.A(n_13841),
.B(n_13725),
.Y(n_14006)
);

NAND2xp5_ASAP7_75t_L g14007 ( 
.A(n_13934),
.B(n_13786),
.Y(n_14007)
);

INVx3_ASAP7_75t_L g14008 ( 
.A(n_13954),
.Y(n_14008)
);

NAND2xp5_ASAP7_75t_L g14009 ( 
.A(n_13849),
.B(n_13943),
.Y(n_14009)
);

NAND2xp5_ASAP7_75t_L g14010 ( 
.A(n_13926),
.B(n_13771),
.Y(n_14010)
);

INVx2_ASAP7_75t_L g14011 ( 
.A(n_13859),
.Y(n_14011)
);

INVx4_ASAP7_75t_L g14012 ( 
.A(n_13918),
.Y(n_14012)
);

INVx1_ASAP7_75t_L g14013 ( 
.A(n_13939),
.Y(n_14013)
);

AND2x4_ASAP7_75t_L g14014 ( 
.A(n_13903),
.B(n_13723),
.Y(n_14014)
);

AND2x2_ASAP7_75t_L g14015 ( 
.A(n_13835),
.B(n_13880),
.Y(n_14015)
);

INVx1_ASAP7_75t_L g14016 ( 
.A(n_13927),
.Y(n_14016)
);

INVx2_ASAP7_75t_L g14017 ( 
.A(n_13933),
.Y(n_14017)
);

INVx1_ASAP7_75t_L g14018 ( 
.A(n_13833),
.Y(n_14018)
);

AND2x2_ASAP7_75t_L g14019 ( 
.A(n_13873),
.B(n_13784),
.Y(n_14019)
);

INVx2_ASAP7_75t_L g14020 ( 
.A(n_13960),
.Y(n_14020)
);

NAND2xp5_ASAP7_75t_L g14021 ( 
.A(n_13910),
.B(n_13773),
.Y(n_14021)
);

HB1xp67_ASAP7_75t_L g14022 ( 
.A(n_13856),
.Y(n_14022)
);

OR2x2_ASAP7_75t_L g14023 ( 
.A(n_13953),
.B(n_13776),
.Y(n_14023)
);

NAND2xp5_ASAP7_75t_L g14024 ( 
.A(n_13922),
.B(n_13790),
.Y(n_14024)
);

INVx2_ASAP7_75t_L g14025 ( 
.A(n_13959),
.Y(n_14025)
);

OR2x2_ASAP7_75t_L g14026 ( 
.A(n_13840),
.B(n_13800),
.Y(n_14026)
);

INVx2_ASAP7_75t_L g14027 ( 
.A(n_13930),
.Y(n_14027)
);

AOI22xp33_ASAP7_75t_L g14028 ( 
.A1(n_13836),
.A2(n_13753),
.B1(n_13797),
.B2(n_13801),
.Y(n_14028)
);

INVx2_ASAP7_75t_L g14029 ( 
.A(n_13955),
.Y(n_14029)
);

OR2x2_ASAP7_75t_L g14030 ( 
.A(n_13832),
.B(n_13782),
.Y(n_14030)
);

INVx2_ASAP7_75t_L g14031 ( 
.A(n_13935),
.Y(n_14031)
);

AND2x2_ASAP7_75t_L g14032 ( 
.A(n_13979),
.B(n_13728),
.Y(n_14032)
);

AND2x2_ASAP7_75t_L g14033 ( 
.A(n_13881),
.B(n_13733),
.Y(n_14033)
);

NAND2xp5_ASAP7_75t_L g14034 ( 
.A(n_13956),
.B(n_13802),
.Y(n_14034)
);

INVx1_ASAP7_75t_L g14035 ( 
.A(n_13839),
.Y(n_14035)
);

AND2x4_ASAP7_75t_L g14036 ( 
.A(n_13875),
.B(n_13734),
.Y(n_14036)
);

INVx1_ASAP7_75t_L g14037 ( 
.A(n_13860),
.Y(n_14037)
);

INVx1_ASAP7_75t_L g14038 ( 
.A(n_13878),
.Y(n_14038)
);

AND2x2_ASAP7_75t_L g14039 ( 
.A(n_13884),
.B(n_13735),
.Y(n_14039)
);

AND2x4_ASAP7_75t_L g14040 ( 
.A(n_13898),
.B(n_13736),
.Y(n_14040)
);

HB1xp67_ASAP7_75t_L g14041 ( 
.A(n_13938),
.Y(n_14041)
);

OR2x2_ASAP7_75t_L g14042 ( 
.A(n_13844),
.B(n_13793),
.Y(n_14042)
);

CKINVDCx20_ASAP7_75t_R g14043 ( 
.A(n_13882),
.Y(n_14043)
);

INVx1_ASAP7_75t_L g14044 ( 
.A(n_13924),
.Y(n_14044)
);

AND2x2_ASAP7_75t_L g14045 ( 
.A(n_13964),
.B(n_13737),
.Y(n_14045)
);

INVx1_ASAP7_75t_L g14046 ( 
.A(n_13928),
.Y(n_14046)
);

NAND2xp5_ASAP7_75t_L g14047 ( 
.A(n_13868),
.B(n_13809),
.Y(n_14047)
);

INVx4_ASAP7_75t_L g14048 ( 
.A(n_13961),
.Y(n_14048)
);

NAND2xp5_ASAP7_75t_SL g14049 ( 
.A(n_13830),
.B(n_13807),
.Y(n_14049)
);

OR2x2_ASAP7_75t_L g14050 ( 
.A(n_13929),
.B(n_13740),
.Y(n_14050)
);

INVx2_ASAP7_75t_L g14051 ( 
.A(n_13966),
.Y(n_14051)
);

INVx2_ASAP7_75t_L g14052 ( 
.A(n_13919),
.Y(n_14052)
);

NOR2xp67_ASAP7_75t_L g14053 ( 
.A(n_13940),
.B(n_13744),
.Y(n_14053)
);

NAND2xp5_ASAP7_75t_L g14054 ( 
.A(n_13862),
.B(n_13748),
.Y(n_14054)
);

NAND2xp5_ASAP7_75t_L g14055 ( 
.A(n_13865),
.B(n_13750),
.Y(n_14055)
);

AND2x2_ASAP7_75t_L g14056 ( 
.A(n_13887),
.B(n_13803),
.Y(n_14056)
);

INVx1_ASAP7_75t_L g14057 ( 
.A(n_13925),
.Y(n_14057)
);

HB1xp67_ASAP7_75t_L g14058 ( 
.A(n_13946),
.Y(n_14058)
);

INVxp67_ASAP7_75t_L g14059 ( 
.A(n_13923),
.Y(n_14059)
);

INVxp67_ASAP7_75t_L g14060 ( 
.A(n_13913),
.Y(n_14060)
);

NAND2xp5_ASAP7_75t_L g14061 ( 
.A(n_13885),
.B(n_13808),
.Y(n_14061)
);

BUFx6f_ASAP7_75t_L g14062 ( 
.A(n_13963),
.Y(n_14062)
);

INVx1_ASAP7_75t_L g14063 ( 
.A(n_13870),
.Y(n_14063)
);

AND2x2_ASAP7_75t_L g14064 ( 
.A(n_13888),
.B(n_13789),
.Y(n_14064)
);

NAND2xp5_ASAP7_75t_L g14065 ( 
.A(n_13837),
.B(n_13775),
.Y(n_14065)
);

AND2x2_ASAP7_75t_L g14066 ( 
.A(n_13942),
.B(n_2335),
.Y(n_14066)
);

AND2x2_ASAP7_75t_L g14067 ( 
.A(n_13861),
.B(n_2336),
.Y(n_14067)
);

INVx2_ASAP7_75t_L g14068 ( 
.A(n_13893),
.Y(n_14068)
);

BUFx3_ASAP7_75t_L g14069 ( 
.A(n_13932),
.Y(n_14069)
);

AND2x4_ASAP7_75t_L g14070 ( 
.A(n_13895),
.B(n_2336),
.Y(n_14070)
);

BUFx3_ASAP7_75t_L g14071 ( 
.A(n_13937),
.Y(n_14071)
);

HB1xp67_ASAP7_75t_L g14072 ( 
.A(n_13912),
.Y(n_14072)
);

AND2x2_ASAP7_75t_L g14073 ( 
.A(n_13920),
.B(n_2337),
.Y(n_14073)
);

INVx1_ASAP7_75t_L g14074 ( 
.A(n_13886),
.Y(n_14074)
);

AND2x4_ASAP7_75t_SL g14075 ( 
.A(n_13907),
.B(n_2337),
.Y(n_14075)
);

INVx1_ASAP7_75t_SL g14076 ( 
.A(n_13962),
.Y(n_14076)
);

AND2x4_ASAP7_75t_L g14077 ( 
.A(n_13908),
.B(n_2338),
.Y(n_14077)
);

INVx1_ASAP7_75t_L g14078 ( 
.A(n_13883),
.Y(n_14078)
);

INVx1_ASAP7_75t_L g14079 ( 
.A(n_13871),
.Y(n_14079)
);

AND2x2_ASAP7_75t_L g14080 ( 
.A(n_13890),
.B(n_2339),
.Y(n_14080)
);

NAND2xp5_ASAP7_75t_L g14081 ( 
.A(n_13906),
.B(n_2340),
.Y(n_14081)
);

AND2x4_ASAP7_75t_L g14082 ( 
.A(n_13874),
.B(n_2341),
.Y(n_14082)
);

INVxp67_ASAP7_75t_L g14083 ( 
.A(n_13825),
.Y(n_14083)
);

AND2x2_ASAP7_75t_L g14084 ( 
.A(n_13863),
.B(n_2341),
.Y(n_14084)
);

INVx1_ASAP7_75t_L g14085 ( 
.A(n_13965),
.Y(n_14085)
);

INVx1_ASAP7_75t_L g14086 ( 
.A(n_13827),
.Y(n_14086)
);

OR2x2_ASAP7_75t_L g14087 ( 
.A(n_13931),
.B(n_2342),
.Y(n_14087)
);

INVx2_ASAP7_75t_L g14088 ( 
.A(n_13948),
.Y(n_14088)
);

AND2x4_ASAP7_75t_L g14089 ( 
.A(n_13877),
.B(n_2343),
.Y(n_14089)
);

NAND2xp5_ASAP7_75t_L g14090 ( 
.A(n_13848),
.B(n_2343),
.Y(n_14090)
);

AND2x2_ASAP7_75t_L g14091 ( 
.A(n_13915),
.B(n_2344),
.Y(n_14091)
);

INVx1_ASAP7_75t_L g14092 ( 
.A(n_13896),
.Y(n_14092)
);

INVx1_ASAP7_75t_L g14093 ( 
.A(n_13973),
.Y(n_14093)
);

AND2x2_ASAP7_75t_L g14094 ( 
.A(n_13916),
.B(n_2344),
.Y(n_14094)
);

INVx1_ASAP7_75t_L g14095 ( 
.A(n_13978),
.Y(n_14095)
);

INVx2_ASAP7_75t_L g14096 ( 
.A(n_13952),
.Y(n_14096)
);

INVx2_ASAP7_75t_L g14097 ( 
.A(n_13866),
.Y(n_14097)
);

NAND2xp5_ASAP7_75t_L g14098 ( 
.A(n_13975),
.B(n_2345),
.Y(n_14098)
);

HB1xp67_ASAP7_75t_L g14099 ( 
.A(n_13944),
.Y(n_14099)
);

INVx1_ASAP7_75t_L g14100 ( 
.A(n_13949),
.Y(n_14100)
);

OR2x2_ASAP7_75t_L g14101 ( 
.A(n_13936),
.B(n_2346),
.Y(n_14101)
);

INVx1_ASAP7_75t_SL g14102 ( 
.A(n_13950),
.Y(n_14102)
);

OR2x2_ASAP7_75t_L g14103 ( 
.A(n_13899),
.B(n_2346),
.Y(n_14103)
);

INVx1_ASAP7_75t_L g14104 ( 
.A(n_13947),
.Y(n_14104)
);

AND2x4_ASAP7_75t_L g14105 ( 
.A(n_13905),
.B(n_13914),
.Y(n_14105)
);

OR2x2_ASAP7_75t_L g14106 ( 
.A(n_13879),
.B(n_2347),
.Y(n_14106)
);

INVx1_ASAP7_75t_L g14107 ( 
.A(n_13917),
.Y(n_14107)
);

OR2x2_ASAP7_75t_L g14108 ( 
.A(n_13847),
.B(n_2347),
.Y(n_14108)
);

AND2x2_ASAP7_75t_L g14109 ( 
.A(n_13904),
.B(n_2348),
.Y(n_14109)
);

AND2x4_ASAP7_75t_L g14110 ( 
.A(n_13967),
.B(n_2348),
.Y(n_14110)
);

INVx1_ASAP7_75t_L g14111 ( 
.A(n_13968),
.Y(n_14111)
);

AND2x4_ASAP7_75t_L g14112 ( 
.A(n_13977),
.B(n_2349),
.Y(n_14112)
);

OAI22xp33_ASAP7_75t_L g14113 ( 
.A1(n_13994),
.A2(n_13876),
.B1(n_13894),
.B2(n_13834),
.Y(n_14113)
);

NAND2xp5_ASAP7_75t_L g14114 ( 
.A(n_13983),
.B(n_13891),
.Y(n_14114)
);

INVx1_ASAP7_75t_L g14115 ( 
.A(n_13997),
.Y(n_14115)
);

AND2x2_ASAP7_75t_L g14116 ( 
.A(n_14004),
.B(n_13981),
.Y(n_14116)
);

NAND2xp5_ASAP7_75t_L g14117 ( 
.A(n_14015),
.B(n_13984),
.Y(n_14117)
);

AND2x2_ASAP7_75t_L g14118 ( 
.A(n_14001),
.B(n_13957),
.Y(n_14118)
);

INVx1_ASAP7_75t_L g14119 ( 
.A(n_14072),
.Y(n_14119)
);

AOI22xp33_ASAP7_75t_L g14120 ( 
.A1(n_14049),
.A2(n_13851),
.B1(n_13902),
.B2(n_13869),
.Y(n_14120)
);

AND2x2_ASAP7_75t_L g14121 ( 
.A(n_13993),
.B(n_13900),
.Y(n_14121)
);

BUFx3_ASAP7_75t_L g14122 ( 
.A(n_14062),
.Y(n_14122)
);

INVx3_ASAP7_75t_L g14123 ( 
.A(n_14012),
.Y(n_14123)
);

AND2x2_ASAP7_75t_L g14124 ( 
.A(n_14033),
.B(n_13872),
.Y(n_14124)
);

AND2x2_ASAP7_75t_L g14125 ( 
.A(n_14056),
.B(n_13921),
.Y(n_14125)
);

AOI21xp5_ASAP7_75t_L g14126 ( 
.A1(n_13982),
.A2(n_13909),
.B(n_13945),
.Y(n_14126)
);

OR2x2_ASAP7_75t_L g14127 ( 
.A(n_13987),
.B(n_13958),
.Y(n_14127)
);

INVx1_ASAP7_75t_L g14128 ( 
.A(n_14022),
.Y(n_14128)
);

AOI221xp5_ASAP7_75t_L g14129 ( 
.A1(n_14028),
.A2(n_13969),
.B1(n_13976),
.B2(n_13974),
.C(n_13970),
.Y(n_14129)
);

AND2x2_ASAP7_75t_L g14130 ( 
.A(n_13989),
.B(n_13972),
.Y(n_14130)
);

AND2x2_ASAP7_75t_L g14131 ( 
.A(n_14084),
.B(n_13941),
.Y(n_14131)
);

OAI321xp33_ASAP7_75t_L g14132 ( 
.A1(n_14000),
.A2(n_2351),
.A3(n_2353),
.B1(n_2349),
.B2(n_2350),
.C(n_2352),
.Y(n_14132)
);

AND2x2_ASAP7_75t_L g14133 ( 
.A(n_14064),
.B(n_2350),
.Y(n_14133)
);

NAND2x1p5_ASAP7_75t_SL g14134 ( 
.A(n_13998),
.B(n_14006),
.Y(n_14134)
);

INVx1_ASAP7_75t_L g14135 ( 
.A(n_14058),
.Y(n_14135)
);

AND2x2_ASAP7_75t_SL g14136 ( 
.A(n_14019),
.B(n_2352),
.Y(n_14136)
);

BUFx2_ASAP7_75t_L g14137 ( 
.A(n_14041),
.Y(n_14137)
);

AND2x2_ASAP7_75t_L g14138 ( 
.A(n_14109),
.B(n_2353),
.Y(n_14138)
);

BUFx2_ASAP7_75t_L g14139 ( 
.A(n_14062),
.Y(n_14139)
);

AND2x2_ASAP7_75t_L g14140 ( 
.A(n_14067),
.B(n_13980),
.Y(n_14140)
);

AOI211xp5_ASAP7_75t_SL g14141 ( 
.A1(n_14060),
.A2(n_2356),
.B(n_2354),
.C(n_2355),
.Y(n_14141)
);

OR2x2_ASAP7_75t_L g14142 ( 
.A(n_14023),
.B(n_2354),
.Y(n_14142)
);

INVx2_ASAP7_75t_L g14143 ( 
.A(n_14008),
.Y(n_14143)
);

INVx1_ASAP7_75t_L g14144 ( 
.A(n_13986),
.Y(n_14144)
);

BUFx2_ASAP7_75t_L g14145 ( 
.A(n_14048),
.Y(n_14145)
);

AND2x2_ASAP7_75t_L g14146 ( 
.A(n_14005),
.B(n_2355),
.Y(n_14146)
);

AND2x2_ASAP7_75t_L g14147 ( 
.A(n_14025),
.B(n_2356),
.Y(n_14147)
);

OAI22xp5_ASAP7_75t_L g14148 ( 
.A1(n_14043),
.A2(n_2359),
.B1(n_2357),
.B2(n_2358),
.Y(n_14148)
);

NOR2xp33_ASAP7_75t_L g14149 ( 
.A(n_14007),
.B(n_2358),
.Y(n_14149)
);

HB1xp67_ASAP7_75t_L g14150 ( 
.A(n_14053),
.Y(n_14150)
);

NAND2xp5_ASAP7_75t_L g14151 ( 
.A(n_13996),
.B(n_2360),
.Y(n_14151)
);

INVx1_ASAP7_75t_L g14152 ( 
.A(n_14099),
.Y(n_14152)
);

INVx4_ASAP7_75t_L g14153 ( 
.A(n_13985),
.Y(n_14153)
);

INVx2_ASAP7_75t_L g14154 ( 
.A(n_14075),
.Y(n_14154)
);

INVx2_ASAP7_75t_L g14155 ( 
.A(n_14069),
.Y(n_14155)
);

HB1xp67_ASAP7_75t_L g14156 ( 
.A(n_13988),
.Y(n_14156)
);

INVx1_ASAP7_75t_L g14157 ( 
.A(n_14066),
.Y(n_14157)
);

OAI22xp33_ASAP7_75t_L g14158 ( 
.A1(n_13999),
.A2(n_2363),
.B1(n_2361),
.B2(n_2362),
.Y(n_14158)
);

INVx2_ASAP7_75t_L g14159 ( 
.A(n_14071),
.Y(n_14159)
);

INVx1_ASAP7_75t_L g14160 ( 
.A(n_14017),
.Y(n_14160)
);

OR2x2_ASAP7_75t_L g14161 ( 
.A(n_14010),
.B(n_2361),
.Y(n_14161)
);

AND2x2_ASAP7_75t_L g14162 ( 
.A(n_14080),
.B(n_2362),
.Y(n_14162)
);

INVx2_ASAP7_75t_L g14163 ( 
.A(n_14029),
.Y(n_14163)
);

OR2x2_ASAP7_75t_L g14164 ( 
.A(n_14002),
.B(n_2363),
.Y(n_14164)
);

AOI33xp33_ASAP7_75t_L g14165 ( 
.A1(n_14102),
.A2(n_2366),
.A3(n_2368),
.B1(n_2364),
.B2(n_2365),
.B3(n_2367),
.Y(n_14165)
);

INVx1_ASAP7_75t_L g14166 ( 
.A(n_14046),
.Y(n_14166)
);

NAND2xp5_ASAP7_75t_L g14167 ( 
.A(n_14091),
.B(n_2365),
.Y(n_14167)
);

INVxp67_ASAP7_75t_L g14168 ( 
.A(n_14009),
.Y(n_14168)
);

INVx1_ASAP7_75t_L g14169 ( 
.A(n_14039),
.Y(n_14169)
);

AND2x2_ASAP7_75t_L g14170 ( 
.A(n_14094),
.B(n_14073),
.Y(n_14170)
);

INVx1_ASAP7_75t_L g14171 ( 
.A(n_14032),
.Y(n_14171)
);

INVx2_ASAP7_75t_SL g14172 ( 
.A(n_14082),
.Y(n_14172)
);

NAND3xp33_ASAP7_75t_L g14173 ( 
.A(n_14013),
.B(n_2366),
.C(n_2367),
.Y(n_14173)
);

INVxp67_ASAP7_75t_L g14174 ( 
.A(n_13991),
.Y(n_14174)
);

OAI21xp5_ASAP7_75t_L g14175 ( 
.A1(n_14059),
.A2(n_14024),
.B(n_14090),
.Y(n_14175)
);

AND2x2_ASAP7_75t_L g14176 ( 
.A(n_14031),
.B(n_2369),
.Y(n_14176)
);

BUFx2_ASAP7_75t_L g14177 ( 
.A(n_14016),
.Y(n_14177)
);

INVx2_ASAP7_75t_L g14178 ( 
.A(n_14020),
.Y(n_14178)
);

OR2x2_ASAP7_75t_L g14179 ( 
.A(n_14026),
.B(n_2369),
.Y(n_14179)
);

OR2x2_ASAP7_75t_L g14180 ( 
.A(n_14042),
.B(n_2370),
.Y(n_14180)
);

AND2x2_ASAP7_75t_L g14181 ( 
.A(n_14044),
.B(n_2370),
.Y(n_14181)
);

OA21x2_ASAP7_75t_L g14182 ( 
.A1(n_14061),
.A2(n_2371),
.B(n_2372),
.Y(n_14182)
);

BUFx3_ASAP7_75t_L g14183 ( 
.A(n_14036),
.Y(n_14183)
);

AND2x2_ASAP7_75t_L g14184 ( 
.A(n_14011),
.B(n_2371),
.Y(n_14184)
);

BUFx2_ASAP7_75t_L g14185 ( 
.A(n_14014),
.Y(n_14185)
);

INVx1_ASAP7_75t_L g14186 ( 
.A(n_14045),
.Y(n_14186)
);

INVx1_ASAP7_75t_L g14187 ( 
.A(n_13995),
.Y(n_14187)
);

OR2x2_ASAP7_75t_L g14188 ( 
.A(n_14103),
.B(n_2372),
.Y(n_14188)
);

INVx2_ASAP7_75t_L g14189 ( 
.A(n_14070),
.Y(n_14189)
);

OR2x2_ASAP7_75t_L g14190 ( 
.A(n_14030),
.B(n_13990),
.Y(n_14190)
);

INVx2_ASAP7_75t_L g14191 ( 
.A(n_14077),
.Y(n_14191)
);

INVx1_ASAP7_75t_L g14192 ( 
.A(n_14003),
.Y(n_14192)
);

OAI211xp5_ASAP7_75t_L g14193 ( 
.A1(n_14055),
.A2(n_2376),
.B(n_2373),
.C(n_2375),
.Y(n_14193)
);

AOI31xp33_ASAP7_75t_L g14194 ( 
.A1(n_14076),
.A2(n_2377),
.A3(n_2375),
.B(n_2376),
.Y(n_14194)
);

NAND2xp5_ASAP7_75t_L g14195 ( 
.A(n_14085),
.B(n_2378),
.Y(n_14195)
);

AND2x2_ASAP7_75t_L g14196 ( 
.A(n_14051),
.B(n_2379),
.Y(n_14196)
);

AND2x2_ASAP7_75t_L g14197 ( 
.A(n_14027),
.B(n_2379),
.Y(n_14197)
);

INVx2_ASAP7_75t_L g14198 ( 
.A(n_14110),
.Y(n_14198)
);

INVx1_ASAP7_75t_L g14199 ( 
.A(n_14074),
.Y(n_14199)
);

NAND2xp5_ASAP7_75t_L g14200 ( 
.A(n_14078),
.B(n_2380),
.Y(n_14200)
);

AND2x2_ASAP7_75t_L g14201 ( 
.A(n_14093),
.B(n_2380),
.Y(n_14201)
);

HB1xp67_ASAP7_75t_L g14202 ( 
.A(n_14037),
.Y(n_14202)
);

HB1xp67_ASAP7_75t_L g14203 ( 
.A(n_14095),
.Y(n_14203)
);

AOI221xp5_ASAP7_75t_L g14204 ( 
.A1(n_14083),
.A2(n_2383),
.B1(n_2381),
.B2(n_2382),
.C(n_2384),
.Y(n_14204)
);

HB1xp67_ASAP7_75t_L g14205 ( 
.A(n_14040),
.Y(n_14205)
);

AO21x2_ASAP7_75t_L g14206 ( 
.A1(n_14081),
.A2(n_2381),
.B(n_2385),
.Y(n_14206)
);

INVxp67_ASAP7_75t_L g14207 ( 
.A(n_14065),
.Y(n_14207)
);

INVx2_ASAP7_75t_L g14208 ( 
.A(n_14089),
.Y(n_14208)
);

INVx1_ASAP7_75t_L g14209 ( 
.A(n_14050),
.Y(n_14209)
);

AND2x4_ASAP7_75t_L g14210 ( 
.A(n_14052),
.B(n_2385),
.Y(n_14210)
);

AND2x4_ASAP7_75t_L g14211 ( 
.A(n_14068),
.B(n_2386),
.Y(n_14211)
);

INVx2_ASAP7_75t_L g14212 ( 
.A(n_14112),
.Y(n_14212)
);

AND2x4_ASAP7_75t_L g14213 ( 
.A(n_14063),
.B(n_2386),
.Y(n_14213)
);

INVx5_ASAP7_75t_L g14214 ( 
.A(n_14105),
.Y(n_14214)
);

INVx1_ASAP7_75t_L g14215 ( 
.A(n_14018),
.Y(n_14215)
);

AND2x2_ASAP7_75t_L g14216 ( 
.A(n_14100),
.B(n_2387),
.Y(n_14216)
);

INVxp67_ASAP7_75t_SL g14217 ( 
.A(n_14021),
.Y(n_14217)
);

BUFx3_ASAP7_75t_L g14218 ( 
.A(n_14057),
.Y(n_14218)
);

INVx1_ASAP7_75t_L g14219 ( 
.A(n_14035),
.Y(n_14219)
);

AND2x2_ASAP7_75t_L g14220 ( 
.A(n_14104),
.B(n_2387),
.Y(n_14220)
);

AND2x2_ASAP7_75t_L g14221 ( 
.A(n_14108),
.B(n_2388),
.Y(n_14221)
);

OR2x2_ASAP7_75t_L g14222 ( 
.A(n_14047),
.B(n_2389),
.Y(n_14222)
);

INVx2_ASAP7_75t_SL g14223 ( 
.A(n_14097),
.Y(n_14223)
);

INVx1_ASAP7_75t_L g14224 ( 
.A(n_14038),
.Y(n_14224)
);

AO21x2_ASAP7_75t_L g14225 ( 
.A1(n_14098),
.A2(n_2390),
.B(n_2391),
.Y(n_14225)
);

AND2x2_ASAP7_75t_L g14226 ( 
.A(n_14054),
.B(n_2390),
.Y(n_14226)
);

OR2x2_ASAP7_75t_L g14227 ( 
.A(n_14034),
.B(n_2391),
.Y(n_14227)
);

AND2x2_ASAP7_75t_L g14228 ( 
.A(n_14116),
.B(n_14088),
.Y(n_14228)
);

AND2x2_ASAP7_75t_L g14229 ( 
.A(n_14125),
.B(n_14096),
.Y(n_14229)
);

INVx2_ASAP7_75t_L g14230 ( 
.A(n_14214),
.Y(n_14230)
);

INVx1_ASAP7_75t_L g14231 ( 
.A(n_14205),
.Y(n_14231)
);

OR2x2_ASAP7_75t_L g14232 ( 
.A(n_14185),
.B(n_14101),
.Y(n_14232)
);

AND2x2_ASAP7_75t_L g14233 ( 
.A(n_14123),
.B(n_14106),
.Y(n_14233)
);

INVx1_ASAP7_75t_L g14234 ( 
.A(n_14150),
.Y(n_14234)
);

AND2x2_ASAP7_75t_L g14235 ( 
.A(n_14170),
.B(n_14087),
.Y(n_14235)
);

NOR2xp33_ASAP7_75t_L g14236 ( 
.A(n_14153),
.B(n_14214),
.Y(n_14236)
);

INVx1_ASAP7_75t_L g14237 ( 
.A(n_14137),
.Y(n_14237)
);

INVx2_ASAP7_75t_L g14238 ( 
.A(n_14122),
.Y(n_14238)
);

AND2x2_ASAP7_75t_L g14239 ( 
.A(n_14139),
.B(n_14079),
.Y(n_14239)
);

INVx1_ASAP7_75t_L g14240 ( 
.A(n_14115),
.Y(n_14240)
);

INVx1_ASAP7_75t_L g14241 ( 
.A(n_14145),
.Y(n_14241)
);

INVxp67_ASAP7_75t_L g14242 ( 
.A(n_14117),
.Y(n_14242)
);

INVx1_ASAP7_75t_L g14243 ( 
.A(n_14133),
.Y(n_14243)
);

AND2x2_ASAP7_75t_L g14244 ( 
.A(n_14140),
.B(n_14111),
.Y(n_14244)
);

OR2x2_ASAP7_75t_L g14245 ( 
.A(n_14134),
.B(n_14092),
.Y(n_14245)
);

INVxp67_ASAP7_75t_L g14246 ( 
.A(n_14203),
.Y(n_14246)
);

NAND2xp5_ASAP7_75t_L g14247 ( 
.A(n_14136),
.B(n_14086),
.Y(n_14247)
);

INVx1_ASAP7_75t_L g14248 ( 
.A(n_14156),
.Y(n_14248)
);

INVx1_ASAP7_75t_L g14249 ( 
.A(n_14177),
.Y(n_14249)
);

INVx1_ASAP7_75t_L g14250 ( 
.A(n_14142),
.Y(n_14250)
);

AND2x2_ASAP7_75t_L g14251 ( 
.A(n_14118),
.B(n_14107),
.Y(n_14251)
);

HB1xp67_ASAP7_75t_L g14252 ( 
.A(n_14182),
.Y(n_14252)
);

NAND2xp5_ASAP7_75t_L g14253 ( 
.A(n_14124),
.B(n_13992),
.Y(n_14253)
);

NAND2xp5_ASAP7_75t_L g14254 ( 
.A(n_14141),
.B(n_2394),
.Y(n_14254)
);

AND2x2_ASAP7_75t_L g14255 ( 
.A(n_14121),
.B(n_2394),
.Y(n_14255)
);

INVx1_ASAP7_75t_L g14256 ( 
.A(n_14138),
.Y(n_14256)
);

NOR2xp67_ASAP7_75t_SL g14257 ( 
.A(n_14183),
.B(n_2395),
.Y(n_14257)
);

CKINVDCx11_ASAP7_75t_R g14258 ( 
.A(n_14155),
.Y(n_14258)
);

INVx1_ASAP7_75t_L g14259 ( 
.A(n_14162),
.Y(n_14259)
);

AND2x2_ASAP7_75t_L g14260 ( 
.A(n_14154),
.B(n_2395),
.Y(n_14260)
);

NAND2xp5_ASAP7_75t_L g14261 ( 
.A(n_14172),
.B(n_2396),
.Y(n_14261)
);

INVx1_ASAP7_75t_L g14262 ( 
.A(n_14135),
.Y(n_14262)
);

INVx2_ASAP7_75t_L g14263 ( 
.A(n_14188),
.Y(n_14263)
);

INVx1_ASAP7_75t_L g14264 ( 
.A(n_14146),
.Y(n_14264)
);

NAND2xp5_ASAP7_75t_L g14265 ( 
.A(n_14128),
.B(n_14169),
.Y(n_14265)
);

OR2x2_ASAP7_75t_L g14266 ( 
.A(n_14114),
.B(n_2396),
.Y(n_14266)
);

AND2x4_ASAP7_75t_L g14267 ( 
.A(n_14159),
.B(n_2397),
.Y(n_14267)
);

AND2x2_ASAP7_75t_L g14268 ( 
.A(n_14143),
.B(n_2398),
.Y(n_14268)
);

INVx3_ASAP7_75t_L g14269 ( 
.A(n_14218),
.Y(n_14269)
);

NAND2xp5_ASAP7_75t_L g14270 ( 
.A(n_14119),
.B(n_2398),
.Y(n_14270)
);

NOR2xp33_ASAP7_75t_L g14271 ( 
.A(n_14168),
.B(n_2399),
.Y(n_14271)
);

NAND2xp5_ASAP7_75t_L g14272 ( 
.A(n_14152),
.B(n_2399),
.Y(n_14272)
);

INVx1_ASAP7_75t_L g14273 ( 
.A(n_14147),
.Y(n_14273)
);

AND2x2_ASAP7_75t_L g14274 ( 
.A(n_14163),
.B(n_2400),
.Y(n_14274)
);

AND2x2_ASAP7_75t_L g14275 ( 
.A(n_14208),
.B(n_2400),
.Y(n_14275)
);

INVx1_ASAP7_75t_L g14276 ( 
.A(n_14180),
.Y(n_14276)
);

HB1xp67_ASAP7_75t_L g14277 ( 
.A(n_14206),
.Y(n_14277)
);

INVx1_ASAP7_75t_L g14278 ( 
.A(n_14202),
.Y(n_14278)
);

NAND2xp5_ASAP7_75t_SL g14279 ( 
.A(n_14113),
.B(n_2401),
.Y(n_14279)
);

AND2x2_ASAP7_75t_L g14280 ( 
.A(n_14212),
.B(n_2401),
.Y(n_14280)
);

INVx1_ASAP7_75t_L g14281 ( 
.A(n_14164),
.Y(n_14281)
);

AND2x2_ASAP7_75t_L g14282 ( 
.A(n_14171),
.B(n_2402),
.Y(n_14282)
);

AND2x2_ASAP7_75t_L g14283 ( 
.A(n_14186),
.B(n_2402),
.Y(n_14283)
);

INVx1_ASAP7_75t_L g14284 ( 
.A(n_14181),
.Y(n_14284)
);

AND2x2_ASAP7_75t_L g14285 ( 
.A(n_14189),
.B(n_2403),
.Y(n_14285)
);

AND2x4_ASAP7_75t_L g14286 ( 
.A(n_14191),
.B(n_2403),
.Y(n_14286)
);

AND2x2_ASAP7_75t_L g14287 ( 
.A(n_14198),
.B(n_2404),
.Y(n_14287)
);

INVx1_ASAP7_75t_L g14288 ( 
.A(n_14179),
.Y(n_14288)
);

INVx2_ASAP7_75t_L g14289 ( 
.A(n_14221),
.Y(n_14289)
);

INVx1_ASAP7_75t_L g14290 ( 
.A(n_14176),
.Y(n_14290)
);

INVx1_ASAP7_75t_L g14291 ( 
.A(n_14201),
.Y(n_14291)
);

INVxp67_ASAP7_75t_L g14292 ( 
.A(n_14149),
.Y(n_14292)
);

OR2x2_ASAP7_75t_L g14293 ( 
.A(n_14151),
.B(n_14161),
.Y(n_14293)
);

OR2x2_ASAP7_75t_L g14294 ( 
.A(n_14157),
.B(n_2404),
.Y(n_14294)
);

INVx1_ASAP7_75t_L g14295 ( 
.A(n_14167),
.Y(n_14295)
);

INVx1_ASAP7_75t_L g14296 ( 
.A(n_14196),
.Y(n_14296)
);

INVxp67_ASAP7_75t_L g14297 ( 
.A(n_14194),
.Y(n_14297)
);

INVx2_ASAP7_75t_SL g14298 ( 
.A(n_14213),
.Y(n_14298)
);

AND2x2_ASAP7_75t_L g14299 ( 
.A(n_14130),
.B(n_2405),
.Y(n_14299)
);

NAND2xp5_ASAP7_75t_L g14300 ( 
.A(n_14131),
.B(n_2405),
.Y(n_14300)
);

AND2x2_ASAP7_75t_L g14301 ( 
.A(n_14178),
.B(n_2406),
.Y(n_14301)
);

NAND2xp5_ASAP7_75t_L g14302 ( 
.A(n_14165),
.B(n_2406),
.Y(n_14302)
);

INVx1_ASAP7_75t_L g14303 ( 
.A(n_14197),
.Y(n_14303)
);

INVx1_ASAP7_75t_L g14304 ( 
.A(n_14184),
.Y(n_14304)
);

AND2x2_ASAP7_75t_L g14305 ( 
.A(n_14217),
.B(n_2407),
.Y(n_14305)
);

INVx2_ASAP7_75t_L g14306 ( 
.A(n_14211),
.Y(n_14306)
);

AND2x2_ASAP7_75t_L g14307 ( 
.A(n_14160),
.B(n_2407),
.Y(n_14307)
);

INVx2_ASAP7_75t_SL g14308 ( 
.A(n_14210),
.Y(n_14308)
);

INVx1_ASAP7_75t_L g14309 ( 
.A(n_14216),
.Y(n_14309)
);

INVx1_ASAP7_75t_L g14310 ( 
.A(n_14226),
.Y(n_14310)
);

INVx2_ASAP7_75t_L g14311 ( 
.A(n_14225),
.Y(n_14311)
);

NOR2xp33_ASAP7_75t_L g14312 ( 
.A(n_14207),
.B(n_14144),
.Y(n_14312)
);

HB1xp67_ASAP7_75t_L g14313 ( 
.A(n_14209),
.Y(n_14313)
);

INVx4_ASAP7_75t_L g14314 ( 
.A(n_14223),
.Y(n_14314)
);

INVx1_ASAP7_75t_L g14315 ( 
.A(n_14166),
.Y(n_14315)
);

INVx2_ASAP7_75t_L g14316 ( 
.A(n_14127),
.Y(n_14316)
);

OR2x2_ASAP7_75t_L g14317 ( 
.A(n_14190),
.B(n_2408),
.Y(n_14317)
);

INVx1_ASAP7_75t_L g14318 ( 
.A(n_14227),
.Y(n_14318)
);

NAND2xp5_ASAP7_75t_L g14319 ( 
.A(n_14120),
.B(n_2408),
.Y(n_14319)
);

HB1xp67_ASAP7_75t_L g14320 ( 
.A(n_14222),
.Y(n_14320)
);

AND2x2_ASAP7_75t_L g14321 ( 
.A(n_14175),
.B(n_2409),
.Y(n_14321)
);

INVx1_ASAP7_75t_L g14322 ( 
.A(n_14220),
.Y(n_14322)
);

AND2x2_ASAP7_75t_SL g14323 ( 
.A(n_14129),
.B(n_2410),
.Y(n_14323)
);

INVx2_ASAP7_75t_L g14324 ( 
.A(n_14199),
.Y(n_14324)
);

BUFx2_ASAP7_75t_L g14325 ( 
.A(n_14224),
.Y(n_14325)
);

INVx2_ASAP7_75t_L g14326 ( 
.A(n_14187),
.Y(n_14326)
);

INVx1_ASAP7_75t_L g14327 ( 
.A(n_14200),
.Y(n_14327)
);

AND2x2_ASAP7_75t_L g14328 ( 
.A(n_14174),
.B(n_2410),
.Y(n_14328)
);

AND2x2_ASAP7_75t_L g14329 ( 
.A(n_14192),
.B(n_2411),
.Y(n_14329)
);

OR2x2_ASAP7_75t_L g14330 ( 
.A(n_14195),
.B(n_2412),
.Y(n_14330)
);

OAI21xp5_ASAP7_75t_L g14331 ( 
.A1(n_14126),
.A2(n_2412),
.B(n_2413),
.Y(n_14331)
);

AND2x2_ASAP7_75t_L g14332 ( 
.A(n_14215),
.B(n_2413),
.Y(n_14332)
);

NAND2xp5_ASAP7_75t_L g14333 ( 
.A(n_14158),
.B(n_2414),
.Y(n_14333)
);

AND2x2_ASAP7_75t_L g14334 ( 
.A(n_14219),
.B(n_2414),
.Y(n_14334)
);

AND2x2_ASAP7_75t_L g14335 ( 
.A(n_14148),
.B(n_2415),
.Y(n_14335)
);

AND2x2_ASAP7_75t_L g14336 ( 
.A(n_14173),
.B(n_2416),
.Y(n_14336)
);

AND2x4_ASAP7_75t_L g14337 ( 
.A(n_14193),
.B(n_2416),
.Y(n_14337)
);

INVx2_ASAP7_75t_L g14338 ( 
.A(n_14132),
.Y(n_14338)
);

INVx1_ASAP7_75t_L g14339 ( 
.A(n_14204),
.Y(n_14339)
);

OR2x2_ASAP7_75t_L g14340 ( 
.A(n_14185),
.B(n_2417),
.Y(n_14340)
);

AND2x2_ASAP7_75t_L g14341 ( 
.A(n_14116),
.B(n_2417),
.Y(n_14341)
);

NAND2xp5_ASAP7_75t_L g14342 ( 
.A(n_14214),
.B(n_2418),
.Y(n_14342)
);

AND2x4_ASAP7_75t_SL g14343 ( 
.A(n_14123),
.B(n_2418),
.Y(n_14343)
);

OR2x2_ASAP7_75t_L g14344 ( 
.A(n_14185),
.B(n_2419),
.Y(n_14344)
);

AND2x2_ASAP7_75t_L g14345 ( 
.A(n_14116),
.B(n_2419),
.Y(n_14345)
);

OR2x2_ASAP7_75t_L g14346 ( 
.A(n_14185),
.B(n_2420),
.Y(n_14346)
);

INVx2_ASAP7_75t_L g14347 ( 
.A(n_14214),
.Y(n_14347)
);

INVx2_ASAP7_75t_L g14348 ( 
.A(n_14214),
.Y(n_14348)
);

INVx1_ASAP7_75t_L g14349 ( 
.A(n_14205),
.Y(n_14349)
);

NAND2xp5_ASAP7_75t_L g14350 ( 
.A(n_14214),
.B(n_2420),
.Y(n_14350)
);

INVx1_ASAP7_75t_L g14351 ( 
.A(n_14205),
.Y(n_14351)
);

INVx1_ASAP7_75t_L g14352 ( 
.A(n_14205),
.Y(n_14352)
);

AND2x2_ASAP7_75t_L g14353 ( 
.A(n_14229),
.B(n_2421),
.Y(n_14353)
);

AND2x2_ASAP7_75t_L g14354 ( 
.A(n_14228),
.B(n_14235),
.Y(n_14354)
);

AND2x2_ASAP7_75t_L g14355 ( 
.A(n_14255),
.B(n_2421),
.Y(n_14355)
);

NAND2xp5_ASAP7_75t_L g14356 ( 
.A(n_14230),
.B(n_2422),
.Y(n_14356)
);

NAND2xp5_ASAP7_75t_L g14357 ( 
.A(n_14347),
.B(n_14348),
.Y(n_14357)
);

AND2x4_ASAP7_75t_L g14358 ( 
.A(n_14231),
.B(n_2423),
.Y(n_14358)
);

INVx1_ASAP7_75t_L g14359 ( 
.A(n_14277),
.Y(n_14359)
);

NAND2xp5_ASAP7_75t_L g14360 ( 
.A(n_14236),
.B(n_2424),
.Y(n_14360)
);

AND2x2_ASAP7_75t_L g14361 ( 
.A(n_14349),
.B(n_2424),
.Y(n_14361)
);

BUFx2_ASAP7_75t_L g14362 ( 
.A(n_14252),
.Y(n_14362)
);

AND2x2_ASAP7_75t_L g14363 ( 
.A(n_14351),
.B(n_2425),
.Y(n_14363)
);

NAND2xp5_ASAP7_75t_L g14364 ( 
.A(n_14352),
.B(n_2425),
.Y(n_14364)
);

NAND2xp5_ASAP7_75t_L g14365 ( 
.A(n_14297),
.B(n_2426),
.Y(n_14365)
);

OR2x2_ASAP7_75t_L g14366 ( 
.A(n_14232),
.B(n_2426),
.Y(n_14366)
);

OAI21xp5_ASAP7_75t_L g14367 ( 
.A1(n_14246),
.A2(n_2427),
.B(n_2428),
.Y(n_14367)
);

NAND2xp5_ASAP7_75t_L g14368 ( 
.A(n_14341),
.B(n_2427),
.Y(n_14368)
);

INVx1_ASAP7_75t_L g14369 ( 
.A(n_14350),
.Y(n_14369)
);

INVx1_ASAP7_75t_L g14370 ( 
.A(n_14342),
.Y(n_14370)
);

INVx1_ASAP7_75t_L g14371 ( 
.A(n_14340),
.Y(n_14371)
);

AND2x2_ASAP7_75t_L g14372 ( 
.A(n_14260),
.B(n_2429),
.Y(n_14372)
);

INVx1_ASAP7_75t_L g14373 ( 
.A(n_14344),
.Y(n_14373)
);

AND2x2_ASAP7_75t_L g14374 ( 
.A(n_14244),
.B(n_2430),
.Y(n_14374)
);

INVx2_ASAP7_75t_L g14375 ( 
.A(n_14346),
.Y(n_14375)
);

NAND2xp5_ASAP7_75t_L g14376 ( 
.A(n_14345),
.B(n_14257),
.Y(n_14376)
);

INVx1_ASAP7_75t_L g14377 ( 
.A(n_14313),
.Y(n_14377)
);

NOR2xp33_ASAP7_75t_L g14378 ( 
.A(n_14314),
.B(n_2430),
.Y(n_14378)
);

AND2x2_ASAP7_75t_L g14379 ( 
.A(n_14251),
.B(n_2431),
.Y(n_14379)
);

INVx2_ASAP7_75t_L g14380 ( 
.A(n_14258),
.Y(n_14380)
);

NAND2xp5_ASAP7_75t_L g14381 ( 
.A(n_14298),
.B(n_2431),
.Y(n_14381)
);

AND2x2_ASAP7_75t_L g14382 ( 
.A(n_14233),
.B(n_2432),
.Y(n_14382)
);

NAND2xp5_ASAP7_75t_SL g14383 ( 
.A(n_14249),
.B(n_2432),
.Y(n_14383)
);

AND2x2_ASAP7_75t_L g14384 ( 
.A(n_14299),
.B(n_14241),
.Y(n_14384)
);

INVx2_ASAP7_75t_L g14385 ( 
.A(n_14343),
.Y(n_14385)
);

INVx1_ASAP7_75t_SL g14386 ( 
.A(n_14245),
.Y(n_14386)
);

NAND3xp33_ASAP7_75t_L g14387 ( 
.A(n_14237),
.B(n_2433),
.C(n_2434),
.Y(n_14387)
);

OR2x2_ASAP7_75t_L g14388 ( 
.A(n_14234),
.B(n_2433),
.Y(n_14388)
);

OR2x2_ASAP7_75t_L g14389 ( 
.A(n_14247),
.B(n_2434),
.Y(n_14389)
);

INVx2_ASAP7_75t_L g14390 ( 
.A(n_14269),
.Y(n_14390)
);

NOR2x1_ASAP7_75t_L g14391 ( 
.A(n_14311),
.B(n_2435),
.Y(n_14391)
);

INVx1_ASAP7_75t_L g14392 ( 
.A(n_14275),
.Y(n_14392)
);

AND2x2_ASAP7_75t_L g14393 ( 
.A(n_14264),
.B(n_2435),
.Y(n_14393)
);

NAND2x1_ASAP7_75t_SL g14394 ( 
.A(n_14305),
.B(n_14320),
.Y(n_14394)
);

NOR2xp33_ASAP7_75t_L g14395 ( 
.A(n_14243),
.B(n_2436),
.Y(n_14395)
);

NAND2xp5_ASAP7_75t_L g14396 ( 
.A(n_14337),
.B(n_2436),
.Y(n_14396)
);

INVxp33_ASAP7_75t_SL g14397 ( 
.A(n_14239),
.Y(n_14397)
);

AND2x2_ASAP7_75t_L g14398 ( 
.A(n_14280),
.B(n_2437),
.Y(n_14398)
);

AND2x2_ASAP7_75t_L g14399 ( 
.A(n_14256),
.B(n_2437),
.Y(n_14399)
);

NOR2x1p5_ASAP7_75t_L g14400 ( 
.A(n_14253),
.B(n_2438),
.Y(n_14400)
);

OR2x2_ASAP7_75t_L g14401 ( 
.A(n_14308),
.B(n_2438),
.Y(n_14401)
);

INVx2_ASAP7_75t_L g14402 ( 
.A(n_14286),
.Y(n_14402)
);

INVx1_ASAP7_75t_L g14403 ( 
.A(n_14285),
.Y(n_14403)
);

AND2x2_ASAP7_75t_L g14404 ( 
.A(n_14259),
.B(n_2439),
.Y(n_14404)
);

INVx3_ASAP7_75t_L g14405 ( 
.A(n_14267),
.Y(n_14405)
);

AND2x4_ASAP7_75t_L g14406 ( 
.A(n_14287),
.B(n_14289),
.Y(n_14406)
);

AND3x2_ASAP7_75t_L g14407 ( 
.A(n_14325),
.B(n_14248),
.C(n_14242),
.Y(n_14407)
);

AND2x2_ASAP7_75t_L g14408 ( 
.A(n_14306),
.B(n_2439),
.Y(n_14408)
);

AND2x2_ASAP7_75t_L g14409 ( 
.A(n_14238),
.B(n_2440),
.Y(n_14409)
);

INVx1_ASAP7_75t_L g14410 ( 
.A(n_14282),
.Y(n_14410)
);

AND2x2_ASAP7_75t_L g14411 ( 
.A(n_14284),
.B(n_2440),
.Y(n_14411)
);

NAND4xp75_ASAP7_75t_L g14412 ( 
.A(n_14323),
.B(n_2443),
.C(n_2441),
.D(n_2442),
.Y(n_14412)
);

NAND2xp5_ASAP7_75t_L g14413 ( 
.A(n_14240),
.B(n_2441),
.Y(n_14413)
);

AND2x2_ASAP7_75t_L g14414 ( 
.A(n_14291),
.B(n_2442),
.Y(n_14414)
);

OR2x2_ASAP7_75t_L g14415 ( 
.A(n_14317),
.B(n_2443),
.Y(n_14415)
);

NAND2xp5_ASAP7_75t_L g14416 ( 
.A(n_14283),
.B(n_2444),
.Y(n_14416)
);

INVx1_ASAP7_75t_L g14417 ( 
.A(n_14261),
.Y(n_14417)
);

NAND2xp5_ASAP7_75t_L g14418 ( 
.A(n_14274),
.B(n_2444),
.Y(n_14418)
);

NAND2xp5_ASAP7_75t_L g14419 ( 
.A(n_14268),
.B(n_2445),
.Y(n_14419)
);

INVx1_ASAP7_75t_L g14420 ( 
.A(n_14294),
.Y(n_14420)
);

INVx1_ASAP7_75t_L g14421 ( 
.A(n_14307),
.Y(n_14421)
);

NAND2xp5_ASAP7_75t_L g14422 ( 
.A(n_14278),
.B(n_2446),
.Y(n_14422)
);

INVx2_ASAP7_75t_SL g14423 ( 
.A(n_14301),
.Y(n_14423)
);

AND2x2_ASAP7_75t_L g14424 ( 
.A(n_14273),
.B(n_2446),
.Y(n_14424)
);

NAND2xp5_ASAP7_75t_L g14425 ( 
.A(n_14250),
.B(n_2447),
.Y(n_14425)
);

AND2x2_ASAP7_75t_L g14426 ( 
.A(n_14309),
.B(n_2447),
.Y(n_14426)
);

OR2x2_ASAP7_75t_L g14427 ( 
.A(n_14300),
.B(n_2448),
.Y(n_14427)
);

INVx2_ASAP7_75t_L g14428 ( 
.A(n_14330),
.Y(n_14428)
);

INVx2_ASAP7_75t_SL g14429 ( 
.A(n_14329),
.Y(n_14429)
);

HB1xp67_ASAP7_75t_L g14430 ( 
.A(n_14288),
.Y(n_14430)
);

AND2x2_ASAP7_75t_L g14431 ( 
.A(n_14322),
.B(n_2448),
.Y(n_14431)
);

NAND2xp5_ASAP7_75t_L g14432 ( 
.A(n_14335),
.B(n_2449),
.Y(n_14432)
);

INVx1_ASAP7_75t_L g14433 ( 
.A(n_14332),
.Y(n_14433)
);

INVx1_ASAP7_75t_L g14434 ( 
.A(n_14334),
.Y(n_14434)
);

INVx2_ASAP7_75t_L g14435 ( 
.A(n_14293),
.Y(n_14435)
);

NAND2xp5_ASAP7_75t_L g14436 ( 
.A(n_14276),
.B(n_14290),
.Y(n_14436)
);

INVx1_ASAP7_75t_L g14437 ( 
.A(n_14321),
.Y(n_14437)
);

INVx1_ASAP7_75t_SL g14438 ( 
.A(n_14254),
.Y(n_14438)
);

AND2x4_ASAP7_75t_L g14439 ( 
.A(n_14263),
.B(n_2449),
.Y(n_14439)
);

INVx2_ASAP7_75t_L g14440 ( 
.A(n_14296),
.Y(n_14440)
);

INVx1_ASAP7_75t_L g14441 ( 
.A(n_14265),
.Y(n_14441)
);

AND2x2_ASAP7_75t_L g14442 ( 
.A(n_14303),
.B(n_2450),
.Y(n_14442)
);

INVx2_ASAP7_75t_L g14443 ( 
.A(n_14304),
.Y(n_14443)
);

INVx2_ASAP7_75t_L g14444 ( 
.A(n_14328),
.Y(n_14444)
);

INVx1_ASAP7_75t_L g14445 ( 
.A(n_14270),
.Y(n_14445)
);

HB1xp67_ASAP7_75t_L g14446 ( 
.A(n_14316),
.Y(n_14446)
);

INVx1_ASAP7_75t_L g14447 ( 
.A(n_14272),
.Y(n_14447)
);

AND2x2_ASAP7_75t_L g14448 ( 
.A(n_14310),
.B(n_2450),
.Y(n_14448)
);

NAND2xp5_ASAP7_75t_L g14449 ( 
.A(n_14338),
.B(n_14262),
.Y(n_14449)
);

INVxp67_ASAP7_75t_L g14450 ( 
.A(n_14271),
.Y(n_14450)
);

AND2x4_ASAP7_75t_L g14451 ( 
.A(n_14281),
.B(n_2451),
.Y(n_14451)
);

INVx1_ASAP7_75t_L g14452 ( 
.A(n_14266),
.Y(n_14452)
);

AND2x2_ASAP7_75t_L g14453 ( 
.A(n_14331),
.B(n_2451),
.Y(n_14453)
);

AND2x2_ASAP7_75t_L g14454 ( 
.A(n_14336),
.B(n_2452),
.Y(n_14454)
);

INVx1_ASAP7_75t_L g14455 ( 
.A(n_14333),
.Y(n_14455)
);

INVx1_ASAP7_75t_L g14456 ( 
.A(n_14315),
.Y(n_14456)
);

NAND2xp5_ASAP7_75t_L g14457 ( 
.A(n_14318),
.B(n_2452),
.Y(n_14457)
);

INVx1_ASAP7_75t_L g14458 ( 
.A(n_14324),
.Y(n_14458)
);

INVx2_ASAP7_75t_L g14459 ( 
.A(n_14326),
.Y(n_14459)
);

INVx1_ASAP7_75t_L g14460 ( 
.A(n_14312),
.Y(n_14460)
);

AND2x2_ASAP7_75t_L g14461 ( 
.A(n_14292),
.B(n_2453),
.Y(n_14461)
);

INVx2_ASAP7_75t_L g14462 ( 
.A(n_14295),
.Y(n_14462)
);

INVx1_ASAP7_75t_L g14463 ( 
.A(n_14319),
.Y(n_14463)
);

INVx2_ASAP7_75t_L g14464 ( 
.A(n_14327),
.Y(n_14464)
);

INVx1_ASAP7_75t_L g14465 ( 
.A(n_14302),
.Y(n_14465)
);

AND2x2_ASAP7_75t_L g14466 ( 
.A(n_14279),
.B(n_2453),
.Y(n_14466)
);

NAND4xp75_ASAP7_75t_L g14467 ( 
.A(n_14339),
.B(n_2457),
.C(n_2454),
.D(n_2455),
.Y(n_14467)
);

INVx2_ASAP7_75t_L g14468 ( 
.A(n_14230),
.Y(n_14468)
);

NAND2xp5_ASAP7_75t_L g14469 ( 
.A(n_14230),
.B(n_2454),
.Y(n_14469)
);

NAND2xp5_ASAP7_75t_L g14470 ( 
.A(n_14230),
.B(n_2455),
.Y(n_14470)
);

INVx1_ASAP7_75t_SL g14471 ( 
.A(n_14258),
.Y(n_14471)
);

OAI33xp33_ASAP7_75t_L g14472 ( 
.A1(n_14249),
.A2(n_2459),
.A3(n_2461),
.B1(n_2457),
.B2(n_2458),
.B3(n_2460),
.Y(n_14472)
);

INVx1_ASAP7_75t_L g14473 ( 
.A(n_14277),
.Y(n_14473)
);

OR2x2_ASAP7_75t_L g14474 ( 
.A(n_14230),
.B(n_2458),
.Y(n_14474)
);

INVx1_ASAP7_75t_L g14475 ( 
.A(n_14277),
.Y(n_14475)
);

INVx1_ASAP7_75t_L g14476 ( 
.A(n_14277),
.Y(n_14476)
);

NAND2xp5_ASAP7_75t_L g14477 ( 
.A(n_14230),
.B(n_2459),
.Y(n_14477)
);

NAND2xp5_ASAP7_75t_L g14478 ( 
.A(n_14230),
.B(n_2460),
.Y(n_14478)
);

INVx1_ASAP7_75t_L g14479 ( 
.A(n_14277),
.Y(n_14479)
);

INVx1_ASAP7_75t_L g14480 ( 
.A(n_14277),
.Y(n_14480)
);

INVx1_ASAP7_75t_L g14481 ( 
.A(n_14277),
.Y(n_14481)
);

INVx1_ASAP7_75t_L g14482 ( 
.A(n_14277),
.Y(n_14482)
);

AND2x4_ASAP7_75t_L g14483 ( 
.A(n_14229),
.B(n_2461),
.Y(n_14483)
);

INVx1_ASAP7_75t_L g14484 ( 
.A(n_14277),
.Y(n_14484)
);

NAND2xp5_ASAP7_75t_L g14485 ( 
.A(n_14230),
.B(n_2462),
.Y(n_14485)
);

INVx1_ASAP7_75t_L g14486 ( 
.A(n_14277),
.Y(n_14486)
);

INVx1_ASAP7_75t_L g14487 ( 
.A(n_14277),
.Y(n_14487)
);

OR2x2_ASAP7_75t_L g14488 ( 
.A(n_14230),
.B(n_2462),
.Y(n_14488)
);

INVx1_ASAP7_75t_L g14489 ( 
.A(n_14277),
.Y(n_14489)
);

INVx1_ASAP7_75t_L g14490 ( 
.A(n_14277),
.Y(n_14490)
);

AND2x2_ASAP7_75t_L g14491 ( 
.A(n_14229),
.B(n_2463),
.Y(n_14491)
);

OR2x2_ASAP7_75t_L g14492 ( 
.A(n_14230),
.B(n_2464),
.Y(n_14492)
);

AND2x2_ASAP7_75t_L g14493 ( 
.A(n_14229),
.B(n_2465),
.Y(n_14493)
);

OR2x2_ASAP7_75t_L g14494 ( 
.A(n_14230),
.B(n_2466),
.Y(n_14494)
);

INVx1_ASAP7_75t_L g14495 ( 
.A(n_14277),
.Y(n_14495)
);

NAND2xp5_ASAP7_75t_L g14496 ( 
.A(n_14230),
.B(n_2466),
.Y(n_14496)
);

AND2x2_ASAP7_75t_L g14497 ( 
.A(n_14229),
.B(n_2467),
.Y(n_14497)
);

AND2x2_ASAP7_75t_SL g14498 ( 
.A(n_14314),
.B(n_2467),
.Y(n_14498)
);

INVx2_ASAP7_75t_L g14499 ( 
.A(n_14230),
.Y(n_14499)
);

NOR2x1p5_ASAP7_75t_SL g14500 ( 
.A(n_14245),
.B(n_2468),
.Y(n_14500)
);

AND2x2_ASAP7_75t_L g14501 ( 
.A(n_14229),
.B(n_2468),
.Y(n_14501)
);

NAND2xp5_ASAP7_75t_L g14502 ( 
.A(n_14230),
.B(n_2469),
.Y(n_14502)
);

AND2x2_ASAP7_75t_L g14503 ( 
.A(n_14471),
.B(n_2469),
.Y(n_14503)
);

INVx1_ASAP7_75t_L g14504 ( 
.A(n_14394),
.Y(n_14504)
);

OR2x2_ASAP7_75t_L g14505 ( 
.A(n_14386),
.B(n_14376),
.Y(n_14505)
);

INVx1_ASAP7_75t_L g14506 ( 
.A(n_14362),
.Y(n_14506)
);

AND2x2_ASAP7_75t_L g14507 ( 
.A(n_14380),
.B(n_2470),
.Y(n_14507)
);

INVx1_ASAP7_75t_L g14508 ( 
.A(n_14354),
.Y(n_14508)
);

NAND2xp5_ASAP7_75t_L g14509 ( 
.A(n_14498),
.B(n_2470),
.Y(n_14509)
);

INVx2_ASAP7_75t_L g14510 ( 
.A(n_14407),
.Y(n_14510)
);

INVx1_ASAP7_75t_L g14511 ( 
.A(n_14500),
.Y(n_14511)
);

AND2x2_ASAP7_75t_L g14512 ( 
.A(n_14384),
.B(n_2471),
.Y(n_14512)
);

INVx2_ASAP7_75t_L g14513 ( 
.A(n_14353),
.Y(n_14513)
);

INVxp67_ASAP7_75t_L g14514 ( 
.A(n_14430),
.Y(n_14514)
);

NOR2xp33_ASAP7_75t_L g14515 ( 
.A(n_14397),
.B(n_2471),
.Y(n_14515)
);

INVx1_ASAP7_75t_L g14516 ( 
.A(n_14491),
.Y(n_14516)
);

NOR2x1_ASAP7_75t_L g14517 ( 
.A(n_14391),
.B(n_2472),
.Y(n_14517)
);

AND2x2_ASAP7_75t_L g14518 ( 
.A(n_14385),
.B(n_2472),
.Y(n_14518)
);

AND2x2_ASAP7_75t_L g14519 ( 
.A(n_14405),
.B(n_2473),
.Y(n_14519)
);

A2O1A1Ixp33_ASAP7_75t_L g14520 ( 
.A1(n_14378),
.A2(n_2475),
.B(n_2473),
.C(n_2474),
.Y(n_14520)
);

HB1xp67_ASAP7_75t_L g14521 ( 
.A(n_14400),
.Y(n_14521)
);

INVxp33_ASAP7_75t_L g14522 ( 
.A(n_14446),
.Y(n_14522)
);

OR2x2_ASAP7_75t_L g14523 ( 
.A(n_14401),
.B(n_14366),
.Y(n_14523)
);

NOR2x1_ASAP7_75t_L g14524 ( 
.A(n_14467),
.B(n_2475),
.Y(n_14524)
);

AOI21xp5_ASAP7_75t_L g14525 ( 
.A1(n_14357),
.A2(n_2476),
.B(n_2477),
.Y(n_14525)
);

INVx1_ASAP7_75t_L g14526 ( 
.A(n_14493),
.Y(n_14526)
);

BUFx2_ASAP7_75t_L g14527 ( 
.A(n_14377),
.Y(n_14527)
);

AOI22xp33_ASAP7_75t_SL g14528 ( 
.A1(n_14468),
.A2(n_2479),
.B1(n_2476),
.B2(n_2478),
.Y(n_14528)
);

INVx2_ASAP7_75t_L g14529 ( 
.A(n_14497),
.Y(n_14529)
);

NAND2xp5_ASAP7_75t_L g14530 ( 
.A(n_14501),
.B(n_2478),
.Y(n_14530)
);

OR2x2_ASAP7_75t_L g14531 ( 
.A(n_14499),
.B(n_2479),
.Y(n_14531)
);

AND2x2_ASAP7_75t_L g14532 ( 
.A(n_14406),
.B(n_2480),
.Y(n_14532)
);

INVx1_ASAP7_75t_L g14533 ( 
.A(n_14374),
.Y(n_14533)
);

AND2x2_ASAP7_75t_L g14534 ( 
.A(n_14402),
.B(n_2481),
.Y(n_14534)
);

INVx1_ASAP7_75t_L g14535 ( 
.A(n_14355),
.Y(n_14535)
);

NAND2xp5_ASAP7_75t_L g14536 ( 
.A(n_14379),
.B(n_2481),
.Y(n_14536)
);

INVx2_ASAP7_75t_L g14537 ( 
.A(n_14415),
.Y(n_14537)
);

INVx1_ASAP7_75t_L g14538 ( 
.A(n_14382),
.Y(n_14538)
);

INVx1_ASAP7_75t_SL g14539 ( 
.A(n_14372),
.Y(n_14539)
);

AND2x2_ASAP7_75t_L g14540 ( 
.A(n_14408),
.B(n_2482),
.Y(n_14540)
);

NOR2xp67_ASAP7_75t_SL g14541 ( 
.A(n_14412),
.B(n_2482),
.Y(n_14541)
);

INVx2_ASAP7_75t_L g14542 ( 
.A(n_14483),
.Y(n_14542)
);

INVx1_ASAP7_75t_L g14543 ( 
.A(n_14398),
.Y(n_14543)
);

AOI22xp33_ASAP7_75t_L g14544 ( 
.A1(n_14390),
.A2(n_14435),
.B1(n_14443),
.B2(n_14440),
.Y(n_14544)
);

INVx1_ASAP7_75t_L g14545 ( 
.A(n_14361),
.Y(n_14545)
);

INVx2_ASAP7_75t_SL g14546 ( 
.A(n_14358),
.Y(n_14546)
);

AND2x2_ASAP7_75t_L g14547 ( 
.A(n_14409),
.B(n_2483),
.Y(n_14547)
);

INVx1_ASAP7_75t_L g14548 ( 
.A(n_14363),
.Y(n_14548)
);

INVx1_ASAP7_75t_L g14549 ( 
.A(n_14393),
.Y(n_14549)
);

INVx1_ASAP7_75t_L g14550 ( 
.A(n_14399),
.Y(n_14550)
);

INVx1_ASAP7_75t_L g14551 ( 
.A(n_14404),
.Y(n_14551)
);

AND2x2_ASAP7_75t_L g14552 ( 
.A(n_14375),
.B(n_2483),
.Y(n_14552)
);

AND2x2_ASAP7_75t_L g14553 ( 
.A(n_14429),
.B(n_14410),
.Y(n_14553)
);

BUFx2_ASAP7_75t_SL g14554 ( 
.A(n_14451),
.Y(n_14554)
);

INVx1_ASAP7_75t_SL g14555 ( 
.A(n_14389),
.Y(n_14555)
);

OR2x2_ASAP7_75t_L g14556 ( 
.A(n_14365),
.B(n_2484),
.Y(n_14556)
);

INVxp67_ASAP7_75t_SL g14557 ( 
.A(n_14359),
.Y(n_14557)
);

INVx2_ASAP7_75t_L g14558 ( 
.A(n_14474),
.Y(n_14558)
);

INVxp67_ASAP7_75t_L g14559 ( 
.A(n_14395),
.Y(n_14559)
);

NAND2xp5_ASAP7_75t_L g14560 ( 
.A(n_14439),
.B(n_2484),
.Y(n_14560)
);

INVx1_ASAP7_75t_L g14561 ( 
.A(n_14488),
.Y(n_14561)
);

NAND2xp5_ASAP7_75t_L g14562 ( 
.A(n_14411),
.B(n_2485),
.Y(n_14562)
);

OR2x2_ASAP7_75t_L g14563 ( 
.A(n_14381),
.B(n_14360),
.Y(n_14563)
);

INVx1_ASAP7_75t_L g14564 ( 
.A(n_14492),
.Y(n_14564)
);

INVx3_ASAP7_75t_L g14565 ( 
.A(n_14494),
.Y(n_14565)
);

INVx1_ASAP7_75t_L g14566 ( 
.A(n_14388),
.Y(n_14566)
);

OR2x2_ASAP7_75t_L g14567 ( 
.A(n_14371),
.B(n_2486),
.Y(n_14567)
);

NOR2x1_ASAP7_75t_L g14568 ( 
.A(n_14387),
.B(n_2486),
.Y(n_14568)
);

AOI22xp33_ASAP7_75t_L g14569 ( 
.A1(n_14465),
.A2(n_2489),
.B1(n_2487),
.B2(n_2488),
.Y(n_14569)
);

INVx1_ASAP7_75t_L g14570 ( 
.A(n_14414),
.Y(n_14570)
);

OR2x2_ASAP7_75t_L g14571 ( 
.A(n_14373),
.B(n_2487),
.Y(n_14571)
);

INVx1_ASAP7_75t_L g14572 ( 
.A(n_14426),
.Y(n_14572)
);

INVx1_ASAP7_75t_L g14573 ( 
.A(n_14431),
.Y(n_14573)
);

AND2x2_ASAP7_75t_L g14574 ( 
.A(n_14392),
.B(n_2488),
.Y(n_14574)
);

AOI22xp5_ASAP7_75t_L g14575 ( 
.A1(n_14460),
.A2(n_2491),
.B1(n_2489),
.B2(n_2490),
.Y(n_14575)
);

NAND2xp5_ASAP7_75t_L g14576 ( 
.A(n_14424),
.B(n_2490),
.Y(n_14576)
);

HB1xp67_ASAP7_75t_L g14577 ( 
.A(n_14473),
.Y(n_14577)
);

AND2x2_ASAP7_75t_L g14578 ( 
.A(n_14403),
.B(n_2491),
.Y(n_14578)
);

INVx1_ASAP7_75t_L g14579 ( 
.A(n_14442),
.Y(n_14579)
);

NAND2xp5_ASAP7_75t_L g14580 ( 
.A(n_14448),
.B(n_2492),
.Y(n_14580)
);

INVxp67_ASAP7_75t_SL g14581 ( 
.A(n_14475),
.Y(n_14581)
);

INVx2_ASAP7_75t_L g14582 ( 
.A(n_14427),
.Y(n_14582)
);

NOR2xp33_ASAP7_75t_L g14583 ( 
.A(n_14421),
.B(n_2492),
.Y(n_14583)
);

AND2x2_ASAP7_75t_L g14584 ( 
.A(n_14423),
.B(n_2493),
.Y(n_14584)
);

AND2x2_ASAP7_75t_L g14585 ( 
.A(n_14444),
.B(n_14433),
.Y(n_14585)
);

AND2x2_ASAP7_75t_L g14586 ( 
.A(n_14434),
.B(n_2494),
.Y(n_14586)
);

INVx1_ASAP7_75t_L g14587 ( 
.A(n_14368),
.Y(n_14587)
);

INVx1_ASAP7_75t_L g14588 ( 
.A(n_14396),
.Y(n_14588)
);

INVx2_ASAP7_75t_L g14589 ( 
.A(n_14454),
.Y(n_14589)
);

INVx1_ASAP7_75t_L g14590 ( 
.A(n_14476),
.Y(n_14590)
);

OR2x2_ASAP7_75t_L g14591 ( 
.A(n_14356),
.B(n_2494),
.Y(n_14591)
);

INVx1_ASAP7_75t_L g14592 ( 
.A(n_14479),
.Y(n_14592)
);

INVx1_ASAP7_75t_L g14593 ( 
.A(n_14480),
.Y(n_14593)
);

OR2x2_ASAP7_75t_L g14594 ( 
.A(n_14502),
.B(n_2495),
.Y(n_14594)
);

AND2x2_ASAP7_75t_L g14595 ( 
.A(n_14453),
.B(n_2495),
.Y(n_14595)
);

OR2x2_ASAP7_75t_L g14596 ( 
.A(n_14496),
.B(n_2496),
.Y(n_14596)
);

INVx1_ASAP7_75t_L g14597 ( 
.A(n_14481),
.Y(n_14597)
);

NOR3xp33_ASAP7_75t_L g14598 ( 
.A(n_14449),
.B(n_2496),
.C(n_2497),
.Y(n_14598)
);

INVx2_ASAP7_75t_L g14599 ( 
.A(n_14482),
.Y(n_14599)
);

INVx1_ASAP7_75t_SL g14600 ( 
.A(n_14466),
.Y(n_14600)
);

NAND2xp5_ASAP7_75t_L g14601 ( 
.A(n_14461),
.B(n_2497),
.Y(n_14601)
);

INVxp67_ASAP7_75t_SL g14602 ( 
.A(n_14484),
.Y(n_14602)
);

AND2x2_ASAP7_75t_L g14603 ( 
.A(n_14437),
.B(n_2498),
.Y(n_14603)
);

NAND2xp5_ASAP7_75t_L g14604 ( 
.A(n_14420),
.B(n_2498),
.Y(n_14604)
);

INVxp67_ASAP7_75t_L g14605 ( 
.A(n_14416),
.Y(n_14605)
);

INVx1_ASAP7_75t_L g14606 ( 
.A(n_14486),
.Y(n_14606)
);

AND2x4_ASAP7_75t_L g14607 ( 
.A(n_14459),
.B(n_2499),
.Y(n_14607)
);

INVx1_ASAP7_75t_L g14608 ( 
.A(n_14487),
.Y(n_14608)
);

AND2x2_ASAP7_75t_L g14609 ( 
.A(n_14438),
.B(n_2499),
.Y(n_14609)
);

NAND2x1p5_ASAP7_75t_L g14610 ( 
.A(n_14383),
.B(n_14452),
.Y(n_14610)
);

NOR2x1_ASAP7_75t_L g14611 ( 
.A(n_14489),
.B(n_2500),
.Y(n_14611)
);

AND2x2_ASAP7_75t_L g14612 ( 
.A(n_14428),
.B(n_2500),
.Y(n_14612)
);

AND2x2_ASAP7_75t_L g14613 ( 
.A(n_14369),
.B(n_2501),
.Y(n_14613)
);

OAI22xp33_ASAP7_75t_L g14614 ( 
.A1(n_14432),
.A2(n_2503),
.B1(n_2501),
.B2(n_2502),
.Y(n_14614)
);

NAND2xp5_ASAP7_75t_L g14615 ( 
.A(n_14490),
.B(n_2502),
.Y(n_14615)
);

AND2x2_ASAP7_75t_L g14616 ( 
.A(n_14370),
.B(n_2503),
.Y(n_14616)
);

AND2x4_ASAP7_75t_L g14617 ( 
.A(n_14462),
.B(n_2504),
.Y(n_14617)
);

INVxp67_ASAP7_75t_SL g14618 ( 
.A(n_14495),
.Y(n_14618)
);

NOR2xp33_ASAP7_75t_L g14619 ( 
.A(n_14472),
.B(n_2504),
.Y(n_14619)
);

OAI21xp33_ASAP7_75t_L g14620 ( 
.A1(n_14436),
.A2(n_2505),
.B(n_2506),
.Y(n_14620)
);

INVx1_ASAP7_75t_L g14621 ( 
.A(n_14469),
.Y(n_14621)
);

NAND2xp5_ASAP7_75t_L g14622 ( 
.A(n_14463),
.B(n_2505),
.Y(n_14622)
);

AND2x2_ASAP7_75t_L g14623 ( 
.A(n_14455),
.B(n_2506),
.Y(n_14623)
);

AND2x2_ASAP7_75t_L g14624 ( 
.A(n_14367),
.B(n_2508),
.Y(n_14624)
);

AND2x2_ASAP7_75t_L g14625 ( 
.A(n_14450),
.B(n_2508),
.Y(n_14625)
);

NOR2xp33_ASAP7_75t_L g14626 ( 
.A(n_14419),
.B(n_2509),
.Y(n_14626)
);

OR2x2_ASAP7_75t_L g14627 ( 
.A(n_14485),
.B(n_2509),
.Y(n_14627)
);

AOI22xp5_ASAP7_75t_L g14628 ( 
.A1(n_14441),
.A2(n_2512),
.B1(n_2510),
.B2(n_2511),
.Y(n_14628)
);

INVx1_ASAP7_75t_L g14629 ( 
.A(n_14470),
.Y(n_14629)
);

NAND3xp33_ASAP7_75t_L g14630 ( 
.A(n_14458),
.B(n_2511),
.C(n_2512),
.Y(n_14630)
);

INVx1_ASAP7_75t_L g14631 ( 
.A(n_14477),
.Y(n_14631)
);

INVx1_ASAP7_75t_L g14632 ( 
.A(n_14478),
.Y(n_14632)
);

NOR2xp67_ASAP7_75t_L g14633 ( 
.A(n_14418),
.B(n_2513),
.Y(n_14633)
);

INVx1_ASAP7_75t_L g14634 ( 
.A(n_14364),
.Y(n_14634)
);

INVx2_ASAP7_75t_L g14635 ( 
.A(n_14417),
.Y(n_14635)
);

OR2x2_ASAP7_75t_L g14636 ( 
.A(n_14425),
.B(n_2513),
.Y(n_14636)
);

INVx1_ASAP7_75t_L g14637 ( 
.A(n_14422),
.Y(n_14637)
);

INVx1_ASAP7_75t_L g14638 ( 
.A(n_14413),
.Y(n_14638)
);

NOR2x1p5_ASAP7_75t_L g14639 ( 
.A(n_14457),
.B(n_2514),
.Y(n_14639)
);

AND2x2_ASAP7_75t_L g14640 ( 
.A(n_14464),
.B(n_2514),
.Y(n_14640)
);

NAND2x1p5_ASAP7_75t_L g14641 ( 
.A(n_14456),
.B(n_2515),
.Y(n_14641)
);

INVx1_ASAP7_75t_L g14642 ( 
.A(n_14445),
.Y(n_14642)
);

OAI21xp5_ASAP7_75t_L g14643 ( 
.A1(n_14447),
.A2(n_2515),
.B(n_2516),
.Y(n_14643)
);

AOI221xp5_ASAP7_75t_L g14644 ( 
.A1(n_14362),
.A2(n_2519),
.B1(n_2517),
.B2(n_2518),
.C(n_2520),
.Y(n_14644)
);

AND2x2_ASAP7_75t_L g14645 ( 
.A(n_14471),
.B(n_2517),
.Y(n_14645)
);

INVx2_ASAP7_75t_L g14646 ( 
.A(n_14380),
.Y(n_14646)
);

OR2x2_ASAP7_75t_L g14647 ( 
.A(n_14511),
.B(n_2518),
.Y(n_14647)
);

OAI21xp5_ASAP7_75t_SL g14648 ( 
.A1(n_14522),
.A2(n_2519),
.B(n_2520),
.Y(n_14648)
);

OAI31xp33_ASAP7_75t_L g14649 ( 
.A1(n_14504),
.A2(n_2523),
.A3(n_2521),
.B(n_2522),
.Y(n_14649)
);

INVx1_ASAP7_75t_L g14650 ( 
.A(n_14517),
.Y(n_14650)
);

NAND2xp5_ASAP7_75t_L g14651 ( 
.A(n_14508),
.B(n_2521),
.Y(n_14651)
);

OR2x2_ASAP7_75t_L g14652 ( 
.A(n_14554),
.B(n_2522),
.Y(n_14652)
);

AND2x2_ASAP7_75t_L g14653 ( 
.A(n_14503),
.B(n_2523),
.Y(n_14653)
);

NAND2xp5_ASAP7_75t_L g14654 ( 
.A(n_14645),
.B(n_2524),
.Y(n_14654)
);

AND2x4_ASAP7_75t_L g14655 ( 
.A(n_14646),
.B(n_2524),
.Y(n_14655)
);

AND2x2_ASAP7_75t_L g14656 ( 
.A(n_14507),
.B(n_2525),
.Y(n_14656)
);

NAND2xp5_ASAP7_75t_L g14657 ( 
.A(n_14512),
.B(n_2525),
.Y(n_14657)
);

A2O1A1Ixp33_ASAP7_75t_R g14658 ( 
.A1(n_14553),
.A2(n_2528),
.B(n_2526),
.C(n_2527),
.Y(n_14658)
);

AND2x2_ASAP7_75t_L g14659 ( 
.A(n_14518),
.B(n_14532),
.Y(n_14659)
);

NAND2xp5_ASAP7_75t_L g14660 ( 
.A(n_14519),
.B(n_2526),
.Y(n_14660)
);

INVx1_ASAP7_75t_L g14661 ( 
.A(n_14611),
.Y(n_14661)
);

OR2x6_ASAP7_75t_L g14662 ( 
.A(n_14510),
.B(n_2528),
.Y(n_14662)
);

NAND2xp5_ASAP7_75t_L g14663 ( 
.A(n_14546),
.B(n_2529),
.Y(n_14663)
);

OR2x2_ASAP7_75t_L g14664 ( 
.A(n_14505),
.B(n_2529),
.Y(n_14664)
);

CKINVDCx20_ASAP7_75t_R g14665 ( 
.A(n_14521),
.Y(n_14665)
);

INVx1_ASAP7_75t_L g14666 ( 
.A(n_14527),
.Y(n_14666)
);

AOI21xp5_ASAP7_75t_L g14667 ( 
.A1(n_14509),
.A2(n_2530),
.B(n_2531),
.Y(n_14667)
);

AO22x2_ASAP7_75t_L g14668 ( 
.A1(n_14557),
.A2(n_2532),
.B1(n_2530),
.B2(n_2531),
.Y(n_14668)
);

INVx2_ASAP7_75t_SL g14669 ( 
.A(n_14641),
.Y(n_14669)
);

AND2x2_ASAP7_75t_L g14670 ( 
.A(n_14513),
.B(n_2533),
.Y(n_14670)
);

INVx3_ASAP7_75t_L g14671 ( 
.A(n_14565),
.Y(n_14671)
);

INVx1_ASAP7_75t_L g14672 ( 
.A(n_14577),
.Y(n_14672)
);

INVx1_ASAP7_75t_L g14673 ( 
.A(n_14540),
.Y(n_14673)
);

NAND2xp5_ASAP7_75t_L g14674 ( 
.A(n_14539),
.B(n_2533),
.Y(n_14674)
);

NAND2xp5_ASAP7_75t_L g14675 ( 
.A(n_14547),
.B(n_2535),
.Y(n_14675)
);

INVx1_ASAP7_75t_L g14676 ( 
.A(n_14584),
.Y(n_14676)
);

OAI22xp5_ASAP7_75t_L g14677 ( 
.A1(n_14544),
.A2(n_2537),
.B1(n_2535),
.B2(n_2536),
.Y(n_14677)
);

INVx1_ASAP7_75t_L g14678 ( 
.A(n_14567),
.Y(n_14678)
);

OR2x2_ASAP7_75t_L g14679 ( 
.A(n_14506),
.B(n_2536),
.Y(n_14679)
);

OAI322xp33_ASAP7_75t_L g14680 ( 
.A1(n_14514),
.A2(n_2542),
.A3(n_2541),
.B1(n_2539),
.B2(n_2537),
.C1(n_2538),
.C2(n_2540),
.Y(n_14680)
);

NAND2xp5_ASAP7_75t_L g14681 ( 
.A(n_14617),
.B(n_2539),
.Y(n_14681)
);

NAND2x1_ASAP7_75t_L g14682 ( 
.A(n_14541),
.B(n_2540),
.Y(n_14682)
);

INVx1_ASAP7_75t_L g14683 ( 
.A(n_14571),
.Y(n_14683)
);

AOI31xp33_ASAP7_75t_L g14684 ( 
.A1(n_14524),
.A2(n_2543),
.A3(n_2541),
.B(n_2542),
.Y(n_14684)
);

NAND3xp33_ASAP7_75t_L g14685 ( 
.A(n_14619),
.B(n_2544),
.C(n_2545),
.Y(n_14685)
);

OAI22xp33_ASAP7_75t_L g14686 ( 
.A1(n_14599),
.A2(n_2546),
.B1(n_2544),
.B2(n_2545),
.Y(n_14686)
);

NOR2xp33_ASAP7_75t_L g14687 ( 
.A(n_14538),
.B(n_2547),
.Y(n_14687)
);

INVx1_ASAP7_75t_L g14688 ( 
.A(n_14607),
.Y(n_14688)
);

AND2x2_ASAP7_75t_L g14689 ( 
.A(n_14529),
.B(n_2547),
.Y(n_14689)
);

OR4x1_ASAP7_75t_L g14690 ( 
.A(n_14590),
.B(n_2550),
.C(n_2548),
.D(n_2549),
.Y(n_14690)
);

INVx2_ASAP7_75t_L g14691 ( 
.A(n_14607),
.Y(n_14691)
);

INVx2_ASAP7_75t_L g14692 ( 
.A(n_14523),
.Y(n_14692)
);

NAND2xp5_ASAP7_75t_L g14693 ( 
.A(n_14528),
.B(n_2548),
.Y(n_14693)
);

OR2x2_ASAP7_75t_L g14694 ( 
.A(n_14542),
.B(n_2550),
.Y(n_14694)
);

INVx1_ASAP7_75t_L g14695 ( 
.A(n_14586),
.Y(n_14695)
);

AOI22xp5_ASAP7_75t_L g14696 ( 
.A1(n_14585),
.A2(n_14516),
.B1(n_14526),
.B2(n_14533),
.Y(n_14696)
);

NOR2xp67_ASAP7_75t_SL g14697 ( 
.A(n_14561),
.B(n_2551),
.Y(n_14697)
);

INVx1_ASAP7_75t_L g14698 ( 
.A(n_14531),
.Y(n_14698)
);

INVx1_ASAP7_75t_L g14699 ( 
.A(n_14534),
.Y(n_14699)
);

NAND2xp67_ASAP7_75t_L g14700 ( 
.A(n_14574),
.B(n_2552),
.Y(n_14700)
);

OAI22xp5_ASAP7_75t_L g14701 ( 
.A1(n_14535),
.A2(n_14543),
.B1(n_14610),
.B2(n_14589),
.Y(n_14701)
);

INVx1_ASAP7_75t_L g14702 ( 
.A(n_14578),
.Y(n_14702)
);

INVxp67_ASAP7_75t_L g14703 ( 
.A(n_14515),
.Y(n_14703)
);

NOR2xp33_ASAP7_75t_L g14704 ( 
.A(n_14620),
.B(n_2553),
.Y(n_14704)
);

INVx2_ASAP7_75t_L g14705 ( 
.A(n_14639),
.Y(n_14705)
);

INVx2_ASAP7_75t_L g14706 ( 
.A(n_14591),
.Y(n_14706)
);

INVx1_ASAP7_75t_L g14707 ( 
.A(n_14603),
.Y(n_14707)
);

CKINVDCx16_ASAP7_75t_R g14708 ( 
.A(n_14568),
.Y(n_14708)
);

INVx1_ASAP7_75t_L g14709 ( 
.A(n_14552),
.Y(n_14709)
);

NAND2xp5_ASAP7_75t_L g14710 ( 
.A(n_14581),
.B(n_2554),
.Y(n_14710)
);

INVx1_ASAP7_75t_L g14711 ( 
.A(n_14530),
.Y(n_14711)
);

AND2x2_ASAP7_75t_L g14712 ( 
.A(n_14549),
.B(n_2554),
.Y(n_14712)
);

INVx1_ASAP7_75t_L g14713 ( 
.A(n_14602),
.Y(n_14713)
);

NAND2xp5_ASAP7_75t_L g14714 ( 
.A(n_14618),
.B(n_2555),
.Y(n_14714)
);

INVx1_ASAP7_75t_SL g14715 ( 
.A(n_14612),
.Y(n_14715)
);

NAND2xp5_ASAP7_75t_L g14716 ( 
.A(n_14633),
.B(n_2555),
.Y(n_14716)
);

INVx1_ASAP7_75t_L g14717 ( 
.A(n_14536),
.Y(n_14717)
);

AOI32xp33_ASAP7_75t_L g14718 ( 
.A1(n_14600),
.A2(n_2559),
.A3(n_2556),
.B1(n_2557),
.B2(n_2561),
.Y(n_14718)
);

NAND4xp25_ASAP7_75t_L g14719 ( 
.A(n_14545),
.B(n_2559),
.C(n_2556),
.D(n_2557),
.Y(n_14719)
);

INVx1_ASAP7_75t_L g14720 ( 
.A(n_14595),
.Y(n_14720)
);

AND2x2_ASAP7_75t_L g14721 ( 
.A(n_14550),
.B(n_2561),
.Y(n_14721)
);

NOR2xp33_ASAP7_75t_L g14722 ( 
.A(n_14551),
.B(n_2562),
.Y(n_14722)
);

NOR2xp33_ASAP7_75t_L g14723 ( 
.A(n_14570),
.B(n_2562),
.Y(n_14723)
);

AND2x2_ASAP7_75t_L g14724 ( 
.A(n_14572),
.B(n_2563),
.Y(n_14724)
);

OAI32xp33_ASAP7_75t_L g14725 ( 
.A1(n_14592),
.A2(n_2565),
.A3(n_2563),
.B1(n_2564),
.B2(n_2566),
.Y(n_14725)
);

BUFx2_ASAP7_75t_L g14726 ( 
.A(n_14643),
.Y(n_14726)
);

INVx1_ASAP7_75t_L g14727 ( 
.A(n_14609),
.Y(n_14727)
);

INVx2_ASAP7_75t_L g14728 ( 
.A(n_14594),
.Y(n_14728)
);

INVx2_ASAP7_75t_L g14729 ( 
.A(n_14596),
.Y(n_14729)
);

INVx1_ASAP7_75t_L g14730 ( 
.A(n_14562),
.Y(n_14730)
);

HB1xp67_ASAP7_75t_L g14731 ( 
.A(n_14640),
.Y(n_14731)
);

INVx1_ASAP7_75t_L g14732 ( 
.A(n_14576),
.Y(n_14732)
);

INVx1_ASAP7_75t_L g14733 ( 
.A(n_14580),
.Y(n_14733)
);

OAI22xp5_ASAP7_75t_L g14734 ( 
.A1(n_14573),
.A2(n_2568),
.B1(n_2566),
.B2(n_2567),
.Y(n_14734)
);

INVx1_ASAP7_75t_L g14735 ( 
.A(n_14560),
.Y(n_14735)
);

NAND2xp5_ASAP7_75t_L g14736 ( 
.A(n_14579),
.B(n_2567),
.Y(n_14736)
);

AND2x2_ASAP7_75t_L g14737 ( 
.A(n_14537),
.B(n_2569),
.Y(n_14737)
);

AND2x2_ASAP7_75t_L g14738 ( 
.A(n_14548),
.B(n_2569),
.Y(n_14738)
);

OAI31xp33_ASAP7_75t_L g14739 ( 
.A1(n_14593),
.A2(n_2572),
.A3(n_2570),
.B(n_2571),
.Y(n_14739)
);

AND2x2_ASAP7_75t_L g14740 ( 
.A(n_14558),
.B(n_2570),
.Y(n_14740)
);

INVx1_ASAP7_75t_SL g14741 ( 
.A(n_14613),
.Y(n_14741)
);

INVxp67_ASAP7_75t_SL g14742 ( 
.A(n_14583),
.Y(n_14742)
);

OAI32xp33_ASAP7_75t_L g14743 ( 
.A1(n_14597),
.A2(n_2573),
.A3(n_2571),
.B1(n_2572),
.B2(n_2574),
.Y(n_14743)
);

AOI21x1_ASAP7_75t_L g14744 ( 
.A1(n_14525),
.A2(n_2573),
.B(n_2574),
.Y(n_14744)
);

NAND2xp33_ASAP7_75t_SL g14745 ( 
.A(n_14566),
.B(n_2575),
.Y(n_14745)
);

OAI21xp5_ASAP7_75t_L g14746 ( 
.A1(n_14559),
.A2(n_2575),
.B(n_2576),
.Y(n_14746)
);

INVx2_ASAP7_75t_L g14747 ( 
.A(n_14627),
.Y(n_14747)
);

INVx1_ASAP7_75t_L g14748 ( 
.A(n_14601),
.Y(n_14748)
);

INVx1_ASAP7_75t_L g14749 ( 
.A(n_14616),
.Y(n_14749)
);

OR2x2_ASAP7_75t_L g14750 ( 
.A(n_14604),
.B(n_2576),
.Y(n_14750)
);

INVx1_ASAP7_75t_SL g14751 ( 
.A(n_14555),
.Y(n_14751)
);

INVx1_ASAP7_75t_L g14752 ( 
.A(n_14625),
.Y(n_14752)
);

OAI21xp5_ASAP7_75t_L g14753 ( 
.A1(n_14606),
.A2(n_14608),
.B(n_14622),
.Y(n_14753)
);

NAND2xp5_ASAP7_75t_L g14754 ( 
.A(n_14623),
.B(n_2577),
.Y(n_14754)
);

NAND2x1p5_ASAP7_75t_L g14755 ( 
.A(n_14564),
.B(n_2578),
.Y(n_14755)
);

AND2x4_ASAP7_75t_L g14756 ( 
.A(n_14582),
.B(n_2580),
.Y(n_14756)
);

AOI22xp33_ASAP7_75t_L g14757 ( 
.A1(n_14621),
.A2(n_2582),
.B1(n_2580),
.B2(n_2581),
.Y(n_14757)
);

OAI221xp5_ASAP7_75t_L g14758 ( 
.A1(n_14598),
.A2(n_2583),
.B1(n_2581),
.B2(n_2582),
.C(n_2584),
.Y(n_14758)
);

AND2x2_ASAP7_75t_L g14759 ( 
.A(n_14624),
.B(n_2583),
.Y(n_14759)
);

AOI21xp5_ASAP7_75t_L g14760 ( 
.A1(n_14615),
.A2(n_2584),
.B(n_2585),
.Y(n_14760)
);

INVx1_ASAP7_75t_L g14761 ( 
.A(n_14556),
.Y(n_14761)
);

AOI22xp5_ASAP7_75t_L g14762 ( 
.A1(n_14626),
.A2(n_2587),
.B1(n_2585),
.B2(n_2586),
.Y(n_14762)
);

INVx1_ASAP7_75t_L g14763 ( 
.A(n_14636),
.Y(n_14763)
);

INVx1_ASAP7_75t_L g14764 ( 
.A(n_14630),
.Y(n_14764)
);

INVx1_ASAP7_75t_L g14765 ( 
.A(n_14563),
.Y(n_14765)
);

INVx1_ASAP7_75t_L g14766 ( 
.A(n_14520),
.Y(n_14766)
);

INVx1_ASAP7_75t_L g14767 ( 
.A(n_14628),
.Y(n_14767)
);

INVx1_ASAP7_75t_SL g14768 ( 
.A(n_14635),
.Y(n_14768)
);

INVx1_ASAP7_75t_L g14769 ( 
.A(n_14575),
.Y(n_14769)
);

NAND2xp5_ASAP7_75t_L g14770 ( 
.A(n_14569),
.B(n_14614),
.Y(n_14770)
);

INVx1_ASAP7_75t_L g14771 ( 
.A(n_14587),
.Y(n_14771)
);

AOI22xp5_ASAP7_75t_L g14772 ( 
.A1(n_14605),
.A2(n_2588),
.B1(n_2586),
.B2(n_2587),
.Y(n_14772)
);

INVx1_ASAP7_75t_L g14773 ( 
.A(n_14629),
.Y(n_14773)
);

OAI21xp5_ASAP7_75t_L g14774 ( 
.A1(n_14642),
.A2(n_2588),
.B(n_2589),
.Y(n_14774)
);

INVx1_ASAP7_75t_L g14775 ( 
.A(n_14631),
.Y(n_14775)
);

INVx1_ASAP7_75t_L g14776 ( 
.A(n_14632),
.Y(n_14776)
);

OAI21xp33_ASAP7_75t_L g14777 ( 
.A1(n_14588),
.A2(n_2589),
.B(n_2590),
.Y(n_14777)
);

OR2x2_ASAP7_75t_L g14778 ( 
.A(n_14634),
.B(n_2590),
.Y(n_14778)
);

INVx1_ASAP7_75t_L g14779 ( 
.A(n_14637),
.Y(n_14779)
);

NAND2xp33_ASAP7_75t_SL g14780 ( 
.A(n_14638),
.B(n_2592),
.Y(n_14780)
);

AOI22xp5_ASAP7_75t_L g14781 ( 
.A1(n_14644),
.A2(n_2595),
.B1(n_2593),
.B2(n_2594),
.Y(n_14781)
);

AND2x2_ASAP7_75t_L g14782 ( 
.A(n_14503),
.B(n_2593),
.Y(n_14782)
);

NAND2xp5_ASAP7_75t_L g14783 ( 
.A(n_14653),
.B(n_2594),
.Y(n_14783)
);

AND2x2_ASAP7_75t_L g14784 ( 
.A(n_14782),
.B(n_2596),
.Y(n_14784)
);

INVx1_ASAP7_75t_SL g14785 ( 
.A(n_14652),
.Y(n_14785)
);

INVx1_ASAP7_75t_L g14786 ( 
.A(n_14668),
.Y(n_14786)
);

NAND2x1_ASAP7_75t_L g14787 ( 
.A(n_14661),
.B(n_2596),
.Y(n_14787)
);

NOR2xp33_ASAP7_75t_L g14788 ( 
.A(n_14684),
.B(n_2597),
.Y(n_14788)
);

INVx1_ASAP7_75t_L g14789 ( 
.A(n_14668),
.Y(n_14789)
);

INVx1_ASAP7_75t_L g14790 ( 
.A(n_14700),
.Y(n_14790)
);

INVx1_ASAP7_75t_L g14791 ( 
.A(n_14647),
.Y(n_14791)
);

OAI32xp33_ASAP7_75t_L g14792 ( 
.A1(n_14708),
.A2(n_2600),
.A3(n_2598),
.B1(n_2599),
.B2(n_2601),
.Y(n_14792)
);

NAND2xp33_ASAP7_75t_L g14793 ( 
.A(n_14650),
.B(n_2598),
.Y(n_14793)
);

INVx2_ASAP7_75t_L g14794 ( 
.A(n_14755),
.Y(n_14794)
);

AOI22xp33_ASAP7_75t_L g14795 ( 
.A1(n_14666),
.A2(n_2601),
.B1(n_2599),
.B2(n_2600),
.Y(n_14795)
);

INVx1_ASAP7_75t_L g14796 ( 
.A(n_14679),
.Y(n_14796)
);

A2O1A1Ixp33_ASAP7_75t_L g14797 ( 
.A1(n_14718),
.A2(n_2604),
.B(n_2602),
.C(n_2603),
.Y(n_14797)
);

INVx2_ASAP7_75t_L g14798 ( 
.A(n_14662),
.Y(n_14798)
);

INVx1_ASAP7_75t_L g14799 ( 
.A(n_14656),
.Y(n_14799)
);

AOI22xp5_ASAP7_75t_L g14800 ( 
.A1(n_14665),
.A2(n_2605),
.B1(n_2602),
.B2(n_2603),
.Y(n_14800)
);

OAI221xp5_ASAP7_75t_L g14801 ( 
.A1(n_14696),
.A2(n_2607),
.B1(n_2605),
.B2(n_2606),
.C(n_2608),
.Y(n_14801)
);

INVx1_ASAP7_75t_L g14802 ( 
.A(n_14664),
.Y(n_14802)
);

AOI22xp33_ASAP7_75t_L g14803 ( 
.A1(n_14672),
.A2(n_2608),
.B1(n_2606),
.B2(n_2607),
.Y(n_14803)
);

OR2x2_ASAP7_75t_L g14804 ( 
.A(n_14669),
.B(n_14662),
.Y(n_14804)
);

NOR2xp33_ASAP7_75t_L g14805 ( 
.A(n_14719),
.B(n_2609),
.Y(n_14805)
);

INVxp67_ASAP7_75t_L g14806 ( 
.A(n_14697),
.Y(n_14806)
);

AO221x1_ASAP7_75t_L g14807 ( 
.A1(n_14701),
.A2(n_2611),
.B1(n_2609),
.B2(n_2610),
.C(n_2612),
.Y(n_14807)
);

OAI22xp5_ASAP7_75t_L g14808 ( 
.A1(n_14751),
.A2(n_2612),
.B1(n_2610),
.B2(n_2611),
.Y(n_14808)
);

AOI22xp33_ASAP7_75t_L g14809 ( 
.A1(n_14692),
.A2(n_2615),
.B1(n_2613),
.B2(n_2614),
.Y(n_14809)
);

INVx1_ASAP7_75t_L g14810 ( 
.A(n_14694),
.Y(n_14810)
);

AOI322xp5_ASAP7_75t_L g14811 ( 
.A1(n_14768),
.A2(n_2618),
.A3(n_2617),
.B1(n_2615),
.B2(n_2613),
.C1(n_2614),
.C2(n_2616),
.Y(n_14811)
);

INVx2_ASAP7_75t_L g14812 ( 
.A(n_14690),
.Y(n_14812)
);

BUFx2_ASAP7_75t_L g14813 ( 
.A(n_14745),
.Y(n_14813)
);

NAND2xp5_ASAP7_75t_L g14814 ( 
.A(n_14655),
.B(n_2617),
.Y(n_14814)
);

OR2x2_ASAP7_75t_L g14815 ( 
.A(n_14682),
.B(n_14691),
.Y(n_14815)
);

AND2x2_ASAP7_75t_L g14816 ( 
.A(n_14659),
.B(n_2619),
.Y(n_14816)
);

OR2x2_ASAP7_75t_L g14817 ( 
.A(n_14663),
.B(n_2619),
.Y(n_14817)
);

INVx2_ASAP7_75t_L g14818 ( 
.A(n_14756),
.Y(n_14818)
);

NAND2xp5_ASAP7_75t_L g14819 ( 
.A(n_14712),
.B(n_2620),
.Y(n_14819)
);

INVx1_ASAP7_75t_L g14820 ( 
.A(n_14721),
.Y(n_14820)
);

OAI22xp5_ASAP7_75t_L g14821 ( 
.A1(n_14781),
.A2(n_2622),
.B1(n_2620),
.B2(n_2621),
.Y(n_14821)
);

NAND2xp5_ASAP7_75t_L g14822 ( 
.A(n_14724),
.B(n_2621),
.Y(n_14822)
);

AND2x2_ASAP7_75t_L g14823 ( 
.A(n_14671),
.B(n_2622),
.Y(n_14823)
);

INVx1_ASAP7_75t_L g14824 ( 
.A(n_14738),
.Y(n_14824)
);

NAND2x2_ASAP7_75t_L g14825 ( 
.A(n_14744),
.B(n_2623),
.Y(n_14825)
);

INVx1_ASAP7_75t_SL g14826 ( 
.A(n_14780),
.Y(n_14826)
);

AOI33xp33_ASAP7_75t_L g14827 ( 
.A1(n_14713),
.A2(n_2625),
.A3(n_2627),
.B1(n_2623),
.B2(n_2624),
.B3(n_2626),
.Y(n_14827)
);

INVx1_ASAP7_75t_SL g14828 ( 
.A(n_14737),
.Y(n_14828)
);

AOI22xp5_ASAP7_75t_L g14829 ( 
.A1(n_14741),
.A2(n_2627),
.B1(n_2624),
.B2(n_2625),
.Y(n_14829)
);

OAI21xp5_ASAP7_75t_L g14830 ( 
.A1(n_14685),
.A2(n_2628),
.B(n_2629),
.Y(n_14830)
);

INVx1_ASAP7_75t_L g14831 ( 
.A(n_14670),
.Y(n_14831)
);

INVx2_ASAP7_75t_L g14832 ( 
.A(n_14778),
.Y(n_14832)
);

INVx1_ASAP7_75t_L g14833 ( 
.A(n_14689),
.Y(n_14833)
);

HB1xp67_ASAP7_75t_L g14834 ( 
.A(n_14688),
.Y(n_14834)
);

INVx1_ASAP7_75t_L g14835 ( 
.A(n_14710),
.Y(n_14835)
);

INVxp67_ASAP7_75t_L g14836 ( 
.A(n_14687),
.Y(n_14836)
);

NAND3x2_ASAP7_75t_L g14837 ( 
.A(n_14726),
.B(n_2628),
.C(n_2629),
.Y(n_14837)
);

HB1xp67_ASAP7_75t_L g14838 ( 
.A(n_14716),
.Y(n_14838)
);

AND2x2_ASAP7_75t_L g14839 ( 
.A(n_14673),
.B(n_2630),
.Y(n_14839)
);

INVx2_ASAP7_75t_L g14840 ( 
.A(n_14759),
.Y(n_14840)
);

AND2x2_ASAP7_75t_L g14841 ( 
.A(n_14720),
.B(n_2630),
.Y(n_14841)
);

HB1xp67_ASAP7_75t_L g14842 ( 
.A(n_14731),
.Y(n_14842)
);

INVx1_ASAP7_75t_L g14843 ( 
.A(n_14714),
.Y(n_14843)
);

OR2x2_ASAP7_75t_L g14844 ( 
.A(n_14674),
.B(n_2631),
.Y(n_14844)
);

AOI22xp5_ASAP7_75t_L g14845 ( 
.A1(n_14715),
.A2(n_2633),
.B1(n_2631),
.B2(n_2632),
.Y(n_14845)
);

INVx1_ASAP7_75t_SL g14846 ( 
.A(n_14740),
.Y(n_14846)
);

OAI21xp33_ASAP7_75t_L g14847 ( 
.A1(n_14770),
.A2(n_2632),
.B(n_2633),
.Y(n_14847)
);

OR2x2_ASAP7_75t_L g14848 ( 
.A(n_14651),
.B(n_2634),
.Y(n_14848)
);

AND2x2_ASAP7_75t_L g14849 ( 
.A(n_14676),
.B(n_14695),
.Y(n_14849)
);

INVxp67_ASAP7_75t_L g14850 ( 
.A(n_14722),
.Y(n_14850)
);

INVx2_ASAP7_75t_L g14851 ( 
.A(n_14750),
.Y(n_14851)
);

NAND2xp5_ASAP7_75t_L g14852 ( 
.A(n_14723),
.B(n_2635),
.Y(n_14852)
);

NAND2xp5_ASAP7_75t_L g14853 ( 
.A(n_14649),
.B(n_2636),
.Y(n_14853)
);

INVx4_ASAP7_75t_L g14854 ( 
.A(n_14706),
.Y(n_14854)
);

INVx2_ASAP7_75t_L g14855 ( 
.A(n_14705),
.Y(n_14855)
);

INVx1_ASAP7_75t_L g14856 ( 
.A(n_14657),
.Y(n_14856)
);

INVx1_ASAP7_75t_L g14857 ( 
.A(n_14660),
.Y(n_14857)
);

OAI211xp5_ASAP7_75t_L g14858 ( 
.A1(n_14753),
.A2(n_2638),
.B(n_2636),
.C(n_2637),
.Y(n_14858)
);

NAND2xp5_ASAP7_75t_L g14859 ( 
.A(n_14686),
.B(n_2637),
.Y(n_14859)
);

OR2x2_ASAP7_75t_L g14860 ( 
.A(n_14693),
.B(n_2639),
.Y(n_14860)
);

INVxp33_ASAP7_75t_L g14861 ( 
.A(n_14704),
.Y(n_14861)
);

INVx2_ASAP7_75t_L g14862 ( 
.A(n_14702),
.Y(n_14862)
);

INVx1_ASAP7_75t_L g14863 ( 
.A(n_14654),
.Y(n_14863)
);

AOI211xp5_ASAP7_75t_L g14864 ( 
.A1(n_14648),
.A2(n_2641),
.B(n_2639),
.C(n_2640),
.Y(n_14864)
);

OAI32xp33_ASAP7_75t_L g14865 ( 
.A1(n_14736),
.A2(n_2642),
.A3(n_2640),
.B1(n_2641),
.B2(n_2643),
.Y(n_14865)
);

AOI21xp33_ASAP7_75t_SL g14866 ( 
.A1(n_14677),
.A2(n_2642),
.B(n_2643),
.Y(n_14866)
);

OAI22xp5_ASAP7_75t_L g14867 ( 
.A1(n_14764),
.A2(n_14758),
.B1(n_14766),
.B2(n_14707),
.Y(n_14867)
);

AOI21xp33_ASAP7_75t_L g14868 ( 
.A1(n_14658),
.A2(n_2644),
.B(n_2645),
.Y(n_14868)
);

OAI32xp33_ASAP7_75t_L g14869 ( 
.A1(n_14767),
.A2(n_2646),
.A3(n_2644),
.B1(n_2645),
.B2(n_2647),
.Y(n_14869)
);

AOI22xp5_ASAP7_75t_L g14870 ( 
.A1(n_14765),
.A2(n_2648),
.B1(n_2646),
.B2(n_2647),
.Y(n_14870)
);

INVx1_ASAP7_75t_L g14871 ( 
.A(n_14675),
.Y(n_14871)
);

AO22x1_ASAP7_75t_L g14872 ( 
.A1(n_14742),
.A2(n_2650),
.B1(n_2648),
.B2(n_2649),
.Y(n_14872)
);

INVx2_ASAP7_75t_SL g14873 ( 
.A(n_14678),
.Y(n_14873)
);

INVx1_ASAP7_75t_L g14874 ( 
.A(n_14754),
.Y(n_14874)
);

O2A1O1Ixp33_ASAP7_75t_L g14875 ( 
.A1(n_14725),
.A2(n_2653),
.B(n_2651),
.C(n_2652),
.Y(n_14875)
);

INVx1_ASAP7_75t_L g14876 ( 
.A(n_14681),
.Y(n_14876)
);

OR2x2_ASAP7_75t_L g14877 ( 
.A(n_14699),
.B(n_2651),
.Y(n_14877)
);

OAI33xp33_ASAP7_75t_L g14878 ( 
.A1(n_14769),
.A2(n_2655),
.A3(n_2657),
.B1(n_2653),
.B2(n_2654),
.B3(n_2656),
.Y(n_14878)
);

INVx2_ASAP7_75t_L g14879 ( 
.A(n_14749),
.Y(n_14879)
);

AND2x4_ASAP7_75t_L g14880 ( 
.A(n_14727),
.B(n_2655),
.Y(n_14880)
);

INVx1_ASAP7_75t_L g14881 ( 
.A(n_14709),
.Y(n_14881)
);

NAND2xp5_ASAP7_75t_L g14882 ( 
.A(n_14739),
.B(n_2656),
.Y(n_14882)
);

AOI22xp5_ASAP7_75t_L g14883 ( 
.A1(n_14752),
.A2(n_2660),
.B1(n_2658),
.B2(n_2659),
.Y(n_14883)
);

AND2x2_ASAP7_75t_L g14884 ( 
.A(n_14683),
.B(n_14698),
.Y(n_14884)
);

INVx2_ASAP7_75t_L g14885 ( 
.A(n_14728),
.Y(n_14885)
);

OAI222xp33_ASAP7_75t_L g14886 ( 
.A1(n_14703),
.A2(n_2662),
.B1(n_2664),
.B2(n_2659),
.C1(n_2661),
.C2(n_2663),
.Y(n_14886)
);

OAI22xp33_ASAP7_75t_SL g14887 ( 
.A1(n_14771),
.A2(n_2664),
.B1(n_2661),
.B2(n_2662),
.Y(n_14887)
);

OAI22xp33_ASAP7_75t_L g14888 ( 
.A1(n_14773),
.A2(n_2667),
.B1(n_2665),
.B2(n_2666),
.Y(n_14888)
);

INVxp67_ASAP7_75t_L g14889 ( 
.A(n_14734),
.Y(n_14889)
);

NOR2xp33_ASAP7_75t_SL g14890 ( 
.A(n_14680),
.B(n_14777),
.Y(n_14890)
);

INVx1_ASAP7_75t_L g14891 ( 
.A(n_14774),
.Y(n_14891)
);

INVx1_ASAP7_75t_L g14892 ( 
.A(n_14746),
.Y(n_14892)
);

INVx2_ASAP7_75t_L g14893 ( 
.A(n_14729),
.Y(n_14893)
);

INVx2_ASAP7_75t_SL g14894 ( 
.A(n_14747),
.Y(n_14894)
);

NOR2xp33_ASAP7_75t_SL g14895 ( 
.A(n_14763),
.B(n_14761),
.Y(n_14895)
);

NAND2xp5_ASAP7_75t_L g14896 ( 
.A(n_14667),
.B(n_2666),
.Y(n_14896)
);

INVx1_ASAP7_75t_L g14897 ( 
.A(n_14762),
.Y(n_14897)
);

NAND2xp33_ASAP7_75t_SL g14898 ( 
.A(n_14775),
.B(n_14776),
.Y(n_14898)
);

OAI32xp33_ASAP7_75t_L g14899 ( 
.A1(n_14779),
.A2(n_2669),
.A3(n_2667),
.B1(n_2668),
.B2(n_2670),
.Y(n_14899)
);

INVx1_ASAP7_75t_L g14900 ( 
.A(n_14772),
.Y(n_14900)
);

AOI31xp33_ASAP7_75t_L g14901 ( 
.A1(n_14760),
.A2(n_2672),
.A3(n_2670),
.B(n_2671),
.Y(n_14901)
);

OAI32xp33_ASAP7_75t_L g14902 ( 
.A1(n_14735),
.A2(n_2674),
.A3(n_2671),
.B1(n_2673),
.B2(n_2675),
.Y(n_14902)
);

OAI22xp5_ASAP7_75t_L g14903 ( 
.A1(n_14711),
.A2(n_2676),
.B1(n_2674),
.B2(n_2675),
.Y(n_14903)
);

INVx1_ASAP7_75t_L g14904 ( 
.A(n_14717),
.Y(n_14904)
);

OAI322xp33_ASAP7_75t_L g14905 ( 
.A1(n_14748),
.A2(n_14732),
.A3(n_14733),
.B1(n_14730),
.B2(n_14743),
.C1(n_14757),
.C2(n_2678),
.Y(n_14905)
);

INVx1_ASAP7_75t_L g14906 ( 
.A(n_14668),
.Y(n_14906)
);

NAND4xp25_ASAP7_75t_L g14907 ( 
.A(n_14696),
.B(n_2679),
.C(n_2676),
.D(n_2677),
.Y(n_14907)
);

OR2x2_ASAP7_75t_L g14908 ( 
.A(n_14652),
.B(n_2677),
.Y(n_14908)
);

AOI22xp5_ASAP7_75t_L g14909 ( 
.A1(n_14895),
.A2(n_2681),
.B1(n_2679),
.B2(n_2680),
.Y(n_14909)
);

OR2x2_ASAP7_75t_L g14910 ( 
.A(n_14787),
.B(n_2680),
.Y(n_14910)
);

AOI322xp5_ASAP7_75t_L g14911 ( 
.A1(n_14826),
.A2(n_2688),
.A3(n_2687),
.B1(n_2685),
.B2(n_2681),
.C1(n_2682),
.C2(n_2686),
.Y(n_14911)
);

OAI321xp33_ASAP7_75t_L g14912 ( 
.A1(n_14806),
.A2(n_2687),
.A3(n_2689),
.B1(n_2682),
.B2(n_2685),
.C(n_2688),
.Y(n_14912)
);

OAI22xp33_ASAP7_75t_L g14913 ( 
.A1(n_14825),
.A2(n_14890),
.B1(n_14901),
.B2(n_14804),
.Y(n_14913)
);

INVx1_ASAP7_75t_L g14914 ( 
.A(n_14786),
.Y(n_14914)
);

AOI221xp5_ASAP7_75t_L g14915 ( 
.A1(n_14868),
.A2(n_2691),
.B1(n_2689),
.B2(n_2690),
.C(n_2692),
.Y(n_14915)
);

OAI221xp5_ASAP7_75t_L g14916 ( 
.A1(n_14898),
.A2(n_2693),
.B1(n_2690),
.B2(n_2692),
.C(n_2694),
.Y(n_14916)
);

OAI21xp33_ASAP7_75t_L g14917 ( 
.A1(n_14861),
.A2(n_2693),
.B(n_2694),
.Y(n_14917)
);

OAI322xp33_ASAP7_75t_L g14918 ( 
.A1(n_14789),
.A2(n_2700),
.A3(n_2699),
.B1(n_2697),
.B2(n_2695),
.C1(n_2696),
.C2(n_2698),
.Y(n_14918)
);

OAI22xp33_ASAP7_75t_SL g14919 ( 
.A1(n_14906),
.A2(n_2699),
.B1(n_2697),
.B2(n_2698),
.Y(n_14919)
);

OAI21xp5_ASAP7_75t_L g14920 ( 
.A1(n_14797),
.A2(n_2700),
.B(n_2701),
.Y(n_14920)
);

OAI21xp5_ASAP7_75t_L g14921 ( 
.A1(n_14834),
.A2(n_2701),
.B(n_2702),
.Y(n_14921)
);

HB1xp67_ASAP7_75t_L g14922 ( 
.A(n_14872),
.Y(n_14922)
);

INVx1_ASAP7_75t_L g14923 ( 
.A(n_14816),
.Y(n_14923)
);

NAND2xp33_ASAP7_75t_L g14924 ( 
.A(n_14842),
.B(n_2702),
.Y(n_14924)
);

OAI33xp33_ASAP7_75t_L g14925 ( 
.A1(n_14867),
.A2(n_2705),
.A3(n_2707),
.B1(n_2703),
.B2(n_2704),
.B3(n_2706),
.Y(n_14925)
);

AOI221xp5_ASAP7_75t_L g14926 ( 
.A1(n_14905),
.A2(n_2705),
.B1(n_2703),
.B2(n_2704),
.C(n_2706),
.Y(n_14926)
);

NAND3xp33_ASAP7_75t_SL g14927 ( 
.A(n_14785),
.B(n_2707),
.C(n_2708),
.Y(n_14927)
);

AOI22xp5_ASAP7_75t_L g14928 ( 
.A1(n_14873),
.A2(n_2710),
.B1(n_2708),
.B2(n_2709),
.Y(n_14928)
);

OAI22xp5_ASAP7_75t_L g14929 ( 
.A1(n_14837),
.A2(n_2711),
.B1(n_2709),
.B2(n_2710),
.Y(n_14929)
);

INVx1_ASAP7_75t_L g14930 ( 
.A(n_14839),
.Y(n_14930)
);

AOI22xp5_ASAP7_75t_L g14931 ( 
.A1(n_14894),
.A2(n_2713),
.B1(n_2711),
.B2(n_2712),
.Y(n_14931)
);

INVx1_ASAP7_75t_L g14932 ( 
.A(n_14841),
.Y(n_14932)
);

AOI32xp33_ASAP7_75t_L g14933 ( 
.A1(n_14813),
.A2(n_2714),
.A3(n_2712),
.B1(n_2713),
.B2(n_2715),
.Y(n_14933)
);

NOR2xp33_ASAP7_75t_L g14934 ( 
.A(n_14907),
.B(n_2714),
.Y(n_14934)
);

OAI22xp5_ASAP7_75t_L g14935 ( 
.A1(n_14889),
.A2(n_14815),
.B1(n_14855),
.B2(n_14798),
.Y(n_14935)
);

OAI22xp5_ASAP7_75t_L g14936 ( 
.A1(n_14812),
.A2(n_2718),
.B1(n_2716),
.B2(n_2717),
.Y(n_14936)
);

AOI21xp5_ASAP7_75t_L g14937 ( 
.A1(n_14793),
.A2(n_2716),
.B(n_2717),
.Y(n_14937)
);

AOI211x1_ASAP7_75t_L g14938 ( 
.A1(n_14830),
.A2(n_2720),
.B(n_2718),
.C(n_2719),
.Y(n_14938)
);

AOI22xp5_ASAP7_75t_L g14939 ( 
.A1(n_14805),
.A2(n_2722),
.B1(n_2719),
.B2(n_2721),
.Y(n_14939)
);

OAI22xp5_ASAP7_75t_L g14940 ( 
.A1(n_14862),
.A2(n_2723),
.B1(n_2721),
.B2(n_2722),
.Y(n_14940)
);

OAI22xp5_ASAP7_75t_L g14941 ( 
.A1(n_14879),
.A2(n_2726),
.B1(n_2724),
.B2(n_2725),
.Y(n_14941)
);

NAND3xp33_ASAP7_75t_L g14942 ( 
.A(n_14864),
.B(n_2724),
.C(n_2725),
.Y(n_14942)
);

INVx1_ASAP7_75t_L g14943 ( 
.A(n_14784),
.Y(n_14943)
);

OAI221xp5_ASAP7_75t_L g14944 ( 
.A1(n_14788),
.A2(n_2728),
.B1(n_2726),
.B2(n_2727),
.C(n_2729),
.Y(n_14944)
);

OAI22xp5_ASAP7_75t_L g14945 ( 
.A1(n_14881),
.A2(n_2729),
.B1(n_2727),
.B2(n_2728),
.Y(n_14945)
);

AOI221xp5_ASAP7_75t_L g14946 ( 
.A1(n_14866),
.A2(n_2732),
.B1(n_2730),
.B2(n_2731),
.C(n_2733),
.Y(n_14946)
);

INVx1_ASAP7_75t_L g14947 ( 
.A(n_14823),
.Y(n_14947)
);

INVx1_ASAP7_75t_L g14948 ( 
.A(n_14880),
.Y(n_14948)
);

AOI22xp5_ASAP7_75t_L g14949 ( 
.A1(n_14849),
.A2(n_2732),
.B1(n_2730),
.B2(n_2731),
.Y(n_14949)
);

OAI22xp33_ASAP7_75t_SL g14950 ( 
.A1(n_14790),
.A2(n_2736),
.B1(n_2734),
.B2(n_2735),
.Y(n_14950)
);

AND2x2_ASAP7_75t_L g14951 ( 
.A(n_14884),
.B(n_2735),
.Y(n_14951)
);

INVx1_ASAP7_75t_L g14952 ( 
.A(n_14880),
.Y(n_14952)
);

AOI222xp33_ASAP7_75t_SL g14953 ( 
.A1(n_14828),
.A2(n_2738),
.B1(n_2740),
.B2(n_2736),
.C1(n_2737),
.C2(n_2739),
.Y(n_14953)
);

NAND2xp5_ASAP7_75t_SL g14954 ( 
.A(n_14887),
.B(n_2737),
.Y(n_14954)
);

NOR2x1_ASAP7_75t_L g14955 ( 
.A(n_14854),
.B(n_2738),
.Y(n_14955)
);

AOI222xp33_ASAP7_75t_L g14956 ( 
.A1(n_14900),
.A2(n_2741),
.B1(n_2743),
.B2(n_2739),
.C1(n_2740),
.C2(n_2742),
.Y(n_14956)
);

NOR4xp25_ASAP7_75t_L g14957 ( 
.A(n_14875),
.B(n_2744),
.C(n_2741),
.D(n_2743),
.Y(n_14957)
);

OAI21xp5_ASAP7_75t_L g14958 ( 
.A1(n_14853),
.A2(n_14882),
.B(n_14850),
.Y(n_14958)
);

INVx2_ASAP7_75t_L g14959 ( 
.A(n_14908),
.Y(n_14959)
);

NOR3xp33_ASAP7_75t_L g14960 ( 
.A(n_14854),
.B(n_2744),
.C(n_2745),
.Y(n_14960)
);

AOI21xp5_ASAP7_75t_L g14961 ( 
.A1(n_14896),
.A2(n_2745),
.B(n_2746),
.Y(n_14961)
);

AOI222xp33_ASAP7_75t_L g14962 ( 
.A1(n_14846),
.A2(n_14891),
.B1(n_14892),
.B2(n_14897),
.C1(n_14799),
.C2(n_14904),
.Y(n_14962)
);

OAI22xp5_ASAP7_75t_L g14963 ( 
.A1(n_14885),
.A2(n_2749),
.B1(n_2747),
.B2(n_2748),
.Y(n_14963)
);

AND2x2_ASAP7_75t_L g14964 ( 
.A(n_14840),
.B(n_2747),
.Y(n_14964)
);

AND2x4_ASAP7_75t_L g14965 ( 
.A(n_14794),
.B(n_2749),
.Y(n_14965)
);

AOI31xp33_ASAP7_75t_L g14966 ( 
.A1(n_14802),
.A2(n_2752),
.A3(n_2750),
.B(n_2751),
.Y(n_14966)
);

HB1xp67_ASAP7_75t_L g14967 ( 
.A(n_14877),
.Y(n_14967)
);

INVx1_ASAP7_75t_L g14968 ( 
.A(n_14807),
.Y(n_14968)
);

NAND2xp5_ASAP7_75t_L g14969 ( 
.A(n_14827),
.B(n_14888),
.Y(n_14969)
);

AOI22xp5_ASAP7_75t_L g14970 ( 
.A1(n_14893),
.A2(n_2752),
.B1(n_2750),
.B2(n_2751),
.Y(n_14970)
);

NAND2xp5_ASAP7_75t_L g14971 ( 
.A(n_14845),
.B(n_2753),
.Y(n_14971)
);

AOI21xp5_ASAP7_75t_L g14972 ( 
.A1(n_14783),
.A2(n_2753),
.B(n_2754),
.Y(n_14972)
);

AOI21xp33_ASAP7_75t_L g14973 ( 
.A1(n_14860),
.A2(n_2755),
.B(n_2756),
.Y(n_14973)
);

INVx2_ASAP7_75t_L g14974 ( 
.A(n_14844),
.Y(n_14974)
);

NOR3xp33_ASAP7_75t_L g14975 ( 
.A(n_14791),
.B(n_2755),
.C(n_2757),
.Y(n_14975)
);

AOI221xp5_ASAP7_75t_L g14976 ( 
.A1(n_14820),
.A2(n_2759),
.B1(n_2757),
.B2(n_2758),
.C(n_2760),
.Y(n_14976)
);

OAI22xp33_ASAP7_75t_SL g14977 ( 
.A1(n_14824),
.A2(n_2761),
.B1(n_2758),
.B2(n_2760),
.Y(n_14977)
);

INVx2_ASAP7_75t_L g14978 ( 
.A(n_14817),
.Y(n_14978)
);

OAI21xp5_ASAP7_75t_L g14979 ( 
.A1(n_14836),
.A2(n_2762),
.B(n_2763),
.Y(n_14979)
);

AOI22xp33_ASAP7_75t_L g14980 ( 
.A1(n_14832),
.A2(n_14796),
.B1(n_14818),
.B2(n_14810),
.Y(n_14980)
);

OAI221xp5_ASAP7_75t_L g14981 ( 
.A1(n_14847),
.A2(n_2764),
.B1(n_2762),
.B2(n_2763),
.C(n_2765),
.Y(n_14981)
);

OAI22xp33_ASAP7_75t_L g14982 ( 
.A1(n_14859),
.A2(n_2767),
.B1(n_2764),
.B2(n_2766),
.Y(n_14982)
);

OAI221xp5_ASAP7_75t_SL g14983 ( 
.A1(n_14831),
.A2(n_2769),
.B1(n_2766),
.B2(n_2768),
.C(n_2770),
.Y(n_14983)
);

O2A1O1Ixp33_ASAP7_75t_L g14984 ( 
.A1(n_14792),
.A2(n_14869),
.B(n_14821),
.C(n_14865),
.Y(n_14984)
);

OAI22xp5_ASAP7_75t_L g14985 ( 
.A1(n_14801),
.A2(n_2770),
.B1(n_2768),
.B2(n_2769),
.Y(n_14985)
);

INVx1_ASAP7_75t_L g14986 ( 
.A(n_14819),
.Y(n_14986)
);

INVx1_ASAP7_75t_L g14987 ( 
.A(n_14822),
.Y(n_14987)
);

NAND2xp5_ASAP7_75t_L g14988 ( 
.A(n_14829),
.B(n_2771),
.Y(n_14988)
);

AOI22xp5_ASAP7_75t_L g14989 ( 
.A1(n_14833),
.A2(n_2773),
.B1(n_2771),
.B2(n_2772),
.Y(n_14989)
);

INVx1_ASAP7_75t_L g14990 ( 
.A(n_14814),
.Y(n_14990)
);

BUFx2_ASAP7_75t_L g14991 ( 
.A(n_14848),
.Y(n_14991)
);

INVx1_ASAP7_75t_L g14992 ( 
.A(n_14852),
.Y(n_14992)
);

AOI21xp33_ASAP7_75t_L g14993 ( 
.A1(n_14835),
.A2(n_2772),
.B(n_2773),
.Y(n_14993)
);

OAI22xp5_ASAP7_75t_L g14994 ( 
.A1(n_14809),
.A2(n_2776),
.B1(n_2774),
.B2(n_2775),
.Y(n_14994)
);

O2A1O1Ixp33_ASAP7_75t_L g14995 ( 
.A1(n_14899),
.A2(n_2777),
.B(n_2775),
.C(n_2776),
.Y(n_14995)
);

INVx1_ASAP7_75t_L g14996 ( 
.A(n_14858),
.Y(n_14996)
);

NAND3xp33_ASAP7_75t_L g14997 ( 
.A(n_14838),
.B(n_2778),
.C(n_2779),
.Y(n_14997)
);

OAI211xp5_ASAP7_75t_L g14998 ( 
.A1(n_14795),
.A2(n_2781),
.B(n_2778),
.C(n_2780),
.Y(n_14998)
);

INVx2_ASAP7_75t_L g14999 ( 
.A(n_14851),
.Y(n_14999)
);

NAND2xp5_ASAP7_75t_L g15000 ( 
.A(n_14803),
.B(n_2780),
.Y(n_15000)
);

OAI221xp5_ASAP7_75t_L g15001 ( 
.A1(n_14876),
.A2(n_14843),
.B1(n_14871),
.B2(n_14856),
.C(n_14857),
.Y(n_15001)
);

AND2x4_ASAP7_75t_L g15002 ( 
.A(n_14863),
.B(n_2781),
.Y(n_15002)
);

BUFx2_ASAP7_75t_L g15003 ( 
.A(n_14808),
.Y(n_15003)
);

OAI22xp5_ASAP7_75t_L g15004 ( 
.A1(n_14874),
.A2(n_14800),
.B1(n_14870),
.B2(n_14883),
.Y(n_15004)
);

AOI21xp5_ASAP7_75t_L g15005 ( 
.A1(n_14878),
.A2(n_2782),
.B(n_2784),
.Y(n_15005)
);

AO22x1_ASAP7_75t_L g15006 ( 
.A1(n_14903),
.A2(n_2786),
.B1(n_2782),
.B2(n_2785),
.Y(n_15006)
);

OAI21xp33_ASAP7_75t_L g15007 ( 
.A1(n_14811),
.A2(n_2785),
.B(n_2787),
.Y(n_15007)
);

INVx1_ASAP7_75t_L g15008 ( 
.A(n_14902),
.Y(n_15008)
);

INVx1_ASAP7_75t_L g15009 ( 
.A(n_14886),
.Y(n_15009)
);

INVx1_ASAP7_75t_L g15010 ( 
.A(n_14786),
.Y(n_15010)
);

INVx1_ASAP7_75t_L g15011 ( 
.A(n_14786),
.Y(n_15011)
);

INVx1_ASAP7_75t_L g15012 ( 
.A(n_14786),
.Y(n_15012)
);

AOI21xp5_ASAP7_75t_L g15013 ( 
.A1(n_14842),
.A2(n_2787),
.B(n_2788),
.Y(n_15013)
);

AOI22xp5_ASAP7_75t_L g15014 ( 
.A1(n_14895),
.A2(n_2791),
.B1(n_2789),
.B2(n_2790),
.Y(n_15014)
);

OAI222xp33_ASAP7_75t_L g15015 ( 
.A1(n_14826),
.A2(n_2792),
.B1(n_2794),
.B2(n_2790),
.C1(n_2791),
.C2(n_2793),
.Y(n_15015)
);

AOI222xp33_ASAP7_75t_L g15016 ( 
.A1(n_14898),
.A2(n_2795),
.B1(n_2797),
.B2(n_2792),
.C1(n_2793),
.C2(n_2796),
.Y(n_15016)
);

AOI221xp5_ASAP7_75t_L g15017 ( 
.A1(n_14868),
.A2(n_2797),
.B1(n_2795),
.B2(n_2796),
.C(n_2798),
.Y(n_15017)
);

AOI22xp33_ASAP7_75t_L g15018 ( 
.A1(n_14834),
.A2(n_2800),
.B1(n_2798),
.B2(n_2799),
.Y(n_15018)
);

INVx1_ASAP7_75t_L g15019 ( 
.A(n_14786),
.Y(n_15019)
);

INVx2_ASAP7_75t_L g15020 ( 
.A(n_14880),
.Y(n_15020)
);

OAI221xp5_ASAP7_75t_L g15021 ( 
.A1(n_14898),
.A2(n_2802),
.B1(n_2800),
.B2(n_2801),
.C(n_2803),
.Y(n_15021)
);

AND3x1_ASAP7_75t_L g15022 ( 
.A(n_14890),
.B(n_2801),
.C(n_2802),
.Y(n_15022)
);

AO21x1_ASAP7_75t_L g15023 ( 
.A1(n_14786),
.A2(n_2803),
.B(n_2804),
.Y(n_15023)
);

INVx2_ASAP7_75t_L g15024 ( 
.A(n_14880),
.Y(n_15024)
);

INVxp67_ASAP7_75t_SL g15025 ( 
.A(n_14787),
.Y(n_15025)
);

OAI22xp5_ASAP7_75t_L g15026 ( 
.A1(n_14806),
.A2(n_2806),
.B1(n_2804),
.B2(n_2805),
.Y(n_15026)
);

OA33x2_ASAP7_75t_L g15027 ( 
.A1(n_14867),
.A2(n_2808),
.A3(n_2810),
.B1(n_2805),
.B2(n_2807),
.B3(n_2809),
.Y(n_15027)
);

OAI31xp33_ASAP7_75t_L g15028 ( 
.A1(n_14898),
.A2(n_2809),
.A3(n_2807),
.B(n_2808),
.Y(n_15028)
);

AOI22xp5_ASAP7_75t_L g15029 ( 
.A1(n_14895),
.A2(n_2812),
.B1(n_2810),
.B2(n_2811),
.Y(n_15029)
);

OAI21xp5_ASAP7_75t_SL g15030 ( 
.A1(n_14826),
.A2(n_2811),
.B(n_2812),
.Y(n_15030)
);

INVx2_ASAP7_75t_L g15031 ( 
.A(n_14880),
.Y(n_15031)
);

OR2x2_ASAP7_75t_L g15032 ( 
.A(n_14787),
.B(n_2813),
.Y(n_15032)
);

AOI222xp33_ASAP7_75t_L g15033 ( 
.A1(n_14898),
.A2(n_2815),
.B1(n_2817),
.B2(n_2813),
.C1(n_2814),
.C2(n_2816),
.Y(n_15033)
);

OAI222xp33_ASAP7_75t_L g15034 ( 
.A1(n_14826),
.A2(n_2816),
.B1(n_2818),
.B2(n_2814),
.C1(n_2815),
.C2(n_2817),
.Y(n_15034)
);

OAI22xp5_ASAP7_75t_L g15035 ( 
.A1(n_14806),
.A2(n_2820),
.B1(n_2818),
.B2(n_2819),
.Y(n_15035)
);

O2A1O1Ixp33_ASAP7_75t_L g15036 ( 
.A1(n_14786),
.A2(n_2821),
.B(n_2819),
.C(n_2820),
.Y(n_15036)
);

A2O1A1Ixp33_ASAP7_75t_L g15037 ( 
.A1(n_14875),
.A2(n_2823),
.B(n_2821),
.C(n_2822),
.Y(n_15037)
);

AOI22xp5_ASAP7_75t_L g15038 ( 
.A1(n_14895),
.A2(n_2825),
.B1(n_2822),
.B2(n_2824),
.Y(n_15038)
);

AOI22xp5_ASAP7_75t_L g15039 ( 
.A1(n_14895),
.A2(n_2827),
.B1(n_2824),
.B2(n_2826),
.Y(n_15039)
);

INVx2_ASAP7_75t_L g15040 ( 
.A(n_14910),
.Y(n_15040)
);

OAI32xp33_ASAP7_75t_L g15041 ( 
.A1(n_14914),
.A2(n_2829),
.A3(n_2827),
.B1(n_2828),
.B2(n_2830),
.Y(n_15041)
);

NOR2xp33_ASAP7_75t_L g15042 ( 
.A(n_14948),
.B(n_2828),
.Y(n_15042)
);

OAI221xp5_ASAP7_75t_L g15043 ( 
.A1(n_15027),
.A2(n_2831),
.B1(n_2829),
.B2(n_2830),
.C(n_2832),
.Y(n_15043)
);

INVx1_ASAP7_75t_L g15044 ( 
.A(n_15023),
.Y(n_15044)
);

INVx1_ASAP7_75t_L g15045 ( 
.A(n_14955),
.Y(n_15045)
);

INVx1_ASAP7_75t_L g15046 ( 
.A(n_14951),
.Y(n_15046)
);

INVx1_ASAP7_75t_L g15047 ( 
.A(n_15032),
.Y(n_15047)
);

NAND3xp33_ASAP7_75t_L g15048 ( 
.A(n_15028),
.B(n_2832),
.C(n_2833),
.Y(n_15048)
);

OAI31xp33_ASAP7_75t_L g15049 ( 
.A1(n_14922),
.A2(n_2835),
.A3(n_2833),
.B(n_2834),
.Y(n_15049)
);

NAND2xp5_ASAP7_75t_L g15050 ( 
.A(n_15025),
.B(n_2834),
.Y(n_15050)
);

INVx2_ASAP7_75t_SL g15051 ( 
.A(n_15020),
.Y(n_15051)
);

INVx1_ASAP7_75t_L g15052 ( 
.A(n_14964),
.Y(n_15052)
);

AOI21xp33_ASAP7_75t_L g15053 ( 
.A1(n_15010),
.A2(n_2835),
.B(n_2836),
.Y(n_15053)
);

INVxp67_ASAP7_75t_L g15054 ( 
.A(n_14953),
.Y(n_15054)
);

INVx1_ASAP7_75t_L g15055 ( 
.A(n_14965),
.Y(n_15055)
);

AND2x2_ASAP7_75t_SL g15056 ( 
.A(n_15022),
.B(n_2837),
.Y(n_15056)
);

INVx2_ASAP7_75t_L g15057 ( 
.A(n_14965),
.Y(n_15057)
);

OR2x2_ASAP7_75t_L g15058 ( 
.A(n_14957),
.B(n_2837),
.Y(n_15058)
);

NAND2xp5_ASAP7_75t_L g15059 ( 
.A(n_15006),
.B(n_2838),
.Y(n_15059)
);

INVx1_ASAP7_75t_L g15060 ( 
.A(n_15002),
.Y(n_15060)
);

INVx1_ASAP7_75t_L g15061 ( 
.A(n_15002),
.Y(n_15061)
);

AOI22xp5_ASAP7_75t_L g15062 ( 
.A1(n_14935),
.A2(n_2840),
.B1(n_2838),
.B2(n_2839),
.Y(n_15062)
);

INVx2_ASAP7_75t_L g15063 ( 
.A(n_15024),
.Y(n_15063)
);

OR2x2_ASAP7_75t_L g15064 ( 
.A(n_14927),
.B(n_2839),
.Y(n_15064)
);

INVx1_ASAP7_75t_L g15065 ( 
.A(n_14952),
.Y(n_15065)
);

INVx1_ASAP7_75t_L g15066 ( 
.A(n_15031),
.Y(n_15066)
);

AOI221xp5_ASAP7_75t_L g15067 ( 
.A1(n_14913),
.A2(n_2842),
.B1(n_2840),
.B2(n_2841),
.C(n_2843),
.Y(n_15067)
);

INVx1_ASAP7_75t_L g15068 ( 
.A(n_14924),
.Y(n_15068)
);

AOI22xp5_ASAP7_75t_L g15069 ( 
.A1(n_15009),
.A2(n_14968),
.B1(n_15008),
.B2(n_14934),
.Y(n_15069)
);

AOI22xp5_ASAP7_75t_L g15070 ( 
.A1(n_14996),
.A2(n_14999),
.B1(n_14923),
.B2(n_15011),
.Y(n_15070)
);

INVx1_ASAP7_75t_L g15071 ( 
.A(n_14919),
.Y(n_15071)
);

INVx1_ASAP7_75t_L g15072 ( 
.A(n_14966),
.Y(n_15072)
);

OAI321xp33_ASAP7_75t_L g15073 ( 
.A1(n_15012),
.A2(n_2844),
.A3(n_2846),
.B1(n_2841),
.B2(n_2843),
.C(n_2845),
.Y(n_15073)
);

OAI22xp5_ASAP7_75t_L g15074 ( 
.A1(n_14980),
.A2(n_2847),
.B1(n_2844),
.B2(n_2845),
.Y(n_15074)
);

AOI21xp33_ASAP7_75t_SL g15075 ( 
.A1(n_15016),
.A2(n_2848),
.B(n_2849),
.Y(n_15075)
);

O2A1O1Ixp33_ASAP7_75t_SL g15076 ( 
.A1(n_15037),
.A2(n_2850),
.B(n_2848),
.C(n_2849),
.Y(n_15076)
);

OAI22xp33_ASAP7_75t_L g15077 ( 
.A1(n_15019),
.A2(n_2853),
.B1(n_2850),
.B2(n_2852),
.Y(n_15077)
);

AOI222xp33_ASAP7_75t_L g15078 ( 
.A1(n_15007),
.A2(n_2855),
.B1(n_2857),
.B2(n_2852),
.C1(n_2854),
.C2(n_2856),
.Y(n_15078)
);

AOI21xp5_ASAP7_75t_L g15079 ( 
.A1(n_14954),
.A2(n_14961),
.B(n_14937),
.Y(n_15079)
);

NOR2x1_ASAP7_75t_SL g15080 ( 
.A(n_14998),
.B(n_2855),
.Y(n_15080)
);

INVx1_ASAP7_75t_L g15081 ( 
.A(n_14967),
.Y(n_15081)
);

OAI322xp33_ASAP7_75t_L g15082 ( 
.A1(n_14969),
.A2(n_2861),
.A3(n_2860),
.B1(n_2858),
.B2(n_2856),
.C1(n_2857),
.C2(n_2859),
.Y(n_15082)
);

INVx1_ASAP7_75t_L g15083 ( 
.A(n_14943),
.Y(n_15083)
);

INVx1_ASAP7_75t_SL g15084 ( 
.A(n_14991),
.Y(n_15084)
);

INVx2_ASAP7_75t_L g15085 ( 
.A(n_14959),
.Y(n_15085)
);

AOI22xp33_ASAP7_75t_SL g15086 ( 
.A1(n_15003),
.A2(n_14947),
.B1(n_14942),
.B2(n_14932),
.Y(n_15086)
);

NAND3xp33_ASAP7_75t_L g15087 ( 
.A(n_14915),
.B(n_2858),
.C(n_2859),
.Y(n_15087)
);

A2O1A1Ixp33_ASAP7_75t_L g15088 ( 
.A1(n_15036),
.A2(n_2862),
.B(n_2860),
.C(n_2861),
.Y(n_15088)
);

INVx1_ASAP7_75t_L g15089 ( 
.A(n_14997),
.Y(n_15089)
);

O2A1O1Ixp33_ASAP7_75t_L g15090 ( 
.A1(n_15030),
.A2(n_14929),
.B(n_15034),
.C(n_15015),
.Y(n_15090)
);

OAI22xp5_ASAP7_75t_L g15091 ( 
.A1(n_14939),
.A2(n_2864),
.B1(n_2862),
.B2(n_2863),
.Y(n_15091)
);

INVx1_ASAP7_75t_L g15092 ( 
.A(n_14971),
.Y(n_15092)
);

AOI22xp5_ASAP7_75t_L g15093 ( 
.A1(n_14962),
.A2(n_2865),
.B1(n_2863),
.B2(n_2864),
.Y(n_15093)
);

INVx1_ASAP7_75t_L g15094 ( 
.A(n_14988),
.Y(n_15094)
);

AOI21xp5_ASAP7_75t_SL g15095 ( 
.A1(n_14977),
.A2(n_2865),
.B(n_2866),
.Y(n_15095)
);

INVx1_ASAP7_75t_L g15096 ( 
.A(n_14995),
.Y(n_15096)
);

INVx1_ASAP7_75t_L g15097 ( 
.A(n_15000),
.Y(n_15097)
);

INVxp67_ASAP7_75t_SL g15098 ( 
.A(n_14950),
.Y(n_15098)
);

INVx1_ASAP7_75t_L g15099 ( 
.A(n_14917),
.Y(n_15099)
);

INVx2_ASAP7_75t_SL g15100 ( 
.A(n_14930),
.Y(n_15100)
);

AOI321xp33_ASAP7_75t_L g15101 ( 
.A1(n_14984),
.A2(n_2868),
.A3(n_2870),
.B1(n_2866),
.B2(n_2867),
.C(n_2869),
.Y(n_15101)
);

NAND2xp5_ASAP7_75t_L g15102 ( 
.A(n_14933),
.B(n_2867),
.Y(n_15102)
);

AOI221xp5_ASAP7_75t_L g15103 ( 
.A1(n_14926),
.A2(n_2872),
.B1(n_2869),
.B2(n_2871),
.C(n_2873),
.Y(n_15103)
);

INVx2_ASAP7_75t_L g15104 ( 
.A(n_14938),
.Y(n_15104)
);

OAI222xp33_ASAP7_75t_L g15105 ( 
.A1(n_15001),
.A2(n_2873),
.B1(n_2875),
.B2(n_2871),
.C1(n_2872),
.C2(n_2874),
.Y(n_15105)
);

INVx1_ASAP7_75t_L g15106 ( 
.A(n_14921),
.Y(n_15106)
);

AND2x2_ASAP7_75t_L g15107 ( 
.A(n_14920),
.B(n_2874),
.Y(n_15107)
);

AOI22xp5_ASAP7_75t_L g15108 ( 
.A1(n_14925),
.A2(n_2878),
.B1(n_2876),
.B2(n_2877),
.Y(n_15108)
);

OR2x2_ASAP7_75t_L g15109 ( 
.A(n_14994),
.B(n_2876),
.Y(n_15109)
);

AOI221xp5_ASAP7_75t_L g15110 ( 
.A1(n_15004),
.A2(n_2880),
.B1(n_2878),
.B2(n_2879),
.C(n_2881),
.Y(n_15110)
);

INVx1_ASAP7_75t_L g15111 ( 
.A(n_14960),
.Y(n_15111)
);

INVxp67_ASAP7_75t_SL g15112 ( 
.A(n_15033),
.Y(n_15112)
);

INVx1_ASAP7_75t_L g15113 ( 
.A(n_14944),
.Y(n_15113)
);

INVx1_ASAP7_75t_L g15114 ( 
.A(n_14981),
.Y(n_15114)
);

AOI22xp33_ASAP7_75t_L g15115 ( 
.A1(n_14974),
.A2(n_2883),
.B1(n_2879),
.B2(n_2882),
.Y(n_15115)
);

INVx1_ASAP7_75t_L g15116 ( 
.A(n_14979),
.Y(n_15116)
);

OAI21xp33_ASAP7_75t_SL g15117 ( 
.A1(n_15017),
.A2(n_2882),
.B(n_2883),
.Y(n_15117)
);

INVx1_ASAP7_75t_L g15118 ( 
.A(n_14975),
.Y(n_15118)
);

XNOR2x2_ASAP7_75t_L g15119 ( 
.A(n_14916),
.B(n_2884),
.Y(n_15119)
);

OAI21xp33_ASAP7_75t_L g15120 ( 
.A1(n_14958),
.A2(n_2884),
.B(n_2885),
.Y(n_15120)
);

INVx1_ASAP7_75t_L g15121 ( 
.A(n_15021),
.Y(n_15121)
);

AOI21xp33_ASAP7_75t_L g15122 ( 
.A1(n_14985),
.A2(n_2885),
.B(n_2886),
.Y(n_15122)
);

OAI22xp5_ASAP7_75t_L g15123 ( 
.A1(n_14909),
.A2(n_2888),
.B1(n_2886),
.B2(n_2887),
.Y(n_15123)
);

INVx1_ASAP7_75t_SL g15124 ( 
.A(n_15013),
.Y(n_15124)
);

OR2x2_ASAP7_75t_L g15125 ( 
.A(n_15005),
.B(n_2887),
.Y(n_15125)
);

NOR2xp33_ASAP7_75t_R g15126 ( 
.A(n_14986),
.B(n_2888),
.Y(n_15126)
);

OAI221xp5_ASAP7_75t_L g15127 ( 
.A1(n_14946),
.A2(n_14972),
.B1(n_14973),
.B2(n_15029),
.C(n_15014),
.Y(n_15127)
);

AOI221xp5_ASAP7_75t_L g15128 ( 
.A1(n_14982),
.A2(n_2891),
.B1(n_2889),
.B2(n_2890),
.C(n_2892),
.Y(n_15128)
);

NAND3xp33_ASAP7_75t_L g15129 ( 
.A(n_14956),
.B(n_2889),
.C(n_2890),
.Y(n_15129)
);

INVx1_ASAP7_75t_L g15130 ( 
.A(n_15038),
.Y(n_15130)
);

OR2x2_ASAP7_75t_L g15131 ( 
.A(n_14978),
.B(n_2891),
.Y(n_15131)
);

AOI22xp33_ASAP7_75t_L g15132 ( 
.A1(n_14987),
.A2(n_2895),
.B1(n_2893),
.B2(n_2894),
.Y(n_15132)
);

AND2x2_ASAP7_75t_L g15133 ( 
.A(n_14990),
.B(n_2893),
.Y(n_15133)
);

AOI211xp5_ASAP7_75t_L g15134 ( 
.A1(n_14983),
.A2(n_2896),
.B(n_2894),
.C(n_2895),
.Y(n_15134)
);

NAND2xp5_ASAP7_75t_L g15135 ( 
.A(n_15039),
.B(n_2896),
.Y(n_15135)
);

AOI222xp33_ASAP7_75t_L g15136 ( 
.A1(n_14992),
.A2(n_2899),
.B1(n_2901),
.B2(n_2897),
.C1(n_2898),
.C2(n_2900),
.Y(n_15136)
);

INVx2_ASAP7_75t_L g15137 ( 
.A(n_14928),
.Y(n_15137)
);

INVx1_ASAP7_75t_L g15138 ( 
.A(n_14918),
.Y(n_15138)
);

AOI22xp5_ASAP7_75t_L g15139 ( 
.A1(n_14936),
.A2(n_2900),
.B1(n_2897),
.B2(n_2898),
.Y(n_15139)
);

NAND2xp5_ASAP7_75t_L g15140 ( 
.A(n_14911),
.B(n_2901),
.Y(n_15140)
);

OAI21xp5_ASAP7_75t_L g15141 ( 
.A1(n_14912),
.A2(n_2902),
.B(n_2903),
.Y(n_15141)
);

AND2x2_ASAP7_75t_L g15142 ( 
.A(n_14993),
.B(n_2902),
.Y(n_15142)
);

NAND2xp5_ASAP7_75t_L g15143 ( 
.A(n_15018),
.B(n_2903),
.Y(n_15143)
);

INVx1_ASAP7_75t_L g15144 ( 
.A(n_14931),
.Y(n_15144)
);

NAND2xp5_ASAP7_75t_L g15145 ( 
.A(n_14989),
.B(n_2904),
.Y(n_15145)
);

AND2x2_ASAP7_75t_L g15146 ( 
.A(n_14970),
.B(n_2904),
.Y(n_15146)
);

OAI31xp33_ASAP7_75t_L g15147 ( 
.A1(n_15026),
.A2(n_2907),
.A3(n_2905),
.B(n_2906),
.Y(n_15147)
);

OAI22xp5_ASAP7_75t_L g15148 ( 
.A1(n_14949),
.A2(n_2907),
.B1(n_2905),
.B2(n_2906),
.Y(n_15148)
);

INVx1_ASAP7_75t_L g15149 ( 
.A(n_15035),
.Y(n_15149)
);

INVx2_ASAP7_75t_L g15150 ( 
.A(n_14945),
.Y(n_15150)
);

NAND2xp5_ASAP7_75t_L g15151 ( 
.A(n_14976),
.B(n_2908),
.Y(n_15151)
);

AND2x2_ASAP7_75t_L g15152 ( 
.A(n_14963),
.B(n_2908),
.Y(n_15152)
);

OAI221xp5_ASAP7_75t_L g15153 ( 
.A1(n_14940),
.A2(n_2911),
.B1(n_2909),
.B2(n_2910),
.C(n_2912),
.Y(n_15153)
);

OR2x2_ASAP7_75t_L g15154 ( 
.A(n_15058),
.B(n_15050),
.Y(n_15154)
);

INVx1_ASAP7_75t_L g15155 ( 
.A(n_15133),
.Y(n_15155)
);

AOI21xp33_ASAP7_75t_L g15156 ( 
.A1(n_15051),
.A2(n_15084),
.B(n_15045),
.Y(n_15156)
);

NAND2xp5_ASAP7_75t_L g15157 ( 
.A(n_15056),
.B(n_14941),
.Y(n_15157)
);

NOR3xp33_ASAP7_75t_L g15158 ( 
.A(n_15066),
.B(n_2909),
.C(n_2911),
.Y(n_15158)
);

OAI211xp5_ASAP7_75t_L g15159 ( 
.A1(n_15093),
.A2(n_2914),
.B(n_2912),
.C(n_2913),
.Y(n_15159)
);

NAND2xp5_ASAP7_75t_SL g15160 ( 
.A(n_15101),
.B(n_2913),
.Y(n_15160)
);

INVx1_ASAP7_75t_L g15161 ( 
.A(n_15131),
.Y(n_15161)
);

A2O1A1Ixp33_ASAP7_75t_SL g15162 ( 
.A1(n_15063),
.A2(n_2916),
.B(n_2914),
.C(n_2915),
.Y(n_15162)
);

NAND3xp33_ASAP7_75t_SL g15163 ( 
.A(n_15049),
.B(n_2915),
.C(n_2916),
.Y(n_15163)
);

INVxp67_ASAP7_75t_SL g15164 ( 
.A(n_15059),
.Y(n_15164)
);

OAI31xp33_ASAP7_75t_L g15165 ( 
.A1(n_15044),
.A2(n_2919),
.A3(n_2917),
.B(n_2918),
.Y(n_15165)
);

O2A1O1Ixp33_ASAP7_75t_L g15166 ( 
.A1(n_15088),
.A2(n_2919),
.B(n_2917),
.C(n_2918),
.Y(n_15166)
);

OAI21xp5_ASAP7_75t_L g15167 ( 
.A1(n_15048),
.A2(n_2920),
.B(n_2921),
.Y(n_15167)
);

AOI22x1_ASAP7_75t_L g15168 ( 
.A1(n_15078),
.A2(n_2922),
.B1(n_2920),
.B2(n_2921),
.Y(n_15168)
);

AOI222xp33_ASAP7_75t_L g15169 ( 
.A1(n_15054),
.A2(n_15112),
.B1(n_15065),
.B2(n_15098),
.C1(n_15081),
.C2(n_15117),
.Y(n_15169)
);

INVx1_ASAP7_75t_L g15170 ( 
.A(n_15064),
.Y(n_15170)
);

INVx1_ASAP7_75t_L g15171 ( 
.A(n_15125),
.Y(n_15171)
);

OAI211xp5_ASAP7_75t_L g15172 ( 
.A1(n_15070),
.A2(n_2924),
.B(n_2922),
.C(n_2923),
.Y(n_15172)
);

NAND2xp5_ASAP7_75t_L g15173 ( 
.A(n_15042),
.B(n_2923),
.Y(n_15173)
);

AOI222xp33_ASAP7_75t_L g15174 ( 
.A1(n_15071),
.A2(n_2927),
.B1(n_2929),
.B2(n_2925),
.C1(n_2926),
.C2(n_2928),
.Y(n_15174)
);

AOI221xp5_ASAP7_75t_L g15175 ( 
.A1(n_15075),
.A2(n_2928),
.B1(n_2925),
.B2(n_2927),
.C(n_2930),
.Y(n_15175)
);

INVx1_ASAP7_75t_L g15176 ( 
.A(n_15080),
.Y(n_15176)
);

AOI22xp33_ASAP7_75t_L g15177 ( 
.A1(n_15085),
.A2(n_2932),
.B1(n_2930),
.B2(n_2931),
.Y(n_15177)
);

AOI22x1_ASAP7_75t_L g15178 ( 
.A1(n_15057),
.A2(n_15061),
.B1(n_15060),
.B2(n_15055),
.Y(n_15178)
);

INVx1_ASAP7_75t_L g15179 ( 
.A(n_15140),
.Y(n_15179)
);

OAI221xp5_ASAP7_75t_L g15180 ( 
.A1(n_15147),
.A2(n_2934),
.B1(n_2931),
.B2(n_2933),
.C(n_2935),
.Y(n_15180)
);

OAI21xp5_ASAP7_75t_L g15181 ( 
.A1(n_15129),
.A2(n_2933),
.B(n_2935),
.Y(n_15181)
);

AOI221xp5_ASAP7_75t_L g15182 ( 
.A1(n_15122),
.A2(n_2938),
.B1(n_2936),
.B2(n_2937),
.C(n_2939),
.Y(n_15182)
);

NAND3xp33_ASAP7_75t_L g15183 ( 
.A(n_15134),
.B(n_2936),
.C(n_2937),
.Y(n_15183)
);

NOR3xp33_ASAP7_75t_L g15184 ( 
.A(n_15086),
.B(n_2938),
.C(n_2940),
.Y(n_15184)
);

AOI221xp5_ASAP7_75t_L g15185 ( 
.A1(n_15076),
.A2(n_2942),
.B1(n_2940),
.B2(n_2941),
.C(n_2943),
.Y(n_15185)
);

NAND2xp5_ASAP7_75t_L g15186 ( 
.A(n_15062),
.B(n_2941),
.Y(n_15186)
);

OAI21xp33_ASAP7_75t_L g15187 ( 
.A1(n_15069),
.A2(n_2942),
.B(n_2943),
.Y(n_15187)
);

OAI211xp5_ASAP7_75t_L g15188 ( 
.A1(n_15103),
.A2(n_2947),
.B(n_2945),
.C(n_2946),
.Y(n_15188)
);

AOI22xp5_ASAP7_75t_L g15189 ( 
.A1(n_15100),
.A2(n_2947),
.B1(n_2945),
.B2(n_2946),
.Y(n_15189)
);

OAI21xp33_ASAP7_75t_L g15190 ( 
.A1(n_15138),
.A2(n_2948),
.B(n_2949),
.Y(n_15190)
);

AOI21xp5_ASAP7_75t_L g15191 ( 
.A1(n_15095),
.A2(n_2948),
.B(n_2949),
.Y(n_15191)
);

OAI322xp33_ASAP7_75t_L g15192 ( 
.A1(n_15096),
.A2(n_2955),
.A3(n_2954),
.B1(n_2952),
.B2(n_2950),
.C1(n_2951),
.C2(n_2953),
.Y(n_15192)
);

NAND3xp33_ASAP7_75t_SL g15193 ( 
.A(n_15124),
.B(n_15141),
.C(n_15067),
.Y(n_15193)
);

AOI21xp5_ASAP7_75t_L g15194 ( 
.A1(n_15090),
.A2(n_15079),
.B(n_15102),
.Y(n_15194)
);

OAI31xp33_ASAP7_75t_L g15195 ( 
.A1(n_15043),
.A2(n_2952),
.A3(n_2950),
.B(n_2951),
.Y(n_15195)
);

INVx1_ASAP7_75t_L g15196 ( 
.A(n_15108),
.Y(n_15196)
);

OAI221xp5_ASAP7_75t_L g15197 ( 
.A1(n_15120),
.A2(n_2957),
.B1(n_2954),
.B2(n_2956),
.C(n_2958),
.Y(n_15197)
);

AOI221xp5_ASAP7_75t_L g15198 ( 
.A1(n_15127),
.A2(n_2959),
.B1(n_2956),
.B2(n_2958),
.C(n_2960),
.Y(n_15198)
);

OAI221xp5_ASAP7_75t_L g15199 ( 
.A1(n_15083),
.A2(n_2961),
.B1(n_2959),
.B2(n_2960),
.C(n_2963),
.Y(n_15199)
);

NAND3xp33_ASAP7_75t_SL g15200 ( 
.A(n_15072),
.B(n_2961),
.C(n_2963),
.Y(n_15200)
);

NAND2xp5_ASAP7_75t_L g15201 ( 
.A(n_15046),
.B(n_2964),
.Y(n_15201)
);

OAI22x1_ASAP7_75t_SL g15202 ( 
.A1(n_15047),
.A2(n_2966),
.B1(n_2964),
.B2(n_2965),
.Y(n_15202)
);

OAI22xp33_ASAP7_75t_L g15203 ( 
.A1(n_15139),
.A2(n_2967),
.B1(n_2965),
.B2(n_2966),
.Y(n_15203)
);

INVxp67_ASAP7_75t_L g15204 ( 
.A(n_15142),
.Y(n_15204)
);

INVx1_ASAP7_75t_L g15205 ( 
.A(n_15119),
.Y(n_15205)
);

AOI21xp5_ASAP7_75t_L g15206 ( 
.A1(n_15151),
.A2(n_2967),
.B(n_2968),
.Y(n_15206)
);

AOI22xp5_ASAP7_75t_L g15207 ( 
.A1(n_15149),
.A2(n_2970),
.B1(n_2968),
.B2(n_2969),
.Y(n_15207)
);

OAI221xp5_ASAP7_75t_L g15208 ( 
.A1(n_15128),
.A2(n_2972),
.B1(n_2970),
.B2(n_2971),
.C(n_2973),
.Y(n_15208)
);

INVx2_ASAP7_75t_SL g15209 ( 
.A(n_15126),
.Y(n_15209)
);

AOI221x1_ASAP7_75t_L g15210 ( 
.A1(n_15068),
.A2(n_2974),
.B1(n_2971),
.B2(n_2973),
.C(n_2975),
.Y(n_15210)
);

AOI222xp33_ASAP7_75t_L g15211 ( 
.A1(n_15089),
.A2(n_2976),
.B1(n_2978),
.B2(n_2974),
.C1(n_2975),
.C2(n_2977),
.Y(n_15211)
);

OAI22xp33_ASAP7_75t_L g15212 ( 
.A1(n_15109),
.A2(n_2979),
.B1(n_2976),
.B2(n_2977),
.Y(n_15212)
);

AOI221x1_ASAP7_75t_L g15213 ( 
.A1(n_15111),
.A2(n_2983),
.B1(n_2979),
.B2(n_2980),
.C(n_2984),
.Y(n_15213)
);

AOI21xp5_ASAP7_75t_L g15214 ( 
.A1(n_15135),
.A2(n_2980),
.B(n_2983),
.Y(n_15214)
);

NOR2xp67_ASAP7_75t_L g15215 ( 
.A(n_15073),
.B(n_2985),
.Y(n_15215)
);

NAND2xp5_ASAP7_75t_L g15216 ( 
.A(n_15077),
.B(n_2985),
.Y(n_15216)
);

INVx1_ASAP7_75t_L g15217 ( 
.A(n_15107),
.Y(n_15217)
);

O2A1O1Ixp33_ASAP7_75t_L g15218 ( 
.A1(n_15105),
.A2(n_2988),
.B(n_2986),
.C(n_2987),
.Y(n_15218)
);

NAND2xp5_ASAP7_75t_L g15219 ( 
.A(n_15074),
.B(n_2986),
.Y(n_15219)
);

NAND3xp33_ASAP7_75t_L g15220 ( 
.A(n_15087),
.B(n_2987),
.C(n_2988),
.Y(n_15220)
);

AND2x2_ASAP7_75t_L g15221 ( 
.A(n_15040),
.B(n_2989),
.Y(n_15221)
);

NAND4xp25_ASAP7_75t_L g15222 ( 
.A(n_15121),
.B(n_15114),
.C(n_15099),
.D(n_15130),
.Y(n_15222)
);

OAI221xp5_ASAP7_75t_L g15223 ( 
.A1(n_15143),
.A2(n_2991),
.B1(n_2989),
.B2(n_2990),
.C(n_2992),
.Y(n_15223)
);

OAI21xp33_ASAP7_75t_L g15224 ( 
.A1(n_15113),
.A2(n_2990),
.B(n_2992),
.Y(n_15224)
);

OA22x2_ASAP7_75t_L g15225 ( 
.A1(n_15104),
.A2(n_2995),
.B1(n_2993),
.B2(n_2994),
.Y(n_15225)
);

OAI32xp33_ASAP7_75t_L g15226 ( 
.A1(n_15145),
.A2(n_2995),
.A3(n_2993),
.B1(n_2994),
.B2(n_2996),
.Y(n_15226)
);

INVx1_ASAP7_75t_L g15227 ( 
.A(n_15152),
.Y(n_15227)
);

AOI211x1_ASAP7_75t_L g15228 ( 
.A1(n_15118),
.A2(n_2998),
.B(n_2996),
.C(n_2997),
.Y(n_15228)
);

INVx1_ASAP7_75t_SL g15229 ( 
.A(n_15146),
.Y(n_15229)
);

INVx1_ASAP7_75t_L g15230 ( 
.A(n_15052),
.Y(n_15230)
);

NOR2x1_ASAP7_75t_L g15231 ( 
.A(n_15082),
.B(n_2997),
.Y(n_15231)
);

NOR2xp33_ASAP7_75t_SL g15232 ( 
.A(n_15153),
.B(n_2998),
.Y(n_15232)
);

NOR2x1_ASAP7_75t_L g15233 ( 
.A(n_15106),
.B(n_2999),
.Y(n_15233)
);

OAI32xp33_ASAP7_75t_L g15234 ( 
.A1(n_15150),
.A2(n_3001),
.A3(n_2999),
.B1(n_3000),
.B2(n_3003),
.Y(n_15234)
);

OA22x2_ASAP7_75t_L g15235 ( 
.A1(n_15144),
.A2(n_3003),
.B1(n_3000),
.B2(n_3001),
.Y(n_15235)
);

NAND2xp5_ASAP7_75t_L g15236 ( 
.A(n_15115),
.B(n_3004),
.Y(n_15236)
);

AOI221xp5_ASAP7_75t_L g15237 ( 
.A1(n_15116),
.A2(n_3006),
.B1(n_3004),
.B2(n_3005),
.C(n_3008),
.Y(n_15237)
);

AOI221xp5_ASAP7_75t_L g15238 ( 
.A1(n_15137),
.A2(n_3009),
.B1(n_3005),
.B2(n_3008),
.C(n_3010),
.Y(n_15238)
);

AOI211xp5_ASAP7_75t_L g15239 ( 
.A1(n_15091),
.A2(n_3011),
.B(n_3009),
.C(n_3010),
.Y(n_15239)
);

AOI21xp33_ASAP7_75t_L g15240 ( 
.A1(n_15097),
.A2(n_3012),
.B(n_3013),
.Y(n_15240)
);

AOI322xp5_ASAP7_75t_L g15241 ( 
.A1(n_15092),
.A2(n_3017),
.A3(n_3016),
.B1(n_3014),
.B2(n_3012),
.C1(n_3013),
.C2(n_3015),
.Y(n_15241)
);

OAI221xp5_ASAP7_75t_L g15242 ( 
.A1(n_15123),
.A2(n_3016),
.B1(n_3014),
.B2(n_3015),
.C(n_3017),
.Y(n_15242)
);

NOR2xp33_ASAP7_75t_L g15243 ( 
.A(n_15053),
.B(n_3018),
.Y(n_15243)
);

INVx1_ASAP7_75t_L g15244 ( 
.A(n_15148),
.Y(n_15244)
);

NAND2xp5_ASAP7_75t_L g15245 ( 
.A(n_15136),
.B(n_3018),
.Y(n_15245)
);

AOI21xp5_ASAP7_75t_L g15246 ( 
.A1(n_15094),
.A2(n_3019),
.B(n_3020),
.Y(n_15246)
);

INVx2_ASAP7_75t_L g15247 ( 
.A(n_15041),
.Y(n_15247)
);

OAI21xp5_ASAP7_75t_L g15248 ( 
.A1(n_15110),
.A2(n_3020),
.B(n_3021),
.Y(n_15248)
);

AOI22xp33_ASAP7_75t_L g15249 ( 
.A1(n_15132),
.A2(n_3023),
.B1(n_3021),
.B2(n_3022),
.Y(n_15249)
);

NAND3xp33_ASAP7_75t_L g15250 ( 
.A(n_15101),
.B(n_3022),
.C(n_3023),
.Y(n_15250)
);

A2O1A1Ixp33_ASAP7_75t_L g15251 ( 
.A1(n_15049),
.A2(n_3027),
.B(n_3025),
.C(n_3026),
.Y(n_15251)
);

A2O1A1Ixp33_ASAP7_75t_L g15252 ( 
.A1(n_15049),
.A2(n_3028),
.B(n_3026),
.C(n_3027),
.Y(n_15252)
);

NAND2xp5_ASAP7_75t_L g15253 ( 
.A(n_15133),
.B(n_3029),
.Y(n_15253)
);

AOI22xp5_ASAP7_75t_L g15254 ( 
.A1(n_15051),
.A2(n_3033),
.B1(n_3030),
.B2(n_3032),
.Y(n_15254)
);

NOR2xp33_ASAP7_75t_SL g15255 ( 
.A(n_15056),
.B(n_3030),
.Y(n_15255)
);

NAND2xp5_ASAP7_75t_L g15256 ( 
.A(n_15221),
.B(n_3034),
.Y(n_15256)
);

AOI322xp5_ASAP7_75t_L g15257 ( 
.A1(n_15205),
.A2(n_3039),
.A3(n_3038),
.B1(n_3036),
.B2(n_3034),
.C1(n_3035),
.C2(n_3037),
.Y(n_15257)
);

AOI221xp5_ASAP7_75t_L g15258 ( 
.A1(n_15156),
.A2(n_3037),
.B1(n_3035),
.B2(n_3036),
.C(n_3038),
.Y(n_15258)
);

OAI21xp33_ASAP7_75t_SL g15259 ( 
.A1(n_15195),
.A2(n_3039),
.B(n_3040),
.Y(n_15259)
);

AOI221xp5_ASAP7_75t_L g15260 ( 
.A1(n_15187),
.A2(n_3042),
.B1(n_3040),
.B2(n_3041),
.C(n_3043),
.Y(n_15260)
);

AOI21xp5_ASAP7_75t_L g15261 ( 
.A1(n_15191),
.A2(n_3041),
.B(n_3042),
.Y(n_15261)
);

AOI211xp5_ASAP7_75t_SL g15262 ( 
.A1(n_15190),
.A2(n_3046),
.B(n_3044),
.C(n_3045),
.Y(n_15262)
);

NAND2xp5_ASAP7_75t_L g15263 ( 
.A(n_15228),
.B(n_3044),
.Y(n_15263)
);

OAI322xp33_ASAP7_75t_L g15264 ( 
.A1(n_15255),
.A2(n_3052),
.A3(n_3051),
.B1(n_3049),
.B2(n_3047),
.C1(n_3048),
.C2(n_3050),
.Y(n_15264)
);

AOI22xp5_ASAP7_75t_L g15265 ( 
.A1(n_15184),
.A2(n_3049),
.B1(n_3047),
.B2(n_3048),
.Y(n_15265)
);

OAI22xp5_ASAP7_75t_L g15266 ( 
.A1(n_15249),
.A2(n_3052),
.B1(n_3050),
.B2(n_3051),
.Y(n_15266)
);

OA21x2_ASAP7_75t_L g15267 ( 
.A1(n_15194),
.A2(n_15178),
.B(n_15230),
.Y(n_15267)
);

NAND2xp5_ASAP7_75t_SL g15268 ( 
.A(n_15185),
.B(n_3053),
.Y(n_15268)
);

NOR3xp33_ASAP7_75t_L g15269 ( 
.A(n_15193),
.B(n_3053),
.C(n_3054),
.Y(n_15269)
);

NOR3xp33_ASAP7_75t_L g15270 ( 
.A(n_15222),
.B(n_3054),
.C(n_3055),
.Y(n_15270)
);

A2O1A1Ixp33_ASAP7_75t_L g15271 ( 
.A1(n_15218),
.A2(n_3057),
.B(n_3055),
.C(n_3056),
.Y(n_15271)
);

XOR2x2_ASAP7_75t_L g15272 ( 
.A(n_15250),
.B(n_15160),
.Y(n_15272)
);

AND2x2_ASAP7_75t_L g15273 ( 
.A(n_15176),
.B(n_3056),
.Y(n_15273)
);

NAND2xp5_ASAP7_75t_L g15274 ( 
.A(n_15165),
.B(n_3058),
.Y(n_15274)
);

OAI21xp5_ASAP7_75t_L g15275 ( 
.A1(n_15183),
.A2(n_3058),
.B(n_3059),
.Y(n_15275)
);

INVx2_ASAP7_75t_L g15276 ( 
.A(n_15225),
.Y(n_15276)
);

INVx1_ASAP7_75t_L g15277 ( 
.A(n_15235),
.Y(n_15277)
);

NAND2xp5_ASAP7_75t_L g15278 ( 
.A(n_15158),
.B(n_3059),
.Y(n_15278)
);

AOI21xp5_ASAP7_75t_L g15279 ( 
.A1(n_15157),
.A2(n_3060),
.B(n_3062),
.Y(n_15279)
);

AOI221xp5_ASAP7_75t_L g15280 ( 
.A1(n_15163),
.A2(n_3065),
.B1(n_3060),
.B2(n_3063),
.C(n_3066),
.Y(n_15280)
);

INVx1_ASAP7_75t_L g15281 ( 
.A(n_15233),
.Y(n_15281)
);

NAND4xp25_ASAP7_75t_SL g15282 ( 
.A(n_15169),
.B(n_3066),
.C(n_3063),
.D(n_3065),
.Y(n_15282)
);

NOR2xp33_ASAP7_75t_L g15283 ( 
.A(n_15224),
.B(n_3067),
.Y(n_15283)
);

OAI22xp5_ASAP7_75t_L g15284 ( 
.A1(n_15220),
.A2(n_3069),
.B1(n_3067),
.B2(n_3068),
.Y(n_15284)
);

AOI221x1_ASAP7_75t_L g15285 ( 
.A1(n_15196),
.A2(n_3070),
.B1(n_3068),
.B2(n_3069),
.C(n_3071),
.Y(n_15285)
);

AOI211xp5_ASAP7_75t_L g15286 ( 
.A1(n_15159),
.A2(n_3073),
.B(n_3071),
.C(n_3072),
.Y(n_15286)
);

A2O1A1Ixp33_ASAP7_75t_L g15287 ( 
.A1(n_15166),
.A2(n_3075),
.B(n_3072),
.C(n_3074),
.Y(n_15287)
);

OAI21xp5_ASAP7_75t_SL g15288 ( 
.A1(n_15175),
.A2(n_3074),
.B(n_3076),
.Y(n_15288)
);

AOI211xp5_ASAP7_75t_L g15289 ( 
.A1(n_15180),
.A2(n_3078),
.B(n_3076),
.C(n_3077),
.Y(n_15289)
);

AOI21xp33_ASAP7_75t_SL g15290 ( 
.A1(n_15212),
.A2(n_3077),
.B(n_3078),
.Y(n_15290)
);

NAND3xp33_ASAP7_75t_L g15291 ( 
.A(n_15182),
.B(n_3079),
.C(n_3080),
.Y(n_15291)
);

NAND2xp5_ASAP7_75t_L g15292 ( 
.A(n_15246),
.B(n_3079),
.Y(n_15292)
);

OAI21xp33_ASAP7_75t_L g15293 ( 
.A1(n_15232),
.A2(n_3081),
.B(n_3082),
.Y(n_15293)
);

OAI211xp5_ASAP7_75t_SL g15294 ( 
.A1(n_15231),
.A2(n_3083),
.B(n_3081),
.C(n_3082),
.Y(n_15294)
);

AOI221xp5_ASAP7_75t_L g15295 ( 
.A1(n_15167),
.A2(n_3085),
.B1(n_3083),
.B2(n_3084),
.C(n_3086),
.Y(n_15295)
);

OAI21xp33_ASAP7_75t_L g15296 ( 
.A1(n_15247),
.A2(n_3084),
.B(n_3085),
.Y(n_15296)
);

INVx1_ASAP7_75t_L g15297 ( 
.A(n_15201),
.Y(n_15297)
);

NOR3xp33_ASAP7_75t_L g15298 ( 
.A(n_15173),
.B(n_3087),
.C(n_3088),
.Y(n_15298)
);

AOI222xp33_ASAP7_75t_L g15299 ( 
.A1(n_15215),
.A2(n_3089),
.B1(n_3091),
.B2(n_3087),
.C1(n_3088),
.C2(n_3090),
.Y(n_15299)
);

INVx1_ASAP7_75t_L g15300 ( 
.A(n_15253),
.Y(n_15300)
);

OAI221xp5_ASAP7_75t_L g15301 ( 
.A1(n_15162),
.A2(n_15252),
.B1(n_15251),
.B2(n_15181),
.C(n_15168),
.Y(n_15301)
);

AOI22xp5_ASAP7_75t_L g15302 ( 
.A1(n_15200),
.A2(n_3092),
.B1(n_3089),
.B2(n_3091),
.Y(n_15302)
);

NOR3xp33_ASAP7_75t_SL g15303 ( 
.A(n_15245),
.B(n_3092),
.C(n_3093),
.Y(n_15303)
);

OAI211xp5_ASAP7_75t_L g15304 ( 
.A1(n_15172),
.A2(n_3095),
.B(n_3093),
.C(n_3094),
.Y(n_15304)
);

NOR3xp33_ASAP7_75t_L g15305 ( 
.A(n_15209),
.B(n_3094),
.C(n_3095),
.Y(n_15305)
);

AOI221xp5_ASAP7_75t_L g15306 ( 
.A1(n_15188),
.A2(n_3098),
.B1(n_3096),
.B2(n_3097),
.C(n_3099),
.Y(n_15306)
);

AOI22xp5_ASAP7_75t_L g15307 ( 
.A1(n_15243),
.A2(n_3098),
.B1(n_3096),
.B2(n_3097),
.Y(n_15307)
);

XOR2xp5_ASAP7_75t_L g15308 ( 
.A(n_15202),
.B(n_4080),
.Y(n_15308)
);

NOR4xp25_ASAP7_75t_L g15309 ( 
.A(n_15229),
.B(n_4090),
.C(n_4081),
.D(n_3102),
.Y(n_15309)
);

NAND3xp33_ASAP7_75t_L g15310 ( 
.A(n_15239),
.B(n_15174),
.C(n_15198),
.Y(n_15310)
);

NOR2xp33_ASAP7_75t_L g15311 ( 
.A(n_15197),
.B(n_3100),
.Y(n_15311)
);

O2A1O1Ixp33_ASAP7_75t_L g15312 ( 
.A1(n_15219),
.A2(n_3102),
.B(n_3100),
.C(n_3101),
.Y(n_15312)
);

NAND2xp5_ASAP7_75t_SL g15313 ( 
.A(n_15203),
.B(n_3101),
.Y(n_15313)
);

NOR3xp33_ASAP7_75t_L g15314 ( 
.A(n_15155),
.B(n_3103),
.C(n_3104),
.Y(n_15314)
);

AOI321xp33_ASAP7_75t_L g15315 ( 
.A1(n_15164),
.A2(n_3129),
.A3(n_3112),
.B1(n_3137),
.B2(n_3121),
.C(n_3103),
.Y(n_15315)
);

AOI22xp5_ASAP7_75t_L g15316 ( 
.A1(n_15171),
.A2(n_3107),
.B1(n_3105),
.B2(n_3106),
.Y(n_15316)
);

NOR2xp67_ASAP7_75t_L g15317 ( 
.A(n_15242),
.B(n_15223),
.Y(n_15317)
);

AOI221xp5_ASAP7_75t_L g15318 ( 
.A1(n_15248),
.A2(n_3109),
.B1(n_3107),
.B2(n_3108),
.C(n_3110),
.Y(n_15318)
);

AOI221xp5_ASAP7_75t_L g15319 ( 
.A1(n_15208),
.A2(n_3112),
.B1(n_3109),
.B2(n_3111),
.C(n_3113),
.Y(n_15319)
);

AND2x2_ASAP7_75t_L g15320 ( 
.A(n_15227),
.B(n_3113),
.Y(n_15320)
);

OAI21xp33_ASAP7_75t_SL g15321 ( 
.A1(n_15216),
.A2(n_3111),
.B(n_3114),
.Y(n_15321)
);

NOR3xp33_ASAP7_75t_L g15322 ( 
.A(n_15179),
.B(n_15244),
.C(n_15170),
.Y(n_15322)
);

AOI221xp5_ASAP7_75t_L g15323 ( 
.A1(n_15206),
.A2(n_3117),
.B1(n_3114),
.B2(n_3115),
.C(n_3118),
.Y(n_15323)
);

AND2x2_ASAP7_75t_L g15324 ( 
.A(n_15161),
.B(n_3118),
.Y(n_15324)
);

O2A1O1Ixp5_ASAP7_75t_SL g15325 ( 
.A1(n_15204),
.A2(n_3120),
.B(n_3117),
.C(n_3119),
.Y(n_15325)
);

AOI21xp5_ASAP7_75t_L g15326 ( 
.A1(n_15214),
.A2(n_3120),
.B(n_3121),
.Y(n_15326)
);

INVx1_ASAP7_75t_L g15327 ( 
.A(n_15186),
.Y(n_15327)
);

AOI21xp5_ASAP7_75t_L g15328 ( 
.A1(n_15236),
.A2(n_3122),
.B(n_3123),
.Y(n_15328)
);

INVx1_ASAP7_75t_L g15329 ( 
.A(n_15154),
.Y(n_15329)
);

OAI21xp33_ASAP7_75t_L g15330 ( 
.A1(n_15217),
.A2(n_3122),
.B(n_3123),
.Y(n_15330)
);

NAND2xp5_ASAP7_75t_L g15331 ( 
.A(n_15207),
.B(n_3124),
.Y(n_15331)
);

AOI221x1_ASAP7_75t_L g15332 ( 
.A1(n_15240),
.A2(n_3126),
.B1(n_3124),
.B2(n_3125),
.C(n_3127),
.Y(n_15332)
);

XNOR2xp5_ASAP7_75t_L g15333 ( 
.A(n_15189),
.B(n_3126),
.Y(n_15333)
);

AOI222xp33_ASAP7_75t_L g15334 ( 
.A1(n_15238),
.A2(n_3129),
.B1(n_3131),
.B2(n_3125),
.C1(n_3128),
.C2(n_3130),
.Y(n_15334)
);

NAND4xp75_ASAP7_75t_L g15335 ( 
.A(n_15210),
.B(n_15213),
.C(n_15237),
.D(n_15254),
.Y(n_15335)
);

AOI211xp5_ASAP7_75t_L g15336 ( 
.A1(n_15226),
.A2(n_3131),
.B(n_3128),
.C(n_3130),
.Y(n_15336)
);

AOI21xp33_ASAP7_75t_L g15337 ( 
.A1(n_15211),
.A2(n_3132),
.B(n_3133),
.Y(n_15337)
);

AOI22xp33_ASAP7_75t_SL g15338 ( 
.A1(n_15234),
.A2(n_3135),
.B1(n_3133),
.B2(n_3134),
.Y(n_15338)
);

INVx1_ASAP7_75t_SL g15339 ( 
.A(n_15192),
.Y(n_15339)
);

INVx1_ASAP7_75t_L g15340 ( 
.A(n_15199),
.Y(n_15340)
);

AOI221x1_ASAP7_75t_L g15341 ( 
.A1(n_15241),
.A2(n_3136),
.B1(n_3134),
.B2(n_3135),
.C(n_3138),
.Y(n_15341)
);

NAND2xp5_ASAP7_75t_L g15342 ( 
.A(n_15177),
.B(n_3136),
.Y(n_15342)
);

A2O1A1Ixp33_ASAP7_75t_L g15343 ( 
.A1(n_15218),
.A2(n_3140),
.B(n_3138),
.C(n_3139),
.Y(n_15343)
);

INVxp67_ASAP7_75t_L g15344 ( 
.A(n_15202),
.Y(n_15344)
);

OAI21xp33_ASAP7_75t_L g15345 ( 
.A1(n_15156),
.A2(n_3139),
.B(n_3140),
.Y(n_15345)
);

OAI21xp33_ASAP7_75t_L g15346 ( 
.A1(n_15156),
.A2(n_3141),
.B(n_3142),
.Y(n_15346)
);

NOR2xp33_ASAP7_75t_L g15347 ( 
.A(n_15255),
.B(n_3142),
.Y(n_15347)
);

AND2x2_ASAP7_75t_L g15348 ( 
.A(n_15176),
.B(n_3144),
.Y(n_15348)
);

INVxp67_ASAP7_75t_SL g15349 ( 
.A(n_15202),
.Y(n_15349)
);

AOI21xp5_ASAP7_75t_L g15350 ( 
.A1(n_15156),
.A2(n_3143),
.B(n_3144),
.Y(n_15350)
);

HB1xp67_ASAP7_75t_L g15351 ( 
.A(n_15233),
.Y(n_15351)
);

AOI22x1_ASAP7_75t_L g15352 ( 
.A1(n_15169),
.A2(n_3146),
.B1(n_3143),
.B2(n_3145),
.Y(n_15352)
);

NAND2xp5_ASAP7_75t_L g15353 ( 
.A(n_15273),
.B(n_3145),
.Y(n_15353)
);

AND2x2_ASAP7_75t_L g15354 ( 
.A(n_15349),
.B(n_15344),
.Y(n_15354)
);

NOR2xp67_ASAP7_75t_L g15355 ( 
.A(n_15282),
.B(n_3147),
.Y(n_15355)
);

OAI322xp33_ASAP7_75t_L g15356 ( 
.A1(n_15308),
.A2(n_3152),
.A3(n_3151),
.B1(n_3149),
.B2(n_3146),
.C1(n_3148),
.C2(n_3150),
.Y(n_15356)
);

AOI322xp5_ASAP7_75t_L g15357 ( 
.A1(n_15339),
.A2(n_3153),
.A3(n_3152),
.B1(n_3150),
.B2(n_3148),
.C1(n_3149),
.C2(n_3151),
.Y(n_15357)
);

NAND4xp25_ASAP7_75t_L g15358 ( 
.A(n_15299),
.B(n_3156),
.C(n_3154),
.D(n_3155),
.Y(n_15358)
);

AOI21xp5_ASAP7_75t_L g15359 ( 
.A1(n_15351),
.A2(n_3154),
.B(n_3156),
.Y(n_15359)
);

NAND3xp33_ASAP7_75t_L g15360 ( 
.A(n_15270),
.B(n_3157),
.C(n_3158),
.Y(n_15360)
);

INVx1_ASAP7_75t_L g15361 ( 
.A(n_15348),
.Y(n_15361)
);

INVx1_ASAP7_75t_L g15362 ( 
.A(n_15263),
.Y(n_15362)
);

INVx2_ASAP7_75t_SL g15363 ( 
.A(n_15324),
.Y(n_15363)
);

AOI221xp5_ASAP7_75t_L g15364 ( 
.A1(n_15290),
.A2(n_3159),
.B1(n_3157),
.B2(n_3158),
.C(n_3160),
.Y(n_15364)
);

NAND2xp5_ASAP7_75t_L g15365 ( 
.A(n_15305),
.B(n_3159),
.Y(n_15365)
);

NOR2xp33_ASAP7_75t_L g15366 ( 
.A(n_15294),
.B(n_3160),
.Y(n_15366)
);

NAND4xp25_ASAP7_75t_L g15367 ( 
.A(n_15341),
.B(n_3163),
.C(n_3161),
.D(n_3162),
.Y(n_15367)
);

NAND3xp33_ASAP7_75t_L g15368 ( 
.A(n_15269),
.B(n_3161),
.C(n_3163),
.Y(n_15368)
);

NAND2xp5_ASAP7_75t_L g15369 ( 
.A(n_15314),
.B(n_3164),
.Y(n_15369)
);

NAND4xp25_ASAP7_75t_L g15370 ( 
.A(n_15322),
.B(n_3166),
.C(n_3164),
.D(n_3165),
.Y(n_15370)
);

INVx1_ASAP7_75t_L g15371 ( 
.A(n_15352),
.Y(n_15371)
);

NAND2xp5_ASAP7_75t_L g15372 ( 
.A(n_15262),
.B(n_3166),
.Y(n_15372)
);

AO22x2_ASAP7_75t_L g15373 ( 
.A1(n_15281),
.A2(n_3169),
.B1(n_3167),
.B2(n_3168),
.Y(n_15373)
);

NAND2xp5_ASAP7_75t_SL g15374 ( 
.A(n_15309),
.B(n_3167),
.Y(n_15374)
);

AOI22xp5_ASAP7_75t_L g15375 ( 
.A1(n_15296),
.A2(n_3170),
.B1(n_3168),
.B2(n_3169),
.Y(n_15375)
);

NOR2xp33_ASAP7_75t_L g15376 ( 
.A(n_15345),
.B(n_3170),
.Y(n_15376)
);

AOI31xp33_ASAP7_75t_L g15377 ( 
.A1(n_15277),
.A2(n_15347),
.A3(n_15286),
.B(n_15336),
.Y(n_15377)
);

NAND2xp5_ASAP7_75t_L g15378 ( 
.A(n_15330),
.B(n_15279),
.Y(n_15378)
);

INVx1_ASAP7_75t_L g15379 ( 
.A(n_15256),
.Y(n_15379)
);

INVx1_ASAP7_75t_L g15380 ( 
.A(n_15320),
.Y(n_15380)
);

AOI221xp5_ASAP7_75t_L g15381 ( 
.A1(n_15337),
.A2(n_15293),
.B1(n_15301),
.B2(n_15259),
.C(n_15280),
.Y(n_15381)
);

NAND2xp5_ASAP7_75t_SL g15382 ( 
.A(n_15306),
.B(n_3171),
.Y(n_15382)
);

NAND2xp5_ASAP7_75t_L g15383 ( 
.A(n_15338),
.B(n_15302),
.Y(n_15383)
);

INVx1_ASAP7_75t_L g15384 ( 
.A(n_15274),
.Y(n_15384)
);

INVx2_ASAP7_75t_L g15385 ( 
.A(n_15267),
.Y(n_15385)
);

AOI21xp5_ASAP7_75t_L g15386 ( 
.A1(n_15313),
.A2(n_3171),
.B(n_3172),
.Y(n_15386)
);

AOI21xp5_ASAP7_75t_L g15387 ( 
.A1(n_15261),
.A2(n_3172),
.B(n_3173),
.Y(n_15387)
);

AOI211xp5_ASAP7_75t_L g15388 ( 
.A1(n_15304),
.A2(n_3175),
.B(n_3173),
.C(n_3174),
.Y(n_15388)
);

INVx1_ASAP7_75t_L g15389 ( 
.A(n_15292),
.Y(n_15389)
);

INVx1_ASAP7_75t_L g15390 ( 
.A(n_15346),
.Y(n_15390)
);

NAND3xp33_ASAP7_75t_L g15391 ( 
.A(n_15318),
.B(n_3174),
.C(n_3175),
.Y(n_15391)
);

INVx1_ASAP7_75t_L g15392 ( 
.A(n_15267),
.Y(n_15392)
);

NOR2xp33_ASAP7_75t_L g15393 ( 
.A(n_15321),
.B(n_3176),
.Y(n_15393)
);

INVx1_ASAP7_75t_SL g15394 ( 
.A(n_15335),
.Y(n_15394)
);

NOR3xp33_ASAP7_75t_L g15395 ( 
.A(n_15329),
.B(n_4096),
.C(n_4094),
.Y(n_15395)
);

INVx1_ASAP7_75t_L g15396 ( 
.A(n_15278),
.Y(n_15396)
);

AOI22xp5_ASAP7_75t_L g15397 ( 
.A1(n_15276),
.A2(n_3178),
.B1(n_3176),
.B2(n_3177),
.Y(n_15397)
);

INVx1_ASAP7_75t_L g15398 ( 
.A(n_15333),
.Y(n_15398)
);

NOR2xp33_ASAP7_75t_L g15399 ( 
.A(n_15288),
.B(n_3177),
.Y(n_15399)
);

INVx1_ASAP7_75t_L g15400 ( 
.A(n_15312),
.Y(n_15400)
);

NAND3xp33_ASAP7_75t_L g15401 ( 
.A(n_15258),
.B(n_15323),
.C(n_15334),
.Y(n_15401)
);

NAND3xp33_ASAP7_75t_L g15402 ( 
.A(n_15295),
.B(n_3179),
.C(n_3180),
.Y(n_15402)
);

AOI21xp5_ASAP7_75t_L g15403 ( 
.A1(n_15268),
.A2(n_3179),
.B(n_3181),
.Y(n_15403)
);

NAND3xp33_ASAP7_75t_L g15404 ( 
.A(n_15303),
.B(n_3181),
.C(n_3182),
.Y(n_15404)
);

AND2x4_ASAP7_75t_SL g15405 ( 
.A(n_15300),
.B(n_3182),
.Y(n_15405)
);

AOI22xp33_ASAP7_75t_L g15406 ( 
.A1(n_15311),
.A2(n_3185),
.B1(n_3183),
.B2(n_3184),
.Y(n_15406)
);

NOR2xp33_ASAP7_75t_L g15407 ( 
.A(n_15284),
.B(n_3184),
.Y(n_15407)
);

INVx1_ASAP7_75t_L g15408 ( 
.A(n_15271),
.Y(n_15408)
);

OAI211xp5_ASAP7_75t_L g15409 ( 
.A1(n_15350),
.A2(n_4087),
.B(n_4089),
.C(n_4086),
.Y(n_15409)
);

INVx2_ASAP7_75t_L g15410 ( 
.A(n_15272),
.Y(n_15410)
);

OAI211xp5_ASAP7_75t_L g15411 ( 
.A1(n_15265),
.A2(n_4087),
.B(n_4089),
.C(n_4086),
.Y(n_15411)
);

NOR4xp25_ASAP7_75t_L g15412 ( 
.A(n_15343),
.B(n_3187),
.C(n_3185),
.D(n_3186),
.Y(n_15412)
);

INVx1_ASAP7_75t_SL g15413 ( 
.A(n_15342),
.Y(n_15413)
);

XNOR2xp5_ASAP7_75t_L g15414 ( 
.A(n_15289),
.B(n_4090),
.Y(n_15414)
);

NAND3xp33_ASAP7_75t_L g15415 ( 
.A(n_15298),
.B(n_3186),
.C(n_3187),
.Y(n_15415)
);

NAND2x1_ASAP7_75t_L g15416 ( 
.A(n_15326),
.B(n_3189),
.Y(n_15416)
);

INVx1_ASAP7_75t_L g15417 ( 
.A(n_15331),
.Y(n_15417)
);

INVx1_ASAP7_75t_L g15418 ( 
.A(n_15283),
.Y(n_15418)
);

NOR3xp33_ASAP7_75t_L g15419 ( 
.A(n_15340),
.B(n_4096),
.C(n_4094),
.Y(n_15419)
);

AOI21xp5_ASAP7_75t_L g15420 ( 
.A1(n_15328),
.A2(n_3189),
.B(n_3190),
.Y(n_15420)
);

AOI31xp33_ASAP7_75t_L g15421 ( 
.A1(n_15275),
.A2(n_3192),
.A3(n_3190),
.B(n_3191),
.Y(n_15421)
);

AOI322xp5_ASAP7_75t_L g15422 ( 
.A1(n_15327),
.A2(n_3196),
.A3(n_3195),
.B1(n_3193),
.B2(n_3191),
.C1(n_3192),
.C2(n_3194),
.Y(n_15422)
);

NOR3xp33_ASAP7_75t_L g15423 ( 
.A(n_15297),
.B(n_4079),
.C(n_4078),
.Y(n_15423)
);

NAND2xp5_ASAP7_75t_L g15424 ( 
.A(n_15260),
.B(n_3193),
.Y(n_15424)
);

AOI211xp5_ASAP7_75t_L g15425 ( 
.A1(n_15266),
.A2(n_3198),
.B(n_3195),
.C(n_3197),
.Y(n_15425)
);

INVx1_ASAP7_75t_L g15426 ( 
.A(n_15332),
.Y(n_15426)
);

INVxp67_ASAP7_75t_SL g15427 ( 
.A(n_15307),
.Y(n_15427)
);

INVx1_ASAP7_75t_L g15428 ( 
.A(n_15315),
.Y(n_15428)
);

AOI221x1_ASAP7_75t_L g15429 ( 
.A1(n_15287),
.A2(n_3200),
.B1(n_3197),
.B2(n_3199),
.C(n_3201),
.Y(n_15429)
);

INVx1_ASAP7_75t_L g15430 ( 
.A(n_15285),
.Y(n_15430)
);

OA22x2_ASAP7_75t_L g15431 ( 
.A1(n_15316),
.A2(n_3201),
.B1(n_3199),
.B2(n_3200),
.Y(n_15431)
);

NAND2xp5_ASAP7_75t_L g15432 ( 
.A(n_15257),
.B(n_3202),
.Y(n_15432)
);

NAND3xp33_ASAP7_75t_L g15433 ( 
.A(n_15319),
.B(n_3202),
.C(n_3203),
.Y(n_15433)
);

NAND2xp5_ASAP7_75t_SL g15434 ( 
.A(n_15291),
.B(n_3204),
.Y(n_15434)
);

OA22x2_ASAP7_75t_L g15435 ( 
.A1(n_15325),
.A2(n_3206),
.B1(n_3204),
.B2(n_3205),
.Y(n_15435)
);

INVxp67_ASAP7_75t_SL g15436 ( 
.A(n_15317),
.Y(n_15436)
);

NOR3xp33_ASAP7_75t_L g15437 ( 
.A(n_15310),
.B(n_15264),
.C(n_3205),
.Y(n_15437)
);

XNOR2xp5_ASAP7_75t_L g15438 ( 
.A(n_15308),
.B(n_4071),
.Y(n_15438)
);

INVx1_ASAP7_75t_L g15439 ( 
.A(n_15308),
.Y(n_15439)
);

INVx1_ASAP7_75t_L g15440 ( 
.A(n_15308),
.Y(n_15440)
);

INVx1_ASAP7_75t_L g15441 ( 
.A(n_15308),
.Y(n_15441)
);

NAND3xp33_ASAP7_75t_L g15442 ( 
.A(n_15299),
.B(n_3206),
.C(n_3208),
.Y(n_15442)
);

OAI311xp33_ASAP7_75t_L g15443 ( 
.A1(n_15301),
.A2(n_3211),
.A3(n_3209),
.B1(n_3210),
.C1(n_3212),
.Y(n_15443)
);

NOR2x1_ASAP7_75t_L g15444 ( 
.A(n_15282),
.B(n_3209),
.Y(n_15444)
);

NOR2xp33_ASAP7_75t_L g15445 ( 
.A(n_15294),
.B(n_3211),
.Y(n_15445)
);

NOR3xp33_ASAP7_75t_SL g15446 ( 
.A(n_15282),
.B(n_3212),
.C(n_3213),
.Y(n_15446)
);

NAND4xp25_ASAP7_75t_L g15447 ( 
.A(n_15299),
.B(n_3215),
.C(n_3213),
.D(n_3214),
.Y(n_15447)
);

NAND2xp5_ASAP7_75t_L g15448 ( 
.A(n_15273),
.B(n_3215),
.Y(n_15448)
);

NAND4xp75_ASAP7_75t_L g15449 ( 
.A(n_15267),
.B(n_3219),
.C(n_3216),
.D(n_3218),
.Y(n_15449)
);

NOR3xp33_ASAP7_75t_L g15450 ( 
.A(n_15282),
.B(n_4093),
.C(n_4092),
.Y(n_15450)
);

AOI221x1_ASAP7_75t_SL g15451 ( 
.A1(n_15355),
.A2(n_3221),
.B1(n_3219),
.B2(n_3220),
.C(n_3222),
.Y(n_15451)
);

NAND3xp33_ASAP7_75t_L g15452 ( 
.A(n_15419),
.B(n_3221),
.C(n_3222),
.Y(n_15452)
);

NAND3xp33_ASAP7_75t_SL g15453 ( 
.A(n_15394),
.B(n_3223),
.C(n_3224),
.Y(n_15453)
);

NOR2xp33_ASAP7_75t_L g15454 ( 
.A(n_15358),
.B(n_15447),
.Y(n_15454)
);

NOR2x1_ASAP7_75t_SL g15455 ( 
.A(n_15449),
.B(n_3223),
.Y(n_15455)
);

AOI21xp5_ASAP7_75t_L g15456 ( 
.A1(n_15416),
.A2(n_3224),
.B(n_3225),
.Y(n_15456)
);

INVx1_ASAP7_75t_L g15457 ( 
.A(n_15435),
.Y(n_15457)
);

NAND2xp5_ASAP7_75t_L g15458 ( 
.A(n_15405),
.B(n_3225),
.Y(n_15458)
);

INVx1_ASAP7_75t_L g15459 ( 
.A(n_15438),
.Y(n_15459)
);

NAND3xp33_ASAP7_75t_L g15460 ( 
.A(n_15406),
.B(n_3226),
.C(n_3227),
.Y(n_15460)
);

AOI22xp33_ASAP7_75t_L g15461 ( 
.A1(n_15450),
.A2(n_3229),
.B1(n_3227),
.B2(n_3228),
.Y(n_15461)
);

NAND4xp25_ASAP7_75t_L g15462 ( 
.A(n_15381),
.B(n_3230),
.C(n_3228),
.D(n_3229),
.Y(n_15462)
);

NAND4xp25_ASAP7_75t_L g15463 ( 
.A(n_15388),
.B(n_3232),
.C(n_3230),
.D(n_3231),
.Y(n_15463)
);

NAND3xp33_ASAP7_75t_L g15464 ( 
.A(n_15364),
.B(n_3231),
.C(n_3232),
.Y(n_15464)
);

OAI211xp5_ASAP7_75t_SL g15465 ( 
.A1(n_15432),
.A2(n_15428),
.B(n_15371),
.C(n_15426),
.Y(n_15465)
);

NAND2xp5_ASAP7_75t_L g15466 ( 
.A(n_15357),
.B(n_3233),
.Y(n_15466)
);

NOR2xp33_ASAP7_75t_L g15467 ( 
.A(n_15421),
.B(n_3233),
.Y(n_15467)
);

NOR3xp33_ASAP7_75t_L g15468 ( 
.A(n_15377),
.B(n_3234),
.C(n_3235),
.Y(n_15468)
);

INVx1_ASAP7_75t_L g15469 ( 
.A(n_15353),
.Y(n_15469)
);

NOR3xp33_ASAP7_75t_L g15470 ( 
.A(n_15436),
.B(n_3234),
.C(n_3235),
.Y(n_15470)
);

AOI221xp5_ASAP7_75t_L g15471 ( 
.A1(n_15412),
.A2(n_3238),
.B1(n_3236),
.B2(n_3237),
.C(n_3239),
.Y(n_15471)
);

CKINVDCx5p33_ASAP7_75t_R g15472 ( 
.A(n_15354),
.Y(n_15472)
);

NAND4xp25_ASAP7_75t_L g15473 ( 
.A(n_15366),
.B(n_3239),
.C(n_3236),
.D(n_3237),
.Y(n_15473)
);

NOR2x1_ASAP7_75t_L g15474 ( 
.A(n_15392),
.B(n_3240),
.Y(n_15474)
);

NAND2xp5_ASAP7_75t_SL g15475 ( 
.A(n_15375),
.B(n_15430),
.Y(n_15475)
);

NAND3xp33_ASAP7_75t_L g15476 ( 
.A(n_15437),
.B(n_3240),
.C(n_3241),
.Y(n_15476)
);

AOI211xp5_ASAP7_75t_L g15477 ( 
.A1(n_15409),
.A2(n_15411),
.B(n_15367),
.C(n_15443),
.Y(n_15477)
);

NAND2xp33_ASAP7_75t_L g15478 ( 
.A(n_15395),
.B(n_3242),
.Y(n_15478)
);

NOR2xp67_ASAP7_75t_L g15479 ( 
.A(n_15370),
.B(n_3242),
.Y(n_15479)
);

NOR2xp33_ASAP7_75t_L g15480 ( 
.A(n_15448),
.B(n_3243),
.Y(n_15480)
);

NOR2xp33_ASAP7_75t_L g15481 ( 
.A(n_15372),
.B(n_3243),
.Y(n_15481)
);

AOI221xp5_ASAP7_75t_L g15482 ( 
.A1(n_15445),
.A2(n_3247),
.B1(n_3245),
.B2(n_3246),
.C(n_3248),
.Y(n_15482)
);

OAI211xp5_ASAP7_75t_SL g15483 ( 
.A1(n_15446),
.A2(n_3249),
.B(n_3246),
.C(n_3248),
.Y(n_15483)
);

NOR3xp33_ASAP7_75t_L g15484 ( 
.A(n_15410),
.B(n_3249),
.C(n_3250),
.Y(n_15484)
);

INVx1_ASAP7_75t_L g15485 ( 
.A(n_15431),
.Y(n_15485)
);

HB1xp67_ASAP7_75t_L g15486 ( 
.A(n_15444),
.Y(n_15486)
);

NAND3xp33_ASAP7_75t_L g15487 ( 
.A(n_15425),
.B(n_3251),
.C(n_3252),
.Y(n_15487)
);

INVx1_ASAP7_75t_L g15488 ( 
.A(n_15365),
.Y(n_15488)
);

INVx1_ASAP7_75t_L g15489 ( 
.A(n_15393),
.Y(n_15489)
);

NAND2xp5_ASAP7_75t_L g15490 ( 
.A(n_15359),
.B(n_3251),
.Y(n_15490)
);

NOR2xp33_ASAP7_75t_L g15491 ( 
.A(n_15404),
.B(n_3252),
.Y(n_15491)
);

NOR3xp33_ASAP7_75t_L g15492 ( 
.A(n_15439),
.B(n_3253),
.C(n_3254),
.Y(n_15492)
);

NOR2x1_ASAP7_75t_L g15493 ( 
.A(n_15385),
.B(n_3255),
.Y(n_15493)
);

INVx1_ASAP7_75t_L g15494 ( 
.A(n_15369),
.Y(n_15494)
);

OAI211xp5_ASAP7_75t_SL g15495 ( 
.A1(n_15403),
.A2(n_15434),
.B(n_15441),
.C(n_15440),
.Y(n_15495)
);

NAND2xp5_ASAP7_75t_L g15496 ( 
.A(n_15423),
.B(n_3255),
.Y(n_15496)
);

NAND2xp5_ASAP7_75t_SL g15497 ( 
.A(n_15360),
.B(n_3256),
.Y(n_15497)
);

AOI21xp5_ASAP7_75t_L g15498 ( 
.A1(n_15374),
.A2(n_3256),
.B(n_3257),
.Y(n_15498)
);

NOR3x1_ASAP7_75t_L g15499 ( 
.A(n_15415),
.B(n_3258),
.C(n_3259),
.Y(n_15499)
);

OR2x2_ASAP7_75t_L g15500 ( 
.A(n_15368),
.B(n_4074),
.Y(n_15500)
);

A2O1A1Ixp33_ASAP7_75t_L g15501 ( 
.A1(n_15376),
.A2(n_3260),
.B(n_3258),
.C(n_3259),
.Y(n_15501)
);

NAND2xp5_ASAP7_75t_SL g15502 ( 
.A(n_15442),
.B(n_3260),
.Y(n_15502)
);

INVx1_ASAP7_75t_L g15503 ( 
.A(n_15414),
.Y(n_15503)
);

OAI21xp33_ASAP7_75t_L g15504 ( 
.A1(n_15399),
.A2(n_3261),
.B(n_3263),
.Y(n_15504)
);

HB1xp67_ASAP7_75t_L g15505 ( 
.A(n_15373),
.Y(n_15505)
);

AOI21xp5_ASAP7_75t_L g15506 ( 
.A1(n_15382),
.A2(n_15420),
.B(n_15387),
.Y(n_15506)
);

NOR3x1_ASAP7_75t_L g15507 ( 
.A(n_15433),
.B(n_3261),
.C(n_3263),
.Y(n_15507)
);

INVx1_ASAP7_75t_L g15508 ( 
.A(n_15424),
.Y(n_15508)
);

NAND3xp33_ASAP7_75t_L g15509 ( 
.A(n_15386),
.B(n_3264),
.C(n_3266),
.Y(n_15509)
);

AOI21xp5_ASAP7_75t_L g15510 ( 
.A1(n_15383),
.A2(n_3264),
.B(n_3266),
.Y(n_15510)
);

AOI322xp5_ASAP7_75t_L g15511 ( 
.A1(n_15407),
.A2(n_3273),
.A3(n_3272),
.B1(n_3270),
.B2(n_3267),
.C1(n_3269),
.C2(n_3271),
.Y(n_15511)
);

OAI21xp33_ASAP7_75t_SL g15512 ( 
.A1(n_15363),
.A2(n_3267),
.B(n_3271),
.Y(n_15512)
);

INVx1_ASAP7_75t_L g15513 ( 
.A(n_15373),
.Y(n_15513)
);

INVx1_ASAP7_75t_L g15514 ( 
.A(n_15361),
.Y(n_15514)
);

NAND4xp25_ASAP7_75t_L g15515 ( 
.A(n_15401),
.B(n_15429),
.C(n_15391),
.D(n_15402),
.Y(n_15515)
);

NOR2xp33_ASAP7_75t_L g15516 ( 
.A(n_15380),
.B(n_3272),
.Y(n_15516)
);

NOR2xp33_ASAP7_75t_L g15517 ( 
.A(n_15356),
.B(n_3274),
.Y(n_15517)
);

INVx2_ASAP7_75t_L g15518 ( 
.A(n_15362),
.Y(n_15518)
);

INVxp67_ASAP7_75t_L g15519 ( 
.A(n_15397),
.Y(n_15519)
);

AOI21xp5_ASAP7_75t_L g15520 ( 
.A1(n_15378),
.A2(n_3275),
.B(n_3276),
.Y(n_15520)
);

INVx1_ASAP7_75t_L g15521 ( 
.A(n_15408),
.Y(n_15521)
);

NOR3xp33_ASAP7_75t_SL g15522 ( 
.A(n_15400),
.B(n_3275),
.C(n_3276),
.Y(n_15522)
);

A2O1A1Ixp33_ASAP7_75t_L g15523 ( 
.A1(n_15390),
.A2(n_3279),
.B(n_3277),
.C(n_3278),
.Y(n_15523)
);

AND2x2_ASAP7_75t_L g15524 ( 
.A(n_15427),
.B(n_3277),
.Y(n_15524)
);

NOR3x1_ASAP7_75t_L g15525 ( 
.A(n_15398),
.B(n_3278),
.C(n_3279),
.Y(n_15525)
);

NOR3xp33_ASAP7_75t_SL g15526 ( 
.A(n_15384),
.B(n_3280),
.C(n_3281),
.Y(n_15526)
);

AND2x2_ASAP7_75t_L g15527 ( 
.A(n_15413),
.B(n_3281),
.Y(n_15527)
);

NAND2xp5_ASAP7_75t_L g15528 ( 
.A(n_15379),
.B(n_3282),
.Y(n_15528)
);

AOI21xp33_ASAP7_75t_L g15529 ( 
.A1(n_15389),
.A2(n_3283),
.B(n_3284),
.Y(n_15529)
);

INVx1_ASAP7_75t_L g15530 ( 
.A(n_15418),
.Y(n_15530)
);

INVx2_ASAP7_75t_SL g15531 ( 
.A(n_15417),
.Y(n_15531)
);

CKINVDCx6p67_ASAP7_75t_R g15532 ( 
.A(n_15396),
.Y(n_15532)
);

INVx1_ASAP7_75t_L g15533 ( 
.A(n_15422),
.Y(n_15533)
);

NOR2xp67_ASAP7_75t_L g15534 ( 
.A(n_15367),
.B(n_3283),
.Y(n_15534)
);

OAI321xp33_ASAP7_75t_L g15535 ( 
.A1(n_15367),
.A2(n_3286),
.A3(n_3288),
.B1(n_3289),
.B2(n_3285),
.C(n_3287),
.Y(n_15535)
);

NAND2xp5_ASAP7_75t_L g15536 ( 
.A(n_15524),
.B(n_4083),
.Y(n_15536)
);

NAND4xp75_ASAP7_75t_L g15537 ( 
.A(n_15493),
.B(n_3286),
.C(n_3284),
.D(n_3285),
.Y(n_15537)
);

NOR3xp33_ASAP7_75t_L g15538 ( 
.A(n_15465),
.B(n_15495),
.C(n_15476),
.Y(n_15538)
);

OA22x2_ASAP7_75t_L g15539 ( 
.A1(n_15472),
.A2(n_3289),
.B1(n_3287),
.B2(n_3288),
.Y(n_15539)
);

NOR2x1_ASAP7_75t_L g15540 ( 
.A(n_15474),
.B(n_15513),
.Y(n_15540)
);

AOI211xp5_ASAP7_75t_L g15541 ( 
.A1(n_15453),
.A2(n_15483),
.B(n_15535),
.C(n_15512),
.Y(n_15541)
);

OAI22xp33_ASAP7_75t_L g15542 ( 
.A1(n_15473),
.A2(n_3294),
.B1(n_3292),
.B2(n_3293),
.Y(n_15542)
);

AND2x2_ASAP7_75t_L g15543 ( 
.A(n_15526),
.B(n_3292),
.Y(n_15543)
);

NOR3xp33_ASAP7_75t_L g15544 ( 
.A(n_15475),
.B(n_3293),
.C(n_3294),
.Y(n_15544)
);

OA22x2_ASAP7_75t_L g15545 ( 
.A1(n_15457),
.A2(n_3297),
.B1(n_3295),
.B2(n_3296),
.Y(n_15545)
);

NOR2x1_ASAP7_75t_L g15546 ( 
.A(n_15462),
.B(n_3295),
.Y(n_15546)
);

AND5x1_ASAP7_75t_L g15547 ( 
.A(n_15454),
.B(n_3299),
.C(n_3296),
.D(n_3297),
.E(n_3300),
.Y(n_15547)
);

NAND2xp5_ASAP7_75t_SL g15548 ( 
.A(n_15482),
.B(n_3300),
.Y(n_15548)
);

INVx1_ASAP7_75t_L g15549 ( 
.A(n_15505),
.Y(n_15549)
);

AND2x2_ASAP7_75t_L g15550 ( 
.A(n_15522),
.B(n_3301),
.Y(n_15550)
);

NOR2x1_ASAP7_75t_L g15551 ( 
.A(n_15458),
.B(n_3301),
.Y(n_15551)
);

NOR2xp67_ASAP7_75t_L g15552 ( 
.A(n_15456),
.B(n_3302),
.Y(n_15552)
);

NAND2xp5_ASAP7_75t_L g15553 ( 
.A(n_15527),
.B(n_4082),
.Y(n_15553)
);

INVx2_ASAP7_75t_L g15554 ( 
.A(n_15525),
.Y(n_15554)
);

NOR3xp33_ASAP7_75t_L g15555 ( 
.A(n_15514),
.B(n_3302),
.C(n_3303),
.Y(n_15555)
);

NOR3x1_ASAP7_75t_L g15556 ( 
.A(n_15452),
.B(n_3303),
.C(n_3304),
.Y(n_15556)
);

NAND2xp5_ASAP7_75t_L g15557 ( 
.A(n_15451),
.B(n_4084),
.Y(n_15557)
);

AND2x4_ASAP7_75t_L g15558 ( 
.A(n_15485),
.B(n_3304),
.Y(n_15558)
);

AOI22xp5_ASAP7_75t_L g15559 ( 
.A1(n_15484),
.A2(n_3307),
.B1(n_3305),
.B2(n_3306),
.Y(n_15559)
);

INVxp33_ASAP7_75t_L g15560 ( 
.A(n_15480),
.Y(n_15560)
);

NOR3xp33_ASAP7_75t_L g15561 ( 
.A(n_15521),
.B(n_3305),
.C(n_3306),
.Y(n_15561)
);

INVx1_ASAP7_75t_L g15562 ( 
.A(n_15455),
.Y(n_15562)
);

NAND4xp75_ASAP7_75t_L g15563 ( 
.A(n_15507),
.B(n_3309),
.C(n_3307),
.D(n_3308),
.Y(n_15563)
);

NAND2xp5_ASAP7_75t_L g15564 ( 
.A(n_15468),
.B(n_4093),
.Y(n_15564)
);

AND3x2_ASAP7_75t_L g15565 ( 
.A(n_15486),
.B(n_15470),
.C(n_15492),
.Y(n_15565)
);

NAND3x1_ASAP7_75t_L g15566 ( 
.A(n_15481),
.B(n_3308),
.C(n_3309),
.Y(n_15566)
);

INVx1_ASAP7_75t_L g15567 ( 
.A(n_15466),
.Y(n_15567)
);

NOR2xp33_ASAP7_75t_SL g15568 ( 
.A(n_15516),
.B(n_3310),
.Y(n_15568)
);

NAND2xp5_ASAP7_75t_SL g15569 ( 
.A(n_15471),
.B(n_3311),
.Y(n_15569)
);

INVx1_ASAP7_75t_L g15570 ( 
.A(n_15490),
.Y(n_15570)
);

INVx1_ASAP7_75t_L g15571 ( 
.A(n_15467),
.Y(n_15571)
);

NOR4xp25_ASAP7_75t_L g15572 ( 
.A(n_15515),
.B(n_3314),
.C(n_3312),
.D(n_3313),
.Y(n_15572)
);

AOI211x1_ASAP7_75t_L g15573 ( 
.A1(n_15498),
.A2(n_3314),
.B(n_3312),
.C(n_3313),
.Y(n_15573)
);

NOR2x1_ASAP7_75t_L g15574 ( 
.A(n_15463),
.B(n_3315),
.Y(n_15574)
);

NOR4xp25_ASAP7_75t_SL g15575 ( 
.A(n_15502),
.B(n_3318),
.C(n_3316),
.D(n_3317),
.Y(n_15575)
);

XNOR2x1_ASAP7_75t_SL g15576 ( 
.A(n_15531),
.B(n_3316),
.Y(n_15576)
);

INVx1_ASAP7_75t_L g15577 ( 
.A(n_15534),
.Y(n_15577)
);

NOR2x1_ASAP7_75t_L g15578 ( 
.A(n_15509),
.B(n_3317),
.Y(n_15578)
);

OA21x2_ASAP7_75t_L g15579 ( 
.A1(n_15530),
.A2(n_3329),
.B(n_3319),
.Y(n_15579)
);

NOR2xp33_ASAP7_75t_L g15580 ( 
.A(n_15504),
.B(n_3319),
.Y(n_15580)
);

NAND3xp33_ASAP7_75t_L g15581 ( 
.A(n_15517),
.B(n_3320),
.C(n_3321),
.Y(n_15581)
);

NOR2xp33_ASAP7_75t_SL g15582 ( 
.A(n_15491),
.B(n_3320),
.Y(n_15582)
);

NOR2xp33_ASAP7_75t_L g15583 ( 
.A(n_15487),
.B(n_3321),
.Y(n_15583)
);

OA22x2_ASAP7_75t_L g15584 ( 
.A1(n_15533),
.A2(n_3325),
.B1(n_3322),
.B2(n_3324),
.Y(n_15584)
);

NOR2xp33_ASAP7_75t_L g15585 ( 
.A(n_15460),
.B(n_3322),
.Y(n_15585)
);

NOR2x1p5_ASAP7_75t_L g15586 ( 
.A(n_15496),
.B(n_3325),
.Y(n_15586)
);

INVx1_ASAP7_75t_L g15587 ( 
.A(n_15500),
.Y(n_15587)
);

NAND2xp5_ASAP7_75t_L g15588 ( 
.A(n_15510),
.B(n_4069),
.Y(n_15588)
);

NAND5xp2_ASAP7_75t_L g15589 ( 
.A(n_15477),
.B(n_4073),
.C(n_4074),
.D(n_4070),
.E(n_4069),
.Y(n_15589)
);

NOR2x1p5_ASAP7_75t_SL g15590 ( 
.A(n_15518),
.B(n_3326),
.Y(n_15590)
);

NAND2xp5_ASAP7_75t_L g15591 ( 
.A(n_15520),
.B(n_4070),
.Y(n_15591)
);

INVx1_ASAP7_75t_L g15592 ( 
.A(n_15528),
.Y(n_15592)
);

NAND2xp5_ASAP7_75t_L g15593 ( 
.A(n_15461),
.B(n_15501),
.Y(n_15593)
);

NOR3x1_ASAP7_75t_L g15594 ( 
.A(n_15464),
.B(n_3326),
.C(n_3327),
.Y(n_15594)
);

OAI22xp5_ASAP7_75t_L g15595 ( 
.A1(n_15479),
.A2(n_15519),
.B1(n_15532),
.B2(n_15459),
.Y(n_15595)
);

AND2x2_ASAP7_75t_L g15596 ( 
.A(n_15499),
.B(n_3329),
.Y(n_15596)
);

NAND4xp25_ASAP7_75t_L g15597 ( 
.A(n_15506),
.B(n_15503),
.C(n_15489),
.D(n_15508),
.Y(n_15597)
);

XNOR2xp5_ASAP7_75t_L g15598 ( 
.A(n_15497),
.B(n_3331),
.Y(n_15598)
);

NOR3xp33_ASAP7_75t_L g15599 ( 
.A(n_15469),
.B(n_3330),
.C(n_3331),
.Y(n_15599)
);

NOR2xp67_ASAP7_75t_L g15600 ( 
.A(n_15488),
.B(n_15494),
.Y(n_15600)
);

NOR2x1_ASAP7_75t_L g15601 ( 
.A(n_15523),
.B(n_3330),
.Y(n_15601)
);

NAND5xp2_ASAP7_75t_L g15602 ( 
.A(n_15511),
.B(n_4083),
.C(n_4084),
.D(n_4082),
.E(n_4081),
.Y(n_15602)
);

INVxp67_ASAP7_75t_L g15603 ( 
.A(n_15478),
.Y(n_15603)
);

NOR3xp33_ASAP7_75t_L g15604 ( 
.A(n_15529),
.B(n_3332),
.C(n_3333),
.Y(n_15604)
);

NAND4xp25_ASAP7_75t_L g15605 ( 
.A(n_15477),
.B(n_3334),
.C(n_3332),
.D(n_3333),
.Y(n_15605)
);

AOI211x1_ASAP7_75t_L g15606 ( 
.A1(n_15498),
.A2(n_3337),
.B(n_3334),
.C(n_3336),
.Y(n_15606)
);

AOI21xp5_ASAP7_75t_L g15607 ( 
.A1(n_15478),
.A2(n_3336),
.B(n_3337),
.Y(n_15607)
);

INVx1_ASAP7_75t_L g15608 ( 
.A(n_15524),
.Y(n_15608)
);

NOR2xp33_ASAP7_75t_L g15609 ( 
.A(n_15483),
.B(n_3338),
.Y(n_15609)
);

NAND3xp33_ASAP7_75t_L g15610 ( 
.A(n_15484),
.B(n_3338),
.C(n_3339),
.Y(n_15610)
);

INVx1_ASAP7_75t_L g15611 ( 
.A(n_15524),
.Y(n_15611)
);

NAND3xp33_ASAP7_75t_L g15612 ( 
.A(n_15484),
.B(n_3339),
.C(n_3340),
.Y(n_15612)
);

INVx2_ASAP7_75t_L g15613 ( 
.A(n_15525),
.Y(n_15613)
);

AO22x2_ASAP7_75t_L g15614 ( 
.A1(n_15513),
.A2(n_4079),
.B1(n_4064),
.B2(n_3343),
.Y(n_15614)
);

NAND2xp5_ASAP7_75t_L g15615 ( 
.A(n_15524),
.B(n_4065),
.Y(n_15615)
);

NAND2xp5_ASAP7_75t_L g15616 ( 
.A(n_15524),
.B(n_4065),
.Y(n_15616)
);

NOR4xp75_ASAP7_75t_L g15617 ( 
.A(n_15475),
.B(n_3344),
.C(n_3340),
.D(n_3342),
.Y(n_15617)
);

NOR2x1_ASAP7_75t_L g15618 ( 
.A(n_15493),
.B(n_3342),
.Y(n_15618)
);

NOR3xp33_ASAP7_75t_L g15619 ( 
.A(n_15465),
.B(n_3344),
.C(n_3345),
.Y(n_15619)
);

OAI21x1_ASAP7_75t_L g15620 ( 
.A1(n_15456),
.A2(n_3345),
.B(n_3346),
.Y(n_15620)
);

NAND4xp75_ASAP7_75t_L g15621 ( 
.A(n_15493),
.B(n_3348),
.C(n_3346),
.D(n_3347),
.Y(n_15621)
);

NOR3xp33_ASAP7_75t_L g15622 ( 
.A(n_15465),
.B(n_3347),
.C(n_3349),
.Y(n_15622)
);

NOR2xp33_ASAP7_75t_SL g15623 ( 
.A(n_15524),
.B(n_3349),
.Y(n_15623)
);

NOR3xp33_ASAP7_75t_L g15624 ( 
.A(n_15465),
.B(n_3350),
.C(n_3351),
.Y(n_15624)
);

NAND2xp5_ASAP7_75t_L g15625 ( 
.A(n_15524),
.B(n_4092),
.Y(n_15625)
);

AO22x2_ASAP7_75t_L g15626 ( 
.A1(n_15549),
.A2(n_3352),
.B1(n_3353),
.B2(n_3351),
.Y(n_15626)
);

INVx1_ASAP7_75t_L g15627 ( 
.A(n_15576),
.Y(n_15627)
);

NOR2x1_ASAP7_75t_L g15628 ( 
.A(n_15618),
.B(n_3354),
.Y(n_15628)
);

NOR3xp33_ASAP7_75t_L g15629 ( 
.A(n_15595),
.B(n_3350),
.C(n_3355),
.Y(n_15629)
);

NOR2x1_ASAP7_75t_L g15630 ( 
.A(n_15537),
.B(n_3356),
.Y(n_15630)
);

NOR3xp33_ASAP7_75t_L g15631 ( 
.A(n_15597),
.B(n_3355),
.C(n_3356),
.Y(n_15631)
);

NAND2xp5_ASAP7_75t_L g15632 ( 
.A(n_15558),
.B(n_3358),
.Y(n_15632)
);

NOR2x1_ASAP7_75t_L g15633 ( 
.A(n_15621),
.B(n_3358),
.Y(n_15633)
);

NOR2xp67_ASAP7_75t_L g15634 ( 
.A(n_15589),
.B(n_3359),
.Y(n_15634)
);

NOR2x1_ASAP7_75t_L g15635 ( 
.A(n_15540),
.B(n_3360),
.Y(n_15635)
);

OAI211xp5_ASAP7_75t_L g15636 ( 
.A1(n_15619),
.A2(n_3362),
.B(n_3363),
.C(n_3360),
.Y(n_15636)
);

NOR3xp33_ASAP7_75t_L g15637 ( 
.A(n_15581),
.B(n_3357),
.C(n_3362),
.Y(n_15637)
);

INVx1_ASAP7_75t_L g15638 ( 
.A(n_15590),
.Y(n_15638)
);

NOR2x1_ASAP7_75t_L g15639 ( 
.A(n_15551),
.B(n_3364),
.Y(n_15639)
);

NOR3xp33_ASAP7_75t_L g15640 ( 
.A(n_15538),
.B(n_3357),
.C(n_3364),
.Y(n_15640)
);

NOR3xp33_ASAP7_75t_SL g15641 ( 
.A(n_15557),
.B(n_3365),
.C(n_3366),
.Y(n_15641)
);

AOI21xp33_ASAP7_75t_SL g15642 ( 
.A1(n_15584),
.A2(n_3366),
.B(n_3367),
.Y(n_15642)
);

NOR2xp33_ASAP7_75t_L g15643 ( 
.A(n_15602),
.B(n_4058),
.Y(n_15643)
);

INVx1_ASAP7_75t_L g15644 ( 
.A(n_15536),
.Y(n_15644)
);

NAND2xp5_ASAP7_75t_L g15645 ( 
.A(n_15558),
.B(n_3369),
.Y(n_15645)
);

NOR2x1_ASAP7_75t_L g15646 ( 
.A(n_15562),
.B(n_3369),
.Y(n_15646)
);

NAND3xp33_ASAP7_75t_SL g15647 ( 
.A(n_15622),
.B(n_3368),
.C(n_3370),
.Y(n_15647)
);

NOR2x1_ASAP7_75t_L g15648 ( 
.A(n_15579),
.B(n_3371),
.Y(n_15648)
);

INVx1_ASAP7_75t_L g15649 ( 
.A(n_15615),
.Y(n_15649)
);

NAND3xp33_ASAP7_75t_SL g15650 ( 
.A(n_15624),
.B(n_3368),
.C(n_3372),
.Y(n_15650)
);

OR2x2_ASAP7_75t_L g15651 ( 
.A(n_15572),
.B(n_3372),
.Y(n_15651)
);

INVx1_ASAP7_75t_L g15652 ( 
.A(n_15616),
.Y(n_15652)
);

NOR4xp25_ASAP7_75t_SL g15653 ( 
.A(n_15608),
.B(n_4068),
.C(n_4073),
.D(n_4067),
.Y(n_15653)
);

NOR2x1_ASAP7_75t_L g15654 ( 
.A(n_15579),
.B(n_3374),
.Y(n_15654)
);

NAND2xp5_ASAP7_75t_SL g15655 ( 
.A(n_15542),
.B(n_3373),
.Y(n_15655)
);

NAND3xp33_ASAP7_75t_L g15656 ( 
.A(n_15623),
.B(n_3374),
.C(n_3375),
.Y(n_15656)
);

INVx1_ASAP7_75t_L g15657 ( 
.A(n_15625),
.Y(n_15657)
);

INVx1_ASAP7_75t_L g15658 ( 
.A(n_15553),
.Y(n_15658)
);

NAND3xp33_ASAP7_75t_L g15659 ( 
.A(n_15568),
.B(n_3375),
.C(n_3376),
.Y(n_15659)
);

INVxp67_ASAP7_75t_SL g15660 ( 
.A(n_15566),
.Y(n_15660)
);

NAND4xp25_ASAP7_75t_L g15661 ( 
.A(n_15541),
.B(n_3378),
.C(n_3376),
.D(n_3377),
.Y(n_15661)
);

INVx1_ASAP7_75t_L g15662 ( 
.A(n_15620),
.Y(n_15662)
);

NOR2x1_ASAP7_75t_L g15663 ( 
.A(n_15563),
.B(n_3379),
.Y(n_15663)
);

OAI322xp33_ASAP7_75t_L g15664 ( 
.A1(n_15582),
.A2(n_3403),
.A3(n_3386),
.B1(n_3411),
.B2(n_3420),
.C1(n_3394),
.C2(n_3377),
.Y(n_15664)
);

NOR3xp33_ASAP7_75t_L g15665 ( 
.A(n_15611),
.B(n_3379),
.C(n_3380),
.Y(n_15665)
);

NAND2xp5_ASAP7_75t_L g15666 ( 
.A(n_15561),
.B(n_3381),
.Y(n_15666)
);

NOR3xp33_ASAP7_75t_L g15667 ( 
.A(n_15577),
.B(n_3380),
.C(n_3381),
.Y(n_15667)
);

AOI211xp5_ASAP7_75t_L g15668 ( 
.A1(n_15609),
.A2(n_3384),
.B(n_3382),
.C(n_3383),
.Y(n_15668)
);

NOR2x1_ASAP7_75t_L g15669 ( 
.A(n_15605),
.B(n_3384),
.Y(n_15669)
);

NOR2x1_ASAP7_75t_L g15670 ( 
.A(n_15554),
.B(n_3385),
.Y(n_15670)
);

NOR2x1_ASAP7_75t_L g15671 ( 
.A(n_15613),
.B(n_3385),
.Y(n_15671)
);

NAND2x1p5_ASAP7_75t_SL g15672 ( 
.A(n_15574),
.B(n_4062),
.Y(n_15672)
);

AOI22xp5_ASAP7_75t_L g15673 ( 
.A1(n_15544),
.A2(n_3387),
.B1(n_3383),
.B2(n_3386),
.Y(n_15673)
);

NOR2x1_ASAP7_75t_L g15674 ( 
.A(n_15586),
.B(n_3388),
.Y(n_15674)
);

OR2x2_ASAP7_75t_L g15675 ( 
.A(n_15564),
.B(n_3387),
.Y(n_15675)
);

NOR2xp67_ASAP7_75t_L g15676 ( 
.A(n_15610),
.B(n_3389),
.Y(n_15676)
);

NOR2x1_ASAP7_75t_L g15677 ( 
.A(n_15552),
.B(n_3389),
.Y(n_15677)
);

NOR3x1_ASAP7_75t_L g15678 ( 
.A(n_15612),
.B(n_3388),
.C(n_3390),
.Y(n_15678)
);

INVx1_ASAP7_75t_L g15679 ( 
.A(n_15617),
.Y(n_15679)
);

OAI211xp5_ASAP7_75t_L g15680 ( 
.A1(n_15559),
.A2(n_3392),
.B(n_3393),
.C(n_3391),
.Y(n_15680)
);

NAND2xp5_ASAP7_75t_L g15681 ( 
.A(n_15573),
.B(n_3391),
.Y(n_15681)
);

NAND2xp5_ASAP7_75t_SL g15682 ( 
.A(n_15604),
.B(n_3390),
.Y(n_15682)
);

INVx2_ASAP7_75t_L g15683 ( 
.A(n_15614),
.Y(n_15683)
);

AOI22xp5_ASAP7_75t_L g15684 ( 
.A1(n_15550),
.A2(n_3395),
.B1(n_3392),
.B2(n_3393),
.Y(n_15684)
);

NOR2x1_ASAP7_75t_L g15685 ( 
.A(n_15578),
.B(n_3397),
.Y(n_15685)
);

NOR2x1_ASAP7_75t_SL g15686 ( 
.A(n_15543),
.B(n_3397),
.Y(n_15686)
);

NAND4xp25_ASAP7_75t_L g15687 ( 
.A(n_15594),
.B(n_15556),
.C(n_15606),
.D(n_15580),
.Y(n_15687)
);

NAND3xp33_ASAP7_75t_L g15688 ( 
.A(n_15583),
.B(n_3395),
.C(n_3398),
.Y(n_15688)
);

NAND2xp5_ASAP7_75t_L g15689 ( 
.A(n_15555),
.B(n_3400),
.Y(n_15689)
);

NAND2xp5_ASAP7_75t_SL g15690 ( 
.A(n_15546),
.B(n_3399),
.Y(n_15690)
);

NOR2xp33_ASAP7_75t_L g15691 ( 
.A(n_15588),
.B(n_4059),
.Y(n_15691)
);

NOR2x1p5_ASAP7_75t_L g15692 ( 
.A(n_15591),
.B(n_3400),
.Y(n_15692)
);

NOR2x1p5_ASAP7_75t_L g15693 ( 
.A(n_15593),
.B(n_3401),
.Y(n_15693)
);

NOR3xp33_ASAP7_75t_L g15694 ( 
.A(n_15603),
.B(n_3401),
.C(n_3402),
.Y(n_15694)
);

NAND5xp2_ASAP7_75t_L g15695 ( 
.A(n_15585),
.B(n_3404),
.C(n_3402),
.D(n_3403),
.E(n_3405),
.Y(n_15695)
);

AOI221x1_ASAP7_75t_L g15696 ( 
.A1(n_15567),
.A2(n_3406),
.B1(n_3404),
.B2(n_3405),
.C(n_3407),
.Y(n_15696)
);

NOR3xp33_ASAP7_75t_L g15697 ( 
.A(n_15571),
.B(n_3406),
.C(n_3407),
.Y(n_15697)
);

HB1xp67_ASAP7_75t_L g15698 ( 
.A(n_15539),
.Y(n_15698)
);

AND4x1_ASAP7_75t_L g15699 ( 
.A(n_15587),
.B(n_3410),
.C(n_3408),
.D(n_3409),
.Y(n_15699)
);

NOR3xp33_ASAP7_75t_SL g15700 ( 
.A(n_15607),
.B(n_3408),
.C(n_3409),
.Y(n_15700)
);

INVx2_ASAP7_75t_L g15701 ( 
.A(n_15614),
.Y(n_15701)
);

NAND5xp2_ASAP7_75t_L g15702 ( 
.A(n_15596),
.B(n_3412),
.C(n_3410),
.D(n_3411),
.E(n_3413),
.Y(n_15702)
);

NAND2xp5_ASAP7_75t_L g15703 ( 
.A(n_15599),
.B(n_3414),
.Y(n_15703)
);

NOR3xp33_ASAP7_75t_SL g15704 ( 
.A(n_15569),
.B(n_15598),
.C(n_15548),
.Y(n_15704)
);

NOR2xp67_ASAP7_75t_L g15705 ( 
.A(n_15570),
.B(n_3415),
.Y(n_15705)
);

AND2x4_ASAP7_75t_L g15706 ( 
.A(n_15547),
.B(n_3413),
.Y(n_15706)
);

NAND2xp5_ASAP7_75t_L g15707 ( 
.A(n_15575),
.B(n_3417),
.Y(n_15707)
);

AOI21xp33_ASAP7_75t_L g15708 ( 
.A1(n_15560),
.A2(n_3416),
.B(n_3417),
.Y(n_15708)
);

NAND4xp75_ASAP7_75t_L g15709 ( 
.A(n_15600),
.B(n_3422),
.C(n_3419),
.D(n_3421),
.Y(n_15709)
);

NAND4xp25_ASAP7_75t_L g15710 ( 
.A(n_15601),
.B(n_3423),
.C(n_3419),
.D(n_3422),
.Y(n_15710)
);

NOR3xp33_ASAP7_75t_L g15711 ( 
.A(n_15592),
.B(n_3424),
.C(n_3425),
.Y(n_15711)
);

NOR2x1_ASAP7_75t_L g15712 ( 
.A(n_15545),
.B(n_3425),
.Y(n_15712)
);

NOR2xp33_ASAP7_75t_L g15713 ( 
.A(n_15565),
.B(n_4075),
.Y(n_15713)
);

NAND3xp33_ASAP7_75t_L g15714 ( 
.A(n_15619),
.B(n_3424),
.C(n_3426),
.Y(n_15714)
);

AND2x2_ASAP7_75t_L g15715 ( 
.A(n_15543),
.B(n_3426),
.Y(n_15715)
);

NOR3x1_ASAP7_75t_L g15716 ( 
.A(n_15537),
.B(n_3427),
.C(n_3428),
.Y(n_15716)
);

NOR3xp33_ASAP7_75t_L g15717 ( 
.A(n_15549),
.B(n_3429),
.C(n_3431),
.Y(n_15717)
);

NOR2x1_ASAP7_75t_L g15718 ( 
.A(n_15618),
.B(n_3431),
.Y(n_15718)
);

NAND2xp5_ASAP7_75t_L g15719 ( 
.A(n_15576),
.B(n_3432),
.Y(n_15719)
);

NOR2x1_ASAP7_75t_L g15720 ( 
.A(n_15618),
.B(n_3432),
.Y(n_15720)
);

AND2x4_ASAP7_75t_L g15721 ( 
.A(n_15617),
.B(n_3429),
.Y(n_15721)
);

INVx1_ASAP7_75t_L g15722 ( 
.A(n_15576),
.Y(n_15722)
);

INVx1_ASAP7_75t_L g15723 ( 
.A(n_15576),
.Y(n_15723)
);

NOR2x1_ASAP7_75t_L g15724 ( 
.A(n_15618),
.B(n_3434),
.Y(n_15724)
);

NAND3xp33_ASAP7_75t_L g15725 ( 
.A(n_15619),
.B(n_3433),
.C(n_3434),
.Y(n_15725)
);

NOR2x1_ASAP7_75t_L g15726 ( 
.A(n_15618),
.B(n_3436),
.Y(n_15726)
);

NOR4xp75_ASAP7_75t_L g15727 ( 
.A(n_15557),
.B(n_3438),
.C(n_3433),
.D(n_3437),
.Y(n_15727)
);

NAND3xp33_ASAP7_75t_SL g15728 ( 
.A(n_15619),
.B(n_3437),
.C(n_3439),
.Y(n_15728)
);

NOR2x1_ASAP7_75t_L g15729 ( 
.A(n_15618),
.B(n_3440),
.Y(n_15729)
);

NOR4xp25_ASAP7_75t_L g15730 ( 
.A(n_15549),
.B(n_4091),
.C(n_4063),
.D(n_3441),
.Y(n_15730)
);

NOR3x1_ASAP7_75t_L g15731 ( 
.A(n_15537),
.B(n_3439),
.C(n_3440),
.Y(n_15731)
);

NAND3xp33_ASAP7_75t_L g15732 ( 
.A(n_15619),
.B(n_3441),
.C(n_3442),
.Y(n_15732)
);

AOI21xp5_ASAP7_75t_L g15733 ( 
.A1(n_15660),
.A2(n_3442),
.B(n_3444),
.Y(n_15733)
);

AND4x2_ASAP7_75t_L g15734 ( 
.A(n_15648),
.B(n_3446),
.C(n_3444),
.D(n_3445),
.Y(n_15734)
);

AOI21xp5_ASAP7_75t_L g15735 ( 
.A1(n_15638),
.A2(n_3445),
.B(n_3446),
.Y(n_15735)
);

OAI221xp5_ASAP7_75t_L g15736 ( 
.A1(n_15710),
.A2(n_3449),
.B1(n_3447),
.B2(n_3448),
.C(n_3450),
.Y(n_15736)
);

BUFx3_ASAP7_75t_L g15737 ( 
.A(n_15715),
.Y(n_15737)
);

AOI211xp5_ASAP7_75t_L g15738 ( 
.A1(n_15642),
.A2(n_3450),
.B(n_3447),
.C(n_3448),
.Y(n_15738)
);

OAI21xp33_ASAP7_75t_L g15739 ( 
.A1(n_15643),
.A2(n_3451),
.B(n_3452),
.Y(n_15739)
);

AOI22xp5_ASAP7_75t_L g15740 ( 
.A1(n_15713),
.A2(n_3453),
.B1(n_3451),
.B2(n_3452),
.Y(n_15740)
);

AOI211xp5_ASAP7_75t_L g15741 ( 
.A1(n_15636),
.A2(n_3455),
.B(n_3453),
.C(n_3454),
.Y(n_15741)
);

OAI211xp5_ASAP7_75t_L g15742 ( 
.A1(n_15719),
.A2(n_3456),
.B(n_3457),
.C(n_3455),
.Y(n_15742)
);

NAND2xp5_ASAP7_75t_L g15743 ( 
.A(n_15705),
.B(n_15631),
.Y(n_15743)
);

OAI221xp5_ASAP7_75t_L g15744 ( 
.A1(n_15673),
.A2(n_3457),
.B1(n_3454),
.B2(n_3456),
.C(n_3458),
.Y(n_15744)
);

NOR2x1_ASAP7_75t_L g15745 ( 
.A(n_15654),
.B(n_4075),
.Y(n_15745)
);

AOI222xp33_ASAP7_75t_L g15746 ( 
.A1(n_15647),
.A2(n_3461),
.B1(n_3463),
.B2(n_3459),
.C1(n_3460),
.C2(n_3462),
.Y(n_15746)
);

OAI21xp5_ASAP7_75t_L g15747 ( 
.A1(n_15634),
.A2(n_3459),
.B(n_3460),
.Y(n_15747)
);

OAI211xp5_ASAP7_75t_SL g15748 ( 
.A1(n_15704),
.A2(n_15627),
.B(n_15723),
.C(n_15722),
.Y(n_15748)
);

OAI211xp5_ASAP7_75t_L g15749 ( 
.A1(n_15635),
.A2(n_3464),
.B(n_3465),
.C(n_3463),
.Y(n_15749)
);

NAND3xp33_ASAP7_75t_SL g15750 ( 
.A(n_15653),
.B(n_15668),
.C(n_15727),
.Y(n_15750)
);

AOI221xp5_ASAP7_75t_L g15751 ( 
.A1(n_15650),
.A2(n_3465),
.B1(n_3461),
.B2(n_3464),
.C(n_3466),
.Y(n_15751)
);

OAI211xp5_ASAP7_75t_L g15752 ( 
.A1(n_15646),
.A2(n_3469),
.B(n_3470),
.C(n_3468),
.Y(n_15752)
);

NOR4xp75_ASAP7_75t_L g15753 ( 
.A(n_15690),
.B(n_3469),
.C(n_3467),
.D(n_3468),
.Y(n_15753)
);

NAND4xp25_ASAP7_75t_L g15754 ( 
.A(n_15716),
.B(n_4085),
.C(n_4060),
.D(n_3473),
.Y(n_15754)
);

OAI211xp5_ASAP7_75t_L g15755 ( 
.A1(n_15670),
.A2(n_3473),
.B(n_3474),
.C(n_3471),
.Y(n_15755)
);

AOI221xp5_ASAP7_75t_L g15756 ( 
.A1(n_15728),
.A2(n_3475),
.B1(n_3470),
.B2(n_3474),
.C(n_3476),
.Y(n_15756)
);

NAND2xp5_ASAP7_75t_SL g15757 ( 
.A(n_15721),
.B(n_3476),
.Y(n_15757)
);

NAND2xp5_ASAP7_75t_L g15758 ( 
.A(n_15693),
.B(n_3477),
.Y(n_15758)
);

AOI222xp33_ASAP7_75t_L g15759 ( 
.A1(n_15676),
.A2(n_3480),
.B1(n_3482),
.B2(n_3478),
.C1(n_3479),
.C2(n_3481),
.Y(n_15759)
);

AOI221xp5_ASAP7_75t_L g15760 ( 
.A1(n_15637),
.A2(n_3482),
.B1(n_3478),
.B2(n_3481),
.C(n_3483),
.Y(n_15760)
);

AOI221xp5_ASAP7_75t_L g15761 ( 
.A1(n_15714),
.A2(n_3486),
.B1(n_3484),
.B2(n_3485),
.C(n_3487),
.Y(n_15761)
);

AOI22xp33_ASAP7_75t_L g15762 ( 
.A1(n_15706),
.A2(n_3486),
.B1(n_3484),
.B2(n_3485),
.Y(n_15762)
);

AOI221xp5_ASAP7_75t_L g15763 ( 
.A1(n_15732),
.A2(n_3489),
.B1(n_3487),
.B2(n_3488),
.C(n_3490),
.Y(n_15763)
);

INVx1_ASAP7_75t_L g15764 ( 
.A(n_15671),
.Y(n_15764)
);

NOR3xp33_ASAP7_75t_L g15765 ( 
.A(n_15662),
.B(n_3488),
.C(n_3489),
.Y(n_15765)
);

A2O1A1Ixp33_ASAP7_75t_L g15766 ( 
.A1(n_15691),
.A2(n_4064),
.B(n_3492),
.C(n_3490),
.Y(n_15766)
);

NAND3xp33_ASAP7_75t_L g15767 ( 
.A(n_15629),
.B(n_3491),
.C(n_3492),
.Y(n_15767)
);

NOR2xp33_ASAP7_75t_L g15768 ( 
.A(n_15702),
.B(n_3491),
.Y(n_15768)
);

AOI21xp33_ASAP7_75t_SL g15769 ( 
.A1(n_15672),
.A2(n_3493),
.B(n_3494),
.Y(n_15769)
);

AOI211x1_ASAP7_75t_SL g15770 ( 
.A1(n_15687),
.A2(n_3496),
.B(n_3494),
.C(n_3495),
.Y(n_15770)
);

NOR2xp67_ASAP7_75t_L g15771 ( 
.A(n_15695),
.B(n_4054),
.Y(n_15771)
);

OA22x2_ASAP7_75t_L g15772 ( 
.A1(n_15684),
.A2(n_3498),
.B1(n_3495),
.B2(n_3497),
.Y(n_15772)
);

AOI22xp33_ASAP7_75t_L g15773 ( 
.A1(n_15706),
.A2(n_3500),
.B1(n_3497),
.B2(n_3499),
.Y(n_15773)
);

AOI22xp5_ASAP7_75t_L g15774 ( 
.A1(n_15721),
.A2(n_3502),
.B1(n_3499),
.B2(n_3501),
.Y(n_15774)
);

OAI221xp5_ASAP7_75t_L g15775 ( 
.A1(n_15680),
.A2(n_3503),
.B1(n_3501),
.B2(n_3502),
.C(n_3504),
.Y(n_15775)
);

AO22x2_ASAP7_75t_L g15776 ( 
.A1(n_15683),
.A2(n_3505),
.B1(n_3503),
.B2(n_3504),
.Y(n_15776)
);

AOI21xp33_ASAP7_75t_SL g15777 ( 
.A1(n_15640),
.A2(n_3505),
.B(n_3506),
.Y(n_15777)
);

OAI211xp5_ASAP7_75t_L g15778 ( 
.A1(n_15677),
.A2(n_3508),
.B(n_3509),
.C(n_3507),
.Y(n_15778)
);

OAI211xp5_ASAP7_75t_SL g15779 ( 
.A1(n_15628),
.A2(n_15720),
.B(n_15724),
.C(n_15718),
.Y(n_15779)
);

NOR2x1_ASAP7_75t_L g15780 ( 
.A(n_15701),
.B(n_4076),
.Y(n_15780)
);

BUFx2_ASAP7_75t_L g15781 ( 
.A(n_15639),
.Y(n_15781)
);

NOR2xp67_ASAP7_75t_L g15782 ( 
.A(n_15651),
.B(n_4076),
.Y(n_15782)
);

AND2x2_ASAP7_75t_L g15783 ( 
.A(n_15641),
.B(n_3506),
.Y(n_15783)
);

OAI211xp5_ASAP7_75t_SL g15784 ( 
.A1(n_15726),
.A2(n_3510),
.B(n_3508),
.C(n_3509),
.Y(n_15784)
);

NOR3xp33_ASAP7_75t_L g15785 ( 
.A(n_15644),
.B(n_3510),
.C(n_3511),
.Y(n_15785)
);

AOI21xp5_ASAP7_75t_L g15786 ( 
.A1(n_15707),
.A2(n_3512),
.B(n_3513),
.Y(n_15786)
);

AND5x1_ASAP7_75t_L g15787 ( 
.A(n_15669),
.B(n_3514),
.C(n_3512),
.D(n_3513),
.E(n_3515),
.Y(n_15787)
);

OAI211xp5_ASAP7_75t_SL g15788 ( 
.A1(n_15729),
.A2(n_3517),
.B(n_3514),
.C(n_3516),
.Y(n_15788)
);

AOI211x1_ASAP7_75t_SL g15789 ( 
.A1(n_15655),
.A2(n_3518),
.B(n_3516),
.C(n_3517),
.Y(n_15789)
);

AOI22xp33_ASAP7_75t_L g15790 ( 
.A1(n_15663),
.A2(n_15630),
.B1(n_15633),
.B2(n_15725),
.Y(n_15790)
);

OA22x2_ASAP7_75t_L g15791 ( 
.A1(n_15681),
.A2(n_3520),
.B1(n_3518),
.B2(n_3519),
.Y(n_15791)
);

AOI221xp5_ASAP7_75t_L g15792 ( 
.A1(n_15730),
.A2(n_3522),
.B1(n_3520),
.B2(n_3521),
.C(n_3523),
.Y(n_15792)
);

NAND4xp75_ASAP7_75t_L g15793 ( 
.A(n_15685),
.B(n_15674),
.C(n_15731),
.D(n_15678),
.Y(n_15793)
);

AOI211xp5_ASAP7_75t_L g15794 ( 
.A1(n_15688),
.A2(n_3523),
.B(n_3521),
.C(n_3522),
.Y(n_15794)
);

OAI22xp5_ASAP7_75t_L g15795 ( 
.A1(n_15656),
.A2(n_3526),
.B1(n_3524),
.B2(n_3525),
.Y(n_15795)
);

NOR2xp33_ASAP7_75t_L g15796 ( 
.A(n_15675),
.B(n_15686),
.Y(n_15796)
);

NAND2xp5_ASAP7_75t_SL g15797 ( 
.A(n_15659),
.B(n_15679),
.Y(n_15797)
);

A2O1A1Ixp33_ASAP7_75t_L g15798 ( 
.A1(n_15700),
.A2(n_3528),
.B(n_3526),
.C(n_3527),
.Y(n_15798)
);

OAI211xp5_ASAP7_75t_L g15799 ( 
.A1(n_15698),
.A2(n_3530),
.B(n_3531),
.C(n_3529),
.Y(n_15799)
);

AOI211xp5_ASAP7_75t_L g15800 ( 
.A1(n_15666),
.A2(n_15689),
.B(n_15682),
.C(n_15703),
.Y(n_15800)
);

HB1xp67_ASAP7_75t_L g15801 ( 
.A(n_15699),
.Y(n_15801)
);

AOI221xp5_ASAP7_75t_L g15802 ( 
.A1(n_15649),
.A2(n_3531),
.B1(n_3528),
.B2(n_3530),
.C(n_3532),
.Y(n_15802)
);

INVxp67_ASAP7_75t_L g15803 ( 
.A(n_15632),
.Y(n_15803)
);

OAI211xp5_ASAP7_75t_L g15804 ( 
.A1(n_15712),
.A2(n_3534),
.B(n_3536),
.C(n_3533),
.Y(n_15804)
);

AOI221xp5_ASAP7_75t_L g15805 ( 
.A1(n_15652),
.A2(n_15657),
.B1(n_15658),
.B2(n_15664),
.C(n_15717),
.Y(n_15805)
);

OAI211xp5_ASAP7_75t_L g15806 ( 
.A1(n_15661),
.A2(n_3534),
.B(n_3536),
.C(n_3533),
.Y(n_15806)
);

OAI22xp5_ASAP7_75t_L g15807 ( 
.A1(n_15692),
.A2(n_3538),
.B1(n_3532),
.B2(n_3537),
.Y(n_15807)
);

OAI22xp33_ASAP7_75t_SL g15808 ( 
.A1(n_15645),
.A2(n_3540),
.B1(n_3537),
.B2(n_3539),
.Y(n_15808)
);

INVx1_ASAP7_75t_L g15809 ( 
.A(n_15709),
.Y(n_15809)
);

AOI221xp5_ASAP7_75t_L g15810 ( 
.A1(n_15708),
.A2(n_3543),
.B1(n_3541),
.B2(n_3542),
.C(n_3544),
.Y(n_15810)
);

NAND3xp33_ASAP7_75t_SL g15811 ( 
.A(n_15805),
.B(n_15665),
.C(n_15667),
.Y(n_15811)
);

OR2x2_ASAP7_75t_L g15812 ( 
.A(n_15754),
.B(n_15694),
.Y(n_15812)
);

AND2x4_ASAP7_75t_L g15813 ( 
.A(n_15753),
.B(n_15711),
.Y(n_15813)
);

AOI22xp5_ASAP7_75t_L g15814 ( 
.A1(n_15768),
.A2(n_15697),
.B1(n_15626),
.B2(n_15696),
.Y(n_15814)
);

INVx1_ASAP7_75t_L g15815 ( 
.A(n_15734),
.Y(n_15815)
);

INVx1_ASAP7_75t_L g15816 ( 
.A(n_15791),
.Y(n_15816)
);

AND2x4_ASAP7_75t_L g15817 ( 
.A(n_15787),
.B(n_15626),
.Y(n_15817)
);

NOR3xp33_ASAP7_75t_SL g15818 ( 
.A(n_15748),
.B(n_3544),
.C(n_3545),
.Y(n_15818)
);

NOR2x1_ASAP7_75t_L g15819 ( 
.A(n_15779),
.B(n_3545),
.Y(n_15819)
);

NOR2x1_ASAP7_75t_L g15820 ( 
.A(n_15745),
.B(n_3546),
.Y(n_15820)
);

NAND3xp33_ASAP7_75t_L g15821 ( 
.A(n_15747),
.B(n_3555),
.C(n_3547),
.Y(n_15821)
);

AND3x4_ASAP7_75t_L g15822 ( 
.A(n_15771),
.B(n_3556),
.C(n_3548),
.Y(n_15822)
);

NOR2xp33_ASAP7_75t_L g15823 ( 
.A(n_15739),
.B(n_3548),
.Y(n_15823)
);

NAND2xp5_ASAP7_75t_L g15824 ( 
.A(n_15762),
.B(n_3549),
.Y(n_15824)
);

OAI22xp33_ASAP7_75t_L g15825 ( 
.A1(n_15774),
.A2(n_3551),
.B1(n_3549),
.B2(n_3550),
.Y(n_15825)
);

XOR2x1_ASAP7_75t_L g15826 ( 
.A(n_15764),
.B(n_3552),
.Y(n_15826)
);

NOR3xp33_ASAP7_75t_L g15827 ( 
.A(n_15797),
.B(n_3552),
.C(n_3553),
.Y(n_15827)
);

INVxp33_ASAP7_75t_L g15828 ( 
.A(n_15780),
.Y(n_15828)
);

NOR2x1_ASAP7_75t_L g15829 ( 
.A(n_15793),
.B(n_3554),
.Y(n_15829)
);

NOR2xp33_ASAP7_75t_L g15830 ( 
.A(n_15769),
.B(n_3554),
.Y(n_15830)
);

OAI21xp33_ASAP7_75t_L g15831 ( 
.A1(n_15737),
.A2(n_3555),
.B(n_3556),
.Y(n_15831)
);

INVx1_ASAP7_75t_L g15832 ( 
.A(n_15772),
.Y(n_15832)
);

NAND2xp5_ASAP7_75t_SL g15833 ( 
.A(n_15759),
.B(n_3557),
.Y(n_15833)
);

OAI21xp5_ASAP7_75t_SL g15834 ( 
.A1(n_15770),
.A2(n_3557),
.B(n_3558),
.Y(n_15834)
);

OAI31xp33_ASAP7_75t_L g15835 ( 
.A1(n_15784),
.A2(n_3560),
.A3(n_3558),
.B(n_3559),
.Y(n_15835)
);

NOR2xp33_ASAP7_75t_L g15836 ( 
.A(n_15757),
.B(n_3559),
.Y(n_15836)
);

INVxp67_ASAP7_75t_SL g15837 ( 
.A(n_15782),
.Y(n_15837)
);

INVx2_ASAP7_75t_SL g15838 ( 
.A(n_15783),
.Y(n_15838)
);

NOR2x1_ASAP7_75t_L g15839 ( 
.A(n_15781),
.B(n_3561),
.Y(n_15839)
);

INVx1_ASAP7_75t_L g15840 ( 
.A(n_15758),
.Y(n_15840)
);

AOI31xp33_ASAP7_75t_L g15841 ( 
.A1(n_15790),
.A2(n_3563),
.A3(n_3561),
.B(n_3562),
.Y(n_15841)
);

NAND4xp75_ASAP7_75t_L g15842 ( 
.A(n_15786),
.B(n_15809),
.C(n_15796),
.D(n_15743),
.Y(n_15842)
);

NOR2x1p5_ASAP7_75t_L g15843 ( 
.A(n_15750),
.B(n_3562),
.Y(n_15843)
);

NOR2x1_ASAP7_75t_L g15844 ( 
.A(n_15778),
.B(n_3563),
.Y(n_15844)
);

AOI22xp5_ASAP7_75t_L g15845 ( 
.A1(n_15806),
.A2(n_3566),
.B1(n_3564),
.B2(n_3565),
.Y(n_15845)
);

NOR3x2_ASAP7_75t_L g15846 ( 
.A(n_15789),
.B(n_3573),
.C(n_3564),
.Y(n_15846)
);

INVx1_ASAP7_75t_L g15847 ( 
.A(n_15804),
.Y(n_15847)
);

NOR2xp33_ASAP7_75t_L g15848 ( 
.A(n_15788),
.B(n_3565),
.Y(n_15848)
);

AND2x2_ASAP7_75t_L g15849 ( 
.A(n_15801),
.B(n_3566),
.Y(n_15849)
);

INVx1_ASAP7_75t_L g15850 ( 
.A(n_15767),
.Y(n_15850)
);

OR2x2_ASAP7_75t_L g15851 ( 
.A(n_15773),
.B(n_3567),
.Y(n_15851)
);

NOR2x1_ASAP7_75t_L g15852 ( 
.A(n_15752),
.B(n_3567),
.Y(n_15852)
);

NOR3xp33_ASAP7_75t_L g15853 ( 
.A(n_15803),
.B(n_3569),
.C(n_3570),
.Y(n_15853)
);

NOR2x1_ASAP7_75t_L g15854 ( 
.A(n_15749),
.B(n_3571),
.Y(n_15854)
);

NAND2xp5_ASAP7_75t_L g15855 ( 
.A(n_15792),
.B(n_15738),
.Y(n_15855)
);

NOR2x1_ASAP7_75t_L g15856 ( 
.A(n_15755),
.B(n_3571),
.Y(n_15856)
);

INVx1_ASAP7_75t_L g15857 ( 
.A(n_15798),
.Y(n_15857)
);

NOR3xp33_ASAP7_75t_SL g15858 ( 
.A(n_15775),
.B(n_3572),
.C(n_3573),
.Y(n_15858)
);

NOR3xp33_ASAP7_75t_L g15859 ( 
.A(n_15800),
.B(n_3572),
.C(n_3574),
.Y(n_15859)
);

INVx1_ASAP7_75t_SL g15860 ( 
.A(n_15733),
.Y(n_15860)
);

INVxp33_ASAP7_75t_SL g15861 ( 
.A(n_15777),
.Y(n_15861)
);

NAND4xp75_ASAP7_75t_L g15862 ( 
.A(n_15751),
.B(n_3577),
.C(n_3575),
.D(n_3576),
.Y(n_15862)
);

INVx1_ASAP7_75t_L g15863 ( 
.A(n_15736),
.Y(n_15863)
);

NOR3xp33_ASAP7_75t_SL g15864 ( 
.A(n_15744),
.B(n_3575),
.C(n_3576),
.Y(n_15864)
);

AND2x4_ASAP7_75t_L g15865 ( 
.A(n_15735),
.B(n_3577),
.Y(n_15865)
);

NAND4xp75_ASAP7_75t_L g15866 ( 
.A(n_15756),
.B(n_3580),
.C(n_3578),
.D(n_3579),
.Y(n_15866)
);

AND3x2_ASAP7_75t_L g15867 ( 
.A(n_15765),
.B(n_3580),
.C(n_3579),
.Y(n_15867)
);

NAND4xp75_ASAP7_75t_L g15868 ( 
.A(n_15760),
.B(n_3582),
.C(n_3578),
.D(n_3581),
.Y(n_15868)
);

NOR2x1_ASAP7_75t_L g15869 ( 
.A(n_15742),
.B(n_3581),
.Y(n_15869)
);

AND2x2_ASAP7_75t_L g15870 ( 
.A(n_15746),
.B(n_3582),
.Y(n_15870)
);

NOR2x1_ASAP7_75t_L g15871 ( 
.A(n_15799),
.B(n_3583),
.Y(n_15871)
);

NAND2xp5_ASAP7_75t_L g15872 ( 
.A(n_15741),
.B(n_15794),
.Y(n_15872)
);

NAND2xp5_ASAP7_75t_L g15873 ( 
.A(n_15761),
.B(n_3583),
.Y(n_15873)
);

AOI22xp5_ASAP7_75t_L g15874 ( 
.A1(n_15822),
.A2(n_15795),
.B1(n_15763),
.B2(n_15810),
.Y(n_15874)
);

NAND4xp75_ASAP7_75t_L g15875 ( 
.A(n_15849),
.B(n_15740),
.C(n_15802),
.D(n_15808),
.Y(n_15875)
);

NOR3xp33_ASAP7_75t_L g15876 ( 
.A(n_15811),
.B(n_15807),
.C(n_15785),
.Y(n_15876)
);

XNOR2xp5_ASAP7_75t_L g15877 ( 
.A(n_15846),
.B(n_15776),
.Y(n_15877)
);

INVx2_ASAP7_75t_SL g15878 ( 
.A(n_15820),
.Y(n_15878)
);

OAI22xp5_ASAP7_75t_L g15879 ( 
.A1(n_15845),
.A2(n_15766),
.B1(n_15776),
.B2(n_3586),
.Y(n_15879)
);

OAI22xp5_ASAP7_75t_L g15880 ( 
.A1(n_15821),
.A2(n_3586),
.B1(n_3584),
.B2(n_3585),
.Y(n_15880)
);

OR2x2_ASAP7_75t_L g15881 ( 
.A(n_15851),
.B(n_15824),
.Y(n_15881)
);

AOI22xp5_ASAP7_75t_L g15882 ( 
.A1(n_15843),
.A2(n_15836),
.B1(n_15848),
.B2(n_15830),
.Y(n_15882)
);

NAND4xp75_ASAP7_75t_L g15883 ( 
.A(n_15829),
.B(n_3587),
.C(n_3584),
.D(n_3585),
.Y(n_15883)
);

NAND2xp5_ASAP7_75t_L g15884 ( 
.A(n_15826),
.B(n_3588),
.Y(n_15884)
);

XNOR2xp5_ASAP7_75t_L g15885 ( 
.A(n_15818),
.B(n_3588),
.Y(n_15885)
);

INVx2_ASAP7_75t_L g15886 ( 
.A(n_15867),
.Y(n_15886)
);

OAI221xp5_ASAP7_75t_L g15887 ( 
.A1(n_15835),
.A2(n_3592),
.B1(n_3589),
.B2(n_3591),
.C(n_3593),
.Y(n_15887)
);

INVx2_ASAP7_75t_L g15888 ( 
.A(n_15839),
.Y(n_15888)
);

NOR2x1_ASAP7_75t_L g15889 ( 
.A(n_15819),
.B(n_3589),
.Y(n_15889)
);

XNOR2x1_ASAP7_75t_L g15890 ( 
.A(n_15842),
.B(n_3591),
.Y(n_15890)
);

INVx2_ASAP7_75t_SL g15891 ( 
.A(n_15817),
.Y(n_15891)
);

INVx1_ASAP7_75t_L g15892 ( 
.A(n_15817),
.Y(n_15892)
);

AOI21xp5_ASAP7_75t_L g15893 ( 
.A1(n_15828),
.A2(n_3592),
.B(n_3594),
.Y(n_15893)
);

OR2x2_ASAP7_75t_L g15894 ( 
.A(n_15834),
.B(n_3594),
.Y(n_15894)
);

NAND2xp5_ASAP7_75t_L g15895 ( 
.A(n_15827),
.B(n_3595),
.Y(n_15895)
);

XNOR2xp5_ASAP7_75t_L g15896 ( 
.A(n_15814),
.B(n_3595),
.Y(n_15896)
);

OAI211xp5_ASAP7_75t_SL g15897 ( 
.A1(n_15847),
.A2(n_3600),
.B(n_3596),
.C(n_3597),
.Y(n_15897)
);

INVx4_ASAP7_75t_L g15898 ( 
.A(n_15838),
.Y(n_15898)
);

XNOR2xp5_ASAP7_75t_L g15899 ( 
.A(n_15862),
.B(n_3596),
.Y(n_15899)
);

AOI22xp5_ASAP7_75t_L g15900 ( 
.A1(n_15823),
.A2(n_3602),
.B1(n_3603),
.B2(n_3601),
.Y(n_15900)
);

INVx1_ASAP7_75t_L g15901 ( 
.A(n_15852),
.Y(n_15901)
);

OAI22xp5_ASAP7_75t_SL g15902 ( 
.A1(n_15815),
.A2(n_3602),
.B1(n_3600),
.B2(n_3601),
.Y(n_15902)
);

INVx1_ASAP7_75t_L g15903 ( 
.A(n_15854),
.Y(n_15903)
);

OR2x2_ASAP7_75t_L g15904 ( 
.A(n_15833),
.B(n_15816),
.Y(n_15904)
);

NAND4xp75_ASAP7_75t_L g15905 ( 
.A(n_15832),
.B(n_3607),
.C(n_3605),
.D(n_3606),
.Y(n_15905)
);

NOR2x1_ASAP7_75t_L g15906 ( 
.A(n_15869),
.B(n_3605),
.Y(n_15906)
);

OAI21xp5_ASAP7_75t_L g15907 ( 
.A1(n_15844),
.A2(n_3606),
.B(n_3607),
.Y(n_15907)
);

INVx2_ASAP7_75t_L g15908 ( 
.A(n_15866),
.Y(n_15908)
);

NAND2xp5_ASAP7_75t_L g15909 ( 
.A(n_15859),
.B(n_3608),
.Y(n_15909)
);

NOR2x1p5_ASAP7_75t_L g15910 ( 
.A(n_15868),
.B(n_3608),
.Y(n_15910)
);

OA22x2_ASAP7_75t_L g15911 ( 
.A1(n_15865),
.A2(n_3611),
.B1(n_3609),
.B2(n_3610),
.Y(n_15911)
);

INVx1_ASAP7_75t_L g15912 ( 
.A(n_15856),
.Y(n_15912)
);

INVx1_ASAP7_75t_L g15913 ( 
.A(n_15871),
.Y(n_15913)
);

INVx2_ASAP7_75t_L g15914 ( 
.A(n_15865),
.Y(n_15914)
);

INVx2_ASAP7_75t_L g15915 ( 
.A(n_15813),
.Y(n_15915)
);

OR2x2_ASAP7_75t_L g15916 ( 
.A(n_15873),
.B(n_3609),
.Y(n_15916)
);

INVx1_ASAP7_75t_L g15917 ( 
.A(n_15870),
.Y(n_15917)
);

INVx1_ASAP7_75t_L g15918 ( 
.A(n_15858),
.Y(n_15918)
);

XOR2xp5_ASAP7_75t_L g15919 ( 
.A(n_15812),
.B(n_3612),
.Y(n_15919)
);

INVx1_ASAP7_75t_L g15920 ( 
.A(n_15864),
.Y(n_15920)
);

NAND4xp75_ASAP7_75t_L g15921 ( 
.A(n_15850),
.B(n_3613),
.C(n_3610),
.D(n_3612),
.Y(n_15921)
);

AOI22xp5_ASAP7_75t_L g15922 ( 
.A1(n_15861),
.A2(n_15813),
.B1(n_15825),
.B2(n_15837),
.Y(n_15922)
);

XOR2xp5_ASAP7_75t_L g15923 ( 
.A(n_15863),
.B(n_3614),
.Y(n_15923)
);

INVx2_ASAP7_75t_L g15924 ( 
.A(n_15857),
.Y(n_15924)
);

AOI21xp5_ASAP7_75t_L g15925 ( 
.A1(n_15855),
.A2(n_15872),
.B(n_15860),
.Y(n_15925)
);

NAND4xp75_ASAP7_75t_L g15926 ( 
.A(n_15840),
.B(n_3615),
.C(n_3613),
.D(n_3614),
.Y(n_15926)
);

NAND2xp5_ASAP7_75t_SL g15927 ( 
.A(n_15853),
.B(n_3615),
.Y(n_15927)
);

NOR2xp33_ASAP7_75t_L g15928 ( 
.A(n_15841),
.B(n_3616),
.Y(n_15928)
);

INVx1_ASAP7_75t_L g15929 ( 
.A(n_15831),
.Y(n_15929)
);

NAND2xp33_ASAP7_75t_L g15930 ( 
.A(n_15818),
.B(n_3616),
.Y(n_15930)
);

AOI22xp33_ASAP7_75t_SL g15931 ( 
.A1(n_15891),
.A2(n_3619),
.B1(n_3617),
.B2(n_3618),
.Y(n_15931)
);

AND2x4_ASAP7_75t_L g15932 ( 
.A(n_15892),
.B(n_3618),
.Y(n_15932)
);

INVx1_ASAP7_75t_L g15933 ( 
.A(n_15890),
.Y(n_15933)
);

NOR3xp33_ASAP7_75t_L g15934 ( 
.A(n_15898),
.B(n_15915),
.C(n_15878),
.Y(n_15934)
);

INVx1_ASAP7_75t_L g15935 ( 
.A(n_15884),
.Y(n_15935)
);

INVx2_ASAP7_75t_SL g15936 ( 
.A(n_15910),
.Y(n_15936)
);

OAI21xp5_ASAP7_75t_L g15937 ( 
.A1(n_15885),
.A2(n_15899),
.B(n_15928),
.Y(n_15937)
);

NAND2xp5_ASAP7_75t_L g15938 ( 
.A(n_15896),
.B(n_3620),
.Y(n_15938)
);

AND2x4_ASAP7_75t_L g15939 ( 
.A(n_15908),
.B(n_3619),
.Y(n_15939)
);

INVx1_ASAP7_75t_L g15940 ( 
.A(n_15911),
.Y(n_15940)
);

INVx2_ASAP7_75t_L g15941 ( 
.A(n_15905),
.Y(n_15941)
);

INVx1_ASAP7_75t_L g15942 ( 
.A(n_15883),
.Y(n_15942)
);

AND2x4_ASAP7_75t_L g15943 ( 
.A(n_15914),
.B(n_3620),
.Y(n_15943)
);

NOR2x1_ASAP7_75t_L g15944 ( 
.A(n_15888),
.B(n_3621),
.Y(n_15944)
);

NAND4xp75_ASAP7_75t_L g15945 ( 
.A(n_15906),
.B(n_3624),
.C(n_3621),
.D(n_3622),
.Y(n_15945)
);

INVx1_ASAP7_75t_L g15946 ( 
.A(n_15889),
.Y(n_15946)
);

NOR2xp33_ASAP7_75t_L g15947 ( 
.A(n_15894),
.B(n_3622),
.Y(n_15947)
);

NOR3xp33_ASAP7_75t_L g15948 ( 
.A(n_15924),
.B(n_3625),
.C(n_3626),
.Y(n_15948)
);

XOR2xp5_ASAP7_75t_L g15949 ( 
.A(n_15877),
.B(n_3625),
.Y(n_15949)
);

NOR2x1_ASAP7_75t_L g15950 ( 
.A(n_15886),
.B(n_3626),
.Y(n_15950)
);

OR2x2_ASAP7_75t_L g15951 ( 
.A(n_15880),
.B(n_3627),
.Y(n_15951)
);

NAND4xp75_ASAP7_75t_L g15952 ( 
.A(n_15925),
.B(n_3630),
.C(n_3628),
.D(n_3629),
.Y(n_15952)
);

INVxp67_ASAP7_75t_SL g15953 ( 
.A(n_15916),
.Y(n_15953)
);

INVx2_ASAP7_75t_SL g15954 ( 
.A(n_15895),
.Y(n_15954)
);

NAND2xp5_ASAP7_75t_L g15955 ( 
.A(n_15907),
.B(n_3629),
.Y(n_15955)
);

AND2x2_ASAP7_75t_SL g15956 ( 
.A(n_15876),
.B(n_3628),
.Y(n_15956)
);

INVx1_ASAP7_75t_L g15957 ( 
.A(n_15930),
.Y(n_15957)
);

XNOR2xp5_ASAP7_75t_L g15958 ( 
.A(n_15875),
.B(n_3630),
.Y(n_15958)
);

AND2x4_ASAP7_75t_L g15959 ( 
.A(n_15920),
.B(n_3632),
.Y(n_15959)
);

INVx1_ASAP7_75t_SL g15960 ( 
.A(n_15923),
.Y(n_15960)
);

NAND2xp5_ASAP7_75t_L g15961 ( 
.A(n_15893),
.B(n_3633),
.Y(n_15961)
);

NAND2xp5_ASAP7_75t_L g15962 ( 
.A(n_15900),
.B(n_3633),
.Y(n_15962)
);

INVx1_ASAP7_75t_L g15963 ( 
.A(n_15909),
.Y(n_15963)
);

NOR2xp33_ASAP7_75t_L g15964 ( 
.A(n_15927),
.B(n_3632),
.Y(n_15964)
);

NOR2xp33_ASAP7_75t_L g15965 ( 
.A(n_15879),
.B(n_3634),
.Y(n_15965)
);

NAND4xp75_ASAP7_75t_L g15966 ( 
.A(n_15922),
.B(n_3637),
.C(n_3635),
.D(n_3636),
.Y(n_15966)
);

AND2x2_ASAP7_75t_SL g15967 ( 
.A(n_15904),
.B(n_3635),
.Y(n_15967)
);

HB1xp67_ASAP7_75t_L g15968 ( 
.A(n_15921),
.Y(n_15968)
);

NAND3xp33_ASAP7_75t_SL g15969 ( 
.A(n_15882),
.B(n_3637),
.C(n_3638),
.Y(n_15969)
);

XNOR2xp5_ASAP7_75t_L g15970 ( 
.A(n_15874),
.B(n_15918),
.Y(n_15970)
);

NAND2xp5_ASAP7_75t_L g15971 ( 
.A(n_15929),
.B(n_3641),
.Y(n_15971)
);

AND2x2_ASAP7_75t_L g15972 ( 
.A(n_15901),
.B(n_3639),
.Y(n_15972)
);

INVx1_ASAP7_75t_L g15973 ( 
.A(n_15887),
.Y(n_15973)
);

INVx1_ASAP7_75t_L g15974 ( 
.A(n_15926),
.Y(n_15974)
);

XNOR2xp5_ASAP7_75t_L g15975 ( 
.A(n_15917),
.B(n_3639),
.Y(n_15975)
);

INVx1_ASAP7_75t_L g15976 ( 
.A(n_15903),
.Y(n_15976)
);

AND2x4_ASAP7_75t_L g15977 ( 
.A(n_15912),
.B(n_3641),
.Y(n_15977)
);

OR2x2_ASAP7_75t_L g15978 ( 
.A(n_15913),
.B(n_3642),
.Y(n_15978)
);

AND3x4_ASAP7_75t_L g15979 ( 
.A(n_15881),
.B(n_3645),
.C(n_3644),
.Y(n_15979)
);

NAND3xp33_ASAP7_75t_L g15980 ( 
.A(n_15897),
.B(n_3643),
.C(n_3644),
.Y(n_15980)
);

XNOR2x1_ASAP7_75t_L g15981 ( 
.A(n_15919),
.B(n_3643),
.Y(n_15981)
);

HB1xp67_ASAP7_75t_L g15982 ( 
.A(n_15902),
.Y(n_15982)
);

NAND2xp5_ASAP7_75t_L g15983 ( 
.A(n_15890),
.B(n_3646),
.Y(n_15983)
);

INVx1_ASAP7_75t_L g15984 ( 
.A(n_15890),
.Y(n_15984)
);

INVx1_ASAP7_75t_L g15985 ( 
.A(n_15890),
.Y(n_15985)
);

NAND4xp25_ASAP7_75t_L g15986 ( 
.A(n_15922),
.B(n_3647),
.C(n_3645),
.D(n_3646),
.Y(n_15986)
);

AND2x2_ASAP7_75t_L g15987 ( 
.A(n_15928),
.B(n_3647),
.Y(n_15987)
);

XNOR2xp5_ASAP7_75t_L g15988 ( 
.A(n_15890),
.B(n_3648),
.Y(n_15988)
);

INVx2_ASAP7_75t_L g15989 ( 
.A(n_15905),
.Y(n_15989)
);

AND2x2_ASAP7_75t_L g15990 ( 
.A(n_15928),
.B(n_3648),
.Y(n_15990)
);

NAND2x1p5_ASAP7_75t_L g15991 ( 
.A(n_15906),
.B(n_3649),
.Y(n_15991)
);

OA22x2_ASAP7_75t_L g15992 ( 
.A1(n_15958),
.A2(n_3651),
.B1(n_3649),
.B2(n_3650),
.Y(n_15992)
);

NOR3x1_ASAP7_75t_L g15993 ( 
.A(n_15945),
.B(n_3650),
.C(n_3651),
.Y(n_15993)
);

AOI22xp5_ASAP7_75t_SL g15994 ( 
.A1(n_15988),
.A2(n_15947),
.B1(n_15965),
.B2(n_15987),
.Y(n_15994)
);

OAI22xp5_ASAP7_75t_L g15995 ( 
.A1(n_15938),
.A2(n_3654),
.B1(n_3652),
.B2(n_3653),
.Y(n_15995)
);

NOR4xp25_ASAP7_75t_L g15996 ( 
.A(n_15976),
.B(n_3654),
.C(n_3652),
.D(n_3653),
.Y(n_15996)
);

OAI22xp5_ASAP7_75t_L g15997 ( 
.A1(n_15980),
.A2(n_3657),
.B1(n_3655),
.B2(n_3656),
.Y(n_15997)
);

NOR2x1p5_ASAP7_75t_L g15998 ( 
.A(n_15983),
.B(n_3656),
.Y(n_15998)
);

XNOR2x2_ASAP7_75t_L g15999 ( 
.A(n_15970),
.B(n_3657),
.Y(n_15999)
);

AOI211x1_ASAP7_75t_L g16000 ( 
.A1(n_15961),
.A2(n_3660),
.B(n_3658),
.C(n_3659),
.Y(n_16000)
);

XNOR2xp5_ASAP7_75t_L g16001 ( 
.A(n_15981),
.B(n_3658),
.Y(n_16001)
);

NOR3xp33_ASAP7_75t_SL g16002 ( 
.A(n_15937),
.B(n_3659),
.C(n_3660),
.Y(n_16002)
);

XNOR2xp5_ASAP7_75t_L g16003 ( 
.A(n_15934),
.B(n_3661),
.Y(n_16003)
);

AND2x2_ASAP7_75t_L g16004 ( 
.A(n_15990),
.B(n_3662),
.Y(n_16004)
);

NAND2xp5_ASAP7_75t_SL g16005 ( 
.A(n_15956),
.B(n_3663),
.Y(n_16005)
);

NAND3xp33_ASAP7_75t_SL g16006 ( 
.A(n_15960),
.B(n_3663),
.C(n_3664),
.Y(n_16006)
);

AOI21xp5_ASAP7_75t_L g16007 ( 
.A1(n_15946),
.A2(n_3664),
.B(n_3665),
.Y(n_16007)
);

NAND4xp25_ASAP7_75t_L g16008 ( 
.A(n_15964),
.B(n_3667),
.C(n_3665),
.D(n_3666),
.Y(n_16008)
);

OAI22xp5_ASAP7_75t_L g16009 ( 
.A1(n_15955),
.A2(n_3669),
.B1(n_3666),
.B2(n_3668),
.Y(n_16009)
);

INVx1_ASAP7_75t_L g16010 ( 
.A(n_15950),
.Y(n_16010)
);

AO22x1_ASAP7_75t_L g16011 ( 
.A1(n_15944),
.A2(n_3670),
.B1(n_3668),
.B2(n_3669),
.Y(n_16011)
);

NAND3xp33_ASAP7_75t_SL g16012 ( 
.A(n_15991),
.B(n_3670),
.C(n_3671),
.Y(n_16012)
);

AOI211xp5_ASAP7_75t_L g16013 ( 
.A1(n_15942),
.A2(n_15974),
.B(n_15940),
.C(n_15969),
.Y(n_16013)
);

INVx1_ASAP7_75t_L g16014 ( 
.A(n_15967),
.Y(n_16014)
);

NAND5xp2_ASAP7_75t_L g16015 ( 
.A(n_15933),
.B(n_15984),
.C(n_15985),
.D(n_15957),
.E(n_15973),
.Y(n_16015)
);

XNOR2x1_ASAP7_75t_L g16016 ( 
.A(n_15941),
.B(n_15989),
.Y(n_16016)
);

OA22x2_ASAP7_75t_L g16017 ( 
.A1(n_15979),
.A2(n_3673),
.B1(n_3671),
.B2(n_3672),
.Y(n_16017)
);

OAI222xp33_ASAP7_75t_L g16018 ( 
.A1(n_15951),
.A2(n_3674),
.B1(n_3676),
.B2(n_3672),
.C1(n_3673),
.C2(n_3675),
.Y(n_16018)
);

INVx1_ASAP7_75t_L g16019 ( 
.A(n_15962),
.Y(n_16019)
);

AOI22xp5_ASAP7_75t_L g16020 ( 
.A1(n_15936),
.A2(n_3676),
.B1(n_3674),
.B2(n_3675),
.Y(n_16020)
);

AOI211xp5_ASAP7_75t_SL g16021 ( 
.A1(n_15982),
.A2(n_3686),
.B(n_3694),
.C(n_3677),
.Y(n_16021)
);

NAND3xp33_ASAP7_75t_SL g16022 ( 
.A(n_15935),
.B(n_3677),
.C(n_3678),
.Y(n_16022)
);

OAI322xp33_ASAP7_75t_L g16023 ( 
.A1(n_15963),
.A2(n_3684),
.A3(n_3683),
.B1(n_3681),
.B2(n_3678),
.C1(n_3679),
.C2(n_3682),
.Y(n_16023)
);

NOR2x1p5_ASAP7_75t_L g16024 ( 
.A(n_15953),
.B(n_3679),
.Y(n_16024)
);

AOI22xp5_ASAP7_75t_L g16025 ( 
.A1(n_15948),
.A2(n_15954),
.B1(n_15968),
.B2(n_15952),
.Y(n_16025)
);

NAND3xp33_ASAP7_75t_L g16026 ( 
.A(n_15931),
.B(n_3681),
.C(n_3683),
.Y(n_16026)
);

AOI21xp5_ASAP7_75t_L g16027 ( 
.A1(n_15975),
.A2(n_3684),
.B(n_3685),
.Y(n_16027)
);

INVx1_ASAP7_75t_L g16028 ( 
.A(n_15932),
.Y(n_16028)
);

INVx1_ASAP7_75t_L g16029 ( 
.A(n_15966),
.Y(n_16029)
);

AND2x4_ASAP7_75t_L g16030 ( 
.A(n_15943),
.B(n_4057),
.Y(n_16030)
);

XNOR2x1_ASAP7_75t_L g16031 ( 
.A(n_15949),
.B(n_3687),
.Y(n_16031)
);

NAND3xp33_ASAP7_75t_L g16032 ( 
.A(n_15986),
.B(n_3688),
.C(n_3689),
.Y(n_16032)
);

NOR4xp25_ASAP7_75t_L g16033 ( 
.A(n_15971),
.B(n_3690),
.C(n_3688),
.D(n_3689),
.Y(n_16033)
);

OR2x2_ASAP7_75t_L g16034 ( 
.A(n_15978),
.B(n_3691),
.Y(n_16034)
);

NAND3xp33_ASAP7_75t_L g16035 ( 
.A(n_15939),
.B(n_15972),
.C(n_15977),
.Y(n_16035)
);

OAI22xp5_ASAP7_75t_L g16036 ( 
.A1(n_15959),
.A2(n_3693),
.B1(n_3691),
.B2(n_3692),
.Y(n_16036)
);

INVx1_ASAP7_75t_L g16037 ( 
.A(n_15958),
.Y(n_16037)
);

AND2x4_ASAP7_75t_L g16038 ( 
.A(n_15987),
.B(n_4068),
.Y(n_16038)
);

NAND2xp5_ASAP7_75t_L g16039 ( 
.A(n_15956),
.B(n_3692),
.Y(n_16039)
);

AOI221xp5_ASAP7_75t_L g16040 ( 
.A1(n_15965),
.A2(n_3696),
.B1(n_3694),
.B2(n_3695),
.C(n_3697),
.Y(n_16040)
);

AO22x2_ASAP7_75t_L g16041 ( 
.A1(n_15946),
.A2(n_3703),
.B1(n_3712),
.B2(n_3695),
.Y(n_16041)
);

INVx1_ASAP7_75t_L g16042 ( 
.A(n_15958),
.Y(n_16042)
);

INVx1_ASAP7_75t_L g16043 ( 
.A(n_15958),
.Y(n_16043)
);

AOI211x1_ASAP7_75t_SL g16044 ( 
.A1(n_15937),
.A2(n_3698),
.B(n_3696),
.C(n_3697),
.Y(n_16044)
);

AND2x2_ASAP7_75t_L g16045 ( 
.A(n_15987),
.B(n_3698),
.Y(n_16045)
);

INVx1_ASAP7_75t_L g16046 ( 
.A(n_15958),
.Y(n_16046)
);

INVx2_ASAP7_75t_L g16047 ( 
.A(n_15932),
.Y(n_16047)
);

NAND3xp33_ASAP7_75t_L g16048 ( 
.A(n_15934),
.B(n_3699),
.C(n_3700),
.Y(n_16048)
);

AOI221xp5_ASAP7_75t_L g16049 ( 
.A1(n_15965),
.A2(n_3701),
.B1(n_3699),
.B2(n_3700),
.C(n_3702),
.Y(n_16049)
);

AOI22xp5_ASAP7_75t_L g16050 ( 
.A1(n_15934),
.A2(n_3705),
.B1(n_3702),
.B2(n_3704),
.Y(n_16050)
);

INVx1_ASAP7_75t_L g16051 ( 
.A(n_15958),
.Y(n_16051)
);

INVx1_ASAP7_75t_L g16052 ( 
.A(n_15958),
.Y(n_16052)
);

AND3x2_ASAP7_75t_L g16053 ( 
.A(n_15982),
.B(n_3705),
.C(n_3706),
.Y(n_16053)
);

NAND4xp25_ASAP7_75t_L g16054 ( 
.A(n_15934),
.B(n_3709),
.C(n_3706),
.D(n_3708),
.Y(n_16054)
);

AOI22xp5_ASAP7_75t_L g16055 ( 
.A1(n_15934),
.A2(n_3710),
.B1(n_3708),
.B2(n_3709),
.Y(n_16055)
);

AOI211xp5_ASAP7_75t_SL g16056 ( 
.A1(n_15934),
.A2(n_3718),
.B(n_3727),
.C(n_3710),
.Y(n_16056)
);

INVx1_ASAP7_75t_L g16057 ( 
.A(n_15958),
.Y(n_16057)
);

NOR2xp33_ASAP7_75t_L g16058 ( 
.A(n_15983),
.B(n_3711),
.Y(n_16058)
);

NAND4xp25_ASAP7_75t_L g16059 ( 
.A(n_15934),
.B(n_3713),
.C(n_3711),
.D(n_3712),
.Y(n_16059)
);

INVxp33_ASAP7_75t_SL g16060 ( 
.A(n_15982),
.Y(n_16060)
);

NOR3xp33_ASAP7_75t_L g16061 ( 
.A(n_15934),
.B(n_3713),
.C(n_3714),
.Y(n_16061)
);

OAI22xp5_ASAP7_75t_SL g16062 ( 
.A1(n_16060),
.A2(n_3723),
.B1(n_3732),
.B2(n_3714),
.Y(n_16062)
);

NOR4xp25_ASAP7_75t_L g16063 ( 
.A(n_16010),
.B(n_3717),
.C(n_3715),
.D(n_3716),
.Y(n_16063)
);

OAI221xp5_ASAP7_75t_L g16064 ( 
.A1(n_16001),
.A2(n_3718),
.B1(n_3716),
.B2(n_3717),
.C(n_3719),
.Y(n_16064)
);

INVx1_ASAP7_75t_L g16065 ( 
.A(n_16031),
.Y(n_16065)
);

AND2x4_ASAP7_75t_L g16066 ( 
.A(n_15998),
.B(n_3720),
.Y(n_16066)
);

AOI22xp5_ASAP7_75t_L g16067 ( 
.A1(n_16006),
.A2(n_3723),
.B1(n_3720),
.B2(n_3722),
.Y(n_16067)
);

INVx1_ASAP7_75t_SL g16068 ( 
.A(n_15999),
.Y(n_16068)
);

NAND2xp5_ASAP7_75t_L g16069 ( 
.A(n_16058),
.B(n_4067),
.Y(n_16069)
);

INVx1_ASAP7_75t_L g16070 ( 
.A(n_16039),
.Y(n_16070)
);

AOI22x1_ASAP7_75t_L g16071 ( 
.A1(n_15994),
.A2(n_3726),
.B1(n_3724),
.B2(n_3725),
.Y(n_16071)
);

INVx2_ASAP7_75t_L g16072 ( 
.A(n_16053),
.Y(n_16072)
);

NAND2xp5_ASAP7_75t_L g16073 ( 
.A(n_16000),
.B(n_4050),
.Y(n_16073)
);

BUFx2_ASAP7_75t_L g16074 ( 
.A(n_16017),
.Y(n_16074)
);

INVxp33_ASAP7_75t_SL g16075 ( 
.A(n_16025),
.Y(n_16075)
);

AOI22xp5_ASAP7_75t_L g16076 ( 
.A1(n_16012),
.A2(n_3730),
.B1(n_3728),
.B2(n_3729),
.Y(n_16076)
);

OR2x2_ASAP7_75t_L g16077 ( 
.A(n_16022),
.B(n_3731),
.Y(n_16077)
);

OA21x2_ASAP7_75t_L g16078 ( 
.A1(n_16014),
.A2(n_3731),
.B(n_3733),
.Y(n_16078)
);

AOI22xp33_ASAP7_75t_L g16079 ( 
.A1(n_16032),
.A2(n_3737),
.B1(n_3734),
.B2(n_3735),
.Y(n_16079)
);

INVx1_ASAP7_75t_L g16080 ( 
.A(n_15992),
.Y(n_16080)
);

INVx1_ASAP7_75t_L g16081 ( 
.A(n_16005),
.Y(n_16081)
);

AOI21xp5_ASAP7_75t_L g16082 ( 
.A1(n_16016),
.A2(n_3735),
.B(n_3737),
.Y(n_16082)
);

AOI211xp5_ASAP7_75t_L g16083 ( 
.A1(n_16015),
.A2(n_3740),
.B(n_3738),
.C(n_3739),
.Y(n_16083)
);

OAI22xp5_ASAP7_75t_L g16084 ( 
.A1(n_16026),
.A2(n_3741),
.B1(n_3742),
.B2(n_3740),
.Y(n_16084)
);

NAND2xp5_ASAP7_75t_L g16085 ( 
.A(n_16002),
.B(n_4061),
.Y(n_16085)
);

OAI22xp5_ASAP7_75t_SL g16086 ( 
.A1(n_16029),
.A2(n_16035),
.B1(n_16028),
.B2(n_16047),
.Y(n_16086)
);

NAND2xp5_ASAP7_75t_SL g16087 ( 
.A(n_16027),
.B(n_3739),
.Y(n_16087)
);

OAI22xp5_ASAP7_75t_L g16088 ( 
.A1(n_15997),
.A2(n_3743),
.B1(n_3744),
.B2(n_3742),
.Y(n_16088)
);

O2A1O1Ixp33_ASAP7_75t_L g16089 ( 
.A1(n_16037),
.A2(n_3745),
.B(n_3746),
.C(n_3744),
.Y(n_16089)
);

AOI22x1_ASAP7_75t_L g16090 ( 
.A1(n_16042),
.A2(n_3748),
.B1(n_3741),
.B2(n_3747),
.Y(n_16090)
);

NOR2xp67_ASAP7_75t_L g16091 ( 
.A(n_16043),
.B(n_4052),
.Y(n_16091)
);

INVx2_ASAP7_75t_L g16092 ( 
.A(n_16024),
.Y(n_16092)
);

OAI22xp5_ASAP7_75t_SL g16093 ( 
.A1(n_16046),
.A2(n_3756),
.B1(n_3765),
.B2(n_3747),
.Y(n_16093)
);

XNOR2xp5_ASAP7_75t_L g16094 ( 
.A(n_16013),
.B(n_3748),
.Y(n_16094)
);

NOR3xp33_ASAP7_75t_SL g16095 ( 
.A(n_16051),
.B(n_3758),
.C(n_3749),
.Y(n_16095)
);

NAND2xp5_ASAP7_75t_L g16096 ( 
.A(n_16044),
.B(n_4054),
.Y(n_16096)
);

NAND3xp33_ASAP7_75t_L g16097 ( 
.A(n_16052),
.B(n_3749),
.C(n_3750),
.Y(n_16097)
);

AOI22xp5_ASAP7_75t_L g16098 ( 
.A1(n_16057),
.A2(n_16061),
.B1(n_16019),
.B2(n_16008),
.Y(n_16098)
);

NAND4xp25_ASAP7_75t_L g16099 ( 
.A(n_15993),
.B(n_3754),
.C(n_3752),
.D(n_3753),
.Y(n_16099)
);

INVx1_ASAP7_75t_L g16100 ( 
.A(n_16003),
.Y(n_16100)
);

OAI22xp5_ASAP7_75t_L g16101 ( 
.A1(n_16048),
.A2(n_3754),
.B1(n_3755),
.B2(n_3753),
.Y(n_16101)
);

INVx2_ASAP7_75t_L g16102 ( 
.A(n_16038),
.Y(n_16102)
);

INVx2_ASAP7_75t_L g16103 ( 
.A(n_16038),
.Y(n_16103)
);

NAND2xp5_ASAP7_75t_SL g16104 ( 
.A(n_16033),
.B(n_3752),
.Y(n_16104)
);

BUFx3_ASAP7_75t_L g16105 ( 
.A(n_16030),
.Y(n_16105)
);

OAI21xp33_ASAP7_75t_L g16106 ( 
.A1(n_15996),
.A2(n_16049),
.B(n_16040),
.Y(n_16106)
);

OAI22xp5_ASAP7_75t_SL g16107 ( 
.A1(n_16075),
.A2(n_16034),
.B1(n_16030),
.B2(n_16009),
.Y(n_16107)
);

NAND4xp75_ASAP7_75t_L g16108 ( 
.A(n_16098),
.B(n_16007),
.C(n_16045),
.D(n_16004),
.Y(n_16108)
);

NOR3xp33_ASAP7_75t_SL g16109 ( 
.A(n_16086),
.B(n_16018),
.C(n_16054),
.Y(n_16109)
);

OAI21xp5_ASAP7_75t_L g16110 ( 
.A1(n_16085),
.A2(n_16056),
.B(n_16021),
.Y(n_16110)
);

INVx2_ASAP7_75t_L g16111 ( 
.A(n_16071),
.Y(n_16111)
);

HB1xp67_ASAP7_75t_L g16112 ( 
.A(n_16094),
.Y(n_16112)
);

INVx2_ASAP7_75t_L g16113 ( 
.A(n_16090),
.Y(n_16113)
);

INVx1_ASAP7_75t_SL g16114 ( 
.A(n_16105),
.Y(n_16114)
);

INVx2_ASAP7_75t_SL g16115 ( 
.A(n_16066),
.Y(n_16115)
);

INVx1_ASAP7_75t_L g16116 ( 
.A(n_16066),
.Y(n_16116)
);

NAND2x1_ASAP7_75t_L g16117 ( 
.A(n_16073),
.B(n_16036),
.Y(n_16117)
);

INVx2_ASAP7_75t_L g16118 ( 
.A(n_16078),
.Y(n_16118)
);

INVx1_ASAP7_75t_L g16119 ( 
.A(n_16096),
.Y(n_16119)
);

OA22x2_ASAP7_75t_SL g16120 ( 
.A1(n_16088),
.A2(n_15995),
.B1(n_16011),
.B2(n_16059),
.Y(n_16120)
);

INVx3_ASAP7_75t_L g16121 ( 
.A(n_16077),
.Y(n_16121)
);

INVx1_ASAP7_75t_L g16122 ( 
.A(n_16099),
.Y(n_16122)
);

INVx2_ASAP7_75t_L g16123 ( 
.A(n_16078),
.Y(n_16123)
);

NAND2xp5_ASAP7_75t_L g16124 ( 
.A(n_16083),
.B(n_16050),
.Y(n_16124)
);

NAND2xp5_ASAP7_75t_L g16125 ( 
.A(n_16076),
.B(n_16055),
.Y(n_16125)
);

XNOR2xp5_ASAP7_75t_L g16126 ( 
.A(n_16104),
.B(n_16020),
.Y(n_16126)
);

BUFx2_ASAP7_75t_L g16127 ( 
.A(n_16095),
.Y(n_16127)
);

NOR2x1p5_ASAP7_75t_L g16128 ( 
.A(n_16102),
.B(n_16023),
.Y(n_16128)
);

INVx1_ASAP7_75t_L g16129 ( 
.A(n_16091),
.Y(n_16129)
);

NAND2xp5_ASAP7_75t_L g16130 ( 
.A(n_16067),
.B(n_16041),
.Y(n_16130)
);

XNOR2x1_ASAP7_75t_L g16131 ( 
.A(n_16065),
.B(n_16041),
.Y(n_16131)
);

AO22x2_ASAP7_75t_L g16132 ( 
.A1(n_16103),
.A2(n_3757),
.B1(n_3755),
.B2(n_3756),
.Y(n_16132)
);

XOR2xp5_ASAP7_75t_L g16133 ( 
.A(n_16100),
.B(n_3758),
.Y(n_16133)
);

XNOR2x1_ASAP7_75t_L g16134 ( 
.A(n_16072),
.B(n_3757),
.Y(n_16134)
);

INVx1_ASAP7_75t_L g16135 ( 
.A(n_16087),
.Y(n_16135)
);

XNOR2x1_ASAP7_75t_L g16136 ( 
.A(n_16092),
.B(n_3759),
.Y(n_16136)
);

AO22x2_ASAP7_75t_L g16137 ( 
.A1(n_16108),
.A2(n_16080),
.B1(n_16068),
.B2(n_16081),
.Y(n_16137)
);

INVx1_ASAP7_75t_L g16138 ( 
.A(n_16118),
.Y(n_16138)
);

NOR3xp33_ASAP7_75t_L g16139 ( 
.A(n_16114),
.B(n_16070),
.C(n_16074),
.Y(n_16139)
);

INVx1_ASAP7_75t_L g16140 ( 
.A(n_16123),
.Y(n_16140)
);

HB1xp67_ASAP7_75t_L g16141 ( 
.A(n_16128),
.Y(n_16141)
);

INVx1_ASAP7_75t_L g16142 ( 
.A(n_16130),
.Y(n_16142)
);

INVx1_ASAP7_75t_L g16143 ( 
.A(n_16116),
.Y(n_16143)
);

INVxp67_ASAP7_75t_L g16144 ( 
.A(n_16127),
.Y(n_16144)
);

AO21x2_ASAP7_75t_L g16145 ( 
.A1(n_16119),
.A2(n_16106),
.B(n_16082),
.Y(n_16145)
);

XNOR2xp5_ASAP7_75t_L g16146 ( 
.A(n_16131),
.B(n_16126),
.Y(n_16146)
);

INVx1_ASAP7_75t_L g16147 ( 
.A(n_16124),
.Y(n_16147)
);

INVx3_ASAP7_75t_L g16148 ( 
.A(n_16117),
.Y(n_16148)
);

INVx1_ASAP7_75t_L g16149 ( 
.A(n_16129),
.Y(n_16149)
);

INVx2_ASAP7_75t_L g16150 ( 
.A(n_16134),
.Y(n_16150)
);

AOI211xp5_ASAP7_75t_SL g16151 ( 
.A1(n_16107),
.A2(n_16084),
.B(n_16101),
.C(n_16064),
.Y(n_16151)
);

INVx1_ASAP7_75t_L g16152 ( 
.A(n_16115),
.Y(n_16152)
);

AO22x2_ASAP7_75t_L g16153 ( 
.A1(n_16122),
.A2(n_16135),
.B1(n_16111),
.B2(n_16113),
.Y(n_16153)
);

INVx2_ASAP7_75t_L g16154 ( 
.A(n_16136),
.Y(n_16154)
);

AND2x2_ASAP7_75t_L g16155 ( 
.A(n_16110),
.B(n_16079),
.Y(n_16155)
);

AOI22x1_ASAP7_75t_L g16156 ( 
.A1(n_16112),
.A2(n_16089),
.B1(n_16063),
.B2(n_16097),
.Y(n_16156)
);

OAI22x1_ASAP7_75t_L g16157 ( 
.A1(n_16121),
.A2(n_16069),
.B1(n_16062),
.B2(n_16093),
.Y(n_16157)
);

INVx2_ASAP7_75t_L g16158 ( 
.A(n_16120),
.Y(n_16158)
);

NOR2xp33_ASAP7_75t_L g16159 ( 
.A(n_16148),
.B(n_16125),
.Y(n_16159)
);

OAI22xp5_ASAP7_75t_SL g16160 ( 
.A1(n_16143),
.A2(n_16109),
.B1(n_16133),
.B2(n_16132),
.Y(n_16160)
);

INVx3_ASAP7_75t_L g16161 ( 
.A(n_16158),
.Y(n_16161)
);

INVx1_ASAP7_75t_L g16162 ( 
.A(n_16137),
.Y(n_16162)
);

INVx1_ASAP7_75t_L g16163 ( 
.A(n_16141),
.Y(n_16163)
);

AO22x2_ASAP7_75t_L g16164 ( 
.A1(n_16138),
.A2(n_16140),
.B1(n_16152),
.B2(n_16142),
.Y(n_16164)
);

NAND2xp5_ASAP7_75t_L g16165 ( 
.A(n_16139),
.B(n_16132),
.Y(n_16165)
);

AOI22xp5_ASAP7_75t_SL g16166 ( 
.A1(n_16157),
.A2(n_3761),
.B1(n_3759),
.B2(n_3760),
.Y(n_16166)
);

A2O1A1Ixp33_ASAP7_75t_SL g16167 ( 
.A1(n_16144),
.A2(n_3762),
.B(n_3760),
.C(n_3761),
.Y(n_16167)
);

OAI22xp33_ASAP7_75t_L g16168 ( 
.A1(n_16151),
.A2(n_3766),
.B1(n_3763),
.B2(n_3765),
.Y(n_16168)
);

INVx1_ASAP7_75t_L g16169 ( 
.A(n_16146),
.Y(n_16169)
);

AOI22xp33_ASAP7_75t_L g16170 ( 
.A1(n_16149),
.A2(n_3769),
.B1(n_3767),
.B2(n_3768),
.Y(n_16170)
);

AOI31xp33_ASAP7_75t_L g16171 ( 
.A1(n_16147),
.A2(n_3777),
.A3(n_3785),
.B(n_3767),
.Y(n_16171)
);

AOI22xp5_ASAP7_75t_L g16172 ( 
.A1(n_16153),
.A2(n_3771),
.B1(n_3772),
.B2(n_3769),
.Y(n_16172)
);

AOI31xp33_ASAP7_75t_L g16173 ( 
.A1(n_16154),
.A2(n_3781),
.A3(n_3789),
.B(n_3768),
.Y(n_16173)
);

AOI22xp5_ASAP7_75t_L g16174 ( 
.A1(n_16150),
.A2(n_3774),
.B1(n_3776),
.B2(n_3773),
.Y(n_16174)
);

OAI31xp33_ASAP7_75t_L g16175 ( 
.A1(n_16155),
.A2(n_3776),
.A3(n_3771),
.B(n_3774),
.Y(n_16175)
);

AOI22xp33_ASAP7_75t_SL g16176 ( 
.A1(n_16156),
.A2(n_3780),
.B1(n_3781),
.B2(n_3779),
.Y(n_16176)
);

OAI22xp5_ASAP7_75t_L g16177 ( 
.A1(n_16145),
.A2(n_3780),
.B1(n_3778),
.B2(n_3779),
.Y(n_16177)
);

AO22x2_ASAP7_75t_L g16178 ( 
.A1(n_16138),
.A2(n_3783),
.B1(n_3778),
.B2(n_3782),
.Y(n_16178)
);

AOI22xp5_ASAP7_75t_L g16179 ( 
.A1(n_16139),
.A2(n_3784),
.B1(n_3785),
.B2(n_3783),
.Y(n_16179)
);

OAI22xp5_ASAP7_75t_SL g16180 ( 
.A1(n_16143),
.A2(n_3786),
.B1(n_3782),
.B2(n_3784),
.Y(n_16180)
);

AO22x2_ASAP7_75t_L g16181 ( 
.A1(n_16162),
.A2(n_4057),
.B1(n_4059),
.B2(n_4056),
.Y(n_16181)
);

NAND2xp5_ASAP7_75t_L g16182 ( 
.A(n_16161),
.B(n_3786),
.Y(n_16182)
);

XNOR2xp5_ASAP7_75t_L g16183 ( 
.A(n_16169),
.B(n_3788),
.Y(n_16183)
);

NOR2xp67_ASAP7_75t_L g16184 ( 
.A(n_16163),
.B(n_16165),
.Y(n_16184)
);

OA21x2_ASAP7_75t_L g16185 ( 
.A1(n_16159),
.A2(n_3797),
.B(n_3787),
.Y(n_16185)
);

AOI21xp5_ASAP7_75t_L g16186 ( 
.A1(n_16164),
.A2(n_3787),
.B(n_3788),
.Y(n_16186)
);

NAND4xp25_ASAP7_75t_L g16187 ( 
.A(n_16160),
.B(n_3793),
.C(n_3790),
.D(n_3791),
.Y(n_16187)
);

AOI31xp33_ASAP7_75t_L g16188 ( 
.A1(n_16176),
.A2(n_3794),
.A3(n_3790),
.B(n_3791),
.Y(n_16188)
);

NAND3xp33_ASAP7_75t_SL g16189 ( 
.A(n_16175),
.B(n_3794),
.C(n_3795),
.Y(n_16189)
);

XOR2xp5_ASAP7_75t_L g16190 ( 
.A(n_16177),
.B(n_16166),
.Y(n_16190)
);

OA22x2_ASAP7_75t_L g16191 ( 
.A1(n_16172),
.A2(n_3798),
.B1(n_3795),
.B2(n_3796),
.Y(n_16191)
);

OAI22xp5_ASAP7_75t_L g16192 ( 
.A1(n_16179),
.A2(n_3799),
.B1(n_3796),
.B2(n_3798),
.Y(n_16192)
);

INVx2_ASAP7_75t_L g16193 ( 
.A(n_16178),
.Y(n_16193)
);

AOI21x1_ASAP7_75t_L g16194 ( 
.A1(n_16167),
.A2(n_4063),
.B(n_4051),
.Y(n_16194)
);

NAND3xp33_ASAP7_75t_L g16195 ( 
.A(n_16168),
.B(n_16174),
.C(n_16173),
.Y(n_16195)
);

AOI21xp5_ASAP7_75t_L g16196 ( 
.A1(n_16171),
.A2(n_3799),
.B(n_3800),
.Y(n_16196)
);

INVx2_ASAP7_75t_L g16197 ( 
.A(n_16180),
.Y(n_16197)
);

INVx1_ASAP7_75t_L g16198 ( 
.A(n_16170),
.Y(n_16198)
);

OAI22xp5_ASAP7_75t_L g16199 ( 
.A1(n_16184),
.A2(n_3802),
.B1(n_3800),
.B2(n_3801),
.Y(n_16199)
);

OAI22xp5_ASAP7_75t_SL g16200 ( 
.A1(n_16193),
.A2(n_3803),
.B1(n_3804),
.B2(n_3802),
.Y(n_16200)
);

XOR2xp5_ASAP7_75t_L g16201 ( 
.A(n_16190),
.B(n_3801),
.Y(n_16201)
);

INVx1_ASAP7_75t_L g16202 ( 
.A(n_16195),
.Y(n_16202)
);

OAI22xp5_ASAP7_75t_SL g16203 ( 
.A1(n_16197),
.A2(n_3805),
.B1(n_3806),
.B2(n_3804),
.Y(n_16203)
);

NAND2xp5_ASAP7_75t_L g16204 ( 
.A(n_16198),
.B(n_4060),
.Y(n_16204)
);

OAI22xp5_ASAP7_75t_SL g16205 ( 
.A1(n_16192),
.A2(n_3807),
.B1(n_3808),
.B2(n_3805),
.Y(n_16205)
);

OAI22xp5_ASAP7_75t_L g16206 ( 
.A1(n_16196),
.A2(n_3808),
.B1(n_3803),
.B2(n_3807),
.Y(n_16206)
);

INVx1_ASAP7_75t_L g16207 ( 
.A(n_16189),
.Y(n_16207)
);

OAI22xp5_ASAP7_75t_SL g16208 ( 
.A1(n_16194),
.A2(n_3811),
.B1(n_3813),
.B2(n_3810),
.Y(n_16208)
);

NAND2xp5_ASAP7_75t_L g16209 ( 
.A(n_16188),
.B(n_4047),
.Y(n_16209)
);

INVx3_ASAP7_75t_L g16210 ( 
.A(n_16191),
.Y(n_16210)
);

CKINVDCx16_ASAP7_75t_R g16211 ( 
.A(n_16183),
.Y(n_16211)
);

OAI22xp5_ASAP7_75t_SL g16212 ( 
.A1(n_16185),
.A2(n_3811),
.B1(n_3813),
.B2(n_3810),
.Y(n_16212)
);

AOI22xp5_ASAP7_75t_L g16213 ( 
.A1(n_16202),
.A2(n_16186),
.B1(n_16187),
.B2(n_16181),
.Y(n_16213)
);

INVx2_ASAP7_75t_L g16214 ( 
.A(n_16209),
.Y(n_16214)
);

INVx1_ASAP7_75t_L g16215 ( 
.A(n_16210),
.Y(n_16215)
);

OAI22xp33_ASAP7_75t_L g16216 ( 
.A1(n_16211),
.A2(n_16182),
.B1(n_3815),
.B2(n_3809),
.Y(n_16216)
);

INVx1_ASAP7_75t_L g16217 ( 
.A(n_16210),
.Y(n_16217)
);

AO22x2_ASAP7_75t_L g16218 ( 
.A1(n_16207),
.A2(n_3816),
.B1(n_3814),
.B2(n_3815),
.Y(n_16218)
);

OAI21xp5_ASAP7_75t_L g16219 ( 
.A1(n_16206),
.A2(n_3814),
.B(n_3817),
.Y(n_16219)
);

OAI22x1_ASAP7_75t_L g16220 ( 
.A1(n_16208),
.A2(n_3819),
.B1(n_3817),
.B2(n_3818),
.Y(n_16220)
);

OAI21xp5_ASAP7_75t_L g16221 ( 
.A1(n_16199),
.A2(n_3819),
.B(n_3820),
.Y(n_16221)
);

CKINVDCx5p33_ASAP7_75t_R g16222 ( 
.A(n_16205),
.Y(n_16222)
);

AO21x2_ASAP7_75t_L g16223 ( 
.A1(n_16212),
.A2(n_3829),
.B(n_3820),
.Y(n_16223)
);

INVx3_ASAP7_75t_L g16224 ( 
.A(n_16215),
.Y(n_16224)
);

AOI222xp33_ASAP7_75t_L g16225 ( 
.A1(n_16217),
.A2(n_16200),
.B1(n_16203),
.B2(n_16204),
.C1(n_16201),
.C2(n_3823),
.Y(n_16225)
);

OAI22xp33_ASAP7_75t_L g16226 ( 
.A1(n_16213),
.A2(n_3823),
.B1(n_3821),
.B2(n_3822),
.Y(n_16226)
);

XNOR2xp5_ASAP7_75t_L g16227 ( 
.A(n_16222),
.B(n_3822),
.Y(n_16227)
);

NAND3xp33_ASAP7_75t_L g16228 ( 
.A(n_16214),
.B(n_3821),
.C(n_3824),
.Y(n_16228)
);

OAI21xp5_ASAP7_75t_L g16229 ( 
.A1(n_16221),
.A2(n_3825),
.B(n_3827),
.Y(n_16229)
);

AOI21xp5_ASAP7_75t_L g16230 ( 
.A1(n_16224),
.A2(n_16219),
.B(n_16223),
.Y(n_16230)
);

NAND2xp5_ASAP7_75t_L g16231 ( 
.A(n_16225),
.B(n_16220),
.Y(n_16231)
);

OAI21xp33_ASAP7_75t_L g16232 ( 
.A1(n_16229),
.A2(n_16216),
.B(n_16226),
.Y(n_16232)
);

NAND2xp5_ASAP7_75t_L g16233 ( 
.A(n_16228),
.B(n_16218),
.Y(n_16233)
);

AOI22xp33_ASAP7_75t_L g16234 ( 
.A1(n_16227),
.A2(n_16218),
.B1(n_3830),
.B2(n_3827),
.Y(n_16234)
);

OAI21xp5_ASAP7_75t_L g16235 ( 
.A1(n_16224),
.A2(n_4049),
.B(n_4048),
.Y(n_16235)
);

AOI21xp5_ASAP7_75t_L g16236 ( 
.A1(n_16231),
.A2(n_3828),
.B(n_3830),
.Y(n_16236)
);

AOI222xp33_ASAP7_75t_SL g16237 ( 
.A1(n_16230),
.A2(n_3832),
.B1(n_3834),
.B2(n_3828),
.C1(n_3831),
.C2(n_3833),
.Y(n_16237)
);

OAI222xp33_ASAP7_75t_L g16238 ( 
.A1(n_16233),
.A2(n_3833),
.B1(n_3836),
.B2(n_3837),
.C1(n_3832),
.C2(n_3835),
.Y(n_16238)
);

AOI22xp33_ASAP7_75t_SL g16239 ( 
.A1(n_16232),
.A2(n_3836),
.B1(n_3831),
.B2(n_3835),
.Y(n_16239)
);

AOI21x1_ASAP7_75t_L g16240 ( 
.A1(n_16236),
.A2(n_16234),
.B(n_16235),
.Y(n_16240)
);

A2O1A1Ixp33_ASAP7_75t_L g16241 ( 
.A1(n_16239),
.A2(n_3840),
.B(n_3838),
.C(n_3839),
.Y(n_16241)
);

AOI322xp5_ASAP7_75t_L g16242 ( 
.A1(n_16240),
.A2(n_16237),
.A3(n_16238),
.B1(n_3843),
.B2(n_3840),
.C1(n_3842),
.C2(n_3838),
.Y(n_16242)
);

AOI22xp5_ASAP7_75t_L g16243 ( 
.A1(n_16241),
.A2(n_3842),
.B1(n_3839),
.B2(n_3841),
.Y(n_16243)
);

AOI21xp33_ASAP7_75t_SL g16244 ( 
.A1(n_16243),
.A2(n_3841),
.B(n_3843),
.Y(n_16244)
);

NAND2xp5_ASAP7_75t_L g16245 ( 
.A(n_16242),
.B(n_3844),
.Y(n_16245)
);

AOI22xp5_ASAP7_75t_L g16246 ( 
.A1(n_16245),
.A2(n_16244),
.B1(n_3846),
.B2(n_3844),
.Y(n_16246)
);

AOI22xp5_ASAP7_75t_L g16247 ( 
.A1(n_16245),
.A2(n_3847),
.B1(n_3845),
.B2(n_3846),
.Y(n_16247)
);

AOI22xp33_ASAP7_75t_L g16248 ( 
.A1(n_16246),
.A2(n_3849),
.B1(n_3845),
.B2(n_3848),
.Y(n_16248)
);

AOI211xp5_ASAP7_75t_L g16249 ( 
.A1(n_16248),
.A2(n_16247),
.B(n_3850),
.C(n_3848),
.Y(n_16249)
);


endmodule