module fake_jpeg_13827_n_127 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_127);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_127;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_4),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_27),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_32),
.B(n_34),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_0),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_2),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_38),
.Y(n_41)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_15),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_44),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_50),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_26),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_53),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_26),
.Y(n_53)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_57),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_20),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_19),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_35),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_63),
.A2(n_67),
.B(n_68),
.Y(n_81)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

CKINVDCx10_ASAP7_75t_R g87 ( 
.A(n_65),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVxp33_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

HAxp5_ASAP7_75t_SL g67 ( 
.A(n_54),
.B(n_31),
.CON(n_67),
.SN(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_16),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVxp33_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_72),
.B1(n_73),
.B2(n_55),
.Y(n_77)
);

INVxp33_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_52),
.A2(n_32),
.B1(n_29),
.B2(n_28),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_15),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_74),
.A2(n_16),
.B1(n_19),
.B2(n_17),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_72),
.A2(n_44),
.B1(n_49),
.B2(n_47),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_78),
.B1(n_80),
.B2(n_82),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_79),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_54),
.B1(n_48),
.B2(n_36),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_62),
.A2(n_20),
.B1(n_14),
.B2(n_17),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_62),
.A2(n_73),
.B1(n_66),
.B2(n_64),
.Y(n_82)
);

AND2x6_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_3),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_6),
.Y(n_96)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_60),
.C(n_71),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_92),
.Y(n_103)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_71),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_76),
.B(n_65),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_97),
.Y(n_99)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

AOI21xp33_ASAP7_75t_L g102 ( 
.A1(n_95),
.A2(n_96),
.B(n_6),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_55),
.C(n_61),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_14),
.C(n_45),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_84),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_89),
.A2(n_83),
.B1(n_84),
.B2(n_69),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_100),
.A2(n_94),
.B1(n_98),
.B2(n_21),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_90),
.A2(n_97),
.B(n_93),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_95),
.B(n_59),
.Y(n_111)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_93),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_7),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_88),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_109),
.B(n_105),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_110),
.A2(n_111),
.B(n_99),
.Y(n_114)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_101),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_115),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_114),
.B(n_116),
.Y(n_119)
);

FAx1_ASAP7_75t_SL g115 ( 
.A(n_110),
.B(n_99),
.CI(n_103),
.CON(n_115),
.SN(n_115)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_108),
.Y(n_121)
);

NOR2xp67_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_117),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_10),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_8),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_120),
.B1(n_119),
.B2(n_118),
.Y(n_125)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_123),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_9),
.B(n_124),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_9),
.Y(n_127)
);


endmodule