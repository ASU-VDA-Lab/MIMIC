module fake_jpeg_6531_n_228 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_228);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_11),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_31),
.B(n_32),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_33),
.B(n_35),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_33),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx4f_ASAP7_75t_SL g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx4f_ASAP7_75t_SL g42 ( 
.A(n_38),
.Y(n_42)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

HAxp5_ASAP7_75t_SL g40 ( 
.A(n_20),
.B(n_1),
.CON(n_40),
.SN(n_40)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_41),
.B1(n_27),
.B2(n_25),
.Y(n_60)
);

BUFx12f_ASAP7_75t_SL g41 ( 
.A(n_21),
.Y(n_41)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_46),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_44),
.B(n_54),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_58),
.Y(n_65)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_16),
.B1(n_30),
.B2(n_18),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_31),
.B1(n_37),
.B2(n_58),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_52),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_16),
.B1(n_30),
.B2(n_18),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_53),
.A2(n_61),
.B1(n_15),
.B2(n_19),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_30),
.B1(n_18),
.B2(n_16),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_57),
.B1(n_22),
.B2(n_39),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_22),
.B1(n_27),
.B2(n_19),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_25),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_60),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_15),
.B1(n_19),
.B2(n_26),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_64),
.B(n_63),
.Y(n_93)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_71),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_45),
.B(n_34),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_79),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_69),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_32),
.Y(n_71)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_75),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_39),
.B1(n_31),
.B2(n_28),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_56),
.B(n_20),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_77),
.A2(n_59),
.B1(n_43),
.B2(n_48),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_34),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_51),
.A2(n_31),
.B1(n_24),
.B2(n_23),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_82),
.A2(n_23),
.B1(n_28),
.B2(n_26),
.Y(n_91)
);

MAJx2_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_42),
.C(n_47),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_71),
.C(n_32),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_65),
.B(n_80),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_100),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_80),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_97),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_91),
.A2(n_92),
.B1(n_93),
.B2(n_101),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_68),
.A2(n_56),
.B1(n_62),
.B2(n_54),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_104),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_95),
.A2(n_102),
.B1(n_74),
.B2(n_75),
.Y(n_116)
);

INVx6_ASAP7_75t_SL g96 ( 
.A(n_83),
.Y(n_96)
);

INVxp33_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_63),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_32),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_103),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_61),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_68),
.A2(n_49),
.B1(n_32),
.B2(n_24),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_32),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_114),
.Y(n_146)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_109),
.Y(n_137)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_121),
.C(n_50),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_96),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_111),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_112),
.Y(n_142)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_116),
.A2(n_75),
.B1(n_49),
.B2(n_29),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_78),
.Y(n_117)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_100),
.B(n_73),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_119),
.Y(n_128)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_32),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_123),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_84),
.C(n_90),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_2),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_124),
.A2(n_104),
.B1(n_94),
.B2(n_100),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_127),
.A2(n_134),
.B1(n_135),
.B2(n_147),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_86),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_21),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_87),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_29),
.Y(n_169)
);

NOR2x1_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_102),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_138),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_110),
.A2(n_88),
.B(n_97),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_133),
.A2(n_136),
.B(n_144),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_107),
.A2(n_84),
.B1(n_73),
.B2(n_74),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_122),
.A2(n_74),
.B1(n_78),
.B2(n_89),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_115),
.A2(n_85),
.B(n_52),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_85),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_149),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_66),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_143),
.C(n_121),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_115),
.A2(n_120),
.B(n_118),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_69),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_155),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_160),
.C(n_163),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_132),
.A2(n_123),
.B1(n_109),
.B2(n_105),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_111),
.B1(n_106),
.B2(n_122),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_154),
.A2(n_133),
.B1(n_147),
.B2(n_29),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_145),
.B(n_108),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_157),
.Y(n_174)
);

NOR3xp33_ASAP7_75t_SL g157 ( 
.A(n_130),
.B(n_105),
.C(n_69),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_69),
.C(n_66),
.Y(n_160)
);

MAJx2_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_52),
.C(n_50),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_161),
.B(n_128),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_141),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_81),
.C(n_49),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_144),
.C(n_128),
.Y(n_177)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_169),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_146),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_167),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_137),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_168),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_170),
.A2(n_148),
.B1(n_141),
.B2(n_142),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_131),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_179),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_178),
.C(n_186),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_131),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_158),
.A2(n_127),
.B1(n_130),
.B2(n_138),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_183),
.A2(n_150),
.B1(n_165),
.B2(n_166),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_184),
.Y(n_188)
);

NOR2xp67_ASAP7_75t_SL g185 ( 
.A(n_157),
.B(n_81),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_185),
.A2(n_153),
.B1(n_161),
.B2(n_158),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_29),
.C(n_17),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_187),
.A2(n_189),
.B1(n_195),
.B2(n_198),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_181),
.A2(n_152),
.B(n_159),
.Y(n_189)
);

AND2x4_ASAP7_75t_SL g191 ( 
.A(n_176),
.B(n_152),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_191),
.A2(n_182),
.B1(n_179),
.B2(n_172),
.Y(n_201)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_197),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_159),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_163),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_3),
.Y(n_205)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_181),
.A2(n_160),
.B(n_164),
.Y(n_198)
);

INVx13_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_201),
.A2(n_189),
.B(n_199),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_192),
.A2(n_177),
.B1(n_174),
.B2(n_175),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_192),
.A2(n_178),
.B1(n_186),
.B2(n_5),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_196),
.C(n_190),
.Y(n_213)
);

NOR2x1_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_3),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_L g209 ( 
.A1(n_207),
.A2(n_194),
.B(n_200),
.Y(n_209)
);

NAND3xp33_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_4),
.C(n_5),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_L g212 ( 
.A1(n_208),
.A2(n_7),
.B(n_8),
.Y(n_212)
);

NOR2x1_ASAP7_75t_SL g214 ( 
.A(n_209),
.B(n_195),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_202),
.Y(n_218)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_188),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_204),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_203),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_214),
.A2(n_8),
.B(n_9),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_215),
.B(n_217),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_218),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_206),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_222),
.B(n_218),
.Y(n_223)
);

NAND3xp33_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_224),
.C(n_220),
.Y(n_225)
);

OAI21x1_ASAP7_75t_L g224 ( 
.A1(n_221),
.A2(n_219),
.B(n_12),
.Y(n_224)
);

BUFx24_ASAP7_75t_SL g226 ( 
.A(n_225),
.Y(n_226)
);

INVxp67_ASAP7_75t_SL g227 ( 
.A(n_226),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_227),
.Y(n_228)
);


endmodule