module fake_jpeg_26844_n_92 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_92);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_92;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_62;
wire n_43;
wire n_82;

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_43),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_53),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_1),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_54),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_1),
.Y(n_56)
);

CKINVDCx12_ASAP7_75t_R g68 ( 
.A(n_56),
.Y(n_68)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_44),
.B1(n_49),
.B2(n_45),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_51),
.A2(n_47),
.B1(n_40),
.B2(n_50),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_64),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_68),
.B(n_3),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_70),
.A2(n_62),
.B1(n_60),
.B2(n_66),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_72),
.A2(n_73),
.B1(n_68),
.B2(n_67),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_14),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_15),
.B(n_16),
.Y(n_80)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_77),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_74),
.A2(n_71),
.B(n_59),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_78),
.B(n_79),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_82),
.B(n_80),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_81),
.C(n_18),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_84),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_21),
.C(n_22),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_25),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_26),
.C(n_30),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_31),
.B(n_32),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_36),
.Y(n_92)
);


endmodule