module fake_aes_10233_n_33 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_33);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
BUFx3_ASAP7_75t_L g10 ( .A(n_8), .Y(n_10) );
AND2x6_ASAP7_75t_L g11 ( .A(n_7), .B(n_6), .Y(n_11) );
INVx3_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_5), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
NAND2xp5_ASAP7_75t_SL g15 ( .A(n_0), .B(n_2), .Y(n_15) );
BUFx2_ASAP7_75t_L g16 ( .A(n_1), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_2), .Y(n_17) );
INVx1_ASAP7_75t_SL g18 ( .A(n_16), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_12), .Y(n_19) );
INVx3_ASAP7_75t_L g20 ( .A(n_14), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_13), .B(n_1), .Y(n_21) );
OAI21x1_ASAP7_75t_L g22 ( .A1(n_17), .A2(n_9), .B(n_3), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_19), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_19), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_24), .B(n_18), .Y(n_25) );
AND2x4_ASAP7_75t_L g26 ( .A(n_23), .B(n_20), .Y(n_26) );
NAND4xp25_ASAP7_75t_SL g27 ( .A(n_25), .B(n_21), .C(n_15), .D(n_22), .Y(n_27) );
AOI21xp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_22), .B(n_10), .Y(n_28) );
AOI221xp5_ASAP7_75t_L g29 ( .A1(n_27), .A2(n_3), .B1(n_11), .B2(n_20), .C(n_28), .Y(n_29) );
AND2x4_ASAP7_75t_L g30 ( .A(n_28), .B(n_11), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_30), .Y(n_31) );
BUFx2_ASAP7_75t_L g32 ( .A(n_29), .Y(n_32) );
OA21x2_ASAP7_75t_L g33 ( .A1(n_31), .A2(n_11), .B(n_32), .Y(n_33) );
endmodule