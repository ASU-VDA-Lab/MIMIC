module fake_jpeg_7754_n_109 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_109);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_109;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_26),
.B(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_16),
.B(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_15),
.Y(n_29)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_1),
.Y(n_31)
);

AND2x4_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_1),
.Y(n_32)
);

AO22x1_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_13),
.B1(n_2),
.B2(n_25),
.Y(n_42)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_35),
.A2(n_14),
.B1(n_20),
.B2(n_17),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_32),
.A2(n_23),
.B1(n_24),
.B2(n_14),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_39),
.B1(n_35),
.B2(n_29),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_35),
.B1(n_23),
.B2(n_33),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_33),
.B1(n_29),
.B2(n_34),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_23),
.B(n_24),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_45),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_44),
.B1(n_18),
.B2(n_21),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_32),
.A2(n_20),
.B1(n_21),
.B2(n_19),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_12),
.Y(n_45)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_49),
.A2(n_53),
.B1(n_48),
.B2(n_36),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_26),
.Y(n_50)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_28),
.Y(n_51)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_55),
.Y(n_67)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_19),
.Y(n_56)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_34),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_12),
.Y(n_58)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_17),
.Y(n_61)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_38),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_48),
.Y(n_80)
);

NOR2x1_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_44),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_70),
.B1(n_72),
.B2(n_62),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_75),
.A2(n_53),
.B1(n_63),
.B2(n_42),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_70),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_76),
.B(n_81),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_69),
.A2(n_60),
.B(n_57),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_78),
.C(n_79),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_55),
.C(n_54),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_59),
.Y(n_79)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_82),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_52),
.C(n_53),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_84),
.Y(n_85)
);

XNOR2x1_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_52),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_87),
.A2(n_83),
.B1(n_88),
.B2(n_77),
.Y(n_93)
);

AO221x1_ASAP7_75t_L g88 ( 
.A1(n_84),
.A2(n_64),
.B1(n_36),
.B2(n_40),
.C(n_42),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_89),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_68),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_93),
.A2(n_95),
.B1(n_86),
.B2(n_74),
.Y(n_100)
);

AOI32xp33_ASAP7_75t_SL g95 ( 
.A1(n_87),
.A2(n_53),
.A3(n_79),
.B1(n_78),
.B2(n_44),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_85),
.C(n_89),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_91),
.C(n_85),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_100),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_90),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_98),
.A2(n_99),
.B1(n_94),
.B2(n_64),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_71),
.Y(n_102)
);

OAI31xp33_ASAP7_75t_L g105 ( 
.A1(n_102),
.A2(n_4),
.A3(n_5),
.B(n_8),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_98),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_104),
.B(n_101),
.C(n_11),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_8),
.B(n_10),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_107),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_11),
.Y(n_109)
);


endmodule