module fake_jpeg_27114_n_203 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx4f_ASAP7_75t_SL g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_10),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_17),
.Y(n_34)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_29),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_27),
.Y(n_46)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_39),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_27),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_48),
.B(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_32),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_17),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_33),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_16),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_24),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_62),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_25),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_25),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_64),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_17),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_17),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_66),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_50),
.Y(n_66)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_71),
.Y(n_94)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_75),
.Y(n_105)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_76),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_54),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_40),
.B1(n_42),
.B2(n_37),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_77),
.A2(n_82),
.B1(n_43),
.B2(n_39),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_34),
.B(n_41),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_78),
.Y(n_87)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_79),
.Y(n_100)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_81),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_28),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_40),
.B1(n_43),
.B2(n_42),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_56),
.Y(n_97)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_95),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_26),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_92),
.A2(n_96),
.B(n_101),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_85),
.B(n_30),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_93),
.A2(n_66),
.B(n_75),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_SL g95 ( 
.A(n_68),
.B(n_23),
.C(n_20),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_56),
.B(n_53),
.C(n_49),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_26),
.Y(n_129)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_73),
.Y(n_112)
);

NOR2xp67_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_21),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_69),
.A2(n_23),
.B(n_16),
.C(n_22),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_104),
.A2(n_109),
.B1(n_67),
.B2(n_86),
.Y(n_115)
);

AO22x1_ASAP7_75t_L g108 ( 
.A1(n_77),
.A2(n_20),
.B1(n_19),
.B2(n_23),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_108),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_69),
.A2(n_22),
.B1(n_21),
.B2(n_31),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_111),
.B(n_116),
.Y(n_135)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_72),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_120),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_68),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_83),
.Y(n_117)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_127),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_91),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_119),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_82),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_84),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_125),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_87),
.A2(n_74),
.B(n_73),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_124),
.Y(n_133)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_19),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_129),
.Y(n_146)
);

INVxp33_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_96),
.A2(n_80),
.B1(n_71),
.B2(n_70),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_19),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_105),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_125),
.B(n_114),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_139),
.B(n_141),
.Y(n_161)
);

AOI221xp5_ASAP7_75t_L g140 ( 
.A1(n_128),
.A2(n_101),
.B1(n_90),
.B2(n_89),
.C(n_95),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_144),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_130),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_90),
.C(n_92),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_108),
.Y(n_145)
);

MAJx2_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_122),
.C(n_129),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_110),
.A2(n_107),
.B1(n_106),
.B2(n_21),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_117),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_148),
.A2(n_122),
.B(n_129),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_135),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_150),
.Y(n_166)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_136),
.C(n_144),
.Y(n_167)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_153),
.Y(n_176)
);

NOR3xp33_ASAP7_75t_SL g153 ( 
.A(n_143),
.B(n_126),
.C(n_116),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_137),
.Y(n_154)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_111),
.Y(n_155)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_138),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_157),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_147),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_158),
.A2(n_146),
.B(n_124),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_122),
.Y(n_159)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_159),
.Y(n_171)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_SL g163 ( 
.A1(n_146),
.A2(n_131),
.B(n_128),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_163),
.A2(n_133),
.B1(n_148),
.B2(n_115),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_161),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_152),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_168),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_173),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_136),
.C(n_145),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_159),
.A2(n_134),
.B(n_142),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_158),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

OAI21xp33_ASAP7_75t_L g178 ( 
.A1(n_175),
.A2(n_162),
.B(n_156),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_178),
.A2(n_171),
.B1(n_174),
.B2(n_165),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_164),
.A2(n_169),
.B1(n_170),
.B2(n_153),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_182),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_167),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_0),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_187),
.B(n_188),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_106),
.C(n_118),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_183),
.C(n_180),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_18),
.C(n_1),
.Y(n_193)
);

AOI322xp5_ASAP7_75t_L g191 ( 
.A1(n_186),
.A2(n_178),
.A3(n_31),
.B1(n_11),
.B2(n_9),
.C1(n_18),
.C2(n_5),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_193),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_192),
.A2(n_194),
.B(n_3),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_0),
.C(n_3),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_197),
.Y(n_199)
);

NOR2x1_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_185),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_188),
.C(n_7),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_198),
.Y(n_200)
);

OAI321xp33_ASAP7_75t_L g201 ( 
.A1(n_199),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_176),
.C(n_166),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_201),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_200),
.Y(n_203)
);


endmodule