module fake_netlist_1_8472_n_680 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_680);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_680;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_622;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_39), .Y(n_78) );
BUFx3_ASAP7_75t_L g79 ( .A(n_53), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_46), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_54), .Y(n_81) );
CKINVDCx14_ASAP7_75t_R g82 ( .A(n_62), .Y(n_82) );
BUFx2_ASAP7_75t_L g83 ( .A(n_70), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_57), .Y(n_84) );
CKINVDCx16_ASAP7_75t_R g85 ( .A(n_42), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_71), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_15), .Y(n_87) );
HB1xp67_ASAP7_75t_L g88 ( .A(n_44), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_52), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_29), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_26), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_1), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_25), .Y(n_93) );
INVx3_ASAP7_75t_L g94 ( .A(n_45), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_31), .Y(n_95) );
CKINVDCx14_ASAP7_75t_R g96 ( .A(n_15), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_27), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_1), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_11), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_66), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_74), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_28), .Y(n_102) );
CKINVDCx16_ASAP7_75t_R g103 ( .A(n_14), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_6), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_75), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_65), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_37), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_58), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_30), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_32), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_34), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_72), .Y(n_112) );
INVxp33_ASAP7_75t_SL g113 ( .A(n_2), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_5), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_33), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_51), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_19), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_7), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_38), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g120 ( .A(n_41), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_21), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_50), .Y(n_122) );
INVxp67_ASAP7_75t_SL g123 ( .A(n_5), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_0), .Y(n_124) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_13), .B(n_21), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_105), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_83), .B(n_0), .Y(n_127) );
OAI22xp5_ASAP7_75t_L g128 ( .A1(n_96), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_128) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_103), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_94), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_85), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_94), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_80), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_80), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_101), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_83), .B(n_3), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_120), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_81), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_94), .B(n_4), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_91), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_87), .B(n_6), .Y(n_141) );
AND2x2_ASAP7_75t_L g142 ( .A(n_88), .B(n_7), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_91), .Y(n_143) );
NOR2xp33_ASAP7_75t_SL g144 ( .A(n_100), .B(n_107), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_111), .Y(n_145) );
INVx4_ASAP7_75t_L g146 ( .A(n_79), .Y(n_146) );
NAND2xp33_ASAP7_75t_SL g147 ( .A(n_100), .B(n_8), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_81), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_113), .B(n_8), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_107), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_111), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_87), .B(n_9), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_84), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_110), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_110), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_84), .Y(n_156) );
INVxp67_ASAP7_75t_L g157 ( .A(n_104), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_86), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_86), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_114), .B(n_9), .Y(n_160) );
NAND2xp33_ASAP7_75t_SL g161 ( .A(n_98), .B(n_10), .Y(n_161) );
NAND2xp33_ASAP7_75t_SL g162 ( .A(n_92), .B(n_10), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_89), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_79), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_89), .Y(n_165) );
INVxp67_ASAP7_75t_L g166 ( .A(n_121), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_90), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_132), .Y(n_168) );
AND2x6_ASAP7_75t_L g169 ( .A(n_139), .B(n_90), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_132), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_133), .B(n_82), .Y(n_171) );
NAND3xp33_ASAP7_75t_L g172 ( .A(n_136), .B(n_117), .C(n_124), .Y(n_172) );
BUFx3_ASAP7_75t_L g173 ( .A(n_139), .Y(n_173) );
HB1xp67_ASAP7_75t_L g174 ( .A(n_129), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_133), .B(n_109), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_136), .B(n_92), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_132), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_132), .Y(n_178) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_132), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_140), .Y(n_180) );
AND2x6_ASAP7_75t_L g181 ( .A(n_139), .B(n_95), .Y(n_181) );
AND2x6_ASAP7_75t_L g182 ( .A(n_139), .B(n_95), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_132), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_134), .B(n_78), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_130), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_130), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_167), .Y(n_187) );
OR2x2_ASAP7_75t_L g188 ( .A(n_157), .B(n_117), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_167), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_164), .Y(n_190) );
INVx1_ASAP7_75t_SL g191 ( .A(n_143), .Y(n_191) );
NAND2x1p5_ASAP7_75t_L g192 ( .A(n_141), .B(n_115), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_164), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_141), .A2(n_124), .B1(n_99), .B2(n_118), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_141), .Y(n_195) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_150), .Y(n_196) );
OAI221xp5_ASAP7_75t_L g197 ( .A1(n_166), .A2(n_99), .B1(n_118), .B2(n_123), .C(n_125), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_141), .B(n_97), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_167), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_154), .B(n_122), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_155), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_131), .B(n_108), .Y(n_202) );
BUFx2_ASAP7_75t_L g203 ( .A(n_135), .Y(n_203) );
OR2x2_ASAP7_75t_L g204 ( .A(n_142), .B(n_119), .Y(n_204) );
INVx4_ASAP7_75t_L g205 ( .A(n_146), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_152), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_164), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_142), .B(n_119), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_152), .Y(n_209) );
CKINVDCx16_ASAP7_75t_R g210 ( .A(n_144), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_164), .Y(n_211) );
INVx4_ASAP7_75t_SL g212 ( .A(n_152), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_164), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_151), .Y(n_214) );
INVx2_ASAP7_75t_SL g215 ( .A(n_146), .Y(n_215) );
INVx1_ASAP7_75t_SL g216 ( .A(n_137), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_164), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_134), .B(n_112), .Y(n_218) );
INVx5_ASAP7_75t_L g219 ( .A(n_146), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_138), .B(n_106), .Y(n_220) );
INVx1_ASAP7_75t_SL g221 ( .A(n_126), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_151), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_151), .Y(n_223) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_152), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_163), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_165), .B(n_116), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_163), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_145), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_145), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_138), .Y(n_230) );
NOR2xp33_ASAP7_75t_R g231 ( .A(n_180), .B(n_161), .Y(n_231) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_169), .A2(n_127), .B1(n_149), .B2(n_147), .Y(n_232) );
AND2x4_ASAP7_75t_L g233 ( .A(n_208), .B(n_165), .Y(n_233) );
NOR3xp33_ASAP7_75t_SL g234 ( .A(n_180), .B(n_128), .C(n_162), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_204), .B(n_159), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_187), .Y(n_236) );
XOR2xp5_ASAP7_75t_L g237 ( .A(n_210), .B(n_11), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_187), .Y(n_238) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_174), .Y(n_239) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_221), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_189), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_189), .Y(n_242) );
AND2x4_ASAP7_75t_L g243 ( .A(n_208), .B(n_148), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_171), .B(n_159), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_226), .B(n_158), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_226), .B(n_158), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_199), .Y(n_247) );
BUFx4f_ASAP7_75t_SL g248 ( .A(n_216), .Y(n_248) );
AND2x4_ASAP7_75t_L g249 ( .A(n_212), .B(n_156), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_226), .B(n_156), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_199), .Y(n_251) );
OR2x6_ASAP7_75t_L g252 ( .A(n_192), .B(n_160), .Y(n_252) );
BUFx3_ASAP7_75t_L g253 ( .A(n_169), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_177), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_176), .B(n_153), .Y(n_255) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_224), .Y(n_256) );
NOR2xp67_ASAP7_75t_L g257 ( .A(n_196), .B(n_197), .Y(n_257) );
BUFx4f_ASAP7_75t_SL g258 ( .A(n_191), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_176), .B(n_153), .Y(n_259) );
INVx6_ASAP7_75t_L g260 ( .A(n_224), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_195), .A2(n_148), .B(n_146), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_204), .B(n_93), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_188), .B(n_116), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_214), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_212), .B(n_115), .Y(n_265) );
INVx2_ASAP7_75t_SL g266 ( .A(n_173), .Y(n_266) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_201), .Y(n_267) );
BUFx4f_ASAP7_75t_L g268 ( .A(n_169), .Y(n_268) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_201), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_214), .Y(n_270) );
NOR2xp67_ASAP7_75t_L g271 ( .A(n_172), .B(n_12), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_169), .A2(n_102), .B1(n_97), .B2(n_14), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_198), .B(n_102), .Y(n_273) );
NOR2x1_ASAP7_75t_L g274 ( .A(n_188), .B(n_12), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_198), .B(n_13), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_177), .Y(n_276) );
AND2x4_ASAP7_75t_L g277 ( .A(n_212), .B(n_16), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_230), .Y(n_278) );
AO22x1_ASAP7_75t_L g279 ( .A1(n_169), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_279) );
OAI22xp33_ASAP7_75t_L g280 ( .A1(n_192), .A2(n_17), .B1(n_18), .B2(n_19), .Y(n_280) );
BUFx2_ASAP7_75t_L g281 ( .A(n_169), .Y(n_281) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_224), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_198), .B(n_20), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_200), .B(n_56), .Y(n_284) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_203), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_212), .B(n_55), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_230), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_177), .Y(n_288) );
INVxp67_ASAP7_75t_SL g289 ( .A(n_192), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_177), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_224), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_224), .Y(n_292) );
NOR3xp33_ASAP7_75t_SL g293 ( .A(n_202), .B(n_20), .C(n_22), .Y(n_293) );
INVx3_ASAP7_75t_L g294 ( .A(n_173), .Y(n_294) );
INVx4_ASAP7_75t_L g295 ( .A(n_181), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_203), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_206), .B(n_59), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_295), .B(n_194), .Y(n_298) );
BUFx3_ASAP7_75t_L g299 ( .A(n_253), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_264), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_235), .B(n_181), .Y(n_301) );
AOI22xp5_ASAP7_75t_L g302 ( .A1(n_289), .A2(n_182), .B1(n_181), .B2(n_209), .Y(n_302) );
INVx3_ASAP7_75t_L g303 ( .A(n_249), .Y(n_303) );
INVx5_ASAP7_75t_L g304 ( .A(n_295), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g305 ( .A1(n_233), .A2(n_181), .B1(n_182), .B2(n_227), .Y(n_305) );
INVx5_ASAP7_75t_L g306 ( .A(n_295), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_233), .B(n_181), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_233), .B(n_185), .Y(n_308) );
INVx3_ASAP7_75t_L g309 ( .A(n_249), .Y(n_309) );
INVx2_ASAP7_75t_SL g310 ( .A(n_277), .Y(n_310) );
AND2x6_ASAP7_75t_L g311 ( .A(n_253), .B(n_181), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_278), .A2(n_215), .B(n_205), .Y(n_312) );
OR2x2_ASAP7_75t_L g313 ( .A(n_240), .B(n_220), .Y(n_313) );
CKINVDCx20_ASAP7_75t_R g314 ( .A(n_248), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g315 ( .A1(n_252), .A2(n_175), .B1(n_184), .B2(n_218), .Y(n_315) );
BUFx6f_ASAP7_75t_L g316 ( .A(n_268), .Y(n_316) );
OAI22xp33_ASAP7_75t_L g317 ( .A1(n_258), .A2(n_229), .B1(n_228), .B2(n_186), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_296), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_243), .B(n_185), .Y(n_319) );
BUFx2_ASAP7_75t_L g320 ( .A(n_277), .Y(n_320) );
AOI22xp5_ASAP7_75t_L g321 ( .A1(n_257), .A2(n_182), .B1(n_225), .B2(n_186), .Y(n_321) );
A2O1A1Ixp33_ASAP7_75t_L g322 ( .A1(n_278), .A2(n_229), .B(n_228), .C(n_223), .Y(n_322) );
CKINVDCx20_ASAP7_75t_R g323 ( .A(n_296), .Y(n_323) );
AND2x4_ASAP7_75t_L g324 ( .A(n_252), .B(n_182), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_239), .B(n_182), .Y(n_325) );
INVx3_ASAP7_75t_L g326 ( .A(n_249), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_287), .Y(n_327) );
BUFx3_ASAP7_75t_L g328 ( .A(n_268), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_264), .Y(n_329) );
BUFx10_ASAP7_75t_L g330 ( .A(n_277), .Y(n_330) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_285), .Y(n_331) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_268), .B(n_219), .Y(n_332) );
OAI21x1_ASAP7_75t_L g333 ( .A1(n_286), .A2(n_168), .B(n_178), .Y(n_333) );
INVx2_ASAP7_75t_SL g334 ( .A(n_252), .Y(n_334) );
BUFx2_ASAP7_75t_L g335 ( .A(n_252), .Y(n_335) );
AND2x4_ASAP7_75t_SL g336 ( .A(n_267), .B(n_205), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_243), .A2(n_182), .B1(n_222), .B2(n_223), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_243), .B(n_222), .Y(n_338) );
AOI21xp5_ASAP7_75t_L g339 ( .A1(n_287), .A2(n_215), .B(n_205), .Y(n_339) );
BUFx12f_ASAP7_75t_L g340 ( .A(n_263), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_263), .B(n_219), .Y(n_341) );
BUFx12f_ASAP7_75t_L g342 ( .A(n_281), .Y(n_342) );
NAND3xp33_ASAP7_75t_L g343 ( .A(n_272), .B(n_219), .C(n_170), .Y(n_343) );
INVx2_ASAP7_75t_SL g344 ( .A(n_281), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_270), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_255), .B(n_219), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_259), .B(n_219), .Y(n_347) );
NOR2x1_ASAP7_75t_SL g348 ( .A(n_270), .B(n_170), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_313), .B(n_244), .Y(n_349) );
OR2x6_ASAP7_75t_L g350 ( .A(n_324), .B(n_245), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_340), .B(n_269), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_308), .B(n_236), .Y(n_352) );
OA21x2_ASAP7_75t_L g353 ( .A1(n_333), .A2(n_217), .B(n_190), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_300), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_308), .B(n_236), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_300), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_320), .A2(n_250), .B1(n_246), .B2(n_273), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_329), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_319), .B(n_242), .Y(n_359) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_340), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_313), .B(n_262), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_331), .A2(n_274), .B1(n_275), .B2(n_283), .Y(n_362) );
NAND2xp33_ASAP7_75t_L g363 ( .A(n_311), .B(n_266), .Y(n_363) );
INVx4_ASAP7_75t_L g364 ( .A(n_324), .Y(n_364) );
OR2x6_ASAP7_75t_L g365 ( .A(n_324), .B(n_266), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_329), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_320), .A2(n_232), .B1(n_247), .B2(n_238), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_319), .B(n_242), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_327), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_338), .B(n_241), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_318), .B(n_237), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_338), .B(n_234), .Y(n_372) );
NAND2xp33_ASAP7_75t_R g373 ( .A(n_318), .B(n_231), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_327), .Y(n_374) );
NAND2x1p5_ASAP7_75t_L g375 ( .A(n_304), .B(n_247), .Y(n_375) );
INVx2_ASAP7_75t_SL g376 ( .A(n_330), .Y(n_376) );
AO31x2_ASAP7_75t_L g377 ( .A1(n_315), .A2(n_297), .A3(n_193), .B(n_207), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_345), .Y(n_378) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_304), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_352), .B(n_335), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_352), .B(n_335), .Y(n_381) );
OAI21x1_ASAP7_75t_L g382 ( .A1(n_353), .A2(n_333), .B(n_312), .Y(n_382) );
OAI21x1_ASAP7_75t_L g383 ( .A1(n_353), .A2(n_339), .B(n_211), .Y(n_383) );
AOI21xp5_ASAP7_75t_L g384 ( .A1(n_353), .A2(n_310), .B(n_348), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_372), .A2(n_323), .B1(n_334), .B2(n_237), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_349), .A2(n_323), .B1(n_334), .B2(n_298), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_350), .A2(n_361), .B1(n_357), .B2(n_351), .Y(n_387) );
OAI21xp33_ASAP7_75t_SL g388 ( .A1(n_369), .A2(n_310), .B(n_302), .Y(n_388) );
CKINVDCx11_ASAP7_75t_R g389 ( .A(n_365), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_350), .A2(n_325), .B1(n_317), .B2(n_301), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_369), .A2(n_305), .B1(n_337), .B2(n_321), .Y(n_391) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_374), .Y(n_392) );
AO31x2_ASAP7_75t_L g393 ( .A1(n_367), .A2(n_322), .A3(n_348), .B(n_251), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_374), .B(n_336), .Y(n_394) );
AOI221xp5_ASAP7_75t_L g395 ( .A1(n_378), .A2(n_280), .B1(n_293), .B2(n_279), .C(n_341), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_354), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_354), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_355), .B(n_238), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_355), .B(n_241), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_356), .B(n_251), .Y(n_400) );
AOI22xp33_ASAP7_75t_SL g401 ( .A1(n_364), .A2(n_314), .B1(n_336), .B2(n_330), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_350), .A2(n_307), .B1(n_344), .B2(n_343), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_356), .Y(n_403) );
AO21x2_ASAP7_75t_L g404 ( .A1(n_358), .A2(n_271), .B(n_190), .Y(n_404) );
OAI211xp5_ASAP7_75t_L g405 ( .A1(n_362), .A2(n_314), .B(n_284), .C(n_346), .Y(n_405) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_375), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_389), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_396), .Y(n_408) );
INVxp67_ASAP7_75t_L g409 ( .A(n_406), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_392), .B(n_358), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_399), .B(n_366), .Y(n_411) );
AOI33xp33_ASAP7_75t_L g412 ( .A1(n_385), .A2(n_378), .A3(n_368), .B1(n_359), .B2(n_366), .B3(n_370), .Y(n_412) );
NAND2xp33_ASAP7_75t_R g413 ( .A(n_394), .B(n_371), .Y(n_413) );
BUFx3_ASAP7_75t_L g414 ( .A(n_406), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_387), .B(n_371), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_396), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_399), .B(n_370), .Y(n_417) );
AOI22x1_ASAP7_75t_SL g418 ( .A1(n_397), .A2(n_364), .B1(n_279), .B2(n_373), .Y(n_418) );
NOR4xp25_ASAP7_75t_SL g419 ( .A(n_395), .B(n_265), .C(n_332), .D(n_292), .Y(n_419) );
INVxp67_ASAP7_75t_SL g420 ( .A(n_392), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_401), .Y(n_421) );
OAI221xp5_ASAP7_75t_L g422 ( .A1(n_386), .A2(n_360), .B1(n_350), .B2(n_364), .C(n_365), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_401), .A2(n_350), .B1(n_365), .B2(n_364), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_397), .Y(n_424) );
OAI332xp33_ASAP7_75t_L g425 ( .A1(n_403), .A2(n_347), .A3(n_22), .B1(n_376), .B2(n_193), .B3(n_211), .C1(n_207), .C2(n_213), .Y(n_425) );
AND2x4_ASAP7_75t_L g426 ( .A(n_403), .B(n_399), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_400), .Y(n_427) );
BUFx3_ASAP7_75t_L g428 ( .A(n_398), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_383), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_380), .B(n_359), .Y(n_430) );
AOI222xp33_ASAP7_75t_L g431 ( .A1(n_395), .A2(n_368), .B1(n_346), .B2(n_342), .C1(n_363), .C2(n_330), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_394), .A2(n_365), .B1(n_375), .B2(n_376), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_400), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_390), .A2(n_365), .B1(n_375), .B2(n_344), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_380), .B(n_377), .Y(n_435) );
NOR4xp25_ASAP7_75t_SL g436 ( .A(n_405), .B(n_292), .C(n_291), .D(n_377), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_393), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_380), .A2(n_303), .B1(n_309), .B2(n_326), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_398), .Y(n_439) );
AOI21xp33_ASAP7_75t_SL g440 ( .A1(n_405), .A2(n_23), .B(n_24), .Y(n_440) );
OAI31xp33_ASAP7_75t_L g441 ( .A1(n_391), .A2(n_303), .A3(n_309), .B(n_326), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_393), .Y(n_442) );
INVx2_ASAP7_75t_SL g443 ( .A(n_414), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_420), .B(n_393), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_435), .B(n_393), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_408), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_429), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_435), .B(n_393), .Y(n_448) );
NOR2xp33_ASAP7_75t_R g449 ( .A(n_413), .B(n_342), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_408), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_428), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_416), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_439), .B(n_393), .Y(n_453) );
INVx4_ASAP7_75t_L g454 ( .A(n_414), .Y(n_454) );
OR2x2_ASAP7_75t_SL g455 ( .A(n_410), .B(n_379), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_416), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_429), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_426), .B(n_393), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_417), .B(n_381), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_426), .B(n_417), .Y(n_460) );
OAI33xp33_ASAP7_75t_L g461 ( .A1(n_424), .A2(n_391), .A3(n_402), .B1(n_217), .B2(n_213), .B3(n_168), .Y(n_461) );
OAI33xp33_ASAP7_75t_L g462 ( .A1(n_424), .A2(n_402), .A3(n_178), .B1(n_291), .B2(n_388), .B3(n_404), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_437), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_437), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_411), .B(n_381), .Y(n_465) );
INVx3_ASAP7_75t_L g466 ( .A(n_426), .Y(n_466) );
NAND2x1_ASAP7_75t_L g467 ( .A(n_427), .B(n_384), .Y(n_467) );
INVx3_ASAP7_75t_L g468 ( .A(n_426), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_442), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_411), .B(n_377), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_442), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_410), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_427), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_433), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_428), .B(n_377), .Y(n_475) );
OAI21xp5_ASAP7_75t_L g476 ( .A1(n_415), .A2(n_388), .B(n_384), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_433), .Y(n_477) );
OAI31xp33_ASAP7_75t_L g478 ( .A1(n_423), .A2(n_309), .A3(n_303), .B(n_326), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_430), .B(n_377), .Y(n_479) );
AND2x4_ASAP7_75t_L g480 ( .A(n_409), .B(n_383), .Y(n_480) );
OAI33xp33_ASAP7_75t_L g481 ( .A1(n_421), .A2(n_404), .A3(n_254), .B1(n_290), .B2(n_288), .B3(n_276), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_430), .B(n_404), .Y(n_482) );
AOI221xp5_ASAP7_75t_L g483 ( .A1(n_425), .A2(n_261), .B1(n_404), .B2(n_177), .C(n_179), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_421), .A2(n_379), .B1(n_311), .B2(n_294), .Y(n_484) );
OA33x2_ASAP7_75t_L g485 ( .A1(n_434), .A2(n_35), .A3(n_36), .B1(n_40), .B2(n_43), .B3(n_47), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_412), .B(n_379), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_418), .Y(n_487) );
AOI221xp5_ASAP7_75t_L g488 ( .A1(n_422), .A2(n_183), .B1(n_179), .B2(n_294), .C(n_282), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_436), .B(n_383), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_432), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_418), .Y(n_491) );
AOI33xp33_ASAP7_75t_L g492 ( .A1(n_438), .A2(n_288), .A3(n_276), .B1(n_290), .B2(n_254), .B3(n_63), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_441), .Y(n_493) );
INVxp67_ASAP7_75t_SL g494 ( .A(n_431), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_472), .B(n_407), .Y(n_495) );
NAND2xp33_ASAP7_75t_R g496 ( .A(n_449), .B(n_407), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_470), .B(n_382), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_470), .B(n_382), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_491), .B(n_440), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_472), .B(n_460), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_447), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_450), .Y(n_502) );
AND2x2_ASAP7_75t_SL g503 ( .A(n_454), .B(n_379), .Y(n_503) );
BUFx2_ASAP7_75t_L g504 ( .A(n_455), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_460), .B(n_419), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_466), .B(n_382), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_458), .B(n_353), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_458), .B(n_379), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_456), .Y(n_509) );
OR2x4_ASAP7_75t_L g510 ( .A(n_491), .B(n_316), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_445), .B(n_48), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_447), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_445), .B(n_49), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_494), .A2(n_256), .B1(n_282), .B2(n_260), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_456), .Y(n_515) );
NAND2x1_ASAP7_75t_SL g516 ( .A(n_454), .B(n_294), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_479), .B(n_183), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_446), .Y(n_518) );
CKINVDCx5p33_ASAP7_75t_R g519 ( .A(n_454), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_448), .B(n_60), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_446), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_473), .B(n_282), .Y(n_522) );
OAI21xp33_ASAP7_75t_L g523 ( .A1(n_487), .A2(n_183), .B(n_179), .Y(n_523) );
AND2x2_ASAP7_75t_SL g524 ( .A(n_454), .B(n_316), .Y(n_524) );
INVx4_ASAP7_75t_L g525 ( .A(n_443), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_448), .B(n_61), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_452), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_482), .B(n_64), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_473), .B(n_256), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_452), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_479), .B(n_183), .Y(n_531) );
NOR2xp33_ASAP7_75t_R g532 ( .A(n_443), .B(n_311), .Y(n_532) );
INVxp67_ASAP7_75t_L g533 ( .A(n_451), .Y(n_533) );
NOR2xp33_ASAP7_75t_R g534 ( .A(n_466), .B(n_311), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_474), .B(n_256), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_487), .B(n_67), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_482), .B(n_68), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_477), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_463), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_477), .B(n_465), .Y(n_540) );
INVxp67_ASAP7_75t_SL g541 ( .A(n_475), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_475), .B(n_69), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_463), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_463), .Y(n_544) );
INVxp67_ASAP7_75t_L g545 ( .A(n_485), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_466), .B(n_73), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_459), .B(n_282), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_447), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_457), .Y(n_549) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_455), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_466), .B(n_76), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_519), .B(n_478), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_541), .B(n_468), .Y(n_553) );
OR2x6_ASAP7_75t_L g554 ( .A(n_504), .B(n_467), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_502), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_502), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_508), .B(n_468), .Y(n_557) );
AND2x2_ASAP7_75t_SL g558 ( .A(n_503), .B(n_490), .Y(n_558) );
INVx1_ASAP7_75t_SL g559 ( .A(n_503), .Y(n_559) );
OAI21xp5_ASAP7_75t_SL g560 ( .A1(n_545), .A2(n_483), .B(n_484), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_509), .Y(n_561) );
AOI21xp33_ASAP7_75t_L g562 ( .A1(n_499), .A2(n_486), .B(n_467), .Y(n_562) );
NAND3xp33_ASAP7_75t_L g563 ( .A(n_533), .B(n_492), .C(n_488), .Y(n_563) );
AOI221xp5_ASAP7_75t_L g564 ( .A1(n_540), .A2(n_476), .B1(n_462), .B2(n_469), .C(n_471), .Y(n_564) );
OAI21xp33_ASAP7_75t_L g565 ( .A1(n_550), .A2(n_444), .B(n_453), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_510), .A2(n_484), .B1(n_453), .B2(n_468), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_500), .B(n_468), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_525), .Y(n_568) );
AOI221xp5_ASAP7_75t_L g569 ( .A1(n_495), .A2(n_464), .B1(n_469), .B2(n_471), .C(n_481), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_538), .B(n_444), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_497), .B(n_480), .Y(n_571) );
OAI21xp5_ASAP7_75t_L g572 ( .A1(n_523), .A2(n_493), .B(n_480), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_509), .Y(n_573) );
AND2x4_ASAP7_75t_L g574 ( .A(n_504), .B(n_480), .Y(n_574) );
OAI221xp5_ASAP7_75t_L g575 ( .A1(n_505), .A2(n_493), .B1(n_489), .B2(n_457), .C(n_179), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_515), .B(n_493), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_525), .Y(n_577) );
O2A1O1Ixp33_ASAP7_75t_L g578 ( .A1(n_536), .A2(n_461), .B(n_489), .C(n_457), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_524), .A2(n_306), .B(n_304), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_510), .A2(n_306), .B1(n_304), .B2(n_299), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_515), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_511), .A2(n_256), .B1(n_282), .B2(n_260), .Y(n_582) );
CKINVDCx16_ASAP7_75t_R g583 ( .A(n_496), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_525), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_510), .A2(n_304), .B1(n_306), .B2(n_299), .Y(n_585) );
INVxp67_ASAP7_75t_SL g586 ( .A(n_517), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_508), .B(n_77), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_511), .A2(n_260), .B1(n_311), .B2(n_179), .Y(n_588) );
OAI21xp33_ASAP7_75t_L g589 ( .A1(n_497), .A2(n_183), .B(n_328), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_498), .B(n_316), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_518), .Y(n_591) );
NAND2x1_ASAP7_75t_SL g592 ( .A(n_513), .B(n_311), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_498), .B(n_260), .Y(n_593) );
BUFx2_ASAP7_75t_L g594 ( .A(n_516), .Y(n_594) );
INVx1_ASAP7_75t_SL g595 ( .A(n_516), .Y(n_595) );
OR2x6_ASAP7_75t_L g596 ( .A(n_513), .B(n_316), .Y(n_596) );
OAI21xp33_ASAP7_75t_SL g597 ( .A1(n_524), .A2(n_306), .B(n_316), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_521), .B(n_306), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_586), .B(n_530), .Y(n_599) );
AOI21xp5_ASAP7_75t_L g600 ( .A1(n_597), .A2(n_526), .B(n_520), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_555), .Y(n_601) );
NAND2xp33_ASAP7_75t_L g602 ( .A(n_559), .B(n_532), .Y(n_602) );
INVx2_ASAP7_75t_SL g603 ( .A(n_568), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_576), .B(n_530), .Y(n_604) );
XNOR2xp5_ASAP7_75t_L g605 ( .A(n_583), .B(n_526), .Y(n_605) );
INVx1_ASAP7_75t_SL g606 ( .A(n_559), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_556), .Y(n_607) );
AOI321xp33_ASAP7_75t_L g608 ( .A1(n_552), .A2(n_537), .A3(n_528), .B1(n_542), .B2(n_507), .C(n_506), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_557), .B(n_506), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_561), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_560), .B(n_506), .Y(n_611) );
AND2x4_ASAP7_75t_L g612 ( .A(n_574), .B(n_539), .Y(n_612) );
AOI21xp5_ASAP7_75t_L g613 ( .A1(n_572), .A2(n_558), .B(n_589), .Y(n_613) );
AOI22x1_ASAP7_75t_L g614 ( .A1(n_594), .A2(n_595), .B1(n_577), .B2(n_584), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_573), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_581), .Y(n_616) );
INVx1_ASAP7_75t_SL g617 ( .A(n_553), .Y(n_617) );
XOR2x2_ASAP7_75t_L g618 ( .A(n_592), .B(n_551), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_571), .B(n_543), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_591), .Y(n_620) );
AOI21x1_ASAP7_75t_SL g621 ( .A1(n_574), .A2(n_546), .B(n_547), .Y(n_621) );
XNOR2x1_ASAP7_75t_L g622 ( .A(n_567), .B(n_546), .Y(n_622) );
INVxp67_ASAP7_75t_SL g623 ( .A(n_578), .Y(n_623) );
NAND2xp33_ASAP7_75t_R g624 ( .A(n_596), .B(n_534), .Y(n_624) );
BUFx3_ASAP7_75t_L g625 ( .A(n_595), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_570), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_593), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_617), .B(n_565), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_599), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_602), .A2(n_554), .B(n_572), .Y(n_630) );
AOI211xp5_ASAP7_75t_L g631 ( .A1(n_611), .A2(n_562), .B(n_575), .C(n_566), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_602), .A2(n_554), .B(n_596), .Y(n_632) );
NOR3xp33_ASAP7_75t_L g633 ( .A(n_613), .B(n_563), .C(n_569), .Y(n_633) );
NAND4xp25_ASAP7_75t_SL g634 ( .A(n_600), .B(n_563), .C(n_564), .D(n_588), .Y(n_634) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_603), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_601), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_619), .B(n_554), .Y(n_637) );
BUFx3_ASAP7_75t_L g638 ( .A(n_625), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_607), .Y(n_639) );
NOR3xp33_ASAP7_75t_L g640 ( .A(n_627), .B(n_587), .C(n_585), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_614), .Y(n_641) );
INVx8_ASAP7_75t_L g642 ( .A(n_612), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_619), .B(n_596), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_610), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_615), .Y(n_645) );
OAI321xp33_ASAP7_75t_L g646 ( .A1(n_608), .A2(n_580), .A3(n_582), .B1(n_514), .B2(n_590), .C(n_517), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_622), .A2(n_527), .B1(n_543), .B2(n_544), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_616), .Y(n_648) );
OR2x2_ASAP7_75t_L g649 ( .A(n_626), .B(n_539), .Y(n_649) );
NAND2x1p5_ASAP7_75t_L g650 ( .A(n_638), .B(n_625), .Y(n_650) );
NOR2x1_ASAP7_75t_L g651 ( .A(n_641), .B(n_605), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_642), .A2(n_622), .B1(n_603), .B2(n_612), .Y(n_652) );
INVx1_ASAP7_75t_SL g653 ( .A(n_638), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_635), .Y(n_654) );
NOR4xp25_ASAP7_75t_L g655 ( .A(n_634), .B(n_641), .C(n_646), .D(n_629), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_630), .B(n_618), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_642), .B(n_606), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_642), .A2(n_618), .B(n_604), .Y(n_658) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_633), .A2(n_620), .B1(n_609), .B2(n_544), .C(n_598), .Y(n_659) );
AOI221xp5_ASAP7_75t_L g660 ( .A1(n_628), .A2(n_636), .B1(n_648), .B2(n_639), .C(n_645), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_647), .B(n_531), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_642), .A2(n_624), .B1(n_621), .B2(n_531), .Y(n_662) );
O2A1O1Ixp33_ASAP7_75t_L g663 ( .A1(n_635), .A2(n_579), .B(n_529), .C(n_522), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_631), .A2(n_624), .B1(n_501), .B2(n_512), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g665 ( .A1(n_640), .A2(n_501), .B1(n_512), .B2(n_548), .Y(n_665) );
AO22x2_ASAP7_75t_L g666 ( .A1(n_628), .A2(n_548), .B1(n_549), .B2(n_535), .Y(n_666) );
NAND4xp25_ASAP7_75t_L g667 ( .A(n_632), .B(n_637), .C(n_643), .D(n_644), .Y(n_667) );
O2A1O1Ixp33_ASAP7_75t_L g668 ( .A1(n_649), .A2(n_633), .B(n_641), .C(n_623), .Y(n_668) );
NOR3xp33_ASAP7_75t_SL g669 ( .A(n_667), .B(n_656), .C(n_668), .Y(n_669) );
CKINVDCx5p33_ASAP7_75t_R g670 ( .A(n_653), .Y(n_670) );
XNOR2xp5_ASAP7_75t_L g671 ( .A(n_651), .B(n_655), .Y(n_671) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_664), .A2(n_652), .B1(n_658), .B2(n_657), .Y(n_672) );
AND3x1_ASAP7_75t_L g673 ( .A(n_669), .B(n_660), .C(n_659), .Y(n_673) );
BUFx3_ASAP7_75t_L g674 ( .A(n_670), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g675 ( .A1(n_671), .A2(n_662), .B1(n_654), .B2(n_665), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_674), .Y(n_676) );
XNOR2xp5_ASAP7_75t_L g677 ( .A(n_673), .B(n_672), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_676), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_678), .A2(n_677), .B1(n_675), .B2(n_650), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g680 ( .A1(n_679), .A2(n_677), .B1(n_666), .B2(n_663), .C(n_661), .Y(n_680) );
endmodule