module fake_jpeg_30531_n_503 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_503);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_503;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_4),
.B(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx24_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_50),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_52),
.Y(n_132)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_55),
.Y(n_131)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_56),
.Y(n_136)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_58),
.Y(n_133)
);

CKINVDCx9p33_ASAP7_75t_R g59 ( 
.A(n_49),
.Y(n_59)
);

INVx5_ASAP7_75t_SL g157 ( 
.A(n_59),
.Y(n_157)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_29),
.B(n_8),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_62),
.B(n_69),
.Y(n_139)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_63),
.Y(n_150)
);

CKINVDCx6p67_ASAP7_75t_R g64 ( 
.A(n_27),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g140 ( 
.A(n_64),
.Y(n_140)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_29),
.B(n_8),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_70),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_37),
.B(n_8),
.C(n_14),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_71),
.B(n_26),
.Y(n_154)
);

BUFx24_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_72),
.Y(n_124)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_73),
.Y(n_158)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_74),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_37),
.B(n_8),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_84),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_20),
.B(n_7),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_76),
.B(n_78),
.Y(n_145)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_24),
.B(n_7),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_79),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

BUFx10_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_81),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_83),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_27),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_24),
.B(n_9),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_86),
.B(n_89),
.Y(n_159)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_9),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_20),
.B(n_6),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_97),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_92),
.Y(n_147)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

BUFx10_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_99),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_59),
.A2(n_35),
.B1(n_18),
.B2(n_41),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_104),
.A2(n_105),
.B1(n_118),
.B2(n_119),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_48),
.B1(n_28),
.B2(n_43),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_65),
.A2(n_48),
.B1(n_43),
.B2(n_28),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_117),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_89),
.B1(n_71),
.B2(n_68),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_64),
.A2(n_35),
.B1(n_18),
.B2(n_38),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_64),
.B(n_30),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_120),
.B(n_125),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_64),
.A2(n_35),
.B1(n_18),
.B2(n_38),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_121),
.A2(n_128),
.B1(n_130),
.B2(n_138),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_61),
.B(n_30),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_63),
.A2(n_30),
.B1(n_45),
.B2(n_44),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_85),
.A2(n_36),
.B1(n_38),
.B2(n_41),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_56),
.A2(n_18),
.B1(n_35),
.B2(n_38),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_88),
.A2(n_41),
.B1(n_35),
.B2(n_18),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_141),
.A2(n_149),
.B1(n_99),
.B2(n_67),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_73),
.A2(n_35),
.B1(n_41),
.B2(n_27),
.Y(n_149)
);

AND2x2_ASAP7_75t_SL g151 ( 
.A(n_53),
.B(n_0),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_80),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_94),
.B(n_34),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_19),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_154),
.B(n_21),
.Y(n_201)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_160),
.Y(n_219)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_108),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_161),
.Y(n_246)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_107),
.Y(n_162)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_162),
.Y(n_223)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_163),
.Y(n_226)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_102),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_164),
.Y(n_257)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_165),
.Y(n_225)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_167),
.Y(n_228)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_168),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_126),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_169),
.B(n_172),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_157),
.A2(n_74),
.B1(n_82),
.B2(n_81),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_171),
.A2(n_178),
.B1(n_192),
.B2(n_213),
.Y(n_239)
);

A2O1A1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_159),
.A2(n_72),
.B(n_44),
.C(n_39),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_173),
.B(n_206),
.Y(n_264)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_133),
.Y(n_174)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_174),
.Y(n_233)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_102),
.Y(n_175)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_175),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_L g176 ( 
.A1(n_111),
.A2(n_70),
.B1(n_66),
.B2(n_52),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_176),
.A2(n_183),
.B1(n_212),
.B2(n_141),
.Y(n_236)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_132),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_177),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_157),
.A2(n_79),
.B1(n_96),
.B2(n_93),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_134),
.Y(n_179)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_179),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_132),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_181),
.Y(n_261)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_124),
.Y(n_182)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_182),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_117),
.A2(n_91),
.B1(n_92),
.B2(n_60),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_184),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_135),
.Y(n_185)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_185),
.Y(n_251)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_116),
.Y(n_186)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_186),
.Y(n_253)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_115),
.Y(n_187)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_187),
.Y(n_254)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_116),
.Y(n_188)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_188),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_189),
.B(n_194),
.Y(n_234)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_110),
.Y(n_190)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_190),
.Y(n_260)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_143),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_191),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_128),
.A2(n_77),
.B1(n_55),
.B2(n_58),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_109),
.B(n_95),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_137),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_195),
.B(n_199),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_140),
.A2(n_51),
.B1(n_50),
.B2(n_54),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_196),
.Y(n_240)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_142),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_197),
.A2(n_205),
.B1(n_209),
.B2(n_210),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_100),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_198),
.Y(n_249)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_143),
.Y(n_199)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_100),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_200),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_139),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_126),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_202),
.B(n_204),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_113),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_203),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_135),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_126),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_124),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_SL g207 ( 
.A1(n_145),
.A2(n_72),
.B(n_98),
.Y(n_207)
);

NOR2x1_ASAP7_75t_R g229 ( 
.A(n_207),
.B(n_121),
.Y(n_229)
);

NAND3xp33_ASAP7_75t_L g208 ( 
.A(n_129),
.B(n_39),
.C(n_34),
.Y(n_208)
);

NOR2xp67_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_119),
.Y(n_232)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_140),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_123),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_111),
.A2(n_39),
.B1(n_21),
.B2(n_26),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_211),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_127),
.A2(n_34),
.B1(n_44),
.B2(n_26),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_127),
.A2(n_32),
.B1(n_42),
.B2(n_46),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_214),
.A2(n_57),
.B1(n_42),
.B2(n_32),
.Y(n_218)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_113),
.Y(n_215)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_142),
.Y(n_216)
);

BUFx2_ASAP7_75t_SL g217 ( 
.A(n_112),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_218),
.A2(n_236),
.B1(n_177),
.B2(n_156),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_166),
.A2(n_151),
.B1(n_125),
.B2(n_138),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_220),
.A2(n_224),
.B1(n_243),
.B2(n_255),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_221),
.B(n_112),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_173),
.B(n_154),
.C(n_151),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_222),
.B(n_230),
.C(n_162),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_166),
.A2(n_114),
.B1(n_148),
.B2(n_152),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_229),
.A2(n_104),
.B1(n_204),
.B2(n_185),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_172),
.B(n_139),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_232),
.B(n_206),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_193),
.A2(n_101),
.B(n_146),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_241),
.A2(n_247),
.B(n_182),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_180),
.A2(n_114),
.B1(n_148),
.B2(n_106),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_170),
.A2(n_146),
.B(n_158),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_209),
.A2(n_158),
.B1(n_136),
.B2(n_83),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_248),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_176),
.A2(n_130),
.B1(n_106),
.B2(n_144),
.Y(n_255)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_223),
.Y(n_265)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_265),
.Y(n_321)
);

BUFx2_ASAP7_75t_SL g266 ( 
.A(n_249),
.Y(n_266)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_266),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_250),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_267),
.B(n_268),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_250),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_269),
.B(n_296),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_270),
.B(n_274),
.Y(n_318)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_256),
.Y(n_271)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_271),
.Y(n_343)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_223),
.Y(n_272)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_272),
.Y(n_335)
);

A2O1A1Ixp33_ASAP7_75t_SL g319 ( 
.A1(n_273),
.A2(n_112),
.B(n_252),
.C(n_228),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_167),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_275),
.Y(n_336)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_251),
.Y(n_276)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_276),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_160),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_277),
.B(n_281),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_250),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_278),
.B(n_280),
.Y(n_344)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_235),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_279),
.Y(n_331)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_247),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_221),
.B(n_210),
.Y(n_281)
);

INVx4_ASAP7_75t_SL g283 ( 
.A(n_227),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_283),
.B(n_286),
.Y(n_322)
);

OAI32xp33_ASAP7_75t_L g284 ( 
.A1(n_230),
.A2(n_179),
.A3(n_184),
.B1(n_168),
.B2(n_174),
.Y(n_284)
);

OAI32xp33_ASAP7_75t_L g329 ( 
.A1(n_284),
.A2(n_237),
.A3(n_233),
.B1(n_219),
.B2(n_225),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_165),
.Y(n_286)
);

BUFx12f_ASAP7_75t_L g287 ( 
.A(n_235),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_287),
.A2(n_288),
.B1(n_290),
.B2(n_291),
.Y(n_323)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_235),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_289),
.A2(n_293),
.B1(n_302),
.B2(n_305),
.Y(n_340)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_226),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_219),
.Y(n_291)
);

AOI32xp33_ASAP7_75t_L g292 ( 
.A1(n_229),
.A2(n_149),
.A3(n_203),
.B1(n_136),
.B2(n_215),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_306),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_220),
.A2(n_197),
.B1(n_216),
.B2(n_175),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_222),
.B(n_164),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_299),
.C(n_307),
.Y(n_311)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_226),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_295),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_264),
.B(n_234),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_240),
.A2(n_200),
.B1(n_198),
.B2(n_185),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_297),
.A2(n_304),
.B1(n_262),
.B2(n_252),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_245),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_298),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_264),
.B(n_186),
.Y(n_299)
);

OA22x2_ASAP7_75t_L g312 ( 
.A1(n_300),
.A2(n_256),
.B1(n_242),
.B2(n_258),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_231),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_301),
.A2(n_262),
.B(n_249),
.Y(n_317)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_238),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_241),
.A2(n_155),
.B1(n_144),
.B2(n_191),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_303),
.A2(n_260),
.B1(n_254),
.B2(n_242),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_246),
.B(n_199),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_238),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_260),
.B(n_188),
.C(n_204),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_301),
.A2(n_240),
.B1(n_239),
.B2(n_236),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_308),
.A2(n_310),
.B1(n_324),
.B2(n_332),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_285),
.A2(n_239),
.B1(n_255),
.B2(n_244),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_312),
.A2(n_327),
.B1(n_338),
.B2(n_341),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_315),
.A2(n_316),
.B1(n_328),
.B2(n_330),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_282),
.A2(n_254),
.B1(n_181),
.B2(n_261),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_317),
.A2(n_319),
.B(n_307),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_285),
.A2(n_263),
.B1(n_258),
.B2(n_253),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_294),
.B(n_253),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_325),
.B(n_326),
.C(n_337),
.Y(n_353)
);

MAJx2_ASAP7_75t_L g326 ( 
.A(n_269),
.B(n_228),
.C(n_263),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_282),
.A2(n_237),
.B1(n_233),
.B2(n_227),
.Y(n_328)
);

OAI32xp33_ASAP7_75t_L g364 ( 
.A1(n_329),
.A2(n_287),
.A3(n_19),
.B1(n_6),
.B2(n_12),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_273),
.A2(n_225),
.B1(n_257),
.B2(n_42),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_300),
.A2(n_257),
.B1(n_32),
.B2(n_19),
.Y(n_332)
);

OAI32xp33_ASAP7_75t_L g334 ( 
.A1(n_277),
.A2(n_257),
.A3(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_334)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_334),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_306),
.B(n_19),
.C(n_1),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_303),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_338)
);

OAI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_284),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_314),
.A2(n_286),
.B(n_296),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_347),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_308),
.A2(n_298),
.B1(n_305),
.B2(n_302),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_348),
.A2(n_352),
.B1(n_361),
.B2(n_365),
.Y(n_397)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_321),
.Y(n_349)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_349),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_342),
.B(n_265),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_350),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_322),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_351),
.B(n_375),
.Y(n_395)
);

OAI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_312),
.A2(n_319),
.B1(n_329),
.B2(n_316),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_344),
.A2(n_276),
.B(n_275),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_354),
.A2(n_362),
.B(n_368),
.Y(n_382)
);

AO21x1_ASAP7_75t_L g399 ( 
.A1(n_355),
.A2(n_358),
.B(n_373),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_342),
.B(n_299),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_356),
.B(n_363),
.Y(n_389)
);

AOI322xp5_ASAP7_75t_L g358 ( 
.A1(n_309),
.A2(n_272),
.A3(n_279),
.B1(n_288),
.B2(n_290),
.C1(n_295),
.C2(n_287),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_322),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_359),
.Y(n_384)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_321),
.Y(n_360)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_360),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_310),
.A2(n_271),
.B1(n_283),
.B2(n_291),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_317),
.A2(n_287),
.B(n_19),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_330),
.Y(n_363)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_364),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_340),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_335),
.Y(n_366)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_366),
.Y(n_393)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_335),
.Y(n_367)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_367),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_309),
.A2(n_5),
.B(n_13),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_311),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_369),
.A2(n_370),
.B1(n_313),
.B2(n_315),
.Y(n_400)
);

OAI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_312),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_313),
.B(n_4),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_371),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_319),
.A2(n_5),
.B(n_11),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_325),
.B(n_5),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_374),
.B(n_337),
.C(n_320),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_319),
.A2(n_11),
.B(n_13),
.Y(n_375)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_336),
.Y(n_377)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_377),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_353),
.B(n_311),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_379),
.B(n_381),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_350),
.B(n_318),
.Y(n_380)
);

CKINVDCx14_ASAP7_75t_R g427 ( 
.A(n_380),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_353),
.B(n_333),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_385),
.B(n_387),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_353),
.B(n_333),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_346),
.A2(n_312),
.B1(n_324),
.B2(n_326),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_388),
.A2(n_361),
.B1(n_370),
.B2(n_354),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_374),
.B(n_320),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_390),
.B(n_392),
.C(n_396),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_374),
.B(n_332),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_347),
.B(n_328),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_347),
.B(n_339),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_398),
.B(n_402),
.C(n_405),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_400),
.B(n_357),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_356),
.B(n_339),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_368),
.B(n_336),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_397),
.A2(n_346),
.B1(n_351),
.B2(n_359),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_407),
.A2(n_417),
.B1(n_420),
.B2(n_423),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_391),
.A2(n_357),
.B1(n_352),
.B2(n_348),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_408),
.A2(n_409),
.B1(n_411),
.B2(n_414),
.Y(n_436)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_386),
.Y(n_410)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_410),
.Y(n_438)
);

OAI21x1_ASAP7_75t_L g412 ( 
.A1(n_395),
.A2(n_355),
.B(n_319),
.Y(n_412)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_412),
.Y(n_440)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_386),
.Y(n_413)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_413),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_396),
.A2(n_391),
.B1(n_388),
.B2(n_383),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_378),
.B(n_369),
.Y(n_415)
);

CKINVDCx14_ASAP7_75t_R g432 ( 
.A(n_415),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_397),
.A2(n_372),
.B1(n_376),
.B2(n_364),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_393),
.Y(n_418)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_418),
.Y(n_442)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_393),
.Y(n_419)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_419),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_384),
.A2(n_372),
.B1(n_376),
.B2(n_358),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_401),
.Y(n_421)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_421),
.B(n_422),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_401),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_400),
.A2(n_372),
.B1(n_373),
.B2(n_375),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_399),
.A2(n_362),
.B(n_377),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_424),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_389),
.A2(n_323),
.B1(n_349),
.B2(n_367),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_425),
.B(n_398),
.Y(n_443)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_403),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_428),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_416),
.B(n_379),
.C(n_381),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_430),
.B(n_431),
.C(n_437),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_416),
.B(n_387),
.C(n_402),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_429),
.B(n_385),
.C(n_390),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_443),
.A2(n_417),
.B1(n_412),
.B2(n_421),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_429),
.B(n_389),
.C(n_392),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_444),
.B(n_445),
.C(n_422),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_406),
.B(n_405),
.C(n_382),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_406),
.B(n_426),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_447),
.B(n_448),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_426),
.B(n_399),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_414),
.B(n_382),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_449),
.B(n_423),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_435),
.A2(n_408),
.B1(n_411),
.B2(n_409),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_450),
.A2(n_436),
.B1(n_435),
.B2(n_449),
.Y(n_468)
);

BUFx24_ASAP7_75t_SL g451 ( 
.A(n_432),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_451),
.B(n_453),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_433),
.A2(n_424),
.B(n_420),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_452),
.A2(n_454),
.B(n_460),
.Y(n_466)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_439),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_433),
.A2(n_407),
.B(n_425),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_439),
.B(n_427),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_455),
.B(n_461),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_456),
.B(n_462),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_459),
.B(n_445),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_440),
.A2(n_428),
.B(n_419),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_447),
.B(n_404),
.Y(n_461)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_438),
.Y(n_463)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_463),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_443),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_464),
.B(n_444),
.Y(n_467)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_467),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_468),
.A2(n_450),
.B1(n_452),
.B2(n_454),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_462),
.B(n_448),
.C(n_430),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_470),
.A2(n_473),
.B(n_477),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_471),
.B(n_474),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_457),
.B(n_437),
.C(n_431),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_457),
.B(n_446),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_459),
.A2(n_442),
.B1(n_441),
.B2(n_434),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_475),
.B(n_469),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_458),
.B(n_418),
.C(n_413),
.Y(n_477)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_479),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_471),
.B(n_458),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_482),
.A2(n_484),
.B(n_477),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_468),
.A2(n_460),
.B1(n_410),
.B2(n_403),
.Y(n_483)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_483),
.Y(n_492)
);

OAI321xp33_ASAP7_75t_L g484 ( 
.A1(n_466),
.A2(n_334),
.A3(n_394),
.B1(n_360),
.B2(n_366),
.C(n_371),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_485),
.B(n_486),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_476),
.B(n_331),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_481),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_487),
.B(n_489),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_478),
.A2(n_472),
.B(n_470),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_490),
.A2(n_473),
.B(n_482),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_494),
.B(n_495),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_488),
.B(n_465),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_491),
.A2(n_476),
.B(n_480),
.Y(n_496)
);

A2O1A1O1Ixp25_ASAP7_75t_L g498 ( 
.A1(n_496),
.A2(n_492),
.B(n_480),
.C(n_474),
.D(n_479),
.Y(n_498)
);

OAI31xp33_ASAP7_75t_SL g499 ( 
.A1(n_498),
.A2(n_493),
.A3(n_483),
.B(n_475),
.Y(n_499)
);

OAI321xp33_ASAP7_75t_L g500 ( 
.A1(n_499),
.A2(n_497),
.A3(n_343),
.B1(n_331),
.B2(n_345),
.C(n_365),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_500),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_501),
.A2(n_343),
.B(n_345),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_502),
.A2(n_15),
.B(n_501),
.Y(n_503)
);


endmodule