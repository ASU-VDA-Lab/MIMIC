module fake_ibex_1188_n_4047 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_861, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_840, n_561, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_158, n_859, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_875, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_373, n_854, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_835, n_168, n_526, n_785, n_155, n_824, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_852, n_789, n_654, n_656, n_724, n_437, n_731, n_602, n_842, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_851, n_689, n_793, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_847, n_830, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_869, n_718, n_801, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_803, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_776, n_409, n_582, n_818, n_653, n_214, n_238, n_579, n_843, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_485, n_870, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_572, n_867, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_4047);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_861;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_840;
input n_561;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_158;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_875;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_854;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_852;
input n_789;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_842;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_851;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_847;
input n_830;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_869;
input n_718;
input n_801;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_867;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;

output n_4047;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_3590;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_3812;
wire n_2017;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_2290;
wire n_3750;
wire n_3838;
wire n_957;
wire n_3272;
wire n_3674;
wire n_3255;
wire n_1652;
wire n_969;
wire n_1859;
wire n_2183;
wire n_1954;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_2682;
wire n_3605;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_4004;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_1722;
wire n_3931;
wire n_911;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_3340;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3411;
wire n_3025;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_2230;
wire n_963;
wire n_1782;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_3904;
wire n_3175;
wire n_3729;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_3984;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_1730;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_3211;
wire n_3479;
wire n_1840;
wire n_2837;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_3982;
wire n_2605;
wire n_2343;
wire n_2887;
wire n_1641;
wire n_2565;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_4031;
wire n_3724;
wire n_939;
wire n_1636;
wire n_1687;
wire n_3192;
wire n_3533;
wire n_3753;
wire n_3896;
wire n_2192;
wire n_1766;
wire n_3566;
wire n_3184;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_3890;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_1937;
wire n_2311;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_3839;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3509;
wire n_3472;
wire n_1749;
wire n_1680;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_3976;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_4002;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3987;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_3969;
wire n_1081;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_3996;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_4015;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3881;
wire n_3884;
wire n_3507;
wire n_3949;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_2333;
wire n_2436;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_3699;
wire n_1955;
wire n_3668;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3148;
wire n_3022;
wire n_2822;
wire n_3766;
wire n_4014;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_3973;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3977;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_2215;
wire n_1449;
wire n_1071;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3979;
wire n_3714;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_3943;
wire n_3809;
wire n_979;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3910;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_3667;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_3822;
wire n_1637;
wire n_3310;
wire n_2900;
wire n_3858;
wire n_1401;
wire n_3764;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_1620;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3225;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_1653;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_1296;
wire n_3060;
wire n_971;
wire n_1326;
wire n_1350;
wire n_3627;
wire n_906;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_3777;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_2541;
wire n_2987;
wire n_881;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3808;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_4012;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_3874;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_3652;
wire n_1818;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_3241;
wire n_2746;
wire n_2256;
wire n_3317;
wire n_3800;
wire n_3887;
wire n_3963;
wire n_3461;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_3583;
wire n_2019;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_889;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_3950;
wire n_2070;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_3320;
wire n_3117;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_1964;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_3957;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3634;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3788;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_3626;
wire n_3733;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_3986;
wire n_2853;
wire n_1932;
wire n_3775;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_1189;
wire n_4008;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_4039;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_3815;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1421;
wire n_1203;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_1793;
wire n_2573;
wire n_1237;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_3849;
wire n_965;
wire n_1109;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_4040;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3855;
wire n_3357;
wire n_4033;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_1236;
wire n_3364;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3188;
wire n_3037;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1477;
wire n_1184;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_4005;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_3680;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_3503;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_3568;
wire n_944;
wire n_3312;
wire n_3003;
wire n_1848;
wire n_4009;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_2252;
wire n_1982;
wire n_3932;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_3331;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_4011;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_2991;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1485;
wire n_1069;
wire n_2239;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_1345;
wire n_2434;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3584;
wire n_3470;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3797;
wire n_1115;
wire n_998;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_2823;
wire n_3274;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_4042;
wire n_2525;
wire n_3829;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1523;
wire n_1086;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_4041;
wire n_1836;
wire n_2398;
wire n_3401;
wire n_3032;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_3978;
wire n_2570;
wire n_3123;
wire n_4025;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_3948;
wire n_1599;
wire n_1400;
wire n_1539;
wire n_1806;
wire n_2711;
wire n_3070;
wire n_2842;
wire n_3477;
wire n_2635;
wire n_3646;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3897;
wire n_4024;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_4010;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_1574;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_1746;
wire n_2716;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_3495;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_4035;
wire n_2781;
wire n_3419;
wire n_3629;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_3999;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_3167;
wire n_3687;
wire n_997;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_1428;
wire n_2691;
wire n_4026;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_2463;
wire n_2654;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_3877;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_2439;
wire n_1925;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_1475;
wire n_3337;
wire n_2465;
wire n_1263;
wire n_3316;
wire n_3925;
wire n_1185;
wire n_1683;
wire n_3575;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_3955;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_4030;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1845;
wire n_1104;
wire n_2205;
wire n_1011;
wire n_2875;
wire n_2684;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_3835;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_3902;
wire n_3927;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_1815;
wire n_972;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_920;
wire n_2442;
wire n_3985;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_2997;
wire n_3747;
wire n_1349;
wire n_1331;
wire n_1223;
wire n_961;
wire n_991;
wire n_2127;
wire n_3735;
wire n_1323;
wire n_3891;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_4003;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_996;
wire n_3632;
wire n_3914;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_3372;
wire n_3499;
wire n_3552;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_3990;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_4044;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2187;
wire n_2105;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3269;
wire n_3029;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_2647;
wire n_1626;
wire n_3995;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_4000;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_3908;
wire n_1099;
wire n_2141;
wire n_3696;
wire n_3113;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3960;
wire n_4007;
wire n_3608;
wire n_3190;
wire n_1524;
wire n_1055;
wire n_3878;
wire n_4016;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_4028;
wire n_2210;
wire n_1517;
wire n_3940;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3778;
wire n_3912;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_3993;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_4001;
wire n_1289;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_3356;
wire n_1191;
wire n_2004;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_1942;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_2274;
wire n_2698;
wire n_3899;
wire n_1617;
wire n_1839;
wire n_3930;
wire n_1587;
wire n_2555;
wire n_2330;
wire n_2639;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_3760;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_4021;
wire n_1538;
wire n_2528;
wire n_3773;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3424;
wire n_3462;
wire n_3745;
wire n_2437;
wire n_2351;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_993;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_3314;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_1241;
wire n_3645;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_4019;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_2154;
wire n_1976;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_3162;
wire n_2984;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_1647;
wire n_1901;
wire n_3333;
wire n_3096;
wire n_3705;
wire n_4023;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1415;
wire n_1238;
wire n_3959;
wire n_3743;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_3860;
wire n_2137;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3493;
wire n_2447;
wire n_3044;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_4034;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_3273;
wire n_950;
wire n_2700;
wire n_3139;
wire n_1222;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3647;
wire n_3623;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_4029;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_919;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_3604;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_3649;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_3740;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2576;
wire n_2348;
wire n_2675;
wire n_2417;
wire n_2043;
wire n_3601;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2973;
wire n_3651;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3085;
wire n_3059;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_3994;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3648;
wire n_3234;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_4032;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_2367;
wire n_3236;
wire n_3576;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3062;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_3391;
wire n_4017;
wire n_1542;
wire n_946;
wire n_1547;
wire n_1362;
wire n_1586;
wire n_3497;
wire n_1097;
wire n_3354;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3586;
wire n_3561;
wire n_956;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1887;
wire n_1212;
wire n_1199;
wire n_3400;
wire n_3942;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_1828;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_3774;
wire n_3972;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_4036;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1361;
wire n_1187;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_3173;
wire n_2872;
wire n_3102;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_3998;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_3989;
wire n_2119;
wire n_1010;
wire n_3844;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3305;
wire n_3051;
wire n_1635;
wire n_1572;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_3343;
wire n_3752;
wire n_3786;
wire n_2637;
wire n_1329;
wire n_2409;
wire n_2337;
wire n_4045;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1369;
wire n_1297;
wire n_1912;
wire n_3143;
wire n_3543;
wire n_1734;
wire n_3655;
wire n_3742;
wire n_3791;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_3532;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_3725;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_2914;
wire n_1833;
wire n_3551;
wire n_2371;
wire n_914;
wire n_3992;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_3326;
wire n_1168;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_2942;
wire n_3947;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_2296;
wire n_3782;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_3831;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_2310;
wire n_3223;
wire n_3318;
wire n_4013;
wire n_1397;
wire n_1211;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1193;
wire n_980;
wire n_1488;
wire n_2928;
wire n_3380;
wire n_2227;
wire n_2652;
wire n_3483;
wire n_1074;
wire n_3557;
wire n_3596;
wire n_3207;
wire n_3067;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3369;
wire n_3823;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_1022;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_3124;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3286;
wire n_1092;
wire n_4038;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3837;
wire n_3612;
wire n_3046;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1142;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1516;
wire n_1027;
wire n_3893;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_2357;
wire n_2303;
wire n_2618;
wire n_2653;
wire n_2855;
wire n_3938;
wire n_924;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_2136;
wire n_3617;
wire n_4027;
wire n_3602;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_1450;
wire n_2302;
wire n_2082;
wire n_2560;
wire n_2453;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2802;
wire n_2443;
wire n_3189;
wire n_3052;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_2066;
wire n_1974;
wire n_1158;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_4046;
wire n_2770;
wire n_2961;
wire n_2704;
wire n_2996;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_2168;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_3613;
wire n_1383;
wire n_990;
wire n_3675;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_4018;
wire n_2378;
wire n_888;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_2969;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_3933;
wire n_955;
wire n_1916;
wire n_1333;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_3873;
wire n_3738;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_3793;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_3988;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_1355;
wire n_3691;
wire n_2544;
wire n_3193;
wire n_3501;
wire n_3635;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1780;
wire n_1091;
wire n_1678;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_1525;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_3685;
wire n_3851;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_3768;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_3980;
wire n_2430;
wire n_2676;
wire n_921;
wire n_2673;
wire n_3515;
wire n_3489;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3494;
wire n_3040;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_3677;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;
wire n_2658;

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_208),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_166),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_584),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_177),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_843),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_378),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_851),
.Y(n_885)
);

CKINVDCx20_ASAP7_75t_R g886 ( 
.A(n_824),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_877),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_549),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_825),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_836),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_466),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_469),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_558),
.Y(n_893)
);

BUFx5_ASAP7_75t_L g894 ( 
.A(n_267),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_589),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_830),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_21),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_124),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_809),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_532),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_815),
.Y(n_901)
);

CKINVDCx20_ASAP7_75t_R g902 ( 
.A(n_732),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_854),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_127),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_153),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_223),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_755),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_147),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_869),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_723),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_83),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_261),
.Y(n_912)
);

CKINVDCx20_ASAP7_75t_R g913 ( 
.A(n_61),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_248),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_257),
.Y(n_915)
);

INVx2_ASAP7_75t_SL g916 ( 
.A(n_618),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_783),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_803),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_814),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_377),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_70),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_202),
.Y(n_922)
);

BUFx8_ASAP7_75t_SL g923 ( 
.A(n_292),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_816),
.Y(n_924)
);

CKINVDCx16_ASAP7_75t_R g925 ( 
.A(n_867),
.Y(n_925)
);

CKINVDCx20_ASAP7_75t_R g926 ( 
.A(n_290),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_797),
.Y(n_927)
);

CKINVDCx16_ASAP7_75t_R g928 ( 
.A(n_571),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_874),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_53),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_435),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_844),
.Y(n_932)
);

CKINVDCx20_ASAP7_75t_R g933 ( 
.A(n_812),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_304),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_696),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_262),
.Y(n_936)
);

BUFx5_ASAP7_75t_L g937 ( 
.A(n_783),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_832),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_95),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_278),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_832),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_230),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_117),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_288),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_827),
.Y(n_945)
);

CKINVDCx20_ASAP7_75t_R g946 ( 
.A(n_265),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_801),
.Y(n_947)
);

BUFx10_ASAP7_75t_L g948 ( 
.A(n_299),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_862),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_821),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_280),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_423),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_329),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_142),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_793),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_870),
.Y(n_956)
);

BUFx3_ASAP7_75t_L g957 ( 
.A(n_338),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_108),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_107),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_188),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_438),
.Y(n_961)
);

CKINVDCx20_ASAP7_75t_R g962 ( 
.A(n_690),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_515),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_269),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_90),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_590),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_565),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_399),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_25),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_550),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_560),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_671),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_154),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_286),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_829),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_672),
.Y(n_976)
);

CKINVDCx20_ASAP7_75t_R g977 ( 
.A(n_384),
.Y(n_977)
);

BUFx3_ASAP7_75t_L g978 ( 
.A(n_845),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_805),
.Y(n_979)
);

CKINVDCx20_ASAP7_75t_R g980 ( 
.A(n_817),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_206),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_441),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_373),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_517),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_743),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_10),
.Y(n_986)
);

BUFx2_ASAP7_75t_SL g987 ( 
.A(n_508),
.Y(n_987)
);

BUFx5_ASAP7_75t_L g988 ( 
.A(n_779),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_837),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_17),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_811),
.Y(n_991)
);

CKINVDCx20_ASAP7_75t_R g992 ( 
.A(n_405),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_467),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_875),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_566),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_140),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_807),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_502),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_21),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_871),
.Y(n_1000)
);

CKINVDCx20_ASAP7_75t_R g1001 ( 
.A(n_188),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_670),
.Y(n_1002)
);

CKINVDCx20_ASAP7_75t_R g1003 ( 
.A(n_586),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_654),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_866),
.Y(n_1005)
);

INVx4_ASAP7_75t_R g1006 ( 
.A(n_868),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_254),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_804),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_597),
.Y(n_1009)
);

INVx2_ASAP7_75t_SL g1010 ( 
.A(n_557),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_353),
.Y(n_1011)
);

BUFx5_ASAP7_75t_L g1012 ( 
.A(n_800),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_486),
.Y(n_1013)
);

BUFx10_ASAP7_75t_L g1014 ( 
.A(n_659),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_430),
.Y(n_1015)
);

CKINVDCx16_ASAP7_75t_R g1016 ( 
.A(n_456),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_188),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_864),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_199),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_792),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_772),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_846),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_813),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_853),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_690),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_168),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_840),
.Y(n_1027)
);

BUFx10_ASAP7_75t_L g1028 ( 
.A(n_135),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_859),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_474),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_323),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_362),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_684),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_385),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_634),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_838),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_147),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_92),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_818),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_289),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_469),
.Y(n_1041)
);

CKINVDCx20_ASAP7_75t_R g1042 ( 
.A(n_707),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_675),
.Y(n_1043)
);

CKINVDCx14_ASAP7_75t_R g1044 ( 
.A(n_833),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_207),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_289),
.Y(n_1046)
);

BUFx5_ASAP7_75t_L g1047 ( 
.A(n_495),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_266),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_40),
.Y(n_1049)
);

BUFx3_ASAP7_75t_L g1050 ( 
.A(n_219),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_187),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_277),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_794),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_393),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_645),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_28),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_506),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_481),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_808),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_554),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_476),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_628),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_390),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_430),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_826),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_310),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_265),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_567),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_156),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_561),
.Y(n_1070)
);

BUFx2_ASAP7_75t_SL g1071 ( 
.A(n_751),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_215),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_340),
.Y(n_1073)
);

INVx1_ASAP7_75t_SL g1074 ( 
.A(n_462),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_68),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_238),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_0),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_587),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_564),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_52),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_412),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_125),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_186),
.Y(n_1083)
);

HB1xp67_ASAP7_75t_L g1084 ( 
.A(n_395),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_48),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_652),
.Y(n_1086)
);

INVxp67_ASAP7_75t_L g1087 ( 
.A(n_873),
.Y(n_1087)
);

CKINVDCx20_ASAP7_75t_R g1088 ( 
.A(n_255),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_872),
.Y(n_1089)
);

INVx1_ASAP7_75t_SL g1090 ( 
.A(n_250),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_814),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_138),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_863),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_237),
.Y(n_1094)
);

CKINVDCx16_ASAP7_75t_R g1095 ( 
.A(n_642),
.Y(n_1095)
);

BUFx2_ASAP7_75t_L g1096 ( 
.A(n_552),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_860),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_86),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_865),
.Y(n_1099)
);

INVxp67_ASAP7_75t_L g1100 ( 
.A(n_831),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_828),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_234),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_310),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_735),
.Y(n_1104)
);

BUFx10_ASAP7_75t_L g1105 ( 
.A(n_849),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_90),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_842),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_835),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_850),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_812),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_643),
.Y(n_1111)
);

CKINVDCx20_ASAP7_75t_R g1112 ( 
.A(n_852),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_710),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_615),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_806),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_857),
.Y(n_1116)
);

BUFx3_ASAP7_75t_L g1117 ( 
.A(n_533),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_697),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_498),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_488),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_425),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_453),
.Y(n_1122)
);

CKINVDCx20_ASAP7_75t_R g1123 ( 
.A(n_608),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_119),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_210),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_67),
.Y(n_1126)
);

CKINVDCx20_ASAP7_75t_R g1127 ( 
.A(n_226),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_144),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_677),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_815),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_594),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_854),
.Y(n_1132)
);

BUFx3_ASAP7_75t_L g1133 ( 
.A(n_810),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_616),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_328),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_729),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_712),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_592),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_358),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_93),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_42),
.Y(n_1141)
);

INVx2_ASAP7_75t_SL g1142 ( 
.A(n_272),
.Y(n_1142)
);

INVx2_ASAP7_75t_SL g1143 ( 
.A(n_240),
.Y(n_1143)
);

INVxp67_ASAP7_75t_SL g1144 ( 
.A(n_420),
.Y(n_1144)
);

BUFx10_ASAP7_75t_L g1145 ( 
.A(n_510),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_339),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_101),
.Y(n_1147)
);

BUFx8_ASAP7_75t_SL g1148 ( 
.A(n_780),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_637),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_88),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_590),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_590),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_497),
.Y(n_1153)
);

INVx1_ASAP7_75t_SL g1154 ( 
.A(n_40),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_287),
.Y(n_1155)
);

CKINVDCx20_ASAP7_75t_R g1156 ( 
.A(n_477),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_847),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_563),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_302),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_861),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_754),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_870),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_413),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_575),
.Y(n_1164)
);

BUFx5_ASAP7_75t_L g1165 ( 
.A(n_224),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_376),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_612),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_384),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_457),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_795),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_132),
.Y(n_1171)
);

CKINVDCx20_ASAP7_75t_R g1172 ( 
.A(n_6),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_510),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_841),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_776),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_746),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_155),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_371),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_227),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_868),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_848),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_855),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_518),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_522),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_574),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_17),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_145),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_858),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_311),
.Y(n_1189)
);

CKINVDCx20_ASAP7_75t_R g1190 ( 
.A(n_314),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_613),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_480),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_538),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_555),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_466),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_258),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_823),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_756),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_798),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_799),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_120),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_236),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_820),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_35),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_796),
.Y(n_1205)
);

CKINVDCx14_ASAP7_75t_R g1206 ( 
.A(n_798),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_278),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_29),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_424),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_856),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_386),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_81),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_362),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_775),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_822),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_528),
.Y(n_1216)
);

INVx1_ASAP7_75t_SL g1217 ( 
.A(n_314),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_549),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_231),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_732),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_468),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_665),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_309),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_834),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_517),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_641),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_436),
.Y(n_1227)
);

CKINVDCx16_ASAP7_75t_R g1228 ( 
.A(n_376),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_769),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_40),
.Y(n_1230)
);

INVx2_ASAP7_75t_SL g1231 ( 
.A(n_876),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_160),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_101),
.Y(n_1233)
);

CKINVDCx20_ASAP7_75t_R g1234 ( 
.A(n_330),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_56),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_537),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_153),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_122),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_359),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_618),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_322),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_824),
.Y(n_1242)
);

INVxp67_ASAP7_75t_L g1243 ( 
.A(n_777),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_810),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_186),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_71),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_626),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_664),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_231),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_160),
.Y(n_1250)
);

CKINVDCx20_ASAP7_75t_R g1251 ( 
.A(n_839),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_284),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_423),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_232),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_93),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_463),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_64),
.Y(n_1257)
);

INVx1_ASAP7_75t_SL g1258 ( 
.A(n_736),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_172),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_568),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_82),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_145),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_213),
.Y(n_1263)
);

CKINVDCx20_ASAP7_75t_R g1264 ( 
.A(n_802),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_324),
.Y(n_1265)
);

INVx1_ASAP7_75t_SL g1266 ( 
.A(n_366),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_874),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_398),
.Y(n_1268)
);

BUFx10_ASAP7_75t_L g1269 ( 
.A(n_490),
.Y(n_1269)
);

INVx1_ASAP7_75t_SL g1270 ( 
.A(n_85),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_340),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_819),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_937),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_916),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_937),
.Y(n_1275)
);

INVxp67_ASAP7_75t_SL g1276 ( 
.A(n_1081),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1010),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1142),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1143),
.Y(n_1279)
);

INVxp33_ASAP7_75t_L g1280 ( 
.A(n_892),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_918),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_937),
.Y(n_1282)
);

INVxp33_ASAP7_75t_SL g1283 ( 
.A(n_998),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_937),
.Y(n_1284)
);

INVxp33_ASAP7_75t_SL g1285 ( 
.A(n_1084),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1045),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_923),
.Y(n_1287)
);

INVxp33_ASAP7_75t_L g1288 ( 
.A(n_1096),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1138),
.Y(n_1289)
);

CKINVDCx20_ASAP7_75t_R g1290 ( 
.A(n_904),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1223),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1271),
.Y(n_1292)
);

INVxp67_ASAP7_75t_L g1293 ( 
.A(n_922),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_937),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_913),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_1044),
.Y(n_1296)
);

INVxp67_ASAP7_75t_L g1297 ( 
.A(n_922),
.Y(n_1297)
);

INVxp67_ASAP7_75t_L g1298 ( 
.A(n_951),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_1044),
.Y(n_1299)
);

CKINVDCx16_ASAP7_75t_R g1300 ( 
.A(n_928),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1206),
.Y(n_1301)
);

INVx4_ASAP7_75t_R g1302 ( 
.A(n_951),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1065),
.B(n_1016),
.Y(n_1303)
);

CKINVDCx20_ASAP7_75t_R g1304 ( 
.A(n_926),
.Y(n_1304)
);

CKINVDCx20_ASAP7_75t_R g1305 ( 
.A(n_946),
.Y(n_1305)
);

INVxp67_ASAP7_75t_L g1306 ( 
.A(n_957),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_912),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_1206),
.Y(n_1308)
);

INVxp67_ASAP7_75t_SL g1309 ( 
.A(n_957),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_921),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_1148),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_930),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_931),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_939),
.Y(n_1314)
);

INVxp67_ASAP7_75t_L g1315 ( 
.A(n_986),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_952),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_958),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_960),
.Y(n_1318)
);

NOR2xp67_ASAP7_75t_L g1319 ( 
.A(n_907),
.B(n_0),
.Y(n_1319)
);

INVxp67_ASAP7_75t_SL g1320 ( 
.A(n_986),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_977),
.Y(n_1321)
);

INVxp33_ASAP7_75t_SL g1322 ( 
.A(n_1149),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_937),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_1228),
.Y(n_1324)
);

INVxp67_ASAP7_75t_L g1325 ( 
.A(n_1040),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_988),
.Y(n_1326)
);

INVxp33_ASAP7_75t_SL g1327 ( 
.A(n_1272),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_968),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_971),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_974),
.Y(n_1330)
);

CKINVDCx16_ASAP7_75t_R g1331 ( 
.A(n_925),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_981),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_993),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1007),
.Y(n_1334)
);

CKINVDCx20_ASAP7_75t_R g1335 ( 
.A(n_992),
.Y(n_1335)
);

INVxp67_ASAP7_75t_SL g1336 ( 
.A(n_1050),
.Y(n_1336)
);

CKINVDCx20_ASAP7_75t_R g1337 ( 
.A(n_1001),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1019),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1026),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_978),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1034),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_978),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1048),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1051),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1054),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_988),
.Y(n_1346)
);

INVxp33_ASAP7_75t_SL g1347 ( 
.A(n_879),
.Y(n_1347)
);

CKINVDCx20_ASAP7_75t_R g1348 ( 
.A(n_1003),
.Y(n_1348)
);

INVxp33_ASAP7_75t_L g1349 ( 
.A(n_883),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1064),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1066),
.Y(n_1351)
);

BUFx6f_ASAP7_75t_L g1352 ( 
.A(n_935),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1068),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1073),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_988),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1083),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1094),
.Y(n_1357)
);

INVx3_ASAP7_75t_L g1358 ( 
.A(n_948),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_880),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_882),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_884),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_1015),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_888),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1293),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1293),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1297),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1297),
.Y(n_1367)
);

AND2x6_ASAP7_75t_L g1368 ( 
.A(n_1358),
.B(n_1052),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1298),
.Y(n_1369)
);

BUFx6f_ASAP7_75t_L g1370 ( 
.A(n_1352),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1298),
.Y(n_1371)
);

AOI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1283),
.A2(n_895),
.B1(n_898),
.B2(n_897),
.Y(n_1372)
);

BUFx6f_ASAP7_75t_L g1373 ( 
.A(n_1352),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1340),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1342),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1306),
.B(n_900),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_1274),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1273),
.Y(n_1378)
);

BUFx6f_ASAP7_75t_L g1379 ( 
.A(n_1352),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1275),
.A2(n_996),
.B(n_915),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1315),
.B(n_1325),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1282),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1284),
.Y(n_1383)
);

AOI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1285),
.A2(n_905),
.B1(n_908),
.B2(n_906),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1276),
.B(n_911),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1309),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1320),
.B(n_914),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1336),
.B(n_920),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1294),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1323),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1280),
.B(n_1361),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1277),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1286),
.B(n_1231),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1278),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1288),
.B(n_948),
.Y(n_1395)
);

BUFx6f_ASAP7_75t_L g1396 ( 
.A(n_1326),
.Y(n_1396)
);

OA21x2_ASAP7_75t_L g1397 ( 
.A1(n_1346),
.A2(n_996),
.B(n_915),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1279),
.B(n_1087),
.Y(n_1398)
);

BUFx6f_ASAP7_75t_L g1399 ( 
.A(n_1355),
.Y(n_1399)
);

INVx3_ASAP7_75t_L g1400 ( 
.A(n_1292),
.Y(n_1400)
);

NOR2x1_ASAP7_75t_L g1401 ( 
.A(n_1289),
.B(n_1291),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1296),
.B(n_1043),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1299),
.B(n_1133),
.Y(n_1403)
);

OAI22x1_ASAP7_75t_SL g1404 ( 
.A1(n_1295),
.A2(n_1088),
.B1(n_1123),
.B2(n_1080),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1359),
.Y(n_1405)
);

AND2x6_ASAP7_75t_L g1406 ( 
.A(n_1307),
.B(n_1052),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_SL g1407 ( 
.A1(n_1304),
.A2(n_1156),
.B1(n_1172),
.B2(n_1127),
.Y(n_1407)
);

BUFx6f_ASAP7_75t_L g1408 ( 
.A(n_1310),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1301),
.B(n_1133),
.Y(n_1409)
);

INVx6_ASAP7_75t_L g1410 ( 
.A(n_1331),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1349),
.B(n_1028),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1312),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1360),
.Y(n_1413)
);

INVx3_ASAP7_75t_L g1414 ( 
.A(n_1313),
.Y(n_1414)
);

INVx4_ASAP7_75t_L g1415 ( 
.A(n_1308),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1363),
.Y(n_1416)
);

INVx3_ASAP7_75t_L g1417 ( 
.A(n_1314),
.Y(n_1417)
);

CKINVDCx20_ASAP7_75t_R g1418 ( 
.A(n_1305),
.Y(n_1418)
);

BUFx6f_ASAP7_75t_L g1419 ( 
.A(n_1316),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1317),
.B(n_1318),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1328),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1329),
.Y(n_1422)
);

OA21x2_ASAP7_75t_L g1423 ( 
.A1(n_1330),
.A2(n_1106),
.B(n_1078),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1332),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1324),
.B(n_1061),
.Y(n_1425)
);

CKINVDCx11_ASAP7_75t_R g1426 ( 
.A(n_1321),
.Y(n_1426)
);

BUFx6f_ASAP7_75t_L g1427 ( 
.A(n_1333),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1334),
.B(n_1145),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1338),
.Y(n_1429)
);

AOI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1322),
.A2(n_936),
.B1(n_943),
.B2(n_942),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1339),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1327),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1341),
.Y(n_1433)
);

INVxp33_ASAP7_75t_SL g1434 ( 
.A(n_1311),
.Y(n_1434)
);

AND2x4_ASAP7_75t_L g1435 ( 
.A(n_1319),
.B(n_1061),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1343),
.B(n_1102),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1344),
.Y(n_1437)
);

CKINVDCx11_ASAP7_75t_R g1438 ( 
.A(n_1335),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1345),
.B(n_1100),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1350),
.B(n_1145),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1351),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1353),
.A2(n_953),
.B1(n_954),
.B2(n_944),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1354),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_1337),
.Y(n_1444)
);

INVx3_ASAP7_75t_L g1445 ( 
.A(n_1356),
.Y(n_1445)
);

AOI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1357),
.A2(n_959),
.B1(n_963),
.B2(n_961),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1348),
.Y(n_1447)
);

OA21x2_ASAP7_75t_L g1448 ( 
.A1(n_1302),
.A2(n_1140),
.B(n_1114),
.Y(n_1448)
);

AOI22xp5_ASAP7_75t_SL g1449 ( 
.A1(n_1362),
.A2(n_1219),
.B1(n_1234),
.B2(n_1190),
.Y(n_1449)
);

BUFx2_ASAP7_75t_L g1450 ( 
.A(n_1359),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1281),
.Y(n_1451)
);

INVx3_ASAP7_75t_L g1452 ( 
.A(n_1358),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1293),
.Y(n_1453)
);

BUFx3_ASAP7_75t_L g1454 ( 
.A(n_1358),
.Y(n_1454)
);

BUFx6f_ASAP7_75t_L g1455 ( 
.A(n_1352),
.Y(n_1455)
);

BUFx3_ASAP7_75t_L g1456 ( 
.A(n_1358),
.Y(n_1456)
);

AND2x2_ASAP7_75t_SL g1457 ( 
.A(n_1300),
.B(n_1095),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1293),
.B(n_964),
.Y(n_1458)
);

BUFx6f_ASAP7_75t_L g1459 ( 
.A(n_1352),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1280),
.Y(n_1460)
);

INVx3_ASAP7_75t_L g1461 ( 
.A(n_1358),
.Y(n_1461)
);

AOI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1283),
.A2(n_965),
.B1(n_967),
.B2(n_966),
.Y(n_1462)
);

OA21x2_ASAP7_75t_L g1463 ( 
.A1(n_1273),
.A2(n_1140),
.B(n_1114),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1293),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1280),
.B(n_1269),
.Y(n_1465)
);

INVxp67_ASAP7_75t_L g1466 ( 
.A(n_1361),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1288),
.A2(n_973),
.B1(n_982),
.B2(n_970),
.Y(n_1467)
);

AND2x6_ASAP7_75t_L g1468 ( 
.A(n_1358),
.B(n_1117),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1280),
.B(n_1269),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1293),
.B(n_983),
.Y(n_1470)
);

CKINVDCx6p67_ASAP7_75t_R g1471 ( 
.A(n_1300),
.Y(n_1471)
);

BUFx6f_ASAP7_75t_L g1472 ( 
.A(n_1352),
.Y(n_1472)
);

AOI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1283),
.A2(n_984),
.B1(n_995),
.B2(n_990),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1347),
.Y(n_1474)
);

AND2x6_ASAP7_75t_L g1475 ( 
.A(n_1358),
.B(n_1117),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1293),
.Y(n_1476)
);

INVx3_ASAP7_75t_L g1477 ( 
.A(n_1358),
.Y(n_1477)
);

OAI22x1_ASAP7_75t_R g1478 ( 
.A1(n_1290),
.A2(n_902),
.B1(n_933),
.B2(n_886),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1293),
.Y(n_1479)
);

CKINVDCx8_ASAP7_75t_R g1480 ( 
.A(n_1300),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1293),
.B(n_999),
.Y(n_1481)
);

BUFx12f_ASAP7_75t_L g1482 ( 
.A(n_1287),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1280),
.Y(n_1483)
);

OAI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1273),
.A2(n_1245),
.B(n_1193),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1281),
.Y(n_1485)
);

OAI22x1_ASAP7_75t_L g1486 ( 
.A1(n_1303),
.A2(n_1011),
.B1(n_1013),
.B2(n_1009),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1281),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_L g1488 ( 
.A(n_1274),
.B(n_1243),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1281),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1281),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1280),
.B(n_1241),
.Y(n_1491)
);

NOR2x1_ASAP7_75t_L g1492 ( 
.A(n_1358),
.B(n_1120),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1293),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1281),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1358),
.B(n_890),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1274),
.B(n_1017),
.Y(n_1496)
);

INVx6_ASAP7_75t_L g1497 ( 
.A(n_1281),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_SL g1498 ( 
.A(n_1358),
.B(n_894),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1293),
.Y(n_1499)
);

BUFx8_ASAP7_75t_SL g1500 ( 
.A(n_1290),
.Y(n_1500)
);

OAI21x1_ASAP7_75t_L g1501 ( 
.A1(n_1273),
.A2(n_1265),
.B(n_1247),
.Y(n_1501)
);

BUFx6f_ASAP7_75t_L g1502 ( 
.A(n_1352),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_R g1503 ( 
.A(n_1474),
.B(n_962),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1428),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1500),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_1426),
.Y(n_1506)
);

BUFx6f_ASAP7_75t_L g1507 ( 
.A(n_1423),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1460),
.B(n_1014),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_1438),
.Y(n_1509)
);

CKINVDCx20_ASAP7_75t_R g1510 ( 
.A(n_1483),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1491),
.B(n_1014),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1491),
.B(n_1105),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1411),
.Y(n_1513)
);

CKINVDCx20_ASAP7_75t_R g1514 ( 
.A(n_1418),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1428),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1411),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1440),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1471),
.Y(n_1518)
);

CKINVDCx20_ASAP7_75t_R g1519 ( 
.A(n_1444),
.Y(n_1519)
);

CKINVDCx20_ASAP7_75t_R g1520 ( 
.A(n_1405),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_1413),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_R g1522 ( 
.A(n_1416),
.B(n_980),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_1480),
.Y(n_1523)
);

CKINVDCx20_ASAP7_75t_R g1524 ( 
.A(n_1450),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_1482),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1380),
.A2(n_1265),
.B(n_1247),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_1434),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1447),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1484),
.Y(n_1529)
);

BUFx2_ASAP7_75t_L g1530 ( 
.A(n_1391),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_1404),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1432),
.Y(n_1532)
);

BUFx3_ASAP7_75t_L g1533 ( 
.A(n_1497),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_1410),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1466),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1465),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1414),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1501),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1417),
.Y(n_1539)
);

CKINVDCx20_ASAP7_75t_R g1540 ( 
.A(n_1478),
.Y(n_1540)
);

BUFx2_ASAP7_75t_L g1541 ( 
.A(n_1469),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1397),
.Y(n_1542)
);

CKINVDCx20_ASAP7_75t_R g1543 ( 
.A(n_1449),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_1407),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_R g1545 ( 
.A(n_1457),
.B(n_1025),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1445),
.Y(n_1546)
);

BUFx8_ASAP7_75t_L g1547 ( 
.A(n_1395),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1463),
.Y(n_1548)
);

INVx8_ASAP7_75t_L g1549 ( 
.A(n_1368),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1467),
.Y(n_1550)
);

BUFx3_ASAP7_75t_L g1551 ( 
.A(n_1375),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_1372),
.Y(n_1552)
);

BUFx6f_ASAP7_75t_SL g1553 ( 
.A(n_1425),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1384),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1392),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_1462),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_1473),
.Y(n_1557)
);

INVx3_ASAP7_75t_L g1558 ( 
.A(n_1408),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1394),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1430),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_1442),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_1415),
.Y(n_1562)
);

CKINVDCx20_ASAP7_75t_R g1563 ( 
.A(n_1446),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1452),
.B(n_1030),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1486),
.Y(n_1565)
);

BUFx6f_ASAP7_75t_L g1566 ( 
.A(n_1406),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_1454),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_1456),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_1468),
.Y(n_1569)
);

BUFx2_ASAP7_75t_L g1570 ( 
.A(n_1468),
.Y(n_1570)
);

BUFx6f_ASAP7_75t_L g1571 ( 
.A(n_1406),
.Y(n_1571)
);

CKINVDCx20_ASAP7_75t_R g1572 ( 
.A(n_1376),
.Y(n_1572)
);

INVxp67_ASAP7_75t_SL g1573 ( 
.A(n_1420),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_R g1574 ( 
.A(n_1475),
.B(n_1042),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_1475),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1419),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1461),
.B(n_1031),
.Y(n_1577)
);

AOI21x1_ASAP7_75t_L g1578 ( 
.A1(n_1498),
.A2(n_1131),
.B(n_1126),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_1377),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1385),
.B(n_1032),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1422),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1422),
.Y(n_1582)
);

AOI21x1_ASAP7_75t_L g1583 ( 
.A1(n_1378),
.A2(n_1389),
.B(n_1382),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1495),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_1458),
.Y(n_1585)
);

BUFx2_ASAP7_75t_L g1586 ( 
.A(n_1406),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1470),
.Y(n_1587)
);

INVxp67_ASAP7_75t_SL g1588 ( 
.A(n_1427),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1481),
.B(n_894),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_1387),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_1388),
.Y(n_1591)
);

BUFx10_ASAP7_75t_L g1592 ( 
.A(n_1496),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1402),
.Y(n_1593)
);

BUFx3_ASAP7_75t_L g1594 ( 
.A(n_1448),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_1403),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1441),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_1409),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_1386),
.Y(n_1598)
);

CKINVDCx20_ASAP7_75t_R g1599 ( 
.A(n_1364),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_1477),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1365),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1366),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_1393),
.Y(n_1603)
);

BUFx2_ASAP7_75t_L g1604 ( 
.A(n_1436),
.Y(n_1604)
);

INVxp67_ASAP7_75t_L g1605 ( 
.A(n_1439),
.Y(n_1605)
);

INVx2_ASAP7_75t_SL g1606 ( 
.A(n_1435),
.Y(n_1606)
);

CKINVDCx20_ASAP7_75t_R g1607 ( 
.A(n_1367),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1374),
.Y(n_1608)
);

INVx3_ASAP7_75t_L g1609 ( 
.A(n_1451),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_1369),
.Y(n_1610)
);

AND2x6_ASAP7_75t_L g1611 ( 
.A(n_1492),
.B(n_881),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_1371),
.Y(n_1612)
);

CKINVDCx16_ASAP7_75t_R g1613 ( 
.A(n_1401),
.Y(n_1613)
);

AND2x4_ASAP7_75t_L g1614 ( 
.A(n_1453),
.B(n_1144),
.Y(n_1614)
);

CKINVDCx6p67_ASAP7_75t_R g1615 ( 
.A(n_1464),
.Y(n_1615)
);

INVx4_ASAP7_75t_L g1616 ( 
.A(n_1383),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_1476),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_1479),
.Y(n_1618)
);

CKINVDCx20_ASAP7_75t_R g1619 ( 
.A(n_1493),
.Y(n_1619)
);

BUFx6f_ASAP7_75t_L g1620 ( 
.A(n_1383),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_1499),
.Y(n_1621)
);

NOR2xp67_ASAP7_75t_L g1622 ( 
.A(n_1398),
.B(n_0),
.Y(n_1622)
);

CKINVDCx20_ASAP7_75t_R g1623 ( 
.A(n_1412),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_1488),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1424),
.B(n_1037),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_1485),
.Y(n_1626)
);

BUFx2_ASAP7_75t_L g1627 ( 
.A(n_1431),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_1487),
.Y(n_1628)
);

BUFx6f_ASAP7_75t_L g1629 ( 
.A(n_1396),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_1489),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1490),
.Y(n_1631)
);

CKINVDCx20_ASAP7_75t_R g1632 ( 
.A(n_1421),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_1494),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1429),
.B(n_889),
.Y(n_1634)
);

CKINVDCx20_ASAP7_75t_R g1635 ( 
.A(n_1433),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_1437),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1396),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_R g1638 ( 
.A(n_1443),
.B(n_1112),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_1399),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1390),
.Y(n_1640)
);

CKINVDCx20_ASAP7_75t_R g1641 ( 
.A(n_1370),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_1370),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_1373),
.Y(n_1643)
);

NOR2x1p5_ASAP7_75t_L g1644 ( 
.A(n_1379),
.B(n_1038),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1502),
.Y(n_1645)
);

BUFx3_ASAP7_75t_L g1646 ( 
.A(n_1455),
.Y(n_1646)
);

INVx4_ASAP7_75t_L g1647 ( 
.A(n_1459),
.Y(n_1647)
);

CKINVDCx20_ASAP7_75t_R g1648 ( 
.A(n_1472),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_1472),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1381),
.B(n_894),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_1500),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_1500),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_1500),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_1500),
.Y(n_1654)
);

BUFx2_ASAP7_75t_L g1655 ( 
.A(n_1460),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1460),
.B(n_1041),
.Y(n_1656)
);

CKINVDCx16_ASAP7_75t_R g1657 ( 
.A(n_1460),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_1500),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1428),
.B(n_1046),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_R g1660 ( 
.A(n_1474),
.B(n_1220),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_1500),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_1500),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_1500),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_1500),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1428),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_1500),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_R g1667 ( 
.A(n_1474),
.B(n_1222),
.Y(n_1667)
);

AND3x1_ASAP7_75t_L g1668 ( 
.A(n_1372),
.B(n_901),
.C(n_899),
.Y(n_1668)
);

NAND2xp33_ASAP7_75t_R g1669 ( 
.A(n_1434),
.B(n_1056),
.Y(n_1669)
);

CKINVDCx20_ASAP7_75t_R g1670 ( 
.A(n_1460),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_1500),
.Y(n_1671)
);

INVx3_ASAP7_75t_L g1672 ( 
.A(n_1400),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_R g1673 ( 
.A(n_1474),
.B(n_1251),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1380),
.Y(n_1674)
);

BUFx6f_ASAP7_75t_L g1675 ( 
.A(n_1423),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_1500),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1573),
.Y(n_1677)
);

BUFx6f_ASAP7_75t_L g1678 ( 
.A(n_1566),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1627),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1504),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1515),
.A2(n_987),
.B1(n_1047),
.B2(n_894),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1530),
.B(n_1057),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1535),
.B(n_1264),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1517),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_SL g1685 ( 
.A(n_1566),
.B(n_1058),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1583),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1536),
.B(n_1060),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1513),
.B(n_1062),
.Y(n_1688)
);

INVx4_ASAP7_75t_L g1689 ( 
.A(n_1562),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_SL g1690 ( 
.A(n_1566),
.B(n_1063),
.Y(n_1690)
);

INVx1_ASAP7_75t_SL g1691 ( 
.A(n_1510),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1507),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1516),
.B(n_1067),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1590),
.B(n_1069),
.Y(n_1694)
);

INVx3_ASAP7_75t_L g1695 ( 
.A(n_1657),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1675),
.Y(n_1696)
);

BUFx6f_ASAP7_75t_L g1697 ( 
.A(n_1571),
.Y(n_1697)
);

BUFx6f_ASAP7_75t_L g1698 ( 
.A(n_1571),
.Y(n_1698)
);

NOR2x1p5_ASAP7_75t_L g1699 ( 
.A(n_1527),
.B(n_1070),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_SL g1700 ( 
.A(n_1571),
.B(n_1072),
.Y(n_1700)
);

INVxp33_ASAP7_75t_L g1701 ( 
.A(n_1638),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1670),
.Y(n_1702)
);

CKINVDCx20_ASAP7_75t_R g1703 ( 
.A(n_1520),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1665),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1675),
.Y(n_1705)
);

INVx1_ASAP7_75t_SL g1706 ( 
.A(n_1524),
.Y(n_1706)
);

INVx3_ASAP7_75t_L g1707 ( 
.A(n_1551),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1542),
.Y(n_1708)
);

BUFx6f_ASAP7_75t_L g1709 ( 
.A(n_1620),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1548),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1555),
.Y(n_1711)
);

INVxp67_ASAP7_75t_SL g1712 ( 
.A(n_1623),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1526),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1656),
.B(n_1075),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1580),
.A2(n_1165),
.B1(n_1047),
.B2(n_1077),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_1620),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1541),
.B(n_1076),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1591),
.B(n_1079),
.Y(n_1718)
);

BUFx6f_ASAP7_75t_L g1719 ( 
.A(n_1620),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1559),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1625),
.B(n_1085),
.Y(n_1721)
);

BUFx3_ASAP7_75t_L g1722 ( 
.A(n_1641),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1608),
.Y(n_1723)
);

BUFx6f_ASAP7_75t_L g1724 ( 
.A(n_1629),
.Y(n_1724)
);

AND2x2_ASAP7_75t_SL g1725 ( 
.A(n_1668),
.B(n_1141),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1532),
.B(n_1074),
.Y(n_1726)
);

AO22x2_ASAP7_75t_L g1727 ( 
.A1(n_1634),
.A2(n_1071),
.B1(n_1090),
.B2(n_1082),
.Y(n_1727)
);

AND2x4_ASAP7_75t_L g1728 ( 
.A(n_1634),
.B(n_910),
.Y(n_1728)
);

NAND3x1_ASAP7_75t_L g1729 ( 
.A(n_1540),
.B(n_927),
.C(n_924),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1511),
.B(n_1092),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1585),
.B(n_1587),
.Y(n_1731)
);

AND2x6_ASAP7_75t_L g1732 ( 
.A(n_1594),
.B(n_881),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1512),
.B(n_1098),
.Y(n_1733)
);

BUFx2_ASAP7_75t_L g1734 ( 
.A(n_1632),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1603),
.B(n_1103),
.Y(n_1735)
);

INVx4_ASAP7_75t_L g1736 ( 
.A(n_1579),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1601),
.Y(n_1737)
);

BUFx6f_ASAP7_75t_L g1738 ( 
.A(n_1629),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_L g1739 ( 
.A(n_1624),
.B(n_1119),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1631),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_SL g1741 ( 
.A(n_1521),
.B(n_1121),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1636),
.B(n_1508),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1614),
.B(n_1122),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1602),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1614),
.B(n_1124),
.Y(n_1745)
);

INVx6_ASAP7_75t_L g1746 ( 
.A(n_1547),
.Y(n_1746)
);

INVx4_ASAP7_75t_L g1747 ( 
.A(n_1534),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1529),
.Y(n_1748)
);

BUFx3_ASAP7_75t_L g1749 ( 
.A(n_1648),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1537),
.Y(n_1750)
);

BUFx6f_ASAP7_75t_L g1751 ( 
.A(n_1629),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_1506),
.Y(n_1752)
);

INVx2_ASAP7_75t_SL g1753 ( 
.A(n_1547),
.Y(n_1753)
);

INVx2_ASAP7_75t_SL g1754 ( 
.A(n_1644),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_SL g1755 ( 
.A(n_1570),
.B(n_1125),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1539),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1538),
.Y(n_1757)
);

BUFx3_ASAP7_75t_L g1758 ( 
.A(n_1509),
.Y(n_1758)
);

BUFx6f_ASAP7_75t_L g1759 ( 
.A(n_1549),
.Y(n_1759)
);

INVx2_ASAP7_75t_SL g1760 ( 
.A(n_1615),
.Y(n_1760)
);

AND2x4_ASAP7_75t_L g1761 ( 
.A(n_1518),
.B(n_1258),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1659),
.B(n_1128),
.Y(n_1762)
);

AND2x6_ASAP7_75t_L g1763 ( 
.A(n_1549),
.B(n_881),
.Y(n_1763)
);

CKINVDCx20_ASAP7_75t_R g1764 ( 
.A(n_1519),
.Y(n_1764)
);

INVxp67_ASAP7_75t_L g1765 ( 
.A(n_1669),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1605),
.B(n_1134),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1635),
.B(n_1135),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1546),
.Y(n_1768)
);

BUFx6f_ASAP7_75t_L g1769 ( 
.A(n_1549),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1584),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1640),
.Y(n_1771)
);

CKINVDCx5p33_ASAP7_75t_R g1772 ( 
.A(n_1505),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_SL g1773 ( 
.A(n_1586),
.B(n_1598),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1613),
.B(n_1139),
.Y(n_1774)
);

INVx3_ASAP7_75t_L g1775 ( 
.A(n_1672),
.Y(n_1775)
);

BUFx2_ASAP7_75t_L g1776 ( 
.A(n_1503),
.Y(n_1776)
);

BUFx6f_ASAP7_75t_L g1777 ( 
.A(n_1642),
.Y(n_1777)
);

CKINVDCx20_ASAP7_75t_R g1778 ( 
.A(n_1514),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1660),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1674),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1564),
.B(n_1146),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_SL g1782 ( 
.A(n_1569),
.B(n_1147),
.Y(n_1782)
);

A2O1A1Ixp33_ASAP7_75t_L g1783 ( 
.A1(n_1589),
.A2(n_1622),
.B(n_1650),
.C(n_1577),
.Y(n_1783)
);

INVx1_ASAP7_75t_SL g1784 ( 
.A(n_1667),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1528),
.B(n_1552),
.Y(n_1785)
);

INVx1_ASAP7_75t_SL g1786 ( 
.A(n_1673),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1609),
.Y(n_1787)
);

BUFx3_ASAP7_75t_L g1788 ( 
.A(n_1525),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1610),
.B(n_1150),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1612),
.B(n_1152),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1578),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1609),
.Y(n_1792)
);

INVx6_ASAP7_75t_L g1793 ( 
.A(n_1592),
.Y(n_1793)
);

INVx1_ASAP7_75t_SL g1794 ( 
.A(n_1522),
.Y(n_1794)
);

AND2x4_ASAP7_75t_L g1795 ( 
.A(n_1606),
.B(n_929),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1617),
.B(n_1155),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1618),
.B(n_1159),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1604),
.Y(n_1798)
);

BUFx10_ASAP7_75t_L g1799 ( 
.A(n_1651),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_L g1800 ( 
.A(n_1572),
.B(n_1164),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1558),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_L g1802 ( 
.A(n_1550),
.B(n_1166),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1575),
.B(n_1167),
.Y(n_1803)
);

AND2x4_ASAP7_75t_L g1804 ( 
.A(n_1621),
.B(n_938),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1611),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1611),
.Y(n_1806)
);

INVx3_ASAP7_75t_L g1807 ( 
.A(n_1553),
.Y(n_1807)
);

NOR2xp33_ASAP7_75t_L g1808 ( 
.A(n_1599),
.B(n_1171),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1607),
.B(n_1173),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1554),
.B(n_1154),
.Y(n_1810)
);

INVx2_ASAP7_75t_SL g1811 ( 
.A(n_1574),
.Y(n_1811)
);

INVx2_ASAP7_75t_SL g1812 ( 
.A(n_1567),
.Y(n_1812)
);

BUFx6f_ASAP7_75t_L g1813 ( 
.A(n_1643),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1611),
.Y(n_1814)
);

INVx4_ASAP7_75t_L g1815 ( 
.A(n_1639),
.Y(n_1815)
);

NOR2xp33_ASAP7_75t_L g1816 ( 
.A(n_1619),
.B(n_1177),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1561),
.A2(n_1165),
.B1(n_1047),
.B2(n_1178),
.Y(n_1817)
);

BUFx6f_ASAP7_75t_L g1818 ( 
.A(n_1649),
.Y(n_1818)
);

AND2x4_ASAP7_75t_L g1819 ( 
.A(n_1568),
.B(n_945),
.Y(n_1819)
);

INVx3_ASAP7_75t_L g1820 ( 
.A(n_1553),
.Y(n_1820)
);

AND2x4_ASAP7_75t_L g1821 ( 
.A(n_1626),
.B(n_1628),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1630),
.B(n_1183),
.Y(n_1822)
);

AO22x2_ASAP7_75t_L g1823 ( 
.A1(n_1543),
.A2(n_1266),
.B1(n_1270),
.B2(n_1217),
.Y(n_1823)
);

NOR2xp33_ASAP7_75t_L g1824 ( 
.A(n_1556),
.B(n_1185),
.Y(n_1824)
);

BUFx3_ASAP7_75t_L g1825 ( 
.A(n_1652),
.Y(n_1825)
);

BUFx10_ASAP7_75t_L g1826 ( 
.A(n_1653),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1633),
.Y(n_1827)
);

BUFx3_ASAP7_75t_L g1828 ( 
.A(n_1654),
.Y(n_1828)
);

AND2x6_ASAP7_75t_L g1829 ( 
.A(n_1596),
.B(n_881),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1576),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1557),
.B(n_1187),
.Y(n_1831)
);

INVx8_ASAP7_75t_L g1832 ( 
.A(n_1523),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1588),
.Y(n_1833)
);

AND2x4_ASAP7_75t_L g1834 ( 
.A(n_1600),
.B(n_947),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1581),
.Y(n_1835)
);

BUFx6f_ASAP7_75t_L g1836 ( 
.A(n_1616),
.Y(n_1836)
);

BUFx4_ASAP7_75t_L g1837 ( 
.A(n_1658),
.Y(n_1837)
);

INVx4_ASAP7_75t_L g1838 ( 
.A(n_1661),
.Y(n_1838)
);

AOI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1560),
.A2(n_1165),
.B1(n_1047),
.B2(n_1201),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1582),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_SL g1841 ( 
.A(n_1616),
.B(n_1204),
.Y(n_1841)
);

INVx5_ASAP7_75t_L g1842 ( 
.A(n_1647),
.Y(n_1842)
);

INVxp67_ASAP7_75t_SL g1843 ( 
.A(n_1563),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1637),
.Y(n_1844)
);

BUFx6f_ASAP7_75t_L g1845 ( 
.A(n_1646),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1565),
.Y(n_1846)
);

BUFx4f_ASAP7_75t_L g1847 ( 
.A(n_1662),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1593),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_L g1849 ( 
.A1(n_1595),
.A2(n_1165),
.B1(n_1211),
.B2(n_1208),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_SL g1850 ( 
.A(n_1597),
.B(n_1213),
.Y(n_1850)
);

AND2x2_ASAP7_75t_SL g1851 ( 
.A(n_1545),
.B(n_1151),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1544),
.B(n_1216),
.Y(n_1852)
);

BUFx2_ASAP7_75t_L g1853 ( 
.A(n_1663),
.Y(n_1853)
);

INVxp33_ASAP7_75t_L g1854 ( 
.A(n_1664),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1645),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1531),
.Y(n_1856)
);

BUFx6f_ASAP7_75t_L g1857 ( 
.A(n_1666),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1676),
.Y(n_1858)
);

AND2x6_ASAP7_75t_L g1859 ( 
.A(n_1671),
.B(n_891),
.Y(n_1859)
);

NOR2xp33_ASAP7_75t_L g1860 ( 
.A(n_1530),
.B(n_1218),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1583),
.Y(n_1861)
);

HB1xp67_ASAP7_75t_L g1862 ( 
.A(n_1655),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_L g1863 ( 
.A(n_1530),
.B(n_1225),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1573),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1573),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1583),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_SL g1867 ( 
.A(n_1566),
.B(n_1232),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1573),
.B(n_1268),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1573),
.Y(n_1869)
);

AOI22xp33_ASAP7_75t_L g1870 ( 
.A1(n_1504),
.A2(n_1236),
.B1(n_1238),
.B2(n_1235),
.Y(n_1870)
);

AND2x4_ASAP7_75t_L g1871 ( 
.A(n_1655),
.B(n_955),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1530),
.B(n_1239),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1530),
.B(n_1246),
.Y(n_1873)
);

BUFx3_ASAP7_75t_L g1874 ( 
.A(n_1641),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1573),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_SL g1876 ( 
.A(n_1566),
.B(n_1252),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1573),
.Y(n_1877)
);

BUFx3_ASAP7_75t_L g1878 ( 
.A(n_1641),
.Y(n_1878)
);

AOI22xp33_ASAP7_75t_L g1879 ( 
.A1(n_1504),
.A2(n_1253),
.B1(n_1255),
.B2(n_1250),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_SL g1880 ( 
.A(n_1566),
.B(n_1261),
.Y(n_1880)
);

BUFx6f_ASAP7_75t_L g1881 ( 
.A(n_1566),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1530),
.B(n_1256),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1530),
.B(n_1257),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1530),
.B(n_1260),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1573),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1573),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1573),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1583),
.Y(n_1888)
);

INVx1_ASAP7_75t_SL g1889 ( 
.A(n_1510),
.Y(n_1889)
);

AND2x6_ASAP7_75t_L g1890 ( 
.A(n_1566),
.B(n_891),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1573),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1573),
.Y(n_1892)
);

BUFx3_ASAP7_75t_L g1893 ( 
.A(n_1641),
.Y(n_1893)
);

BUFx6f_ASAP7_75t_L g1894 ( 
.A(n_1566),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1573),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1530),
.B(n_885),
.Y(n_1896)
);

BUFx6f_ASAP7_75t_L g1897 ( 
.A(n_1566),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1573),
.Y(n_1898)
);

INVx3_ASAP7_75t_L g1899 ( 
.A(n_1533),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1573),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_SL g1901 ( 
.A(n_1566),
.B(n_887),
.Y(n_1901)
);

HB1xp67_ASAP7_75t_L g1902 ( 
.A(n_1862),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1677),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1864),
.B(n_1153),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1865),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1869),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1875),
.Y(n_1907)
);

AO22x2_ASAP7_75t_L g1908 ( 
.A1(n_1712),
.A2(n_1163),
.B1(n_1168),
.B2(n_1158),
.Y(n_1908)
);

AND2x4_ASAP7_75t_L g1909 ( 
.A(n_1877),
.B(n_985),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1885),
.B(n_1169),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1886),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1887),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1891),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1892),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1895),
.Y(n_1915)
);

BUFx3_ASAP7_75t_L g1916 ( 
.A(n_1703),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1898),
.Y(n_1917)
);

INVx5_ASAP7_75t_L g1918 ( 
.A(n_1763),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1900),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1711),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1720),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1708),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1710),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1872),
.B(n_1873),
.Y(n_1924)
);

INVx3_ASAP7_75t_L g1925 ( 
.A(n_1746),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1868),
.B(n_1184),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1737),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1882),
.B(n_903),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1741),
.B(n_909),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1744),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1883),
.B(n_919),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1680),
.Y(n_1932)
);

AO22x2_ASAP7_75t_L g1933 ( 
.A1(n_1727),
.A2(n_1192),
.B1(n_1194),
.B2(n_1191),
.Y(n_1933)
);

AO22x2_ASAP7_75t_L g1934 ( 
.A1(n_1706),
.A2(n_1196),
.B1(n_1202),
.B2(n_1195),
.Y(n_1934)
);

AO22x2_ASAP7_75t_L g1935 ( 
.A1(n_1889),
.A2(n_1209),
.B1(n_1212),
.B2(n_1207),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1684),
.Y(n_1936)
);

AND2x4_ASAP7_75t_L g1937 ( 
.A(n_1760),
.B(n_989),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1884),
.B(n_932),
.Y(n_1938)
);

NAND2x1p5_ASAP7_75t_L g1939 ( 
.A(n_1777),
.B(n_891),
.Y(n_1939)
);

NAND3xp33_ASAP7_75t_L g1940 ( 
.A(n_1783),
.B(n_893),
.C(n_891),
.Y(n_1940)
);

BUFx8_ASAP7_75t_L g1941 ( 
.A(n_1857),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1704),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1714),
.B(n_1221),
.Y(n_1943)
);

AND2x6_ASAP7_75t_SL g1944 ( 
.A(n_1856),
.B(n_991),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1679),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1748),
.Y(n_1946)
);

BUFx6f_ASAP7_75t_L g1947 ( 
.A(n_1813),
.Y(n_1947)
);

NOR2xp33_ASAP7_75t_L g1948 ( 
.A(n_1810),
.B(n_1802),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_L g1949 ( 
.A(n_1683),
.B(n_941),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1767),
.B(n_950),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1730),
.B(n_1227),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1757),
.Y(n_1952)
);

AOI22xp33_ASAP7_75t_L g1953 ( 
.A1(n_1831),
.A2(n_975),
.B1(n_976),
.B2(n_956),
.Y(n_1953)
);

AO22x2_ASAP7_75t_L g1954 ( 
.A1(n_1846),
.A2(n_1237),
.B1(n_1240),
.B2(n_1233),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_SL g1955 ( 
.A(n_1821),
.B(n_979),
.Y(n_1955)
);

NOR2xp33_ASAP7_75t_L g1956 ( 
.A(n_1742),
.B(n_1824),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1733),
.B(n_1249),
.Y(n_1957)
);

AO22x2_ASAP7_75t_L g1958 ( 
.A1(n_1794),
.A2(n_1259),
.B1(n_1262),
.B2(n_1254),
.Y(n_1958)
);

BUFx3_ASAP7_75t_L g1959 ( 
.A(n_1722),
.Y(n_1959)
);

OR2x6_ASAP7_75t_L g1960 ( 
.A(n_1832),
.B(n_1753),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1780),
.Y(n_1961)
);

NAND2xp33_ASAP7_75t_L g1962 ( 
.A(n_1732),
.B(n_1012),
.Y(n_1962)
);

NOR2xp33_ASAP7_75t_L g1963 ( 
.A(n_1785),
.B(n_994),
.Y(n_1963)
);

NAND2x1p5_ASAP7_75t_L g1964 ( 
.A(n_1818),
.B(n_893),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1694),
.B(n_1718),
.Y(n_1965)
);

AOI22xp33_ASAP7_75t_L g1966 ( 
.A1(n_1725),
.A2(n_1018),
.B1(n_1020),
.B2(n_1008),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1682),
.B(n_1022),
.Y(n_1967)
);

AND2x6_ASAP7_75t_L g1968 ( 
.A(n_1759),
.B(n_893),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1771),
.Y(n_1969)
);

NAND3xp33_ASAP7_75t_L g1970 ( 
.A(n_1739),
.B(n_940),
.C(n_934),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1860),
.B(n_1024),
.Y(n_1971)
);

AND2x4_ASAP7_75t_L g1972 ( 
.A(n_1736),
.B(n_997),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1863),
.B(n_1036),
.Y(n_1973)
);

OAI22xp5_ASAP7_75t_L g1974 ( 
.A1(n_1715),
.A2(n_1055),
.B1(n_1059),
.B2(n_1053),
.Y(n_1974)
);

AO22x2_ASAP7_75t_L g1975 ( 
.A1(n_1726),
.A2(n_1004),
.B1(n_1005),
.B2(n_1002),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1770),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1750),
.Y(n_1977)
);

BUFx6f_ASAP7_75t_L g1978 ( 
.A(n_1709),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1756),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1717),
.B(n_1896),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1768),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1728),
.Y(n_1982)
);

NAND3x1_ASAP7_75t_L g1983 ( 
.A(n_1837),
.B(n_1248),
.C(n_1244),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1728),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1723),
.Y(n_1985)
);

NAND2x1p5_ASAP7_75t_L g1986 ( 
.A(n_1747),
.B(n_934),
.Y(n_1986)
);

AO22x2_ASAP7_75t_L g1987 ( 
.A1(n_1784),
.A2(n_1027),
.B1(n_1029),
.B2(n_1021),
.Y(n_1987)
);

BUFx2_ASAP7_75t_L g1988 ( 
.A(n_1749),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1740),
.Y(n_1989)
);

BUFx3_ASAP7_75t_L g1990 ( 
.A(n_1874),
.Y(n_1990)
);

AND2x4_ASAP7_75t_L g1991 ( 
.A(n_1878),
.B(n_1033),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1721),
.B(n_1086),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1795),
.Y(n_1993)
);

BUFx6f_ASAP7_75t_L g1994 ( 
.A(n_1709),
.Y(n_1994)
);

NOR2xp33_ASAP7_75t_L g1995 ( 
.A(n_1702),
.B(n_1091),
.Y(n_1995)
);

INVx3_ASAP7_75t_L g1996 ( 
.A(n_1893),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1743),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1745),
.Y(n_1998)
);

AND2x4_ASAP7_75t_L g1999 ( 
.A(n_1788),
.B(n_1089),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1787),
.Y(n_2000)
);

AO22x2_ASAP7_75t_L g2001 ( 
.A1(n_1786),
.A2(n_1097),
.B1(n_1099),
.B2(n_1093),
.Y(n_2001)
);

NAND2x1p5_ASAP7_75t_L g2002 ( 
.A(n_1815),
.B(n_940),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1798),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1686),
.Y(n_2004)
);

AO22x2_ASAP7_75t_L g2005 ( 
.A1(n_1843),
.A2(n_1104),
.B1(n_1108),
.B2(n_1101),
.Y(n_2005)
);

NAND2xp33_ASAP7_75t_L g2006 ( 
.A(n_1732),
.B(n_1763),
.Y(n_2006)
);

INVx2_ASAP7_75t_SL g2007 ( 
.A(n_1793),
.Y(n_2007)
);

AOI22xp5_ASAP7_75t_L g2008 ( 
.A1(n_1800),
.A2(n_1808),
.B1(n_1816),
.B2(n_1809),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1861),
.Y(n_2009)
);

NOR2xp33_ASAP7_75t_L g2010 ( 
.A(n_1734),
.B(n_1107),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1792),
.Y(n_2011)
);

CKINVDCx20_ASAP7_75t_R g2012 ( 
.A(n_1764),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1866),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1766),
.B(n_1110),
.Y(n_2014)
);

AO22x2_ASAP7_75t_L g2015 ( 
.A1(n_1823),
.A2(n_1111),
.B1(n_1113),
.B2(n_1109),
.Y(n_2015)
);

NAND2x1p5_ASAP7_75t_L g2016 ( 
.A(n_1695),
.B(n_969),
.Y(n_2016)
);

AND2x6_ASAP7_75t_L g2017 ( 
.A(n_1759),
.B(n_1769),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1841),
.Y(n_2018)
);

INVx6_ASAP7_75t_L g2019 ( 
.A(n_1799),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1687),
.B(n_1115),
.Y(n_2020)
);

NAND2x1p5_ASAP7_75t_L g2021 ( 
.A(n_1842),
.B(n_969),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1888),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1833),
.Y(n_2023)
);

AND2x4_ASAP7_75t_L g2024 ( 
.A(n_1773),
.B(n_1116),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1688),
.B(n_1693),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_1851),
.B(n_1118),
.Y(n_2026)
);

BUFx6f_ASAP7_75t_L g2027 ( 
.A(n_1716),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1830),
.Y(n_2028)
);

AND2x6_ASAP7_75t_L g2029 ( 
.A(n_1769),
.B(n_1035),
.Y(n_2029)
);

NAND2x1p5_ASAP7_75t_L g2030 ( 
.A(n_1842),
.B(n_1035),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1839),
.B(n_1130),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1835),
.Y(n_2032)
);

AND2x4_ASAP7_75t_L g2033 ( 
.A(n_1775),
.B(n_1129),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1681),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1836),
.Y(n_2035)
);

AO22x2_ASAP7_75t_L g2036 ( 
.A1(n_1823),
.A2(n_1136),
.B1(n_1137),
.B2(n_1132),
.Y(n_2036)
);

NAND2x1p5_ASAP7_75t_L g2037 ( 
.A(n_1776),
.B(n_1035),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1836),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1871),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1840),
.Y(n_2040)
);

INVx3_ASAP7_75t_L g2041 ( 
.A(n_1793),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1827),
.Y(n_2042)
);

INVx5_ASAP7_75t_L g2043 ( 
.A(n_1763),
.Y(n_2043)
);

BUFx6f_ASAP7_75t_L g2044 ( 
.A(n_1716),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1804),
.Y(n_2045)
);

AO22x2_ASAP7_75t_L g2046 ( 
.A1(n_1811),
.A2(n_1834),
.B1(n_1765),
.B2(n_1754),
.Y(n_2046)
);

AND2x6_ASAP7_75t_L g2047 ( 
.A(n_1678),
.B(n_1049),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1685),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1690),
.Y(n_2049)
);

INVx2_ASAP7_75t_SL g2050 ( 
.A(n_1832),
.Y(n_2050)
);

NAND3x1_ASAP7_75t_L g2051 ( 
.A(n_1837),
.B(n_1161),
.C(n_1160),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1700),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1867),
.Y(n_2053)
);

CKINVDCx20_ASAP7_75t_R g2054 ( 
.A(n_1778),
.Y(n_2054)
);

BUFx6f_ASAP7_75t_L g2055 ( 
.A(n_1719),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1781),
.B(n_1162),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1876),
.Y(n_2057)
);

AND2x4_ASAP7_75t_L g2058 ( 
.A(n_1812),
.B(n_1170),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1880),
.Y(n_2059)
);

NOR2xp33_ASAP7_75t_L g2060 ( 
.A(n_1735),
.B(n_1701),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_1870),
.B(n_1879),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1789),
.B(n_1174),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1790),
.B(n_1176),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1762),
.Y(n_2064)
);

NOR2xp33_ASAP7_75t_L g2065 ( 
.A(n_1848),
.B(n_1180),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1796),
.B(n_1181),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1901),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_1852),
.B(n_1797),
.Y(n_2068)
);

INVxp67_ASAP7_75t_L g2069 ( 
.A(n_1776),
.Y(n_2069)
);

NAND3xp33_ASAP7_75t_L g2070 ( 
.A(n_1817),
.B(n_1179),
.C(n_1049),
.Y(n_2070)
);

BUFx2_ASAP7_75t_L g2071 ( 
.A(n_1732),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1801),
.Y(n_2072)
);

OR2x6_ASAP7_75t_L g2073 ( 
.A(n_1838),
.B(n_896),
.Y(n_2073)
);

AO22x2_ASAP7_75t_L g2074 ( 
.A1(n_1834),
.A2(n_1214),
.B1(n_1215),
.B2(n_1210),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1719),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1849),
.B(n_1188),
.Y(n_2076)
);

INVxp67_ASAP7_75t_L g2077 ( 
.A(n_1779),
.Y(n_2077)
);

AND2x6_ASAP7_75t_L g2078 ( 
.A(n_1678),
.B(n_1049),
.Y(n_2078)
);

NOR2xp33_ASAP7_75t_L g2079 ( 
.A(n_1774),
.B(n_1197),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_1724),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1822),
.Y(n_2081)
);

NOR2xp33_ASAP7_75t_L g2082 ( 
.A(n_1850),
.B(n_1198),
.Y(n_2082)
);

BUFx2_ASAP7_75t_L g2083 ( 
.A(n_1890),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_1819),
.B(n_1199),
.Y(n_2084)
);

OAI22x1_ASAP7_75t_L g2085 ( 
.A1(n_1699),
.A2(n_1203),
.B1(n_1205),
.B2(n_1200),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1707),
.Y(n_2086)
);

AO22x2_ASAP7_75t_L g2087 ( 
.A1(n_1713),
.A2(n_1226),
.B1(n_1229),
.B2(n_1224),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1755),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1845),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1845),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1738),
.Y(n_2091)
);

AO22x2_ASAP7_75t_L g2092 ( 
.A1(n_1761),
.A2(n_917),
.B1(n_949),
.B2(n_896),
.Y(n_2092)
);

A2O1A1Ixp33_ASAP7_75t_L g2093 ( 
.A1(n_1791),
.A2(n_1023),
.B(n_1182),
.C(n_1000),
.Y(n_2093)
);

AND2x6_ASAP7_75t_L g2094 ( 
.A(n_1697),
.B(n_1049),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1751),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1805),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1806),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1844),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1814),
.Y(n_2099)
);

INVxp67_ASAP7_75t_L g2100 ( 
.A(n_1859),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_1855),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_1697),
.Y(n_2102)
);

AOI22xp33_ASAP7_75t_L g2103 ( 
.A1(n_1807),
.A2(n_1179),
.B1(n_1189),
.B2(n_1186),
.Y(n_2103)
);

BUFx8_ASAP7_75t_L g2104 ( 
.A(n_1853),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1698),
.Y(n_2105)
);

AND2x4_ASAP7_75t_L g2106 ( 
.A(n_1820),
.B(n_1),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_1782),
.B(n_1012),
.Y(n_2107)
);

INVx4_ASAP7_75t_L g2108 ( 
.A(n_1859),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1899),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1803),
.Y(n_2110)
);

NAND2x1p5_ASAP7_75t_L g2111 ( 
.A(n_1758),
.B(n_1186),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1881),
.Y(n_2112)
);

INVx1_ASAP7_75t_SL g2113 ( 
.A(n_1859),
.Y(n_2113)
);

AND2x4_ASAP7_75t_L g2114 ( 
.A(n_1894),
.B(n_2),
.Y(n_2114)
);

AND2x4_ASAP7_75t_L g2115 ( 
.A(n_1897),
.B(n_2),
.Y(n_2115)
);

OAI221xp5_ASAP7_75t_L g2116 ( 
.A1(n_1858),
.A2(n_1230),
.B1(n_1189),
.B2(n_1263),
.C(n_1039),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1829),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1829),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1829),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1890),
.B(n_3),
.Y(n_2120)
);

AND2x4_ASAP7_75t_L g2121 ( 
.A(n_1825),
.B(n_3),
.Y(n_2121)
);

HB1xp67_ASAP7_75t_L g2122 ( 
.A(n_1828),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_1890),
.B(n_3),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_1692),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1696),
.Y(n_2125)
);

CKINVDCx5p33_ASAP7_75t_R g2126 ( 
.A(n_1772),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1729),
.Y(n_2127)
);

AO22x2_ASAP7_75t_L g2128 ( 
.A1(n_1705),
.A2(n_1006),
.B1(n_6),
.B2(n_4),
.Y(n_2128)
);

AND2x4_ASAP7_75t_L g2129 ( 
.A(n_1826),
.B(n_4),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_1854),
.B(n_5),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_SL g2131 ( 
.A(n_1847),
.B(n_1230),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_1677),
.Y(n_2132)
);

AND2x4_ASAP7_75t_L g2133 ( 
.A(n_1677),
.B(n_5),
.Y(n_2133)
);

AOI22xp33_ASAP7_75t_L g2134 ( 
.A1(n_1831),
.A2(n_972),
.B1(n_1039),
.B2(n_935),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_1677),
.Y(n_2135)
);

NAND2x1p5_ASAP7_75t_L g2136 ( 
.A(n_1689),
.B(n_935),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_1677),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_1872),
.B(n_7),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1677),
.Y(n_2139)
);

NAND3xp33_ASAP7_75t_L g2140 ( 
.A(n_1783),
.B(n_1157),
.C(n_972),
.Y(n_2140)
);

AO22x2_ASAP7_75t_L g2141 ( 
.A1(n_1712),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1677),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1677),
.B(n_8),
.Y(n_2143)
);

AND2x4_ASAP7_75t_L g2144 ( 
.A(n_1677),
.B(n_8),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_1677),
.B(n_9),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1677),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_1677),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1677),
.Y(n_2148)
);

BUFx4f_ASAP7_75t_L g2149 ( 
.A(n_1746),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_1677),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_1677),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_1677),
.B(n_10),
.Y(n_2152)
);

INVx2_ASAP7_75t_SL g2153 ( 
.A(n_1746),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1677),
.Y(n_2154)
);

AND2x4_ASAP7_75t_L g2155 ( 
.A(n_1677),
.B(n_11),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1677),
.Y(n_2156)
);

NAND2x1p5_ASAP7_75t_L g2157 ( 
.A(n_1689),
.B(n_1157),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_1677),
.B(n_11),
.Y(n_2158)
);

AOI22xp33_ASAP7_75t_L g2159 ( 
.A1(n_1831),
.A2(n_1242),
.B1(n_1267),
.B2(n_1175),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1677),
.Y(n_2160)
);

AO22x2_ASAP7_75t_L g2161 ( 
.A1(n_1712),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_1677),
.B(n_12),
.Y(n_2162)
);

HB1xp67_ASAP7_75t_L g2163 ( 
.A(n_1862),
.Y(n_2163)
);

AO22x2_ASAP7_75t_L g2164 ( 
.A1(n_1712),
.A2(n_18),
.B1(n_15),
.B2(n_16),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1677),
.Y(n_2165)
);

BUFx8_ASAP7_75t_L g2166 ( 
.A(n_1857),
.Y(n_2166)
);

NAND2x1p5_ASAP7_75t_L g2167 ( 
.A(n_1689),
.B(n_15),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1677),
.Y(n_2168)
);

AOI22xp5_ASAP7_75t_L g2169 ( 
.A1(n_1731),
.A2(n_19),
.B1(n_15),
.B2(n_18),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1677),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1677),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_1872),
.B(n_18),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_1677),
.Y(n_2173)
);

BUFx6f_ASAP7_75t_L g2174 ( 
.A(n_1777),
.Y(n_2174)
);

BUFx8_ASAP7_75t_L g2175 ( 
.A(n_1857),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1677),
.Y(n_2176)
);

NAND2x1p5_ASAP7_75t_L g2177 ( 
.A(n_1689),
.B(n_20),
.Y(n_2177)
);

CKINVDCx5p33_ASAP7_75t_R g2178 ( 
.A(n_1703),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1677),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_1677),
.Y(n_2180)
);

BUFx6f_ASAP7_75t_L g2181 ( 
.A(n_1777),
.Y(n_2181)
);

CKINVDCx5p33_ASAP7_75t_R g2182 ( 
.A(n_1703),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1677),
.Y(n_2183)
);

OAI22xp33_ASAP7_75t_SL g2184 ( 
.A1(n_1741),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_2184)
);

AND2x4_ASAP7_75t_L g2185 ( 
.A(n_1677),
.B(n_20),
.Y(n_2185)
);

HB1xp67_ASAP7_75t_L g2186 ( 
.A(n_1862),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1677),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1677),
.Y(n_2188)
);

BUFx3_ASAP7_75t_L g2189 ( 
.A(n_1703),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_1677),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_1677),
.Y(n_2191)
);

OR2x2_ASAP7_75t_L g2192 ( 
.A(n_1691),
.B(n_23),
.Y(n_2192)
);

AO22x2_ASAP7_75t_L g2193 ( 
.A1(n_1712),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_2193)
);

AND2x4_ASAP7_75t_L g2194 ( 
.A(n_1760),
.B(n_26),
.Y(n_2194)
);

AND2x4_ASAP7_75t_L g2195 ( 
.A(n_1760),
.B(n_27),
.Y(n_2195)
);

AND2x4_ASAP7_75t_L g2196 ( 
.A(n_1760),
.B(n_27),
.Y(n_2196)
);

BUFx12f_ASAP7_75t_L g2197 ( 
.A(n_1799),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1677),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1677),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1677),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1677),
.Y(n_2201)
);

CKINVDCx5p33_ASAP7_75t_R g2202 ( 
.A(n_1703),
.Y(n_2202)
);

BUFx6f_ASAP7_75t_L g2203 ( 
.A(n_1777),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1677),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1677),
.Y(n_2205)
);

OAI221xp5_ASAP7_75t_L g2206 ( 
.A1(n_1731),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.C(n_32),
.Y(n_2206)
);

BUFx8_ASAP7_75t_L g2207 ( 
.A(n_1857),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_1677),
.Y(n_2208)
);

CKINVDCx20_ASAP7_75t_R g2209 ( 
.A(n_1703),
.Y(n_2209)
);

AND2x4_ASAP7_75t_L g2210 ( 
.A(n_1760),
.B(n_31),
.Y(n_2210)
);

AOI22xp5_ASAP7_75t_L g2211 ( 
.A1(n_1731),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1677),
.Y(n_2212)
);

AO22x2_ASAP7_75t_L g2213 ( 
.A1(n_1712),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_2213)
);

NAND3xp33_ASAP7_75t_L g2214 ( 
.A(n_1783),
.B(n_36),
.C(n_37),
.Y(n_2214)
);

HB1xp67_ASAP7_75t_L g2215 ( 
.A(n_1862),
.Y(n_2215)
);

AND2x4_ASAP7_75t_L g2216 ( 
.A(n_1677),
.B(n_37),
.Y(n_2216)
);

OAI221xp5_ASAP7_75t_L g2217 ( 
.A1(n_1731),
.A2(n_41),
.B1(n_38),
.B2(n_39),
.C(n_42),
.Y(n_2217)
);

AND2x4_ASAP7_75t_L g2218 ( 
.A(n_1677),
.B(n_38),
.Y(n_2218)
);

NOR2xp33_ASAP7_75t_SL g2219 ( 
.A(n_1689),
.B(n_39),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1677),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_1677),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_1677),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1677),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_1677),
.Y(n_2224)
);

AND2x4_ASAP7_75t_L g2225 ( 
.A(n_1677),
.B(n_43),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1677),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_1677),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_1677),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_1872),
.B(n_44),
.Y(n_2229)
);

CKINVDCx5p33_ASAP7_75t_R g2230 ( 
.A(n_1703),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1677),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1677),
.Y(n_2232)
);

OAI22xp5_ASAP7_75t_SL g2233 ( 
.A1(n_1703),
.A2(n_46),
.B1(n_47),
.B2(n_45),
.Y(n_2233)
);

AO22x2_ASAP7_75t_L g2234 ( 
.A1(n_1712),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_1677),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_1677),
.B(n_48),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1677),
.Y(n_2237)
);

BUFx6f_ASAP7_75t_L g2238 ( 
.A(n_1777),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1677),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1677),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1677),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_1677),
.B(n_48),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_1677),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_1677),
.Y(n_2244)
);

INVx1_ASAP7_75t_SL g2245 ( 
.A(n_1691),
.Y(n_2245)
);

AND2x4_ASAP7_75t_L g2246 ( 
.A(n_1677),
.B(n_49),
.Y(n_2246)
);

AND2x4_ASAP7_75t_L g2247 ( 
.A(n_1677),
.B(n_49),
.Y(n_2247)
);

INVxp67_ASAP7_75t_L g2248 ( 
.A(n_1862),
.Y(n_2248)
);

AOI22xp5_ASAP7_75t_L g2249 ( 
.A1(n_1731),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_2249)
);

AO22x2_ASAP7_75t_L g2250 ( 
.A1(n_1712),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_1677),
.Y(n_2251)
);

CKINVDCx20_ASAP7_75t_R g2252 ( 
.A(n_1703),
.Y(n_2252)
);

AO22x2_ASAP7_75t_L g2253 ( 
.A1(n_1712),
.A2(n_53),
.B1(n_50),
.B2(n_51),
.Y(n_2253)
);

AND2x4_ASAP7_75t_L g2254 ( 
.A(n_1677),
.B(n_54),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1677),
.Y(n_2255)
);

INVx2_ASAP7_75t_L g2256 ( 
.A(n_1677),
.Y(n_2256)
);

CKINVDCx5p33_ASAP7_75t_R g2257 ( 
.A(n_1703),
.Y(n_2257)
);

AND2x4_ASAP7_75t_L g2258 ( 
.A(n_1677),
.B(n_54),
.Y(n_2258)
);

OAI22xp5_ASAP7_75t_SL g2259 ( 
.A1(n_1703),
.A2(n_57),
.B1(n_58),
.B2(n_56),
.Y(n_2259)
);

NOR2xp33_ASAP7_75t_L g2260 ( 
.A(n_1731),
.B(n_55),
.Y(n_2260)
);

AND2x4_ASAP7_75t_L g2261 ( 
.A(n_1677),
.B(n_55),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_1677),
.B(n_56),
.Y(n_2262)
);

AND2x4_ASAP7_75t_L g2263 ( 
.A(n_1677),
.B(n_57),
.Y(n_2263)
);

INVxp67_ASAP7_75t_L g2264 ( 
.A(n_1862),
.Y(n_2264)
);

AND2x4_ASAP7_75t_L g2265 ( 
.A(n_1677),
.B(n_59),
.Y(n_2265)
);

BUFx6f_ASAP7_75t_L g2266 ( 
.A(n_1777),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_1872),
.B(n_60),
.Y(n_2267)
);

HB1xp67_ASAP7_75t_L g2268 ( 
.A(n_1862),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_1677),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_1677),
.Y(n_2270)
);

AO22x2_ASAP7_75t_L g2271 ( 
.A1(n_1712),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_2271)
);

AOI22xp33_ASAP7_75t_L g2272 ( 
.A1(n_1831),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_1872),
.B(n_65),
.Y(n_2273)
);

OAI22xp5_ASAP7_75t_L g2274 ( 
.A1(n_1677),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_1677),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_1677),
.Y(n_2276)
);

NOR2xp33_ASAP7_75t_L g2277 ( 
.A(n_1731),
.B(n_65),
.Y(n_2277)
);

AND2x4_ASAP7_75t_L g2278 ( 
.A(n_1677),
.B(n_67),
.Y(n_2278)
);

AO22x2_ASAP7_75t_L g2279 ( 
.A1(n_1712),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_1677),
.Y(n_2280)
);

OR2x6_ASAP7_75t_SL g2281 ( 
.A(n_1752),
.B(n_70),
.Y(n_2281)
);

INVxp67_ASAP7_75t_L g2282 ( 
.A(n_1862),
.Y(n_2282)
);

AND2x4_ASAP7_75t_L g2283 ( 
.A(n_1677),
.B(n_68),
.Y(n_2283)
);

HB1xp67_ASAP7_75t_L g2284 ( 
.A(n_1862),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_1677),
.Y(n_2285)
);

CKINVDCx16_ASAP7_75t_R g2286 ( 
.A(n_1703),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_1677),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_1677),
.B(n_72),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_1677),
.Y(n_2289)
);

BUFx2_ASAP7_75t_L g2290 ( 
.A(n_1862),
.Y(n_2290)
);

O2A1O1Ixp5_ASAP7_75t_L g2291 ( 
.A1(n_1940),
.A2(n_75),
.B(n_73),
.C(n_74),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_1927),
.Y(n_2292)
);

INVx2_ASAP7_75t_L g2293 ( 
.A(n_1903),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2068),
.B(n_75),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_1924),
.B(n_76),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_1948),
.B(n_1980),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_1930),
.Y(n_2297)
);

O2A1O1Ixp33_ASAP7_75t_L g2298 ( 
.A1(n_2025),
.A2(n_79),
.B(n_77),
.C(n_78),
.Y(n_2298)
);

AOI21xp5_ASAP7_75t_L g2299 ( 
.A1(n_2140),
.A2(n_2009),
.B(n_2004),
.Y(n_2299)
);

INVx4_ASAP7_75t_L g2300 ( 
.A(n_2149),
.Y(n_2300)
);

INVx5_ASAP7_75t_L g2301 ( 
.A(n_1968),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_1905),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_1997),
.B(n_78),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_1998),
.B(n_80),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_1945),
.Y(n_2305)
);

INVx4_ASAP7_75t_L g2306 ( 
.A(n_1947),
.Y(n_2306)
);

AOI21x1_ASAP7_75t_L g2307 ( 
.A1(n_2013),
.A2(n_84),
.B(n_85),
.Y(n_2307)
);

INVx2_ASAP7_75t_SL g2308 ( 
.A(n_1947),
.Y(n_2308)
);

AOI21xp5_ASAP7_75t_L g2309 ( 
.A1(n_2022),
.A2(n_84),
.B(n_85),
.Y(n_2309)
);

O2A1O1Ixp5_ASAP7_75t_SL g2310 ( 
.A1(n_2127),
.A2(n_639),
.B(n_640),
.C(n_638),
.Y(n_2310)
);

OAI21xp5_ASAP7_75t_L g2311 ( 
.A1(n_1926),
.A2(n_87),
.B(n_88),
.Y(n_2311)
);

AO32x2_ASAP7_75t_L g2312 ( 
.A1(n_2274),
.A2(n_92),
.A3(n_89),
.B1(n_91),
.B2(n_93),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_1935),
.B(n_89),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_1914),
.Y(n_2314)
);

CKINVDCx8_ASAP7_75t_R g2315 ( 
.A(n_2286),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_1919),
.Y(n_2316)
);

AOI21xp5_ASAP7_75t_L g2317 ( 
.A1(n_2006),
.A2(n_94),
.B(n_95),
.Y(n_2317)
);

NOR2xp33_ASAP7_75t_L g2318 ( 
.A(n_1956),
.B(n_94),
.Y(n_2318)
);

BUFx8_ASAP7_75t_L g2319 ( 
.A(n_2197),
.Y(n_2319)
);

OAI21xp5_ASAP7_75t_L g2320 ( 
.A1(n_2093),
.A2(n_96),
.B(n_97),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_SL g2321 ( 
.A(n_2219),
.B(n_640),
.Y(n_2321)
);

A2O1A1Ixp33_ASAP7_75t_L g2322 ( 
.A1(n_2214),
.A2(n_98),
.B(n_96),
.C(n_97),
.Y(n_2322)
);

AOI21x1_ASAP7_75t_L g2323 ( 
.A1(n_2071),
.A2(n_98),
.B(n_99),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_1932),
.B(n_1936),
.Y(n_2324)
);

AOI21xp5_ASAP7_75t_L g2325 ( 
.A1(n_1962),
.A2(n_1952),
.B(n_1946),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2003),
.Y(n_2326)
);

NAND2x1p5_ASAP7_75t_L g2327 ( 
.A(n_2174),
.B(n_2181),
.Y(n_2327)
);

NOR2xp33_ASAP7_75t_L g2328 ( 
.A(n_1965),
.B(n_100),
.Y(n_2328)
);

AOI21xp5_ASAP7_75t_L g2329 ( 
.A1(n_1961),
.A2(n_102),
.B(n_103),
.Y(n_2329)
);

AOI21xp5_ASAP7_75t_L g2330 ( 
.A1(n_2034),
.A2(n_102),
.B(n_103),
.Y(n_2330)
);

BUFx6f_ASAP7_75t_L g2331 ( 
.A(n_1978),
.Y(n_2331)
);

BUFx4f_ASAP7_75t_L g2332 ( 
.A(n_2019),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_1920),
.Y(n_2333)
);

AOI21xp5_ASAP7_75t_L g2334 ( 
.A1(n_2124),
.A2(n_104),
.B(n_105),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_1942),
.B(n_1906),
.Y(n_2335)
);

OR2x6_ASAP7_75t_L g2336 ( 
.A(n_1960),
.B(n_106),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_1907),
.B(n_107),
.Y(n_2337)
);

HB1xp67_ASAP7_75t_L g2338 ( 
.A(n_2290),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_1921),
.Y(n_2339)
);

AOI21x1_ASAP7_75t_L g2340 ( 
.A1(n_2071),
.A2(n_108),
.B(n_109),
.Y(n_2340)
);

AOI21xp5_ASAP7_75t_L g2341 ( 
.A1(n_2125),
.A2(n_108),
.B(n_109),
.Y(n_2341)
);

HB1xp67_ASAP7_75t_L g2342 ( 
.A(n_1902),
.Y(n_2342)
);

BUFx3_ASAP7_75t_L g2343 ( 
.A(n_2174),
.Y(n_2343)
);

HB1xp67_ASAP7_75t_L g2344 ( 
.A(n_2163),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_1911),
.B(n_110),
.Y(n_2345)
);

BUFx2_ASAP7_75t_L g2346 ( 
.A(n_2209),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_SL g2347 ( 
.A(n_1918),
.B(n_644),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_1912),
.B(n_111),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_2132),
.Y(n_2349)
);

AOI21xp5_ASAP7_75t_L g2350 ( 
.A1(n_1922),
.A2(n_111),
.B(n_112),
.Y(n_2350)
);

BUFx6f_ASAP7_75t_L g2351 ( 
.A(n_1978),
.Y(n_2351)
);

OAI21xp5_ASAP7_75t_L g2352 ( 
.A1(n_2143),
.A2(n_112),
.B(n_113),
.Y(n_2352)
);

BUFx6f_ASAP7_75t_L g2353 ( 
.A(n_1994),
.Y(n_2353)
);

AOI21xp5_ASAP7_75t_L g2354 ( 
.A1(n_1923),
.A2(n_114),
.B(n_115),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_2135),
.Y(n_2355)
);

AND2x2_ASAP7_75t_L g2356 ( 
.A(n_1935),
.B(n_114),
.Y(n_2356)
);

AND2x2_ASAP7_75t_L g2357 ( 
.A(n_1934),
.B(n_115),
.Y(n_2357)
);

INVxp67_ASAP7_75t_SL g2358 ( 
.A(n_2186),
.Y(n_2358)
);

AND2x4_ASAP7_75t_L g2359 ( 
.A(n_1913),
.B(n_116),
.Y(n_2359)
);

OAI21xp5_ASAP7_75t_L g2360 ( 
.A1(n_2145),
.A2(n_116),
.B(n_117),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_1915),
.B(n_118),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_SL g2362 ( 
.A(n_2043),
.B(n_2108),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_1917),
.B(n_121),
.Y(n_2363)
);

HB1xp67_ASAP7_75t_L g2364 ( 
.A(n_2215),
.Y(n_2364)
);

INVxp67_ASAP7_75t_SL g2365 ( 
.A(n_2268),
.Y(n_2365)
);

BUFx6f_ASAP7_75t_L g2366 ( 
.A(n_1994),
.Y(n_2366)
);

BUFx6f_ASAP7_75t_L g2367 ( 
.A(n_2027),
.Y(n_2367)
);

BUFx4f_ASAP7_75t_L g2368 ( 
.A(n_2019),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2133),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2139),
.B(n_123),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2144),
.Y(n_2371)
);

AND2x2_ASAP7_75t_L g2372 ( 
.A(n_1934),
.B(n_126),
.Y(n_2372)
);

HB1xp67_ASAP7_75t_L g2373 ( 
.A(n_2284),
.Y(n_2373)
);

AOI21xp5_ASAP7_75t_L g2374 ( 
.A1(n_2070),
.A2(n_128),
.B(n_129),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2137),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2142),
.B(n_130),
.Y(n_2376)
);

AOI21xp5_ASAP7_75t_L g2377 ( 
.A1(n_1904),
.A2(n_131),
.B(n_132),
.Y(n_2377)
);

AOI22xp5_ASAP7_75t_L g2378 ( 
.A1(n_1949),
.A2(n_2008),
.B1(n_1963),
.B2(n_1933),
.Y(n_2378)
);

O2A1O1Ixp33_ASAP7_75t_L g2379 ( 
.A1(n_2061),
.A2(n_2064),
.B(n_2277),
.C(n_2260),
.Y(n_2379)
);

AOI21xp5_ASAP7_75t_L g2380 ( 
.A1(n_1910),
.A2(n_132),
.B(n_133),
.Y(n_2380)
);

AOI21xp5_ASAP7_75t_L g2381 ( 
.A1(n_2152),
.A2(n_133),
.B(n_134),
.Y(n_2381)
);

AOI21xp5_ASAP7_75t_L g2382 ( 
.A1(n_2158),
.A2(n_136),
.B(n_137),
.Y(n_2382)
);

NOR2xp67_ASAP7_75t_L g2383 ( 
.A(n_2248),
.B(n_136),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2147),
.Y(n_2384)
);

AO21x1_ASAP7_75t_L g2385 ( 
.A1(n_2184),
.A2(n_647),
.B(n_646),
.Y(n_2385)
);

AOI21xp5_ASAP7_75t_L g2386 ( 
.A1(n_2162),
.A2(n_137),
.B(n_138),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2146),
.B(n_139),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_2150),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2155),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2148),
.B(n_141),
.Y(n_2390)
);

NOR3xp33_ASAP7_75t_L g2391 ( 
.A(n_2233),
.B(n_143),
.C(n_144),
.Y(n_2391)
);

AND2x2_ASAP7_75t_L g2392 ( 
.A(n_1908),
.B(n_1958),
.Y(n_2392)
);

AOI21xp5_ASAP7_75t_L g2393 ( 
.A1(n_2236),
.A2(n_146),
.B(n_148),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_2156),
.B(n_146),
.Y(n_2394)
);

OAI21xp5_ASAP7_75t_L g2395 ( 
.A1(n_2242),
.A2(n_148),
.B(n_149),
.Y(n_2395)
);

BUFx3_ASAP7_75t_L g2396 ( 
.A(n_2203),
.Y(n_2396)
);

BUFx6f_ASAP7_75t_L g2397 ( 
.A(n_2027),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2155),
.Y(n_2398)
);

AOI21xp5_ASAP7_75t_L g2399 ( 
.A1(n_2262),
.A2(n_150),
.B(n_151),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_2160),
.B(n_152),
.Y(n_2400)
);

AND2x2_ASAP7_75t_L g2401 ( 
.A(n_2015),
.B(n_152),
.Y(n_2401)
);

CKINVDCx10_ASAP7_75t_R g2402 ( 
.A(n_1960),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2170),
.B(n_2171),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_2176),
.B(n_154),
.Y(n_2404)
);

BUFx12f_ASAP7_75t_L g2405 ( 
.A(n_1941),
.Y(n_2405)
);

INVx2_ASAP7_75t_L g2406 ( 
.A(n_2151),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_2179),
.B(n_155),
.Y(n_2407)
);

AOI22xp5_ASAP7_75t_L g2408 ( 
.A1(n_1950),
.A2(n_158),
.B1(n_156),
.B2(n_157),
.Y(n_2408)
);

BUFx2_ASAP7_75t_SL g2409 ( 
.A(n_2252),
.Y(n_2409)
);

OAI21x1_ASAP7_75t_L g2410 ( 
.A1(n_2096),
.A2(n_157),
.B(n_158),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_SL g2411 ( 
.A(n_2044),
.B(n_647),
.Y(n_2411)
);

NAND3xp33_ASAP7_75t_L g2412 ( 
.A(n_1970),
.B(n_2159),
.C(n_2134),
.Y(n_2412)
);

OAI21xp5_ASAP7_75t_L g2413 ( 
.A1(n_2288),
.A2(n_2056),
.B(n_1943),
.Y(n_2413)
);

NOR2xp33_ASAP7_75t_L g2414 ( 
.A(n_2245),
.B(n_159),
.Y(n_2414)
);

NOR2xp67_ASAP7_75t_L g2415 ( 
.A(n_2264),
.B(n_161),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_2183),
.B(n_161),
.Y(n_2416)
);

AOI21xp5_ASAP7_75t_L g2417 ( 
.A1(n_2097),
.A2(n_162),
.B(n_163),
.Y(n_2417)
);

AOI21xp5_ASAP7_75t_L g2418 ( 
.A1(n_2099),
.A2(n_163),
.B(n_164),
.Y(n_2418)
);

AOI21xp5_ASAP7_75t_L g2419 ( 
.A1(n_2107),
.A2(n_164),
.B(n_165),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2154),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2165),
.Y(n_2421)
);

AND2x4_ASAP7_75t_L g2422 ( 
.A(n_2187),
.B(n_165),
.Y(n_2422)
);

AND2x4_ASAP7_75t_L g2423 ( 
.A(n_2188),
.B(n_167),
.Y(n_2423)
);

O2A1O1Ixp33_ASAP7_75t_L g2424 ( 
.A1(n_2026),
.A2(n_2130),
.B(n_1951),
.C(n_1957),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2185),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_2168),
.Y(n_2426)
);

OAI22xp5_ASAP7_75t_L g2427 ( 
.A1(n_2216),
.A2(n_171),
.B1(n_169),
.B2(n_170),
.Y(n_2427)
);

INVx3_ASAP7_75t_L g2428 ( 
.A(n_2203),
.Y(n_2428)
);

BUFx6f_ASAP7_75t_L g2429 ( 
.A(n_2055),
.Y(n_2429)
);

AOI21xp5_ASAP7_75t_L g2430 ( 
.A1(n_1989),
.A2(n_170),
.B(n_171),
.Y(n_2430)
);

BUFx6f_ASAP7_75t_L g2431 ( 
.A(n_2047),
.Y(n_2431)
);

AOI22xp5_ASAP7_75t_L g2432 ( 
.A1(n_2084),
.A2(n_173),
.B1(n_171),
.B2(n_172),
.Y(n_2432)
);

AOI21xp5_ASAP7_75t_L g2433 ( 
.A1(n_1985),
.A2(n_173),
.B(n_174),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2198),
.B(n_173),
.Y(n_2434)
);

A2O1A1Ixp33_ASAP7_75t_L g2435 ( 
.A1(n_2206),
.A2(n_176),
.B(n_174),
.C(n_175),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_2173),
.Y(n_2436)
);

INVx1_ASAP7_75t_SL g2437 ( 
.A(n_2012),
.Y(n_2437)
);

INVx3_ASAP7_75t_L g2438 ( 
.A(n_2238),
.Y(n_2438)
);

NOR3xp33_ASAP7_75t_L g2439 ( 
.A(n_2259),
.B(n_2060),
.C(n_2217),
.Y(n_2439)
);

INVx1_ASAP7_75t_SL g2440 ( 
.A(n_1916),
.Y(n_2440)
);

A2O1A1Ixp33_ASAP7_75t_L g2441 ( 
.A1(n_2169),
.A2(n_180),
.B(n_178),
.C(n_179),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2218),
.Y(n_2442)
);

OR2x6_ASAP7_75t_L g2443 ( 
.A(n_2167),
.B(n_178),
.Y(n_2443)
);

AOI21xp5_ASAP7_75t_L g2444 ( 
.A1(n_2028),
.A2(n_181),
.B(n_182),
.Y(n_2444)
);

AOI21xp5_ASAP7_75t_L g2445 ( 
.A1(n_2032),
.A2(n_182),
.B(n_183),
.Y(n_2445)
);

OAI22xp5_ASAP7_75t_L g2446 ( 
.A1(n_2218),
.A2(n_185),
.B1(n_183),
.B2(n_184),
.Y(n_2446)
);

INVxp67_ASAP7_75t_L g2447 ( 
.A(n_2225),
.Y(n_2447)
);

AO21x1_ASAP7_75t_L g2448 ( 
.A1(n_2021),
.A2(n_649),
.B(n_648),
.Y(n_2448)
);

BUFx2_ASAP7_75t_L g2449 ( 
.A(n_2054),
.Y(n_2449)
);

AOI21xp5_ASAP7_75t_L g2450 ( 
.A1(n_2040),
.A2(n_2101),
.B(n_2098),
.Y(n_2450)
);

AND2x4_ASAP7_75t_L g2451 ( 
.A(n_2199),
.B(n_183),
.Y(n_2451)
);

AOI22xp5_ASAP7_75t_L g2452 ( 
.A1(n_1928),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_2200),
.B(n_184),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2201),
.B(n_187),
.Y(n_2454)
);

O2A1O1Ixp33_ASAP7_75t_L g2455 ( 
.A1(n_2020),
.A2(n_1967),
.B(n_1973),
.C(n_1971),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2180),
.Y(n_2456)
);

A2O1A1Ixp33_ASAP7_75t_L g2457 ( 
.A1(n_2211),
.A2(n_190),
.B(n_187),
.C(n_189),
.Y(n_2457)
);

NAND2x1p5_ASAP7_75t_L g2458 ( 
.A(n_2238),
.B(n_189),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_2204),
.B(n_2205),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2190),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_2208),
.B(n_2212),
.Y(n_2461)
);

AOI22x1_ASAP7_75t_L g2462 ( 
.A1(n_1986),
.A2(n_191),
.B1(n_189),
.B2(n_190),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2225),
.Y(n_2463)
);

BUFx3_ASAP7_75t_L g2464 ( 
.A(n_2266),
.Y(n_2464)
);

OAI21xp5_ASAP7_75t_L g2465 ( 
.A1(n_2014),
.A2(n_190),
.B(n_191),
.Y(n_2465)
);

AOI21x1_ASAP7_75t_L g2466 ( 
.A1(n_2087),
.A2(n_191),
.B(n_192),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_2191),
.Y(n_2467)
);

AND2x6_ASAP7_75t_L g2468 ( 
.A(n_2246),
.B(n_193),
.Y(n_2468)
);

AO32x1_ASAP7_75t_L g2469 ( 
.A1(n_2117),
.A2(n_196),
.A3(n_194),
.B1(n_195),
.B2(n_197),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_L g2470 ( 
.A(n_2220),
.B(n_195),
.Y(n_2470)
);

AOI21xp5_ASAP7_75t_L g2471 ( 
.A1(n_2223),
.A2(n_196),
.B(n_197),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2246),
.Y(n_2472)
);

INVx4_ASAP7_75t_L g2473 ( 
.A(n_1968),
.Y(n_2473)
);

AOI21xp5_ASAP7_75t_L g2474 ( 
.A1(n_2226),
.A2(n_198),
.B(n_199),
.Y(n_2474)
);

BUFx2_ASAP7_75t_L g2475 ( 
.A(n_2178),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2231),
.B(n_200),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_2232),
.B(n_2237),
.Y(n_2477)
);

AOI21xp5_ASAP7_75t_L g2478 ( 
.A1(n_2239),
.A2(n_200),
.B(n_201),
.Y(n_2478)
);

OAI21x1_ASAP7_75t_L g2479 ( 
.A1(n_2030),
.A2(n_200),
.B(n_201),
.Y(n_2479)
);

AOI21xp5_ASAP7_75t_L g2480 ( 
.A1(n_2240),
.A2(n_201),
.B(n_202),
.Y(n_2480)
);

O2A1O1Ixp5_ASAP7_75t_L g2481 ( 
.A1(n_2131),
.A2(n_205),
.B(n_203),
.C(n_204),
.Y(n_2481)
);

NOR2x1p5_ASAP7_75t_SL g2482 ( 
.A(n_2118),
.B(n_2119),
.Y(n_2482)
);

AOI22xp5_ASAP7_75t_L g2483 ( 
.A1(n_1931),
.A2(n_205),
.B1(n_203),
.B2(n_204),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2241),
.B(n_203),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_L g2485 ( 
.A(n_2244),
.B(n_205),
.Y(n_2485)
);

AND2x2_ASAP7_75t_L g2486 ( 
.A(n_2036),
.B(n_206),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2247),
.Y(n_2487)
);

AOI22xp5_ASAP7_75t_L g2488 ( 
.A1(n_1938),
.A2(n_208),
.B1(n_206),
.B2(n_207),
.Y(n_2488)
);

AOI21xp5_ASAP7_75t_L g2489 ( 
.A1(n_2251),
.A2(n_208),
.B(n_209),
.Y(n_2489)
);

INVx1_ASAP7_75t_SL g2490 ( 
.A(n_2189),
.Y(n_2490)
);

BUFx2_ASAP7_75t_L g2491 ( 
.A(n_2182),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_2255),
.B(n_209),
.Y(n_2492)
);

OAI21xp5_ASAP7_75t_L g2493 ( 
.A1(n_1992),
.A2(n_211),
.B(n_212),
.Y(n_2493)
);

NOR2xp67_ASAP7_75t_L g2494 ( 
.A(n_2282),
.B(n_211),
.Y(n_2494)
);

BUFx2_ASAP7_75t_L g2495 ( 
.A(n_2202),
.Y(n_2495)
);

AOI21x1_ASAP7_75t_L g2496 ( 
.A1(n_2087),
.A2(n_214),
.B(n_215),
.Y(n_2496)
);

AOI21x1_ASAP7_75t_L g2497 ( 
.A1(n_2083),
.A2(n_216),
.B(n_217),
.Y(n_2497)
);

AOI21xp5_ASAP7_75t_L g2498 ( 
.A1(n_2269),
.A2(n_216),
.B(n_217),
.Y(n_2498)
);

AOI21xp5_ASAP7_75t_L g2499 ( 
.A1(n_2270),
.A2(n_218),
.B(n_219),
.Y(n_2499)
);

BUFx2_ASAP7_75t_L g2500 ( 
.A(n_2230),
.Y(n_2500)
);

OAI22xp5_ASAP7_75t_L g2501 ( 
.A1(n_2254),
.A2(n_222),
.B1(n_220),
.B2(n_221),
.Y(n_2501)
);

BUFx6f_ASAP7_75t_L g2502 ( 
.A(n_2047),
.Y(n_2502)
);

OAI21xp5_ASAP7_75t_L g2503 ( 
.A1(n_2062),
.A2(n_222),
.B(n_223),
.Y(n_2503)
);

CKINVDCx5p33_ASAP7_75t_R g2504 ( 
.A(n_2257),
.Y(n_2504)
);

BUFx6f_ASAP7_75t_L g2505 ( 
.A(n_2078),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2285),
.B(n_2287),
.Y(n_2506)
);

AND2x4_ASAP7_75t_L g2507 ( 
.A(n_2289),
.B(n_225),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_2221),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_2222),
.Y(n_2509)
);

OAI22xp5_ASAP7_75t_L g2510 ( 
.A1(n_2258),
.A2(n_2261),
.B1(n_2265),
.B2(n_2263),
.Y(n_2510)
);

AOI21xp5_ASAP7_75t_L g2511 ( 
.A1(n_2224),
.A2(n_228),
.B(n_229),
.Y(n_2511)
);

AOI21xp5_ASAP7_75t_L g2512 ( 
.A1(n_2227),
.A2(n_230),
.B(n_232),
.Y(n_2512)
);

AOI21xp5_ASAP7_75t_L g2513 ( 
.A1(n_2228),
.A2(n_232),
.B(n_233),
.Y(n_2513)
);

AOI21xp5_ASAP7_75t_L g2514 ( 
.A1(n_2235),
.A2(n_233),
.B(n_234),
.Y(n_2514)
);

O2A1O1Ixp33_ASAP7_75t_L g2515 ( 
.A1(n_2031),
.A2(n_237),
.B(n_235),
.C(n_236),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_2138),
.B(n_235),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_2172),
.B(n_237),
.Y(n_2517)
);

INVxp67_ASAP7_75t_L g2518 ( 
.A(n_2258),
.Y(n_2518)
);

AOI21xp33_ASAP7_75t_L g2519 ( 
.A1(n_2079),
.A2(n_239),
.B(n_240),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2261),
.Y(n_2520)
);

OAI22xp5_ASAP7_75t_L g2521 ( 
.A1(n_2263),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.Y(n_2521)
);

AOI21xp5_ASAP7_75t_L g2522 ( 
.A1(n_2243),
.A2(n_241),
.B(n_242),
.Y(n_2522)
);

AOI21xp5_ASAP7_75t_L g2523 ( 
.A1(n_2256),
.A2(n_241),
.B(n_242),
.Y(n_2523)
);

OAI21xp5_ASAP7_75t_L g2524 ( 
.A1(n_2063),
.A2(n_242),
.B(n_243),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_L g2525 ( 
.A(n_2229),
.B(n_243),
.Y(n_2525)
);

AOI21xp5_ASAP7_75t_L g2526 ( 
.A1(n_2275),
.A2(n_244),
.B(n_245),
.Y(n_2526)
);

AND2x4_ASAP7_75t_L g2527 ( 
.A(n_2276),
.B(n_246),
.Y(n_2527)
);

BUFx6f_ASAP7_75t_L g2528 ( 
.A(n_2078),
.Y(n_2528)
);

AND2x4_ASAP7_75t_L g2529 ( 
.A(n_2280),
.B(n_246),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2265),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2267),
.B(n_247),
.Y(n_2531)
);

O2A1O1Ixp33_ASAP7_75t_L g2532 ( 
.A1(n_2066),
.A2(n_250),
.B(n_248),
.C(n_249),
.Y(n_2532)
);

A2O1A1Ixp33_ASAP7_75t_L g2533 ( 
.A1(n_2249),
.A2(n_253),
.B(n_251),
.C(n_252),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2273),
.B(n_253),
.Y(n_2534)
);

INVx3_ASAP7_75t_L g2535 ( 
.A(n_2166),
.Y(n_2535)
);

OAI22xp5_ASAP7_75t_L g2536 ( 
.A1(n_2278),
.A2(n_258),
.B1(n_256),
.B2(n_257),
.Y(n_2536)
);

INVxp67_ASAP7_75t_L g2537 ( 
.A(n_2283),
.Y(n_2537)
);

NAND2xp33_ASAP7_75t_L g2538 ( 
.A(n_2078),
.B(n_256),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2283),
.Y(n_2539)
);

NOR2xp33_ASAP7_75t_L g2540 ( 
.A(n_2045),
.B(n_259),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_SL g2541 ( 
.A(n_2111),
.B(n_650),
.Y(n_2541)
);

BUFx6f_ASAP7_75t_L g2542 ( 
.A(n_2094),
.Y(n_2542)
);

NOR2xp33_ASAP7_75t_L g2543 ( 
.A(n_2039),
.B(n_260),
.Y(n_2543)
);

INVx1_ASAP7_75t_SL g2544 ( 
.A(n_1988),
.Y(n_2544)
);

OAI21xp33_ASAP7_75t_L g2545 ( 
.A1(n_1987),
.A2(n_263),
.B(n_264),
.Y(n_2545)
);

BUFx4f_ASAP7_75t_L g2546 ( 
.A(n_2177),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_L g2547 ( 
.A(n_1976),
.B(n_266),
.Y(n_2547)
);

AOI21xp5_ASAP7_75t_L g2548 ( 
.A1(n_1969),
.A2(n_267),
.B(n_268),
.Y(n_2548)
);

INVx6_ASAP7_75t_L g2549 ( 
.A(n_2175),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_1993),
.B(n_270),
.Y(n_2550)
);

OAI21xp5_ASAP7_75t_L g2551 ( 
.A1(n_2076),
.A2(n_271),
.B(n_272),
.Y(n_2551)
);

INVx4_ASAP7_75t_L g2552 ( 
.A(n_2017),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2042),
.B(n_271),
.Y(n_2553)
);

OAI22xp5_ASAP7_75t_L g2554 ( 
.A1(n_2005),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.Y(n_2554)
);

INVx3_ASAP7_75t_L g2555 ( 
.A(n_2207),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_1977),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_SL g2557 ( 
.A(n_2058),
.B(n_651),
.Y(n_2557)
);

INVx5_ASAP7_75t_L g2558 ( 
.A(n_1968),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_1981),
.Y(n_2559)
);

NOR3xp33_ASAP7_75t_L g2560 ( 
.A(n_1955),
.B(n_276),
.C(n_277),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2023),
.Y(n_2561)
);

AND2x2_ASAP7_75t_L g2562 ( 
.A(n_1975),
.B(n_276),
.Y(n_2562)
);

OAI21xp5_ASAP7_75t_L g2563 ( 
.A1(n_1909),
.A2(n_279),
.B(n_281),
.Y(n_2563)
);

AOI21x1_ASAP7_75t_L g2564 ( 
.A1(n_2128),
.A2(n_282),
.B(n_283),
.Y(n_2564)
);

AND2x2_ASAP7_75t_L g2565 ( 
.A(n_1975),
.B(n_282),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_L g2566 ( 
.A(n_1982),
.B(n_283),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_1984),
.B(n_283),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_1979),
.Y(n_2568)
);

INVx3_ASAP7_75t_L g2569 ( 
.A(n_2104),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_SL g2570 ( 
.A(n_2113),
.B(n_652),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2000),
.Y(n_2571)
);

AOI21xp5_ASAP7_75t_L g2572 ( 
.A1(n_2072),
.A2(n_285),
.B(n_286),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_L g2573 ( 
.A(n_1966),
.B(n_285),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2081),
.B(n_285),
.Y(n_2574)
);

HB1xp67_ASAP7_75t_L g2575 ( 
.A(n_1988),
.Y(n_2575)
);

INVx1_ASAP7_75t_SL g2576 ( 
.A(n_1959),
.Y(n_2576)
);

AOI21xp5_ASAP7_75t_L g2577 ( 
.A1(n_2011),
.A2(n_288),
.B(n_289),
.Y(n_2577)
);

AOI21xp5_ASAP7_75t_L g2578 ( 
.A1(n_2116),
.A2(n_2049),
.B(n_2048),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_L g2579 ( 
.A(n_1954),
.B(n_291),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_SL g2580 ( 
.A(n_2016),
.B(n_653),
.Y(n_2580)
);

AOI21xp5_ASAP7_75t_L g2581 ( 
.A1(n_2052),
.A2(n_292),
.B(n_293),
.Y(n_2581)
);

AOI21xp5_ASAP7_75t_L g2582 ( 
.A1(n_2053),
.A2(n_292),
.B(n_293),
.Y(n_2582)
);

INVxp67_ASAP7_75t_L g2583 ( 
.A(n_2281),
.Y(n_2583)
);

AOI21xp5_ASAP7_75t_L g2584 ( 
.A1(n_2057),
.A2(n_293),
.B(n_294),
.Y(n_2584)
);

INVx1_ASAP7_75t_SL g2585 ( 
.A(n_1990),
.Y(n_2585)
);

BUFx2_ASAP7_75t_L g2586 ( 
.A(n_2073),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2141),
.Y(n_2587)
);

AOI21xp5_ASAP7_75t_L g2588 ( 
.A1(n_2059),
.A2(n_295),
.B(n_296),
.Y(n_2588)
);

AO21x1_ASAP7_75t_L g2589 ( 
.A1(n_2114),
.A2(n_655),
.B(n_654),
.Y(n_2589)
);

AND2x2_ASAP7_75t_SL g2590 ( 
.A(n_2121),
.B(n_297),
.Y(n_2590)
);

INVx2_ASAP7_75t_L g2591 ( 
.A(n_2115),
.Y(n_2591)
);

OAI21xp33_ASAP7_75t_L g2592 ( 
.A1(n_2001),
.A2(n_298),
.B(n_299),
.Y(n_2592)
);

AND2x4_ASAP7_75t_L g2593 ( 
.A(n_2110),
.B(n_298),
.Y(n_2593)
);

OAI21x1_ASAP7_75t_L g2594 ( 
.A1(n_2075),
.A2(n_300),
.B(n_301),
.Y(n_2594)
);

OR2x6_ASAP7_75t_SL g2595 ( 
.A(n_2126),
.B(n_2192),
.Y(n_2595)
);

NOR2xp33_ASAP7_75t_L g2596 ( 
.A(n_2010),
.B(n_303),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2018),
.B(n_303),
.Y(n_2597)
);

AOI21xp5_ASAP7_75t_L g2598 ( 
.A1(n_2080),
.A2(n_304),
.B(n_305),
.Y(n_2598)
);

NAND2x1p5_ASAP7_75t_L g2599 ( 
.A(n_2050),
.B(n_2041),
.Y(n_2599)
);

OAI21xp5_ASAP7_75t_L g2600 ( 
.A1(n_2088),
.A2(n_306),
.B(n_307),
.Y(n_2600)
);

OAI21xp5_ASAP7_75t_L g2601 ( 
.A1(n_2067),
.A2(n_308),
.B(n_311),
.Y(n_2601)
);

NAND3xp33_ASAP7_75t_L g2602 ( 
.A(n_2103),
.B(n_312),
.C(n_313),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2024),
.B(n_2272),
.Y(n_2603)
);

O2A1O1Ixp33_ASAP7_75t_SL g2604 ( 
.A1(n_2100),
.A2(n_2123),
.B(n_2120),
.C(n_1929),
.Y(n_2604)
);

O2A1O1Ixp33_ASAP7_75t_L g2605 ( 
.A1(n_1974),
.A2(n_317),
.B(n_315),
.C(n_316),
.Y(n_2605)
);

BUFx6f_ASAP7_75t_L g2606 ( 
.A(n_2094),
.Y(n_2606)
);

AOI21xp5_ASAP7_75t_L g2607 ( 
.A1(n_2091),
.A2(n_2095),
.B(n_2102),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2105),
.Y(n_2608)
);

BUFx6f_ASAP7_75t_L g2609 ( 
.A(n_2094),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2112),
.Y(n_2610)
);

AND2x2_ASAP7_75t_L g2611 ( 
.A(n_2074),
.B(n_318),
.Y(n_2611)
);

OAI22xp5_ASAP7_75t_L g2612 ( 
.A1(n_2510),
.A2(n_2092),
.B1(n_2164),
.B2(n_2161),
.Y(n_2612)
);

HB1xp67_ASAP7_75t_L g2613 ( 
.A(n_2338),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_L g2614 ( 
.A(n_2296),
.B(n_2439),
.Y(n_2614)
);

AOI21xp5_ASAP7_75t_L g2615 ( 
.A1(n_2299),
.A2(n_2046),
.B(n_1964),
.Y(n_2615)
);

AND2x4_ASAP7_75t_L g2616 ( 
.A(n_2473),
.B(n_2301),
.Y(n_2616)
);

NOR2x1_ASAP7_75t_L g2617 ( 
.A(n_2443),
.B(n_2129),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2292),
.Y(n_2618)
);

OAI22xp5_ASAP7_75t_L g2619 ( 
.A1(n_2590),
.A2(n_2378),
.B1(n_2392),
.B2(n_2603),
.Y(n_2619)
);

BUFx2_ASAP7_75t_L g2620 ( 
.A(n_2327),
.Y(n_2620)
);

OAI22xp5_ASAP7_75t_L g2621 ( 
.A1(n_2447),
.A2(n_2193),
.B1(n_2213),
.B2(n_2164),
.Y(n_2621)
);

CKINVDCx5p33_ASAP7_75t_R g2622 ( 
.A(n_2319),
.Y(n_2622)
);

OR2x2_ASAP7_75t_L g2623 ( 
.A(n_2358),
.B(n_2106),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2297),
.Y(n_2624)
);

INVx3_ASAP7_75t_L g2625 ( 
.A(n_2405),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_2293),
.Y(n_2626)
);

INVxp67_ASAP7_75t_L g2627 ( 
.A(n_2365),
.Y(n_2627)
);

BUFx3_ASAP7_75t_L g2628 ( 
.A(n_2319),
.Y(n_2628)
);

CKINVDCx16_ASAP7_75t_R g2629 ( 
.A(n_2336),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_SL g2630 ( 
.A(n_2301),
.B(n_2002),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2305),
.Y(n_2631)
);

BUFx6f_ASAP7_75t_L g2632 ( 
.A(n_2431),
.Y(n_2632)
);

INVx2_ASAP7_75t_L g2633 ( 
.A(n_2302),
.Y(n_2633)
);

NAND3xp33_ASAP7_75t_SL g2634 ( 
.A(n_2545),
.B(n_2157),
.C(n_2136),
.Y(n_2634)
);

O2A1O1Ixp33_ASAP7_75t_L g2635 ( 
.A1(n_2379),
.A2(n_1995),
.B(n_2077),
.C(n_2069),
.Y(n_2635)
);

OAI21xp5_ASAP7_75t_L g2636 ( 
.A1(n_2424),
.A2(n_1937),
.B(n_2065),
.Y(n_2636)
);

NOR2xp33_ASAP7_75t_L g2637 ( 
.A(n_2437),
.B(n_1944),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_SL g2638 ( 
.A(n_2301),
.B(n_2037),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_SL g2639 ( 
.A(n_2558),
.B(n_2194),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_2328),
.B(n_2195),
.Y(n_2640)
);

A2O1A1Ixp33_ASAP7_75t_L g2641 ( 
.A1(n_2455),
.A2(n_2210),
.B(n_2196),
.C(n_1972),
.Y(n_2641)
);

OAI22xp5_ASAP7_75t_L g2642 ( 
.A1(n_2518),
.A2(n_2234),
.B1(n_2250),
.B2(n_2193),
.Y(n_2642)
);

AND2x6_ASAP7_75t_L g2643 ( 
.A(n_2431),
.B(n_2035),
.Y(n_2643)
);

OAI22xp5_ASAP7_75t_SL g2644 ( 
.A1(n_2583),
.A2(n_2085),
.B1(n_1983),
.B2(n_2051),
.Y(n_2644)
);

OAI22xp5_ASAP7_75t_L g2645 ( 
.A1(n_2537),
.A2(n_2234),
.B1(n_2253),
.B2(n_2250),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2326),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2318),
.B(n_2122),
.Y(n_2647)
);

INVx5_ASAP7_75t_L g2648 ( 
.A(n_2549),
.Y(n_2648)
);

NOR2xp33_ASAP7_75t_L g2649 ( 
.A(n_2440),
.B(n_1996),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2561),
.Y(n_2650)
);

NOR2xp33_ASAP7_75t_L g2651 ( 
.A(n_2490),
.B(n_2346),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2314),
.Y(n_2652)
);

AOI21xp5_ASAP7_75t_L g2653 ( 
.A1(n_2538),
.A2(n_1939),
.B(n_2271),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_2333),
.B(n_1953),
.Y(n_2654)
);

AND2x2_ASAP7_75t_L g2655 ( 
.A(n_2313),
.B(n_2279),
.Y(n_2655)
);

BUFx6f_ASAP7_75t_L g2656 ( 
.A(n_2431),
.Y(n_2656)
);

CKINVDCx16_ASAP7_75t_R g2657 ( 
.A(n_2409),
.Y(n_2657)
);

O2A1O1Ixp33_ASAP7_75t_L g2658 ( 
.A1(n_2435),
.A2(n_1991),
.B(n_1999),
.C(n_2082),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2316),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2339),
.Y(n_2660)
);

NOR2xp33_ASAP7_75t_L g2661 ( 
.A(n_2449),
.B(n_1925),
.Y(n_2661)
);

OR2x6_ASAP7_75t_L g2662 ( 
.A(n_2549),
.B(n_2153),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_SL g2663 ( 
.A(n_2558),
.B(n_2007),
.Y(n_2663)
);

OR2x2_ASAP7_75t_L g2664 ( 
.A(n_2342),
.B(n_2038),
.Y(n_2664)
);

INVx3_ASAP7_75t_L g2665 ( 
.A(n_2332),
.Y(n_2665)
);

HB1xp67_ASAP7_75t_L g2666 ( 
.A(n_2344),
.Y(n_2666)
);

INVx3_ASAP7_75t_L g2667 ( 
.A(n_2368),
.Y(n_2667)
);

A2O1A1Ixp33_ASAP7_75t_L g2668 ( 
.A1(n_2605),
.A2(n_2033),
.B(n_2086),
.C(n_2109),
.Y(n_2668)
);

INVx2_ASAP7_75t_L g2669 ( 
.A(n_2349),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_2335),
.B(n_2089),
.Y(n_2670)
);

AOI21xp5_ASAP7_75t_L g2671 ( 
.A1(n_2325),
.A2(n_2578),
.B(n_2604),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2324),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_L g2673 ( 
.A(n_2403),
.B(n_2090),
.Y(n_2673)
);

AND2x2_ASAP7_75t_L g2674 ( 
.A(n_2356),
.B(n_318),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_L g2675 ( 
.A(n_2459),
.B(n_2017),
.Y(n_2675)
);

NAND2x1p5_ASAP7_75t_L g2676 ( 
.A(n_2300),
.B(n_2029),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_SL g2677 ( 
.A(n_2502),
.B(n_2505),
.Y(n_2677)
);

AND2x2_ASAP7_75t_L g2678 ( 
.A(n_2357),
.B(n_319),
.Y(n_2678)
);

AOI21xp5_ASAP7_75t_L g2679 ( 
.A1(n_2450),
.A2(n_319),
.B(n_320),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_SL g2680 ( 
.A(n_2502),
.B(n_320),
.Y(n_2680)
);

BUFx3_ASAP7_75t_L g2681 ( 
.A(n_2343),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_SL g2682 ( 
.A(n_2505),
.B(n_320),
.Y(n_2682)
);

NOR2xp33_ASAP7_75t_L g2683 ( 
.A(n_2586),
.B(n_2595),
.Y(n_2683)
);

AOI21xp5_ASAP7_75t_L g2684 ( 
.A1(n_2607),
.A2(n_321),
.B(n_322),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2568),
.Y(n_2685)
);

AND2x2_ASAP7_75t_L g2686 ( 
.A(n_2372),
.B(n_325),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2461),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2355),
.Y(n_2688)
);

INVx1_ASAP7_75t_SL g2689 ( 
.A(n_2402),
.Y(n_2689)
);

AOI21xp5_ASAP7_75t_L g2690 ( 
.A1(n_2413),
.A2(n_326),
.B(n_327),
.Y(n_2690)
);

INVx1_ASAP7_75t_SL g2691 ( 
.A(n_2576),
.Y(n_2691)
);

BUFx2_ASAP7_75t_L g2692 ( 
.A(n_2396),
.Y(n_2692)
);

OR2x2_ASAP7_75t_L g2693 ( 
.A(n_2364),
.B(n_331),
.Y(n_2693)
);

BUFx6f_ASAP7_75t_L g2694 ( 
.A(n_2528),
.Y(n_2694)
);

INVx2_ASAP7_75t_L g2695 ( 
.A(n_2375),
.Y(n_2695)
);

O2A1O1Ixp33_ASAP7_75t_L g2696 ( 
.A1(n_2557),
.A2(n_334),
.B(n_332),
.C(n_333),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_2477),
.B(n_332),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2506),
.Y(n_2698)
);

NOR2xp33_ASAP7_75t_L g2699 ( 
.A(n_2475),
.B(n_333),
.Y(n_2699)
);

INVx1_ASAP7_75t_SL g2700 ( 
.A(n_2585),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_L g2701 ( 
.A(n_2294),
.B(n_334),
.Y(n_2701)
);

NAND2x1p5_ASAP7_75t_L g2702 ( 
.A(n_2546),
.B(n_335),
.Y(n_2702)
);

AOI21xp5_ASAP7_75t_L g2703 ( 
.A1(n_2541),
.A2(n_336),
.B(n_337),
.Y(n_2703)
);

BUFx6f_ASAP7_75t_L g2704 ( 
.A(n_2542),
.Y(n_2704)
);

NOR2xp33_ASAP7_75t_L g2705 ( 
.A(n_2491),
.B(n_336),
.Y(n_2705)
);

AOI21xp5_ASAP7_75t_L g2706 ( 
.A1(n_2320),
.A2(n_337),
.B(n_338),
.Y(n_2706)
);

AOI21xp5_ASAP7_75t_L g2707 ( 
.A1(n_2580),
.A2(n_338),
.B(n_339),
.Y(n_2707)
);

AOI21xp5_ASAP7_75t_L g2708 ( 
.A1(n_2412),
.A2(n_2322),
.B(n_2352),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2384),
.Y(n_2709)
);

AOI21xp5_ASAP7_75t_L g2710 ( 
.A1(n_2360),
.A2(n_341),
.B(n_342),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2571),
.B(n_341),
.Y(n_2711)
);

AND2x4_ASAP7_75t_L g2712 ( 
.A(n_2388),
.B(n_342),
.Y(n_2712)
);

INVx3_ASAP7_75t_L g2713 ( 
.A(n_2552),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_2373),
.B(n_343),
.Y(n_2714)
);

INVx4_ASAP7_75t_L g2715 ( 
.A(n_2535),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_SL g2716 ( 
.A(n_2542),
.B(n_344),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_SL g2717 ( 
.A(n_2542),
.B(n_345),
.Y(n_2717)
);

INVx6_ASAP7_75t_L g2718 ( 
.A(n_2306),
.Y(n_2718)
);

INVxp67_ASAP7_75t_L g2719 ( 
.A(n_2468),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2556),
.Y(n_2720)
);

AO22x1_ASAP7_75t_L g2721 ( 
.A1(n_2468),
.A2(n_348),
.B1(n_346),
.B2(n_347),
.Y(n_2721)
);

NOR2xp33_ASAP7_75t_L g2722 ( 
.A(n_2495),
.B(n_346),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2559),
.Y(n_2723)
);

O2A1O1Ixp33_ASAP7_75t_L g2724 ( 
.A1(n_2554),
.A2(n_349),
.B(n_347),
.C(n_348),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_SL g2725 ( 
.A(n_2606),
.B(n_348),
.Y(n_2725)
);

NOR3xp33_ASAP7_75t_L g2726 ( 
.A(n_2592),
.B(n_349),
.C(n_350),
.Y(n_2726)
);

INVx1_ASAP7_75t_SL g2727 ( 
.A(n_2464),
.Y(n_2727)
);

OAI21xp5_ASAP7_75t_L g2728 ( 
.A1(n_2291),
.A2(n_349),
.B(n_350),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_L g2729 ( 
.A(n_2369),
.B(n_350),
.Y(n_2729)
);

BUFx12f_ASAP7_75t_L g2730 ( 
.A(n_2504),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_2406),
.Y(n_2731)
);

INVx2_ASAP7_75t_L g2732 ( 
.A(n_2420),
.Y(n_2732)
);

A2O1A1Ixp33_ASAP7_75t_L g2733 ( 
.A1(n_2311),
.A2(n_354),
.B(n_351),
.C(n_352),
.Y(n_2733)
);

AND2x2_ASAP7_75t_SL g2734 ( 
.A(n_2391),
.B(n_354),
.Y(n_2734)
);

BUFx3_ASAP7_75t_L g2735 ( 
.A(n_2555),
.Y(n_2735)
);

O2A1O1Ixp33_ASAP7_75t_SL g2736 ( 
.A1(n_2321),
.A2(n_357),
.B(n_355),
.C(n_356),
.Y(n_2736)
);

BUFx6f_ASAP7_75t_L g2737 ( 
.A(n_2606),
.Y(n_2737)
);

INVx5_ASAP7_75t_L g2738 ( 
.A(n_2606),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_2371),
.B(n_356),
.Y(n_2739)
);

BUFx3_ASAP7_75t_L g2740 ( 
.A(n_2428),
.Y(n_2740)
);

NOR2xp33_ASAP7_75t_L g2741 ( 
.A(n_2500),
.B(n_359),
.Y(n_2741)
);

HB1xp67_ASAP7_75t_L g2742 ( 
.A(n_2575),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_2421),
.Y(n_2743)
);

INVxp67_ASAP7_75t_SL g2744 ( 
.A(n_2527),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2389),
.B(n_360),
.Y(n_2745)
);

AOI21xp5_ASAP7_75t_L g2746 ( 
.A1(n_2395),
.A2(n_360),
.B(n_361),
.Y(n_2746)
);

NOR2xp33_ASAP7_75t_L g2747 ( 
.A(n_2596),
.B(n_2544),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2359),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_2398),
.B(n_361),
.Y(n_2749)
);

AOI21xp5_ASAP7_75t_L g2750 ( 
.A1(n_2426),
.A2(n_2456),
.B(n_2436),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2422),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2422),
.Y(n_2752)
);

OR2x6_ASAP7_75t_L g2753 ( 
.A(n_2569),
.B(n_363),
.Y(n_2753)
);

AOI21xp5_ASAP7_75t_L g2754 ( 
.A1(n_2460),
.A2(n_364),
.B(n_365),
.Y(n_2754)
);

AND2x2_ASAP7_75t_L g2755 ( 
.A(n_2611),
.B(n_364),
.Y(n_2755)
);

INVx4_ASAP7_75t_L g2756 ( 
.A(n_2609),
.Y(n_2756)
);

INVx2_ASAP7_75t_L g2757 ( 
.A(n_2467),
.Y(n_2757)
);

OAI22xp5_ASAP7_75t_L g2758 ( 
.A1(n_2423),
.A2(n_367),
.B1(n_365),
.B2(n_366),
.Y(n_2758)
);

CKINVDCx5p33_ASAP7_75t_R g2759 ( 
.A(n_2315),
.Y(n_2759)
);

NAND3xp33_ASAP7_75t_SL g2760 ( 
.A(n_2563),
.B(n_368),
.C(n_369),
.Y(n_2760)
);

O2A1O1Ixp33_ASAP7_75t_L g2761 ( 
.A1(n_2441),
.A2(n_371),
.B(n_369),
.C(n_370),
.Y(n_2761)
);

AOI21xp5_ASAP7_75t_L g2762 ( 
.A1(n_2508),
.A2(n_370),
.B(n_371),
.Y(n_2762)
);

HB1xp67_ASAP7_75t_L g2763 ( 
.A(n_2509),
.Y(n_2763)
);

AOI21xp5_ASAP7_75t_L g2764 ( 
.A1(n_2347),
.A2(n_372),
.B(n_373),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_L g2765 ( 
.A(n_2425),
.B(n_2442),
.Y(n_2765)
);

BUFx6f_ASAP7_75t_L g2766 ( 
.A(n_2331),
.Y(n_2766)
);

BUFx3_ASAP7_75t_L g2767 ( 
.A(n_2438),
.Y(n_2767)
);

NOR2xp67_ASAP7_75t_L g2768 ( 
.A(n_2308),
.B(n_374),
.Y(n_2768)
);

BUFx3_ASAP7_75t_L g2769 ( 
.A(n_2599),
.Y(n_2769)
);

AOI21xp5_ASAP7_75t_L g2770 ( 
.A1(n_2465),
.A2(n_374),
.B(n_375),
.Y(n_2770)
);

HB1xp67_ASAP7_75t_L g2771 ( 
.A(n_2529),
.Y(n_2771)
);

BUFx6f_ASAP7_75t_L g2772 ( 
.A(n_2331),
.Y(n_2772)
);

AOI21xp5_ASAP7_75t_L g2773 ( 
.A1(n_2493),
.A2(n_2524),
.B(n_2503),
.Y(n_2773)
);

NAND2xp5_ASAP7_75t_L g2774 ( 
.A(n_2463),
.B(n_377),
.Y(n_2774)
);

NOR2xp33_ASAP7_75t_L g2775 ( 
.A(n_2472),
.B(n_378),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_L g2776 ( 
.A(n_2487),
.B(n_378),
.Y(n_2776)
);

O2A1O1Ixp33_ASAP7_75t_L g2777 ( 
.A1(n_2457),
.A2(n_381),
.B(n_379),
.C(n_380),
.Y(n_2777)
);

AND2x2_ASAP7_75t_L g2778 ( 
.A(n_2562),
.B(n_379),
.Y(n_2778)
);

NOR2xp33_ASAP7_75t_L g2779 ( 
.A(n_2520),
.B(n_2530),
.Y(n_2779)
);

AOI22xp33_ASAP7_75t_L g2780 ( 
.A1(n_2587),
.A2(n_381),
.B1(n_379),
.B2(n_380),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_L g2781 ( 
.A(n_2539),
.B(n_382),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_L g2782 ( 
.A(n_2295),
.B(n_382),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_SL g2783 ( 
.A(n_2529),
.B(n_383),
.Y(n_2783)
);

AOI21xp5_ASAP7_75t_L g2784 ( 
.A1(n_2551),
.A2(n_383),
.B(n_385),
.Y(n_2784)
);

BUFx2_ASAP7_75t_L g2785 ( 
.A(n_2351),
.Y(n_2785)
);

OR2x6_ASAP7_75t_L g2786 ( 
.A(n_2451),
.B(n_386),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2410),
.Y(n_2787)
);

AO22x1_ASAP7_75t_L g2788 ( 
.A1(n_2401),
.A2(n_389),
.B1(n_387),
.B2(n_388),
.Y(n_2788)
);

AOI22xp5_ASAP7_75t_L g2789 ( 
.A1(n_2560),
.A2(n_389),
.B1(n_387),
.B2(n_388),
.Y(n_2789)
);

NOR2x1_ASAP7_75t_SL g2790 ( 
.A(n_2351),
.B(n_390),
.Y(n_2790)
);

BUFx6f_ASAP7_75t_L g2791 ( 
.A(n_2351),
.Y(n_2791)
);

NAND2x1_ASAP7_75t_L g2792 ( 
.A(n_2353),
.B(n_2366),
.Y(n_2792)
);

AOI21xp5_ASAP7_75t_L g2793 ( 
.A1(n_2317),
.A2(n_391),
.B(n_392),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2507),
.Y(n_2794)
);

AND2x4_ASAP7_75t_L g2795 ( 
.A(n_2353),
.B(n_394),
.Y(n_2795)
);

BUFx2_ASAP7_75t_L g2796 ( 
.A(n_2353),
.Y(n_2796)
);

INVx2_ASAP7_75t_L g2797 ( 
.A(n_2307),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2303),
.B(n_396),
.Y(n_2798)
);

BUFx6f_ASAP7_75t_L g2799 ( 
.A(n_2366),
.Y(n_2799)
);

AOI21xp5_ASAP7_75t_L g2800 ( 
.A1(n_2374),
.A2(n_396),
.B(n_397),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_L g2801 ( 
.A(n_2304),
.B(n_397),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_SL g2802 ( 
.A(n_2383),
.B(n_398),
.Y(n_2802)
);

BUFx6f_ASAP7_75t_L g2803 ( 
.A(n_2367),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2594),
.Y(n_2804)
);

INVx4_ASAP7_75t_L g2805 ( 
.A(n_2367),
.Y(n_2805)
);

BUFx2_ASAP7_75t_SL g2806 ( 
.A(n_2397),
.Y(n_2806)
);

AND2x2_ASAP7_75t_L g2807 ( 
.A(n_2565),
.B(n_2486),
.Y(n_2807)
);

AOI21xp5_ASAP7_75t_L g2808 ( 
.A1(n_2601),
.A2(n_400),
.B(n_401),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2553),
.Y(n_2809)
);

AOI21xp5_ASAP7_75t_L g2810 ( 
.A1(n_2600),
.A2(n_402),
.B(n_403),
.Y(n_2810)
);

OAI22xp5_ASAP7_75t_L g2811 ( 
.A1(n_2452),
.A2(n_404),
.B1(n_402),
.B2(n_403),
.Y(n_2811)
);

AND2x2_ASAP7_75t_L g2812 ( 
.A(n_2593),
.B(n_403),
.Y(n_2812)
);

OAI22xp5_ASAP7_75t_L g2813 ( 
.A1(n_2483),
.A2(n_408),
.B1(n_406),
.B2(n_407),
.Y(n_2813)
);

O2A1O1Ixp33_ASAP7_75t_SL g2814 ( 
.A1(n_2533),
.A2(n_410),
.B(n_408),
.C(n_409),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_L g2815 ( 
.A(n_2540),
.B(n_411),
.Y(n_2815)
);

OAI22xp5_ASAP7_75t_L g2816 ( 
.A1(n_2488),
.A2(n_413),
.B1(n_411),
.B2(n_412),
.Y(n_2816)
);

AOI21xp5_ASAP7_75t_L g2817 ( 
.A1(n_2608),
.A2(n_413),
.B(n_414),
.Y(n_2817)
);

INVx2_ASAP7_75t_L g2818 ( 
.A(n_2479),
.Y(n_2818)
);

INVxp67_ASAP7_75t_SL g2819 ( 
.A(n_2591),
.Y(n_2819)
);

AND2x4_ASAP7_75t_L g2820 ( 
.A(n_2429),
.B(n_415),
.Y(n_2820)
);

BUFx12f_ASAP7_75t_L g2821 ( 
.A(n_2429),
.Y(n_2821)
);

NAND2x1p5_ASAP7_75t_L g2822 ( 
.A(n_2462),
.B(n_415),
.Y(n_2822)
);

A2O1A1Ixp33_ASAP7_75t_L g2823 ( 
.A1(n_2298),
.A2(n_418),
.B(n_416),
.C(n_417),
.Y(n_2823)
);

NOR2xp33_ASAP7_75t_R g2824 ( 
.A(n_2564),
.B(n_417),
.Y(n_2824)
);

BUFx12f_ASAP7_75t_L g2825 ( 
.A(n_2458),
.Y(n_2825)
);

BUFx2_ASAP7_75t_L g2826 ( 
.A(n_2593),
.Y(n_2826)
);

CKINVDCx5p33_ASAP7_75t_R g2827 ( 
.A(n_2414),
.Y(n_2827)
);

A2O1A1Ixp33_ASAP7_75t_L g2828 ( 
.A1(n_2532),
.A2(n_421),
.B(n_419),
.C(n_420),
.Y(n_2828)
);

INVx2_ASAP7_75t_L g2829 ( 
.A(n_2610),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_2573),
.B(n_421),
.Y(n_2830)
);

OAI22xp5_ASAP7_75t_L g2831 ( 
.A1(n_2408),
.A2(n_425),
.B1(n_422),
.B2(n_424),
.Y(n_2831)
);

HB1xp67_ASAP7_75t_L g2832 ( 
.A(n_2415),
.Y(n_2832)
);

INVx2_ASAP7_75t_L g2833 ( 
.A(n_2337),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_2543),
.B(n_426),
.Y(n_2834)
);

NOR2xp33_ASAP7_75t_SL g2835 ( 
.A(n_2494),
.B(n_426),
.Y(n_2835)
);

OAI21x1_ASAP7_75t_L g2836 ( 
.A1(n_2362),
.A2(n_428),
.B(n_427),
.Y(n_2836)
);

AOI22xp33_ASAP7_75t_L g2837 ( 
.A1(n_2519),
.A2(n_429),
.B1(n_427),
.B2(n_428),
.Y(n_2837)
);

INVx2_ASAP7_75t_L g2838 ( 
.A(n_2345),
.Y(n_2838)
);

INVx3_ASAP7_75t_L g2839 ( 
.A(n_2497),
.Y(n_2839)
);

INVx2_ASAP7_75t_L g2840 ( 
.A(n_2348),
.Y(n_2840)
);

AND2x4_ASAP7_75t_SL g2841 ( 
.A(n_2432),
.B(n_429),
.Y(n_2841)
);

AOI21xp5_ASAP7_75t_L g2842 ( 
.A1(n_2330),
.A2(n_431),
.B(n_432),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_2361),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_L g2844 ( 
.A(n_2363),
.B(n_433),
.Y(n_2844)
);

INVxp67_ASAP7_75t_L g2845 ( 
.A(n_2516),
.Y(n_2845)
);

INVx1_ASAP7_75t_SL g2846 ( 
.A(n_2517),
.Y(n_2846)
);

NOR2xp67_ASAP7_75t_SL g2847 ( 
.A(n_2579),
.B(n_434),
.Y(n_2847)
);

INVx6_ASAP7_75t_L g2848 ( 
.A(n_2482),
.Y(n_2848)
);

NAND2xp5_ASAP7_75t_L g2849 ( 
.A(n_2370),
.B(n_2376),
.Y(n_2849)
);

INVx4_ASAP7_75t_L g2850 ( 
.A(n_2589),
.Y(n_2850)
);

BUFx2_ASAP7_75t_L g2851 ( 
.A(n_2525),
.Y(n_2851)
);

NAND2xp33_ASAP7_75t_SL g2852 ( 
.A(n_2427),
.B(n_435),
.Y(n_2852)
);

O2A1O1Ixp5_ASAP7_75t_SL g2853 ( 
.A1(n_2411),
.A2(n_657),
.B(n_658),
.C(n_656),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_SL g2854 ( 
.A(n_2448),
.B(n_2323),
.Y(n_2854)
);

NAND2xp33_ASAP7_75t_SL g2855 ( 
.A(n_2446),
.B(n_436),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_SL g2856 ( 
.A(n_2340),
.B(n_437),
.Y(n_2856)
);

AOI21xp5_ASAP7_75t_L g2857 ( 
.A1(n_2469),
.A2(n_2382),
.B(n_2381),
.Y(n_2857)
);

INVx3_ASAP7_75t_L g2858 ( 
.A(n_2466),
.Y(n_2858)
);

INVx2_ASAP7_75t_L g2859 ( 
.A(n_2387),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_L g2860 ( 
.A(n_2390),
.B(n_438),
.Y(n_2860)
);

OAI21xp5_ASAP7_75t_L g2861 ( 
.A1(n_2481),
.A2(n_439),
.B(n_440),
.Y(n_2861)
);

INVx2_ASAP7_75t_L g2862 ( 
.A(n_2394),
.Y(n_2862)
);

NAND3xp33_ASAP7_75t_SL g2863 ( 
.A(n_2385),
.B(n_442),
.C(n_443),
.Y(n_2863)
);

AND2x2_ASAP7_75t_L g2864 ( 
.A(n_2531),
.B(n_442),
.Y(n_2864)
);

NAND2xp5_ASAP7_75t_SL g2865 ( 
.A(n_2496),
.B(n_442),
.Y(n_2865)
);

BUFx2_ASAP7_75t_L g2866 ( 
.A(n_2534),
.Y(n_2866)
);

O2A1O1Ixp5_ASAP7_75t_L g2867 ( 
.A1(n_2570),
.A2(n_445),
.B(n_443),
.C(n_444),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2400),
.B(n_444),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_L g2869 ( 
.A(n_2404),
.B(n_445),
.Y(n_2869)
);

AOI22xp5_ASAP7_75t_L g2870 ( 
.A1(n_2501),
.A2(n_448),
.B1(n_446),
.B2(n_447),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_L g2871 ( 
.A(n_2407),
.B(n_446),
.Y(n_2871)
);

OR2x6_ASAP7_75t_L g2872 ( 
.A(n_2521),
.B(n_447),
.Y(n_2872)
);

BUFx2_ASAP7_75t_L g2873 ( 
.A(n_2416),
.Y(n_2873)
);

NAND2x1p5_ASAP7_75t_L g2874 ( 
.A(n_2377),
.B(n_448),
.Y(n_2874)
);

INVx2_ASAP7_75t_SL g2875 ( 
.A(n_2547),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_SL g2876 ( 
.A(n_2536),
.B(n_449),
.Y(n_2876)
);

INVx2_ASAP7_75t_L g2877 ( 
.A(n_2434),
.Y(n_2877)
);

OAI21x1_ASAP7_75t_L g2878 ( 
.A1(n_2310),
.A2(n_451),
.B(n_450),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_SL g2879 ( 
.A(n_2515),
.B(n_449),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2453),
.Y(n_2880)
);

NOR2xp33_ASAP7_75t_L g2881 ( 
.A(n_2566),
.B(n_450),
.Y(n_2881)
);

INVx3_ASAP7_75t_L g2882 ( 
.A(n_2454),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2470),
.B(n_452),
.Y(n_2883)
);

NOR2xp33_ASAP7_75t_L g2884 ( 
.A(n_2567),
.B(n_452),
.Y(n_2884)
);

AOI21xp5_ASAP7_75t_L g2885 ( 
.A1(n_2386),
.A2(n_453),
.B(n_454),
.Y(n_2885)
);

HB1xp67_ASAP7_75t_L g2886 ( 
.A(n_2476),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_L g2887 ( 
.A(n_2484),
.B(n_453),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2485),
.B(n_454),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2492),
.Y(n_2889)
);

AOI21x1_ASAP7_75t_L g2890 ( 
.A1(n_2597),
.A2(n_659),
.B(n_658),
.Y(n_2890)
);

AND2x2_ASAP7_75t_L g2891 ( 
.A(n_2574),
.B(n_455),
.Y(n_2891)
);

AND2x4_ASAP7_75t_L g2892 ( 
.A(n_2550),
.B(n_458),
.Y(n_2892)
);

INVx2_ASAP7_75t_L g2893 ( 
.A(n_2312),
.Y(n_2893)
);

INVxp67_ASAP7_75t_L g2894 ( 
.A(n_2380),
.Y(n_2894)
);

OR2x6_ASAP7_75t_L g2895 ( 
.A(n_2471),
.B(n_459),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2312),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2312),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_2393),
.B(n_460),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2511),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2512),
.Y(n_2900)
);

A2O1A1Ixp33_ASAP7_75t_L g2901 ( 
.A1(n_2399),
.A2(n_465),
.B(n_461),
.C(n_464),
.Y(n_2901)
);

BUFx6f_ASAP7_75t_L g2902 ( 
.A(n_2602),
.Y(n_2902)
);

AND2x2_ASAP7_75t_L g2903 ( 
.A(n_2474),
.B(n_468),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2478),
.B(n_470),
.Y(n_2904)
);

HB1xp67_ASAP7_75t_L g2905 ( 
.A(n_2513),
.Y(n_2905)
);

INVx2_ASAP7_75t_SL g2906 ( 
.A(n_2514),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2480),
.B(n_471),
.Y(n_2907)
);

BUFx6f_ASAP7_75t_L g2908 ( 
.A(n_2419),
.Y(n_2908)
);

NAND2xp5_ASAP7_75t_L g2909 ( 
.A(n_2489),
.B(n_472),
.Y(n_2909)
);

AOI21xp5_ASAP7_75t_L g2910 ( 
.A1(n_2309),
.A2(n_473),
.B(n_474),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_L g2911 ( 
.A(n_2498),
.B(n_475),
.Y(n_2911)
);

A2O1A1Ixp33_ASAP7_75t_L g2912 ( 
.A1(n_2581),
.A2(n_2584),
.B(n_2588),
.C(n_2582),
.Y(n_2912)
);

INVx2_ASAP7_75t_L g2913 ( 
.A(n_2522),
.Y(n_2913)
);

INVx3_ASAP7_75t_L g2914 ( 
.A(n_2499),
.Y(n_2914)
);

AOI21xp5_ASAP7_75t_L g2915 ( 
.A1(n_2334),
.A2(n_476),
.B(n_477),
.Y(n_2915)
);

NAND2x1p5_ASAP7_75t_L g2916 ( 
.A(n_2523),
.B(n_478),
.Y(n_2916)
);

OAI21xp33_ASAP7_75t_L g2917 ( 
.A1(n_2548),
.A2(n_478),
.B(n_479),
.Y(n_2917)
);

INVx2_ASAP7_75t_L g2918 ( 
.A(n_2526),
.Y(n_2918)
);

CKINVDCx8_ASAP7_75t_R g2919 ( 
.A(n_2417),
.Y(n_2919)
);

INVx2_ASAP7_75t_L g2920 ( 
.A(n_2341),
.Y(n_2920)
);

AOI21xp5_ASAP7_75t_L g2921 ( 
.A1(n_2329),
.A2(n_480),
.B(n_482),
.Y(n_2921)
);

OAI22xp5_ASAP7_75t_L g2922 ( 
.A1(n_2572),
.A2(n_485),
.B1(n_483),
.B2(n_484),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_2418),
.B(n_483),
.Y(n_2923)
);

AND2x4_ASAP7_75t_L g2924 ( 
.A(n_2350),
.B(n_483),
.Y(n_2924)
);

BUFx2_ASAP7_75t_L g2925 ( 
.A(n_2354),
.Y(n_2925)
);

INVx3_ASAP7_75t_L g2926 ( 
.A(n_2577),
.Y(n_2926)
);

OR2x6_ASAP7_75t_L g2927 ( 
.A(n_2433),
.B(n_484),
.Y(n_2927)
);

BUFx6f_ASAP7_75t_L g2928 ( 
.A(n_2598),
.Y(n_2928)
);

INVx2_ASAP7_75t_L g2929 ( 
.A(n_2430),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_SL g2930 ( 
.A(n_2444),
.B(n_486),
.Y(n_2930)
);

NAND2xp5_ASAP7_75t_SL g2931 ( 
.A(n_2445),
.B(n_487),
.Y(n_2931)
);

AND2x4_ASAP7_75t_L g2932 ( 
.A(n_2473),
.B(n_489),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_L g2933 ( 
.A(n_2296),
.B(n_491),
.Y(n_2933)
);

BUFx6f_ASAP7_75t_L g2934 ( 
.A(n_2431),
.Y(n_2934)
);

INVx3_ASAP7_75t_L g2935 ( 
.A(n_2628),
.Y(n_2935)
);

AND2x4_ASAP7_75t_L g2936 ( 
.A(n_2617),
.B(n_492),
.Y(n_2936)
);

CKINVDCx5p33_ASAP7_75t_R g2937 ( 
.A(n_2622),
.Y(n_2937)
);

BUFx2_ASAP7_75t_SL g2938 ( 
.A(n_2648),
.Y(n_2938)
);

CKINVDCx8_ASAP7_75t_R g2939 ( 
.A(n_2629),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2618),
.Y(n_2940)
);

BUFx6f_ASAP7_75t_L g2941 ( 
.A(n_2821),
.Y(n_2941)
);

INVx3_ASAP7_75t_SL g2942 ( 
.A(n_2715),
.Y(n_2942)
);

BUFx3_ASAP7_75t_L g2943 ( 
.A(n_2735),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2624),
.Y(n_2944)
);

BUFx3_ASAP7_75t_L g2945 ( 
.A(n_2715),
.Y(n_2945)
);

AOI22xp33_ASAP7_75t_L g2946 ( 
.A1(n_2619),
.A2(n_493),
.B1(n_491),
.B2(n_492),
.Y(n_2946)
);

BUFx3_ASAP7_75t_L g2947 ( 
.A(n_2681),
.Y(n_2947)
);

BUFx3_ASAP7_75t_L g2948 ( 
.A(n_2662),
.Y(n_2948)
);

INVx3_ASAP7_75t_L g2949 ( 
.A(n_2769),
.Y(n_2949)
);

BUFx6f_ASAP7_75t_L g2950 ( 
.A(n_2766),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2631),
.Y(n_2951)
);

CKINVDCx5p33_ASAP7_75t_R g2952 ( 
.A(n_2730),
.Y(n_2952)
);

INVx8_ASAP7_75t_L g2953 ( 
.A(n_2753),
.Y(n_2953)
);

INVx4_ASAP7_75t_L g2954 ( 
.A(n_2665),
.Y(n_2954)
);

BUFx3_ASAP7_75t_L g2955 ( 
.A(n_2667),
.Y(n_2955)
);

BUFx12f_ASAP7_75t_L g2956 ( 
.A(n_2759),
.Y(n_2956)
);

CKINVDCx20_ASAP7_75t_R g2957 ( 
.A(n_2689),
.Y(n_2957)
);

INVx6_ASAP7_75t_SL g2958 ( 
.A(n_2786),
.Y(n_2958)
);

INVx5_ASAP7_75t_L g2959 ( 
.A(n_2625),
.Y(n_2959)
);

BUFx2_ASAP7_75t_L g2960 ( 
.A(n_2627),
.Y(n_2960)
);

HB1xp67_ASAP7_75t_L g2961 ( 
.A(n_2666),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2646),
.Y(n_2962)
);

INVx5_ASAP7_75t_L g2963 ( 
.A(n_2657),
.Y(n_2963)
);

CKINVDCx11_ASAP7_75t_R g2964 ( 
.A(n_2691),
.Y(n_2964)
);

BUFx3_ASAP7_75t_L g2965 ( 
.A(n_2692),
.Y(n_2965)
);

INVx1_ASAP7_75t_SL g2966 ( 
.A(n_2727),
.Y(n_2966)
);

OR2x2_ASAP7_75t_L g2967 ( 
.A(n_2807),
.B(n_493),
.Y(n_2967)
);

BUFx4_ASAP7_75t_SL g2968 ( 
.A(n_2786),
.Y(n_2968)
);

INVxp67_ASAP7_75t_SL g2969 ( 
.A(n_2744),
.Y(n_2969)
);

INVx8_ASAP7_75t_L g2970 ( 
.A(n_2825),
.Y(n_2970)
);

INVx1_ASAP7_75t_SL g2971 ( 
.A(n_2700),
.Y(n_2971)
);

INVx2_ASAP7_75t_L g2972 ( 
.A(n_2626),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2650),
.Y(n_2973)
);

BUFx4f_ASAP7_75t_L g2974 ( 
.A(n_2702),
.Y(n_2974)
);

INVx6_ASAP7_75t_L g2975 ( 
.A(n_2718),
.Y(n_2975)
);

BUFx2_ASAP7_75t_SL g2976 ( 
.A(n_2768),
.Y(n_2976)
);

AND2x2_ASAP7_75t_L g2977 ( 
.A(n_2655),
.B(n_493),
.Y(n_2977)
);

BUFx6f_ASAP7_75t_L g2978 ( 
.A(n_2772),
.Y(n_2978)
);

BUFx2_ASAP7_75t_L g2979 ( 
.A(n_2805),
.Y(n_2979)
);

BUFx6f_ASAP7_75t_L g2980 ( 
.A(n_2772),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2660),
.Y(n_2981)
);

AOI22xp33_ASAP7_75t_L g2982 ( 
.A1(n_2734),
.A2(n_497),
.B1(n_494),
.B2(n_496),
.Y(n_2982)
);

BUFx6f_ASAP7_75t_L g2983 ( 
.A(n_2772),
.Y(n_2983)
);

AND2x2_ASAP7_75t_L g2984 ( 
.A(n_2896),
.B(n_496),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2720),
.Y(n_2985)
);

INVx4_ASAP7_75t_L g2986 ( 
.A(n_2718),
.Y(n_2986)
);

INVx6_ASAP7_75t_L g2987 ( 
.A(n_2805),
.Y(n_2987)
);

INVx6_ASAP7_75t_SL g2988 ( 
.A(n_2932),
.Y(n_2988)
);

BUFx2_ASAP7_75t_SL g2989 ( 
.A(n_2616),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2723),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2685),
.Y(n_2991)
);

BUFx3_ASAP7_75t_L g2992 ( 
.A(n_2740),
.Y(n_2992)
);

INVx2_ASAP7_75t_L g2993 ( 
.A(n_2633),
.Y(n_2993)
);

BUFx3_ASAP7_75t_L g2994 ( 
.A(n_2767),
.Y(n_2994)
);

INVx2_ASAP7_75t_L g2995 ( 
.A(n_2652),
.Y(n_2995)
);

CKINVDCx8_ASAP7_75t_R g2996 ( 
.A(n_2806),
.Y(n_2996)
);

BUFx12f_ASAP7_75t_L g2997 ( 
.A(n_2676),
.Y(n_2997)
);

BUFx2_ASAP7_75t_SL g2998 ( 
.A(n_2616),
.Y(n_2998)
);

INVx3_ASAP7_75t_L g2999 ( 
.A(n_2713),
.Y(n_2999)
);

INVx2_ASAP7_75t_L g3000 ( 
.A(n_2659),
.Y(n_3000)
);

INVx1_ASAP7_75t_SL g3001 ( 
.A(n_2623),
.Y(n_3001)
);

BUFx2_ASAP7_75t_L g3002 ( 
.A(n_2643),
.Y(n_3002)
);

AND2x4_ASAP7_75t_L g3003 ( 
.A(n_2719),
.B(n_500),
.Y(n_3003)
);

INVx5_ASAP7_75t_L g3004 ( 
.A(n_2791),
.Y(n_3004)
);

INVx1_ASAP7_75t_SL g3005 ( 
.A(n_2664),
.Y(n_3005)
);

INVx5_ASAP7_75t_SL g3006 ( 
.A(n_2872),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2672),
.B(n_499),
.Y(n_3007)
);

NAND2x1p5_ASAP7_75t_L g3008 ( 
.A(n_2738),
.B(n_499),
.Y(n_3008)
);

INVx1_ASAP7_75t_SL g3009 ( 
.A(n_2620),
.Y(n_3009)
);

INVx6_ASAP7_75t_L g3010 ( 
.A(n_2738),
.Y(n_3010)
);

INVx2_ASAP7_75t_L g3011 ( 
.A(n_2669),
.Y(n_3011)
);

BUFx6f_ASAP7_75t_SL g3012 ( 
.A(n_2795),
.Y(n_3012)
);

AND2x2_ASAP7_75t_L g3013 ( 
.A(n_2763),
.B(n_501),
.Y(n_3013)
);

BUFx2_ASAP7_75t_SL g3014 ( 
.A(n_2643),
.Y(n_3014)
);

BUFx6f_ASAP7_75t_L g3015 ( 
.A(n_2791),
.Y(n_3015)
);

BUFx3_ASAP7_75t_L g3016 ( 
.A(n_2649),
.Y(n_3016)
);

INVx5_ASAP7_75t_L g3017 ( 
.A(n_2791),
.Y(n_3017)
);

INVx2_ASAP7_75t_SL g3018 ( 
.A(n_2742),
.Y(n_3018)
);

INVx6_ASAP7_75t_L g3019 ( 
.A(n_2756),
.Y(n_3019)
);

BUFx12f_ASAP7_75t_L g3020 ( 
.A(n_2827),
.Y(n_3020)
);

INVx1_ASAP7_75t_SL g3021 ( 
.A(n_2785),
.Y(n_3021)
);

AND2x2_ASAP7_75t_L g3022 ( 
.A(n_2893),
.B(n_501),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2687),
.Y(n_3023)
);

INVx2_ASAP7_75t_SL g3024 ( 
.A(n_2613),
.Y(n_3024)
);

BUFx12f_ASAP7_75t_L g3025 ( 
.A(n_2693),
.Y(n_3025)
);

BUFx4f_ASAP7_75t_SL g3026 ( 
.A(n_2643),
.Y(n_3026)
);

HB1xp67_ASAP7_75t_L g3027 ( 
.A(n_2771),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2698),
.B(n_501),
.Y(n_3028)
);

BUFx2_ASAP7_75t_R g3029 ( 
.A(n_2614),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2688),
.Y(n_3030)
);

INVx1_ASAP7_75t_SL g3031 ( 
.A(n_2796),
.Y(n_3031)
);

BUFx12f_ASAP7_75t_L g3032 ( 
.A(n_2820),
.Y(n_3032)
);

INVx1_ASAP7_75t_SL g3033 ( 
.A(n_2683),
.Y(n_3033)
);

BUFx6f_ASAP7_75t_SL g3034 ( 
.A(n_2820),
.Y(n_3034)
);

INVx1_ASAP7_75t_SL g3035 ( 
.A(n_2826),
.Y(n_3035)
);

BUFx2_ASAP7_75t_SL g3036 ( 
.A(n_2643),
.Y(n_3036)
);

BUFx3_ASAP7_75t_L g3037 ( 
.A(n_2661),
.Y(n_3037)
);

CKINVDCx5p33_ASAP7_75t_R g3038 ( 
.A(n_2637),
.Y(n_3038)
);

BUFx3_ASAP7_75t_L g3039 ( 
.A(n_2651),
.Y(n_3039)
);

BUFx6f_ASAP7_75t_L g3040 ( 
.A(n_2799),
.Y(n_3040)
);

INVx2_ASAP7_75t_L g3041 ( 
.A(n_2695),
.Y(n_3041)
);

OR2x6_ASAP7_75t_L g3042 ( 
.A(n_2721),
.B(n_503),
.Y(n_3042)
);

CKINVDCx5p33_ASAP7_75t_R g3043 ( 
.A(n_2644),
.Y(n_3043)
);

BUFx8_ASAP7_75t_L g3044 ( 
.A(n_2812),
.Y(n_3044)
);

BUFx8_ASAP7_75t_L g3045 ( 
.A(n_2778),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_L g3046 ( 
.A(n_2809),
.B(n_503),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2709),
.Y(n_3047)
);

AND2x2_ASAP7_75t_L g3048 ( 
.A(n_2897),
.B(n_504),
.Y(n_3048)
);

INVx2_ASAP7_75t_L g3049 ( 
.A(n_2731),
.Y(n_3049)
);

BUFx5_ASAP7_75t_L g3050 ( 
.A(n_2899),
.Y(n_3050)
);

INVx4_ASAP7_75t_L g3051 ( 
.A(n_2799),
.Y(n_3051)
);

BUFx10_ASAP7_75t_L g3052 ( 
.A(n_2699),
.Y(n_3052)
);

OR2x6_ASAP7_75t_L g3053 ( 
.A(n_2788),
.B(n_504),
.Y(n_3053)
);

BUFx3_ASAP7_75t_L g3054 ( 
.A(n_2792),
.Y(n_3054)
);

INVx4_ASAP7_75t_L g3055 ( 
.A(n_2799),
.Y(n_3055)
);

INVx1_ASAP7_75t_SL g3056 ( 
.A(n_2803),
.Y(n_3056)
);

BUFx8_ASAP7_75t_L g3057 ( 
.A(n_2755),
.Y(n_3057)
);

BUFx12f_ASAP7_75t_L g3058 ( 
.A(n_2803),
.Y(n_3058)
);

BUFx6f_ASAP7_75t_L g3059 ( 
.A(n_2803),
.Y(n_3059)
);

BUFx12f_ASAP7_75t_L g3060 ( 
.A(n_2851),
.Y(n_3060)
);

AOI22xp33_ASAP7_75t_L g3061 ( 
.A1(n_2612),
.A2(n_507),
.B1(n_505),
.B2(n_506),
.Y(n_3061)
);

CKINVDCx5p33_ASAP7_75t_R g3062 ( 
.A(n_2705),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2732),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2743),
.Y(n_3064)
);

CKINVDCx5p33_ASAP7_75t_R g3065 ( 
.A(n_2722),
.Y(n_3065)
);

INVx2_ASAP7_75t_SL g3066 ( 
.A(n_2757),
.Y(n_3066)
);

BUFx3_ASAP7_75t_L g3067 ( 
.A(n_2632),
.Y(n_3067)
);

INVx2_ASAP7_75t_SL g3068 ( 
.A(n_2663),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2670),
.Y(n_3069)
);

INVxp67_ASAP7_75t_SL g3070 ( 
.A(n_2839),
.Y(n_3070)
);

BUFx3_ASAP7_75t_L g3071 ( 
.A(n_2656),
.Y(n_3071)
);

CKINVDCx11_ASAP7_75t_R g3072 ( 
.A(n_2919),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2673),
.Y(n_3073)
);

AND2x2_ASAP7_75t_L g3074 ( 
.A(n_2674),
.B(n_507),
.Y(n_3074)
);

BUFx5_ASAP7_75t_L g3075 ( 
.A(n_2900),
.Y(n_3075)
);

INVxp67_ASAP7_75t_SL g3076 ( 
.A(n_2712),
.Y(n_3076)
);

BUFx4f_ASAP7_75t_SL g3077 ( 
.A(n_2630),
.Y(n_3077)
);

BUFx12f_ASAP7_75t_L g3078 ( 
.A(n_2866),
.Y(n_3078)
);

HB1xp67_ASAP7_75t_L g3079 ( 
.A(n_2748),
.Y(n_3079)
);

INVx1_ASAP7_75t_SL g3080 ( 
.A(n_2846),
.Y(n_3080)
);

INVx1_ASAP7_75t_SL g3081 ( 
.A(n_2714),
.Y(n_3081)
);

INVx3_ASAP7_75t_L g3082 ( 
.A(n_2656),
.Y(n_3082)
);

BUFx3_ASAP7_75t_L g3083 ( 
.A(n_2694),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2829),
.Y(n_3084)
);

INVxp33_ASAP7_75t_L g3085 ( 
.A(n_2741),
.Y(n_3085)
);

CKINVDCx20_ASAP7_75t_R g3086 ( 
.A(n_2832),
.Y(n_3086)
);

OR2x6_ASAP7_75t_L g3087 ( 
.A(n_2653),
.B(n_509),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2765),
.Y(n_3088)
);

INVx3_ASAP7_75t_L g3089 ( 
.A(n_2694),
.Y(n_3089)
);

HB1xp67_ASAP7_75t_L g3090 ( 
.A(n_2751),
.Y(n_3090)
);

BUFx12f_ASAP7_75t_L g3091 ( 
.A(n_2873),
.Y(n_3091)
);

BUFx6f_ASAP7_75t_L g3092 ( 
.A(n_2704),
.Y(n_3092)
);

BUFx6f_ASAP7_75t_L g3093 ( 
.A(n_2704),
.Y(n_3093)
);

INVx2_ASAP7_75t_L g3094 ( 
.A(n_2833),
.Y(n_3094)
);

AND2x2_ASAP7_75t_L g3095 ( 
.A(n_2678),
.B(n_511),
.Y(n_3095)
);

BUFx3_ASAP7_75t_L g3096 ( 
.A(n_2704),
.Y(n_3096)
);

BUFx8_ASAP7_75t_L g3097 ( 
.A(n_2686),
.Y(n_3097)
);

BUFx3_ASAP7_75t_L g3098 ( 
.A(n_2737),
.Y(n_3098)
);

BUFx2_ASAP7_75t_SL g3099 ( 
.A(n_2638),
.Y(n_3099)
);

BUFx3_ASAP7_75t_L g3100 ( 
.A(n_2737),
.Y(n_3100)
);

INVx4_ASAP7_75t_L g3101 ( 
.A(n_2737),
.Y(n_3101)
);

BUFx2_ASAP7_75t_R g3102 ( 
.A(n_2640),
.Y(n_3102)
);

BUFx3_ASAP7_75t_L g3103 ( 
.A(n_2934),
.Y(n_3103)
);

BUFx6f_ASAP7_75t_L g3104 ( 
.A(n_2934),
.Y(n_3104)
);

CKINVDCx20_ASAP7_75t_R g3105 ( 
.A(n_2647),
.Y(n_3105)
);

AND2x2_ASAP7_75t_L g3106 ( 
.A(n_2838),
.B(n_512),
.Y(n_3106)
);

CKINVDCx16_ASAP7_75t_R g3107 ( 
.A(n_2835),
.Y(n_3107)
);

BUFx6f_ASAP7_75t_L g3108 ( 
.A(n_2934),
.Y(n_3108)
);

INVx2_ASAP7_75t_L g3109 ( 
.A(n_2840),
.Y(n_3109)
);

BUFx12f_ASAP7_75t_L g3110 ( 
.A(n_2875),
.Y(n_3110)
);

BUFx2_ASAP7_75t_L g3111 ( 
.A(n_2752),
.Y(n_3111)
);

INVxp67_ASAP7_75t_SL g3112 ( 
.A(n_2819),
.Y(n_3112)
);

AND2x2_ASAP7_75t_L g3113 ( 
.A(n_2843),
.B(n_512),
.Y(n_3113)
);

BUFx6f_ASAP7_75t_L g3114 ( 
.A(n_2677),
.Y(n_3114)
);

INVx2_ASAP7_75t_SL g3115 ( 
.A(n_2639),
.Y(n_3115)
);

INVxp67_ASAP7_75t_SL g3116 ( 
.A(n_2783),
.Y(n_3116)
);

CKINVDCx11_ASAP7_75t_R g3117 ( 
.A(n_2794),
.Y(n_3117)
);

INVx4_ASAP7_75t_L g3118 ( 
.A(n_2841),
.Y(n_3118)
);

INVxp67_ASAP7_75t_SL g3119 ( 
.A(n_2886),
.Y(n_3119)
);

INVx3_ASAP7_75t_L g3120 ( 
.A(n_2848),
.Y(n_3120)
);

INVx2_ASAP7_75t_L g3121 ( 
.A(n_2859),
.Y(n_3121)
);

BUFx6f_ASAP7_75t_L g3122 ( 
.A(n_2675),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_2711),
.Y(n_3123)
);

BUFx3_ASAP7_75t_L g3124 ( 
.A(n_2864),
.Y(n_3124)
);

BUFx6f_ASAP7_75t_L g3125 ( 
.A(n_2908),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2779),
.Y(n_3126)
);

BUFx12f_ASAP7_75t_L g3127 ( 
.A(n_2874),
.Y(n_3127)
);

BUFx6f_ASAP7_75t_L g3128 ( 
.A(n_2908),
.Y(n_3128)
);

BUFx2_ASAP7_75t_L g3129 ( 
.A(n_2824),
.Y(n_3129)
);

INVx5_ASAP7_75t_SL g3130 ( 
.A(n_2895),
.Y(n_3130)
);

BUFx3_ASAP7_75t_L g3131 ( 
.A(n_2747),
.Y(n_3131)
);

BUFx6f_ASAP7_75t_L g3132 ( 
.A(n_2908),
.Y(n_3132)
);

INVx2_ASAP7_75t_L g3133 ( 
.A(n_2862),
.Y(n_3133)
);

AOI22xp33_ASAP7_75t_L g3134 ( 
.A1(n_2852),
.A2(n_515),
.B1(n_513),
.B2(n_514),
.Y(n_3134)
);

INVx2_ASAP7_75t_SL g3135 ( 
.A(n_2933),
.Y(n_3135)
);

HB1xp67_ASAP7_75t_L g3136 ( 
.A(n_2621),
.Y(n_3136)
);

INVx2_ASAP7_75t_SL g3137 ( 
.A(n_2892),
.Y(n_3137)
);

INVxp67_ASAP7_75t_SL g3138 ( 
.A(n_2858),
.Y(n_3138)
);

INVx8_ASAP7_75t_L g3139 ( 
.A(n_2895),
.Y(n_3139)
);

INVx2_ASAP7_75t_L g3140 ( 
.A(n_2877),
.Y(n_3140)
);

BUFx12f_ASAP7_75t_L g3141 ( 
.A(n_2924),
.Y(n_3141)
);

BUFx3_ASAP7_75t_L g3142 ( 
.A(n_2924),
.Y(n_3142)
);

BUFx3_ASAP7_75t_L g3143 ( 
.A(n_2822),
.Y(n_3143)
);

INVx3_ASAP7_75t_L g3144 ( 
.A(n_2927),
.Y(n_3144)
);

AND2x2_ASAP7_75t_L g3145 ( 
.A(n_2850),
.B(n_2880),
.Y(n_3145)
);

INVx6_ASAP7_75t_SL g3146 ( 
.A(n_2790),
.Y(n_3146)
);

BUFx4_ASAP7_75t_R g3147 ( 
.A(n_2818),
.Y(n_3147)
);

AND2x2_ASAP7_75t_L g3148 ( 
.A(n_2850),
.B(n_2889),
.Y(n_3148)
);

INVx5_ASAP7_75t_L g3149 ( 
.A(n_2882),
.Y(n_3149)
);

BUFx2_ASAP7_75t_L g3150 ( 
.A(n_2641),
.Y(n_3150)
);

INVx1_ASAP7_75t_L g3151 ( 
.A(n_2750),
.Y(n_3151)
);

BUFx3_ASAP7_75t_L g3152 ( 
.A(n_2697),
.Y(n_3152)
);

INVx1_ASAP7_75t_SL g3153 ( 
.A(n_2654),
.Y(n_3153)
);

INVx2_ASAP7_75t_SL g3154 ( 
.A(n_2802),
.Y(n_3154)
);

BUFx3_ASAP7_75t_L g3155 ( 
.A(n_2836),
.Y(n_3155)
);

BUFx3_ASAP7_75t_L g3156 ( 
.A(n_2916),
.Y(n_3156)
);

INVx2_ASAP7_75t_SL g3157 ( 
.A(n_2680),
.Y(n_3157)
);

INVx3_ASAP7_75t_SL g3158 ( 
.A(n_2682),
.Y(n_3158)
);

BUFx2_ASAP7_75t_L g3159 ( 
.A(n_2845),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_2729),
.Y(n_3160)
);

INVx3_ASAP7_75t_L g3161 ( 
.A(n_2890),
.Y(n_3161)
);

BUFx2_ASAP7_75t_L g3162 ( 
.A(n_2636),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_L g3163 ( 
.A(n_2642),
.B(n_516),
.Y(n_3163)
);

BUFx3_ASAP7_75t_L g3164 ( 
.A(n_2891),
.Y(n_3164)
);

BUFx6f_ASAP7_75t_L g3165 ( 
.A(n_2928),
.Y(n_3165)
);

BUFx6f_ASAP7_75t_L g3166 ( 
.A(n_2928),
.Y(n_3166)
);

INVx4_ASAP7_75t_L g3167 ( 
.A(n_2902),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_2645),
.B(n_519),
.Y(n_3168)
);

NAND2x1p5_ASAP7_75t_L g3169 ( 
.A(n_2847),
.B(n_519),
.Y(n_3169)
);

AND2x2_ASAP7_75t_L g3170 ( 
.A(n_2787),
.B(n_519),
.Y(n_3170)
);

OR2x2_ASAP7_75t_L g3171 ( 
.A(n_2849),
.B(n_520),
.Y(n_3171)
);

BUFx6f_ASAP7_75t_L g3172 ( 
.A(n_2902),
.Y(n_3172)
);

AOI22xp33_ASAP7_75t_L g3173 ( 
.A1(n_2855),
.A2(n_522),
.B1(n_520),
.B2(n_521),
.Y(n_3173)
);

INVx5_ASAP7_75t_L g3174 ( 
.A(n_2903),
.Y(n_3174)
);

INVxp67_ASAP7_75t_SL g3175 ( 
.A(n_2797),
.Y(n_3175)
);

OR2x2_ASAP7_75t_L g3176 ( 
.A(n_2782),
.B(n_521),
.Y(n_3176)
);

INVx1_ASAP7_75t_L g3177 ( 
.A(n_2739),
.Y(n_3177)
);

INVxp67_ASAP7_75t_SL g3178 ( 
.A(n_2905),
.Y(n_3178)
);

BUFx8_ASAP7_75t_L g3179 ( 
.A(n_2925),
.Y(n_3179)
);

INVx3_ASAP7_75t_SL g3180 ( 
.A(n_2716),
.Y(n_3180)
);

BUFx3_ASAP7_75t_L g3181 ( 
.A(n_2745),
.Y(n_3181)
);

INVx1_ASAP7_75t_SL g3182 ( 
.A(n_2717),
.Y(n_3182)
);

BUFx3_ASAP7_75t_L g3183 ( 
.A(n_2749),
.Y(n_3183)
);

BUFx3_ASAP7_75t_L g3184 ( 
.A(n_2774),
.Y(n_3184)
);

BUFx2_ASAP7_75t_R g3185 ( 
.A(n_2701),
.Y(n_3185)
);

INVx2_ASAP7_75t_SL g3186 ( 
.A(n_2725),
.Y(n_3186)
);

INVx4_ASAP7_75t_L g3187 ( 
.A(n_2914),
.Y(n_3187)
);

BUFx2_ASAP7_75t_L g3188 ( 
.A(n_2894),
.Y(n_3188)
);

BUFx4_ASAP7_75t_SL g3189 ( 
.A(n_2634),
.Y(n_3189)
);

BUFx6f_ASAP7_75t_L g3190 ( 
.A(n_2898),
.Y(n_3190)
);

INVx2_ASAP7_75t_L g3191 ( 
.A(n_2878),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_2776),
.Y(n_3192)
);

BUFx2_ASAP7_75t_SL g3193 ( 
.A(n_2758),
.Y(n_3193)
);

BUFx3_ASAP7_75t_L g3194 ( 
.A(n_2781),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_2865),
.Y(n_3195)
);

INVx3_ASAP7_75t_L g3196 ( 
.A(n_2926),
.Y(n_3196)
);

INVx2_ASAP7_75t_L g3197 ( 
.A(n_2913),
.Y(n_3197)
);

CKINVDCx6p67_ASAP7_75t_R g3198 ( 
.A(n_2876),
.Y(n_3198)
);

INVx4_ASAP7_75t_L g3199 ( 
.A(n_2906),
.Y(n_3199)
);

INVx2_ASAP7_75t_SL g3200 ( 
.A(n_2834),
.Y(n_3200)
);

INVx4_ASAP7_75t_L g3201 ( 
.A(n_2918),
.Y(n_3201)
);

INVx2_ASAP7_75t_SL g3202 ( 
.A(n_2815),
.Y(n_3202)
);

AND2x2_ASAP7_75t_L g3203 ( 
.A(n_2804),
.B(n_523),
.Y(n_3203)
);

BUFx2_ASAP7_75t_SL g3204 ( 
.A(n_2856),
.Y(n_3204)
);

BUFx2_ASAP7_75t_SL g3205 ( 
.A(n_2789),
.Y(n_3205)
);

INVx2_ASAP7_75t_L g3206 ( 
.A(n_2920),
.Y(n_3206)
);

BUFx6f_ASAP7_75t_L g3207 ( 
.A(n_2830),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_2844),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_2860),
.Y(n_3209)
);

BUFx6f_ASAP7_75t_L g3210 ( 
.A(n_2904),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_2868),
.Y(n_3211)
);

BUFx3_ASAP7_75t_L g3212 ( 
.A(n_2775),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_2869),
.Y(n_3213)
);

INVx3_ASAP7_75t_L g3214 ( 
.A(n_2907),
.Y(n_3214)
);

INVx6_ASAP7_75t_L g3215 ( 
.A(n_2635),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_2871),
.Y(n_3216)
);

INVx6_ASAP7_75t_L g3217 ( 
.A(n_2658),
.Y(n_3217)
);

BUFx2_ASAP7_75t_L g3218 ( 
.A(n_2861),
.Y(n_3218)
);

AND2x2_ASAP7_75t_L g3219 ( 
.A(n_2929),
.B(n_524),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_2883),
.Y(n_3220)
);

BUFx6f_ASAP7_75t_L g3221 ( 
.A(n_2909),
.Y(n_3221)
);

NOR2x1_ASAP7_75t_L g3222 ( 
.A(n_2863),
.B(n_524),
.Y(n_3222)
);

NAND2x1p5_ASAP7_75t_L g3223 ( 
.A(n_2870),
.B(n_525),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_2887),
.Y(n_3224)
);

BUFx6f_ASAP7_75t_L g3225 ( 
.A(n_2911),
.Y(n_3225)
);

INVx5_ASAP7_75t_L g3226 ( 
.A(n_2760),
.Y(n_3226)
);

AND2x2_ASAP7_75t_L g3227 ( 
.A(n_2708),
.B(n_525),
.Y(n_3227)
);

BUFx12f_ASAP7_75t_L g3228 ( 
.A(n_2736),
.Y(n_3228)
);

AND2x4_ASAP7_75t_L g3229 ( 
.A(n_2668),
.B(n_2726),
.Y(n_3229)
);

BUFx6f_ASAP7_75t_L g3230 ( 
.A(n_2923),
.Y(n_3230)
);

INVxp67_ASAP7_75t_SL g3231 ( 
.A(n_2854),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_2888),
.Y(n_3232)
);

OR2x6_ASAP7_75t_L g3233 ( 
.A(n_2710),
.B(n_526),
.Y(n_3233)
);

BUFx3_ASAP7_75t_L g3234 ( 
.A(n_2798),
.Y(n_3234)
);

INVx2_ASAP7_75t_SL g3235 ( 
.A(n_2945),
.Y(n_3235)
);

NOR2xp33_ASAP7_75t_L g3236 ( 
.A(n_2942),
.B(n_2881),
.Y(n_3236)
);

INVx2_ASAP7_75t_L g3237 ( 
.A(n_3066),
.Y(n_3237)
);

BUFx3_ASAP7_75t_L g3238 ( 
.A(n_2970),
.Y(n_3238)
);

OR2x6_ASAP7_75t_L g3239 ( 
.A(n_3139),
.B(n_2953),
.Y(n_3239)
);

NAND2x1p5_ASAP7_75t_L g3240 ( 
.A(n_2974),
.B(n_2879),
.Y(n_3240)
);

OAI21x1_ASAP7_75t_L g3241 ( 
.A1(n_3161),
.A2(n_2671),
.B(n_2615),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_2940),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_2944),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_2951),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_2962),
.Y(n_3245)
);

OR2x2_ASAP7_75t_L g3246 ( 
.A(n_3005),
.B(n_2801),
.Y(n_3246)
);

NOR2xp33_ASAP7_75t_L g3247 ( 
.A(n_3118),
.B(n_2884),
.Y(n_3247)
);

O2A1O1Ixp33_ASAP7_75t_L g3248 ( 
.A1(n_3154),
.A2(n_2733),
.B(n_2823),
.C(n_2828),
.Y(n_3248)
);

AO32x2_ASAP7_75t_L g3249 ( 
.A1(n_3018),
.A2(n_2811),
.A3(n_2831),
.B1(n_2816),
.B2(n_2813),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_2973),
.Y(n_3250)
);

AND2x2_ASAP7_75t_L g3251 ( 
.A(n_3001),
.B(n_2960),
.Y(n_3251)
);

A2O1A1Ixp33_ASAP7_75t_L g3252 ( 
.A1(n_3129),
.A2(n_2746),
.B(n_2724),
.C(n_2696),
.Y(n_3252)
);

OAI21x1_ASAP7_75t_L g3253 ( 
.A1(n_3120),
.A2(n_2857),
.B(n_2853),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_2981),
.Y(n_3254)
);

AO21x2_ASAP7_75t_L g3255 ( 
.A1(n_3231),
.A2(n_2728),
.B(n_2690),
.Y(n_3255)
);

AOI22xp33_ASAP7_75t_L g3256 ( 
.A1(n_3193),
.A2(n_2773),
.B1(n_2917),
.B2(n_2770),
.Y(n_3256)
);

NOR2x1_ASAP7_75t_SL g3257 ( 
.A(n_2989),
.B(n_2922),
.Y(n_3257)
);

OAI21x1_ASAP7_75t_L g3258 ( 
.A1(n_3196),
.A2(n_2706),
.B(n_2684),
.Y(n_3258)
);

BUFx12f_ASAP7_75t_L g3259 ( 
.A(n_2937),
.Y(n_3259)
);

HB1xp67_ASAP7_75t_L g3260 ( 
.A(n_2961),
.Y(n_3260)
);

INVx2_ASAP7_75t_L g3261 ( 
.A(n_2972),
.Y(n_3261)
);

BUFx6f_ASAP7_75t_L g3262 ( 
.A(n_2941),
.Y(n_3262)
);

AND2x4_ASAP7_75t_L g3263 ( 
.A(n_2965),
.B(n_2764),
.Y(n_3263)
);

AO21x1_ASAP7_75t_L g3264 ( 
.A1(n_3119),
.A2(n_2784),
.B(n_2808),
.Y(n_3264)
);

OR2x2_ASAP7_75t_L g3265 ( 
.A(n_2967),
.B(n_526),
.Y(n_3265)
);

BUFx2_ASAP7_75t_R g3266 ( 
.A(n_2939),
.Y(n_3266)
);

OAI22xp5_ASAP7_75t_L g3267 ( 
.A1(n_3006),
.A2(n_2837),
.B1(n_2810),
.B2(n_2901),
.Y(n_3267)
);

AND2x2_ASAP7_75t_L g3268 ( 
.A(n_3153),
.B(n_2780),
.Y(n_3268)
);

INVx2_ASAP7_75t_L g3269 ( 
.A(n_2993),
.Y(n_3269)
);

OA21x2_ASAP7_75t_L g3270 ( 
.A1(n_3162),
.A2(n_2867),
.B(n_2679),
.Y(n_3270)
);

INVx2_ASAP7_75t_L g3271 ( 
.A(n_2995),
.Y(n_3271)
);

INVx2_ASAP7_75t_SL g3272 ( 
.A(n_2963),
.Y(n_3272)
);

AND2x4_ASAP7_75t_L g3273 ( 
.A(n_3142),
.B(n_2817),
.Y(n_3273)
);

BUFx6f_ASAP7_75t_L g3274 ( 
.A(n_2941),
.Y(n_3274)
);

AO21x2_ASAP7_75t_L g3275 ( 
.A1(n_3138),
.A2(n_2814),
.B(n_2762),
.Y(n_3275)
);

OAI21x1_ASAP7_75t_L g3276 ( 
.A1(n_3191),
.A2(n_2754),
.B(n_2930),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_2985),
.Y(n_3277)
);

INVx3_ASAP7_75t_L g3278 ( 
.A(n_2997),
.Y(n_3278)
);

OAI21x1_ASAP7_75t_L g3279 ( 
.A1(n_3197),
.A2(n_2931),
.B(n_2915),
.Y(n_3279)
);

OAI21x1_ASAP7_75t_L g3280 ( 
.A1(n_3206),
.A2(n_2921),
.B(n_2910),
.Y(n_3280)
);

AO21x2_ASAP7_75t_L g3281 ( 
.A1(n_3070),
.A2(n_2703),
.B(n_2707),
.Y(n_3281)
);

INVx3_ASAP7_75t_L g3282 ( 
.A(n_2943),
.Y(n_3282)
);

NAND2xp5_ASAP7_75t_L g3283 ( 
.A(n_3023),
.B(n_2761),
.Y(n_3283)
);

BUFx12f_ASAP7_75t_L g3284 ( 
.A(n_2964),
.Y(n_3284)
);

BUFx6f_ASAP7_75t_L g3285 ( 
.A(n_2947),
.Y(n_3285)
);

AOI22xp33_ASAP7_75t_L g3286 ( 
.A1(n_3205),
.A2(n_2793),
.B1(n_2842),
.B2(n_2800),
.Y(n_3286)
);

BUFx3_ASAP7_75t_L g3287 ( 
.A(n_2992),
.Y(n_3287)
);

AND2x2_ASAP7_75t_L g3288 ( 
.A(n_2977),
.B(n_526),
.Y(n_3288)
);

INVx8_ASAP7_75t_L g3289 ( 
.A(n_2963),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_2990),
.Y(n_3290)
);

BUFx5_ASAP7_75t_L g3291 ( 
.A(n_3058),
.Y(n_3291)
);

BUFx6f_ASAP7_75t_L g3292 ( 
.A(n_2994),
.Y(n_3292)
);

OAI21x1_ASAP7_75t_L g3293 ( 
.A1(n_3151),
.A2(n_3144),
.B(n_3195),
.Y(n_3293)
);

INVx5_ASAP7_75t_L g3294 ( 
.A(n_2935),
.Y(n_3294)
);

AOI21x1_ASAP7_75t_L g3295 ( 
.A1(n_3087),
.A2(n_2885),
.B(n_2912),
.Y(n_3295)
);

AND2x6_ASAP7_75t_L g3296 ( 
.A(n_3130),
.B(n_2777),
.Y(n_3296)
);

AO31x2_ASAP7_75t_L g3297 ( 
.A1(n_3187),
.A2(n_529),
.A3(n_527),
.B(n_528),
.Y(n_3297)
);

OAI21x1_ASAP7_75t_L g3298 ( 
.A1(n_3082),
.A2(n_3089),
.B(n_3222),
.Y(n_3298)
);

INVx2_ASAP7_75t_L g3299 ( 
.A(n_3000),
.Y(n_3299)
);

OAI22xp5_ASAP7_75t_L g3300 ( 
.A1(n_3107),
.A2(n_529),
.B1(n_527),
.B2(n_528),
.Y(n_3300)
);

OR2x6_ASAP7_75t_L g3301 ( 
.A(n_2998),
.B(n_527),
.Y(n_3301)
);

AND2x2_ASAP7_75t_L g3302 ( 
.A(n_2977),
.B(n_530),
.Y(n_3302)
);

OAI22xp33_ASAP7_75t_L g3303 ( 
.A1(n_3042),
.A2(n_533),
.B1(n_531),
.B2(n_532),
.Y(n_3303)
);

INVx2_ASAP7_75t_L g3304 ( 
.A(n_3011),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_2991),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_3094),
.Y(n_3306)
);

OAI21x1_ASAP7_75t_L g3307 ( 
.A1(n_3178),
.A2(n_661),
.B(n_660),
.Y(n_3307)
);

AO31x2_ASAP7_75t_L g3308 ( 
.A1(n_3199),
.A2(n_536),
.A3(n_534),
.B(n_535),
.Y(n_3308)
);

INVx1_ASAP7_75t_SL g3309 ( 
.A(n_2968),
.Y(n_3309)
);

OAI22xp5_ASAP7_75t_L g3310 ( 
.A1(n_3053),
.A2(n_536),
.B1(n_534),
.B2(n_535),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_3109),
.Y(n_3311)
);

INVx2_ASAP7_75t_SL g3312 ( 
.A(n_2959),
.Y(n_3312)
);

AO21x2_ASAP7_75t_L g3313 ( 
.A1(n_3163),
.A2(n_537),
.B(n_538),
.Y(n_3313)
);

OAI21x1_ASAP7_75t_L g3314 ( 
.A1(n_3175),
.A2(n_663),
.B(n_662),
.Y(n_3314)
);

INVx2_ASAP7_75t_L g3315 ( 
.A(n_3041),
.Y(n_3315)
);

A2O1A1Ixp33_ASAP7_75t_L g3316 ( 
.A1(n_3143),
.A2(n_541),
.B(n_539),
.C(n_540),
.Y(n_3316)
);

AO21x2_ASAP7_75t_L g3317 ( 
.A1(n_3168),
.A2(n_539),
.B(n_540),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3121),
.Y(n_3318)
);

INVx2_ASAP7_75t_L g3319 ( 
.A(n_3049),
.Y(n_3319)
);

HB1xp67_ASAP7_75t_L g3320 ( 
.A(n_3112),
.Y(n_3320)
);

BUFx6f_ASAP7_75t_L g3321 ( 
.A(n_2996),
.Y(n_3321)
);

HB1xp67_ASAP7_75t_L g3322 ( 
.A(n_3080),
.Y(n_3322)
);

INVx2_ASAP7_75t_SL g3323 ( 
.A(n_2975),
.Y(n_3323)
);

BUFx2_ASAP7_75t_L g3324 ( 
.A(n_2988),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_3133),
.Y(n_3325)
);

NAND2x1p5_ASAP7_75t_L g3326 ( 
.A(n_2954),
.B(n_542),
.Y(n_3326)
);

AOI22xp33_ASAP7_75t_L g3327 ( 
.A1(n_3217),
.A2(n_545),
.B1(n_543),
.B2(n_544),
.Y(n_3327)
);

CKINVDCx11_ASAP7_75t_R g3328 ( 
.A(n_2957),
.Y(n_3328)
);

AND2x4_ASAP7_75t_L g3329 ( 
.A(n_2979),
.B(n_3174),
.Y(n_3329)
);

AND2x4_ASAP7_75t_L g3330 ( 
.A(n_3174),
.B(n_544),
.Y(n_3330)
);

CKINVDCx6p67_ASAP7_75t_R g3331 ( 
.A(n_2938),
.Y(n_3331)
);

INVxp67_ASAP7_75t_SL g3332 ( 
.A(n_3179),
.Y(n_3332)
);

INVx1_ASAP7_75t_L g3333 ( 
.A(n_3140),
.Y(n_3333)
);

INVx2_ASAP7_75t_SL g3334 ( 
.A(n_2975),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_3024),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_3030),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_3047),
.Y(n_3337)
);

INVx1_ASAP7_75t_L g3338 ( 
.A(n_3063),
.Y(n_3338)
);

OAI21x1_ASAP7_75t_L g3339 ( 
.A1(n_3219),
.A2(n_667),
.B(n_666),
.Y(n_3339)
);

OAI21x1_ASAP7_75t_L g3340 ( 
.A1(n_3145),
.A2(n_3148),
.B(n_3214),
.Y(n_3340)
);

OAI21x1_ASAP7_75t_L g3341 ( 
.A1(n_3145),
.A2(n_667),
.B(n_666),
.Y(n_3341)
);

CKINVDCx5p33_ASAP7_75t_R g3342 ( 
.A(n_2952),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_3064),
.Y(n_3343)
);

OA21x2_ASAP7_75t_L g3344 ( 
.A1(n_3188),
.A2(n_546),
.B(n_547),
.Y(n_3344)
);

OAI21x1_ASAP7_75t_L g3345 ( 
.A1(n_3148),
.A2(n_669),
.B(n_668),
.Y(n_3345)
);

INVx2_ASAP7_75t_L g3346 ( 
.A(n_3084),
.Y(n_3346)
);

AND2x4_ASAP7_75t_L g3347 ( 
.A(n_2986),
.B(n_548),
.Y(n_3347)
);

INVx1_ASAP7_75t_L g3348 ( 
.A(n_3027),
.Y(n_3348)
);

INVx2_ASAP7_75t_L g3349 ( 
.A(n_3203),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_3079),
.Y(n_3350)
);

INVx2_ASAP7_75t_L g3351 ( 
.A(n_3170),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_SL g3352 ( 
.A(n_3149),
.B(n_3141),
.Y(n_3352)
);

BUFx8_ASAP7_75t_L g3353 ( 
.A(n_2956),
.Y(n_3353)
);

OA21x2_ASAP7_75t_L g3354 ( 
.A1(n_3218),
.A2(n_551),
.B(n_552),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_3090),
.Y(n_3355)
);

NAND2x1p5_ASAP7_75t_L g3356 ( 
.A(n_2955),
.B(n_553),
.Y(n_3356)
);

OAI21x1_ASAP7_75t_L g3357 ( 
.A1(n_3170),
.A2(n_674),
.B(n_673),
.Y(n_3357)
);

OAI21x1_ASAP7_75t_L g3358 ( 
.A1(n_3169),
.A2(n_677),
.B(n_676),
.Y(n_3358)
);

OAI21x1_ASAP7_75t_L g3359 ( 
.A1(n_3116),
.A2(n_678),
.B(n_676),
.Y(n_3359)
);

OAI21xp5_ASAP7_75t_L g3360 ( 
.A1(n_3227),
.A2(n_2946),
.B(n_2982),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_3069),
.B(n_3073),
.Y(n_3361)
);

OAI21x1_ASAP7_75t_L g3362 ( 
.A1(n_3008),
.A2(n_679),
.B(n_678),
.Y(n_3362)
);

A2O1A1Ixp33_ASAP7_75t_L g3363 ( 
.A1(n_3156),
.A2(n_556),
.B(n_554),
.C(n_555),
.Y(n_3363)
);

HB1xp67_ASAP7_75t_L g3364 ( 
.A(n_3021),
.Y(n_3364)
);

OAI21x1_ASAP7_75t_L g3365 ( 
.A1(n_3223),
.A2(n_681),
.B(n_680),
.Y(n_3365)
);

OAI21x1_ASAP7_75t_L g3366 ( 
.A1(n_3076),
.A2(n_682),
.B(n_681),
.Y(n_3366)
);

OR2x6_ASAP7_75t_L g3367 ( 
.A(n_2976),
.B(n_557),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_L g3368 ( 
.A(n_3126),
.B(n_558),
.Y(n_3368)
);

INVx5_ASAP7_75t_L g3369 ( 
.A(n_3127),
.Y(n_3369)
);

OAI21x1_ASAP7_75t_L g3370 ( 
.A1(n_2999),
.A2(n_683),
.B(n_682),
.Y(n_3370)
);

INVx2_ASAP7_75t_L g3371 ( 
.A(n_3088),
.Y(n_3371)
);

BUFx2_ASAP7_75t_L g3372 ( 
.A(n_2958),
.Y(n_3372)
);

OAI21x1_ASAP7_75t_L g3373 ( 
.A1(n_3022),
.A2(n_684),
.B(n_683),
.Y(n_3373)
);

AOI21x1_ASAP7_75t_L g3374 ( 
.A1(n_3150),
.A2(n_3002),
.B(n_3229),
.Y(n_3374)
);

INVx4_ASAP7_75t_L g3375 ( 
.A(n_2949),
.Y(n_3375)
);

A2O1A1Ixp33_ASAP7_75t_L g3376 ( 
.A1(n_3226),
.A2(n_561),
.B(n_559),
.C(n_560),
.Y(n_3376)
);

INVx2_ASAP7_75t_L g3377 ( 
.A(n_3106),
.Y(n_3377)
);

NOR2xp33_ASAP7_75t_L g3378 ( 
.A(n_2966),
.B(n_561),
.Y(n_3378)
);

NOR2xp33_ASAP7_75t_L g3379 ( 
.A(n_3085),
.B(n_562),
.Y(n_3379)
);

OAI21x1_ASAP7_75t_L g3380 ( 
.A1(n_3048),
.A2(n_686),
.B(n_685),
.Y(n_3380)
);

BUFx12f_ASAP7_75t_L g3381 ( 
.A(n_3045),
.Y(n_3381)
);

INVx1_ASAP7_75t_SL g3382 ( 
.A(n_3060),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_3048),
.Y(n_3383)
);

OAI21x1_ASAP7_75t_L g3384 ( 
.A1(n_3123),
.A2(n_686),
.B(n_685),
.Y(n_3384)
);

INVx3_ASAP7_75t_L g3385 ( 
.A(n_2987),
.Y(n_3385)
);

OAI21x1_ASAP7_75t_L g3386 ( 
.A1(n_2969),
.A2(n_3173),
.B(n_3134),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_2984),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_L g3388 ( 
.A(n_3113),
.B(n_569),
.Y(n_3388)
);

INVx2_ASAP7_75t_L g3389 ( 
.A(n_3122),
.Y(n_3389)
);

INVx1_ASAP7_75t_L g3390 ( 
.A(n_3159),
.Y(n_3390)
);

AO31x2_ASAP7_75t_L g3391 ( 
.A1(n_3201),
.A2(n_571),
.A3(n_569),
.B(n_570),
.Y(n_3391)
);

AO21x2_ASAP7_75t_L g3392 ( 
.A1(n_3007),
.A2(n_3028),
.B(n_3046),
.Y(n_3392)
);

INVx2_ASAP7_75t_L g3393 ( 
.A(n_3122),
.Y(n_3393)
);

OAI21x1_ASAP7_75t_L g3394 ( 
.A1(n_3208),
.A2(n_688),
.B(n_687),
.Y(n_3394)
);

OAI21x1_ASAP7_75t_L g3395 ( 
.A1(n_3209),
.A2(n_691),
.B(n_689),
.Y(n_3395)
);

AOI22xp33_ASAP7_75t_L g3396 ( 
.A1(n_3215),
.A2(n_574),
.B1(n_572),
.B2(n_573),
.Y(n_3396)
);

AO31x2_ASAP7_75t_L g3397 ( 
.A1(n_3167),
.A2(n_576),
.A3(n_573),
.B(n_575),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_3111),
.Y(n_3398)
);

INVx2_ASAP7_75t_L g3399 ( 
.A(n_3190),
.Y(n_3399)
);

OAI21xp5_ASAP7_75t_L g3400 ( 
.A1(n_3233),
.A2(n_576),
.B(n_577),
.Y(n_3400)
);

OAI22xp33_ASAP7_75t_L g3401 ( 
.A1(n_3198),
.A2(n_578),
.B1(n_576),
.B2(n_577),
.Y(n_3401)
);

OAI21xp5_ASAP7_75t_L g3402 ( 
.A1(n_3061),
.A2(n_577),
.B(n_578),
.Y(n_3402)
);

BUFx12f_ASAP7_75t_L g3403 ( 
.A(n_3057),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_L g3404 ( 
.A(n_3136),
.B(n_3013),
.Y(n_3404)
);

HB1xp67_ASAP7_75t_L g3405 ( 
.A(n_3031),
.Y(n_3405)
);

INVx2_ASAP7_75t_L g3406 ( 
.A(n_3190),
.Y(n_3406)
);

BUFx2_ASAP7_75t_L g3407 ( 
.A(n_3091),
.Y(n_3407)
);

OAI21x1_ASAP7_75t_L g3408 ( 
.A1(n_3211),
.A2(n_3216),
.B(n_3213),
.Y(n_3408)
);

AND2x2_ASAP7_75t_L g3409 ( 
.A(n_3074),
.B(n_579),
.Y(n_3409)
);

OAI21x1_ASAP7_75t_L g3410 ( 
.A1(n_3220),
.A2(n_3232),
.B(n_3224),
.Y(n_3410)
);

NAND2x1p5_ASAP7_75t_L g3411 ( 
.A(n_2948),
.B(n_580),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_3320),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_3242),
.Y(n_3413)
);

OA21x2_ASAP7_75t_L g3414 ( 
.A1(n_3293),
.A2(n_3177),
.B(n_3160),
.Y(n_3414)
);

NOR2xp33_ASAP7_75t_L g3415 ( 
.A(n_3309),
.B(n_3043),
.Y(n_3415)
);

INVx1_ASAP7_75t_SL g3416 ( 
.A(n_3287),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_3243),
.Y(n_3417)
);

INVx3_ASAP7_75t_L g3418 ( 
.A(n_3331),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_3244),
.Y(n_3419)
);

INVx1_ASAP7_75t_L g3420 ( 
.A(n_3245),
.Y(n_3420)
);

BUFx3_ASAP7_75t_L g3421 ( 
.A(n_3238),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_3250),
.Y(n_3422)
);

AOI21x1_ASAP7_75t_L g3423 ( 
.A1(n_3374),
.A2(n_3186),
.B(n_3157),
.Y(n_3423)
);

BUFx2_ASAP7_75t_L g3424 ( 
.A(n_3340),
.Y(n_3424)
);

INVx2_ASAP7_75t_L g3425 ( 
.A(n_3261),
.Y(n_3425)
);

INVx2_ASAP7_75t_L g3426 ( 
.A(n_3269),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_3254),
.Y(n_3427)
);

OAI21x1_ASAP7_75t_L g3428 ( 
.A1(n_3241),
.A2(n_3189),
.B(n_3147),
.Y(n_3428)
);

HB1xp67_ASAP7_75t_L g3429 ( 
.A(n_3260),
.Y(n_3429)
);

INVx2_ASAP7_75t_L g3430 ( 
.A(n_3271),
.Y(n_3430)
);

NOR2xp33_ASAP7_75t_L g3431 ( 
.A(n_3235),
.B(n_3029),
.Y(n_3431)
);

OR2x6_ASAP7_75t_L g3432 ( 
.A(n_3239),
.B(n_3014),
.Y(n_3432)
);

CKINVDCx6p67_ASAP7_75t_R g3433 ( 
.A(n_3369),
.Y(n_3433)
);

INVx2_ASAP7_75t_SL g3434 ( 
.A(n_3285),
.Y(n_3434)
);

INVx2_ASAP7_75t_L g3435 ( 
.A(n_3299),
.Y(n_3435)
);

INVx2_ASAP7_75t_L g3436 ( 
.A(n_3304),
.Y(n_3436)
);

INVx1_ASAP7_75t_L g3437 ( 
.A(n_3277),
.Y(n_3437)
);

INVx1_ASAP7_75t_L g3438 ( 
.A(n_3290),
.Y(n_3438)
);

INVx2_ASAP7_75t_L g3439 ( 
.A(n_3315),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3305),
.Y(n_3440)
);

INVx2_ASAP7_75t_L g3441 ( 
.A(n_3319),
.Y(n_3441)
);

AOI21x1_ASAP7_75t_L g3442 ( 
.A1(n_3253),
.A2(n_3003),
.B(n_3068),
.Y(n_3442)
);

AND2x4_ASAP7_75t_L g3443 ( 
.A(n_3329),
.B(n_3137),
.Y(n_3443)
);

BUFx5_ASAP7_75t_L g3444 ( 
.A(n_3296),
.Y(n_3444)
);

INVx2_ASAP7_75t_SL g3445 ( 
.A(n_3292),
.Y(n_3445)
);

BUFx4f_ASAP7_75t_SL g3446 ( 
.A(n_3381),
.Y(n_3446)
);

AND2x4_ASAP7_75t_L g3447 ( 
.A(n_3251),
.B(n_3016),
.Y(n_3447)
);

BUFx4f_ASAP7_75t_SL g3448 ( 
.A(n_3403),
.Y(n_3448)
);

AOI21xp5_ASAP7_75t_L g3449 ( 
.A1(n_3257),
.A2(n_3056),
.B(n_3182),
.Y(n_3449)
);

BUFx2_ASAP7_75t_L g3450 ( 
.A(n_3364),
.Y(n_3450)
);

OAI21x1_ASAP7_75t_L g3451 ( 
.A1(n_3295),
.A2(n_3192),
.B(n_3171),
.Y(n_3451)
);

AOI21x1_ASAP7_75t_L g3452 ( 
.A1(n_3264),
.A2(n_2936),
.B(n_3115),
.Y(n_3452)
);

BUFx2_ASAP7_75t_L g3453 ( 
.A(n_3405),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3371),
.Y(n_3454)
);

AND2x2_ASAP7_75t_L g3455 ( 
.A(n_3335),
.B(n_3131),
.Y(n_3455)
);

INVx2_ASAP7_75t_L g3456 ( 
.A(n_3346),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_3350),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3355),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_3408),
.Y(n_3459)
);

BUFx2_ASAP7_75t_L g3460 ( 
.A(n_3237),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_3410),
.Y(n_3461)
);

INVx2_ASAP7_75t_L g3462 ( 
.A(n_3306),
.Y(n_3462)
);

INVx2_ASAP7_75t_L g3463 ( 
.A(n_3311),
.Y(n_3463)
);

OR2x2_ASAP7_75t_L g3464 ( 
.A(n_3348),
.B(n_2971),
.Y(n_3464)
);

INVx2_ASAP7_75t_L g3465 ( 
.A(n_3318),
.Y(n_3465)
);

BUFx6f_ASAP7_75t_L g3466 ( 
.A(n_3262),
.Y(n_3466)
);

AND2x2_ASAP7_75t_L g3467 ( 
.A(n_3390),
.B(n_3124),
.Y(n_3467)
);

INVx2_ASAP7_75t_L g3468 ( 
.A(n_3325),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_3336),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_3337),
.Y(n_3470)
);

OA21x2_ASAP7_75t_L g3471 ( 
.A1(n_3298),
.A2(n_3035),
.B(n_3081),
.Y(n_3471)
);

INVx2_ASAP7_75t_L g3472 ( 
.A(n_3333),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3338),
.Y(n_3473)
);

INVx1_ASAP7_75t_L g3474 ( 
.A(n_3343),
.Y(n_3474)
);

INVx2_ASAP7_75t_L g3475 ( 
.A(n_3349),
.Y(n_3475)
);

HB1xp67_ASAP7_75t_L g3476 ( 
.A(n_3322),
.Y(n_3476)
);

BUFx2_ASAP7_75t_L g3477 ( 
.A(n_3399),
.Y(n_3477)
);

INVx2_ASAP7_75t_L g3478 ( 
.A(n_3351),
.Y(n_3478)
);

OAI21x1_ASAP7_75t_L g3479 ( 
.A1(n_3258),
.A2(n_3095),
.B(n_3176),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_3361),
.Y(n_3480)
);

INVx2_ASAP7_75t_L g3481 ( 
.A(n_3398),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3404),
.Y(n_3482)
);

INVx2_ASAP7_75t_L g3483 ( 
.A(n_3406),
.Y(n_3483)
);

OAI21x1_ASAP7_75t_L g3484 ( 
.A1(n_3276),
.A2(n_3279),
.B(n_3307),
.Y(n_3484)
);

AND2x2_ASAP7_75t_L g3485 ( 
.A(n_3389),
.B(n_3164),
.Y(n_3485)
);

INVx2_ASAP7_75t_L g3486 ( 
.A(n_3377),
.Y(n_3486)
);

AO21x1_ASAP7_75t_SL g3487 ( 
.A1(n_3400),
.A2(n_3036),
.B(n_3026),
.Y(n_3487)
);

INVxp33_ASAP7_75t_L g3488 ( 
.A(n_3328),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3387),
.Y(n_3489)
);

OR2x6_ASAP7_75t_L g3490 ( 
.A(n_3239),
.B(n_3099),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_3383),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_L g3492 ( 
.A(n_3246),
.B(n_3200),
.Y(n_3492)
);

INVx2_ASAP7_75t_L g3493 ( 
.A(n_3393),
.Y(n_3493)
);

AND2x2_ASAP7_75t_L g3494 ( 
.A(n_3282),
.B(n_3409),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_L g3495 ( 
.A(n_3392),
.B(n_3202),
.Y(n_3495)
);

INVx2_ASAP7_75t_L g3496 ( 
.A(n_3344),
.Y(n_3496)
);

INVx2_ASAP7_75t_L g3497 ( 
.A(n_3354),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_L g3498 ( 
.A(n_3288),
.B(n_3135),
.Y(n_3498)
);

INVx2_ASAP7_75t_L g3499 ( 
.A(n_3354),
.Y(n_3499)
);

INVx1_ASAP7_75t_L g3500 ( 
.A(n_3368),
.Y(n_3500)
);

AND2x2_ASAP7_75t_L g3501 ( 
.A(n_3302),
.B(n_3033),
.Y(n_3501)
);

BUFx3_ASAP7_75t_L g3502 ( 
.A(n_3274),
.Y(n_3502)
);

AND2x2_ASAP7_75t_L g3503 ( 
.A(n_3375),
.B(n_3039),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_L g3504 ( 
.A(n_3268),
.B(n_3210),
.Y(n_3504)
);

BUFx3_ASAP7_75t_L g3505 ( 
.A(n_3274),
.Y(n_3505)
);

INVx1_ASAP7_75t_L g3506 ( 
.A(n_3265),
.Y(n_3506)
);

INVx2_ASAP7_75t_SL g3507 ( 
.A(n_3289),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_3391),
.Y(n_3508)
);

BUFx2_ASAP7_75t_L g3509 ( 
.A(n_3385),
.Y(n_3509)
);

OAI222xp33_ASAP7_75t_L g3510 ( 
.A1(n_3301),
.A2(n_3086),
.B1(n_3105),
.B2(n_3077),
.C1(n_3009),
.C2(n_3062),
.Y(n_3510)
);

HB1xp67_ASAP7_75t_L g3511 ( 
.A(n_3301),
.Y(n_3511)
);

INVx2_ASAP7_75t_L g3512 ( 
.A(n_3373),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_3380),
.Y(n_3513)
);

INVx2_ASAP7_75t_SL g3514 ( 
.A(n_3294),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_L g3515 ( 
.A(n_3482),
.B(n_3256),
.Y(n_3515)
);

CKINVDCx16_ASAP7_75t_R g3516 ( 
.A(n_3421),
.Y(n_3516)
);

INVx1_ASAP7_75t_L g3517 ( 
.A(n_3413),
.Y(n_3517)
);

INVx3_ASAP7_75t_L g3518 ( 
.A(n_3433),
.Y(n_3518)
);

INVx2_ASAP7_75t_L g3519 ( 
.A(n_3450),
.Y(n_3519)
);

INVx2_ASAP7_75t_L g3520 ( 
.A(n_3453),
.Y(n_3520)
);

AO31x2_ASAP7_75t_L g3521 ( 
.A1(n_3495),
.A2(n_3407),
.A3(n_3378),
.B(n_3247),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_3417),
.Y(n_3522)
);

INVx2_ASAP7_75t_L g3523 ( 
.A(n_3453),
.Y(n_3523)
);

O2A1O1Ixp33_ASAP7_75t_SL g3524 ( 
.A1(n_3510),
.A2(n_3332),
.B(n_3352),
.C(n_3312),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3419),
.Y(n_3525)
);

HB1xp67_ASAP7_75t_L g3526 ( 
.A(n_3429),
.Y(n_3526)
);

BUFx3_ASAP7_75t_L g3527 ( 
.A(n_3503),
.Y(n_3527)
);

BUFx6f_ASAP7_75t_L g3528 ( 
.A(n_3466),
.Y(n_3528)
);

INVx2_ASAP7_75t_SL g3529 ( 
.A(n_3416),
.Y(n_3529)
);

NAND2xp33_ASAP7_75t_SL g3530 ( 
.A(n_3511),
.B(n_3321),
.Y(n_3530)
);

AND2x4_ASAP7_75t_SL g3531 ( 
.A(n_3490),
.B(n_3321),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_3420),
.Y(n_3532)
);

BUFx3_ASAP7_75t_L g3533 ( 
.A(n_3446),
.Y(n_3533)
);

AND2x2_ASAP7_75t_L g3534 ( 
.A(n_3460),
.B(n_3037),
.Y(n_3534)
);

INVx3_ASAP7_75t_L g3535 ( 
.A(n_3490),
.Y(n_3535)
);

BUFx3_ASAP7_75t_L g3536 ( 
.A(n_3448),
.Y(n_3536)
);

OR2x6_ASAP7_75t_L g3537 ( 
.A(n_3432),
.B(n_3284),
.Y(n_3537)
);

AO31x2_ASAP7_75t_L g3538 ( 
.A1(n_3424),
.A2(n_3372),
.A3(n_3236),
.B(n_3324),
.Y(n_3538)
);

OAI21x1_ASAP7_75t_L g3539 ( 
.A1(n_3423),
.A2(n_3442),
.B(n_3428),
.Y(n_3539)
);

NAND2xp33_ASAP7_75t_R g3540 ( 
.A(n_3418),
.B(n_3367),
.Y(n_3540)
);

AND2x2_ASAP7_75t_L g3541 ( 
.A(n_3476),
.B(n_3382),
.Y(n_3541)
);

AND2x4_ASAP7_75t_L g3542 ( 
.A(n_3447),
.B(n_3294),
.Y(n_3542)
);

INVx1_ASAP7_75t_L g3543 ( 
.A(n_3422),
.Y(n_3543)
);

AND2x4_ASAP7_75t_L g3544 ( 
.A(n_3509),
.B(n_3272),
.Y(n_3544)
);

AO31x2_ASAP7_75t_L g3545 ( 
.A1(n_3424),
.A2(n_3379),
.A3(n_3300),
.B(n_3310),
.Y(n_3545)
);

OR2x6_ASAP7_75t_L g3546 ( 
.A(n_3514),
.B(n_3367),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_3480),
.B(n_3313),
.Y(n_3547)
);

BUFx2_ASAP7_75t_L g3548 ( 
.A(n_3502),
.Y(n_3548)
);

INVx2_ASAP7_75t_L g3549 ( 
.A(n_3425),
.Y(n_3549)
);

INVx2_ASAP7_75t_L g3550 ( 
.A(n_3426),
.Y(n_3550)
);

INVx2_ASAP7_75t_L g3551 ( 
.A(n_3430),
.Y(n_3551)
);

NAND2xp33_ASAP7_75t_SL g3552 ( 
.A(n_3509),
.B(n_3278),
.Y(n_3552)
);

AND2x2_ASAP7_75t_L g3553 ( 
.A(n_3467),
.B(n_3323),
.Y(n_3553)
);

AND2x4_ASAP7_75t_L g3554 ( 
.A(n_3443),
.B(n_3263),
.Y(n_3554)
);

INVx1_ASAP7_75t_L g3555 ( 
.A(n_3427),
.Y(n_3555)
);

NAND2xp33_ASAP7_75t_R g3556 ( 
.A(n_3431),
.B(n_3330),
.Y(n_3556)
);

NOR3xp33_ASAP7_75t_SL g3557 ( 
.A(n_3415),
.B(n_3342),
.C(n_3401),
.Y(n_3557)
);

AND2x2_ASAP7_75t_L g3558 ( 
.A(n_3494),
.B(n_3334),
.Y(n_3558)
);

OR2x6_ASAP7_75t_L g3559 ( 
.A(n_3449),
.B(n_3078),
.Y(n_3559)
);

BUFx2_ASAP7_75t_L g3560 ( 
.A(n_3505),
.Y(n_3560)
);

INVx2_ASAP7_75t_L g3561 ( 
.A(n_3435),
.Y(n_3561)
);

OR2x2_ASAP7_75t_L g3562 ( 
.A(n_3412),
.B(n_3388),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3437),
.Y(n_3563)
);

NOR2xp33_ASAP7_75t_R g3564 ( 
.A(n_3507),
.B(n_3353),
.Y(n_3564)
);

AND2x4_ASAP7_75t_L g3565 ( 
.A(n_3485),
.B(n_3273),
.Y(n_3565)
);

CKINVDCx20_ASAP7_75t_R g3566 ( 
.A(n_3434),
.Y(n_3566)
);

AND2x2_ASAP7_75t_L g3567 ( 
.A(n_3455),
.B(n_3172),
.Y(n_3567)
);

INVx4_ASAP7_75t_L g3568 ( 
.A(n_3466),
.Y(n_3568)
);

CKINVDCx5p33_ASAP7_75t_R g3569 ( 
.A(n_3445),
.Y(n_3569)
);

CKINVDCx16_ASAP7_75t_R g3570 ( 
.A(n_3501),
.Y(n_3570)
);

NAND3xp33_ASAP7_75t_SL g3571 ( 
.A(n_3488),
.B(n_3356),
.C(n_3326),
.Y(n_3571)
);

NAND2xp33_ASAP7_75t_R g3572 ( 
.A(n_3471),
.B(n_3347),
.Y(n_3572)
);

AND2x4_ASAP7_75t_L g3573 ( 
.A(n_3504),
.B(n_3054),
.Y(n_3573)
);

INVx4_ASAP7_75t_L g3574 ( 
.A(n_3444),
.Y(n_3574)
);

HB1xp67_ASAP7_75t_L g3575 ( 
.A(n_3456),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_3475),
.B(n_3317),
.Y(n_3576)
);

NOR2xp33_ASAP7_75t_R g3577 ( 
.A(n_3444),
.B(n_3259),
.Y(n_3577)
);

NOR3xp33_ASAP7_75t_SL g3578 ( 
.A(n_3492),
.B(n_3038),
.C(n_3303),
.Y(n_3578)
);

CKINVDCx16_ASAP7_75t_R g3579 ( 
.A(n_3498),
.Y(n_3579)
);

BUFx2_ASAP7_75t_L g3580 ( 
.A(n_3477),
.Y(n_3580)
);

CKINVDCx5p33_ASAP7_75t_R g3581 ( 
.A(n_3464),
.Y(n_3581)
);

NOR3xp33_ASAP7_75t_SL g3582 ( 
.A(n_3500),
.B(n_3065),
.C(n_3376),
.Y(n_3582)
);

INVx2_ASAP7_75t_L g3583 ( 
.A(n_3436),
.Y(n_3583)
);

BUFx3_ASAP7_75t_L g3584 ( 
.A(n_3454),
.Y(n_3584)
);

AND2x4_ASAP7_75t_L g3585 ( 
.A(n_3481),
.B(n_3210),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3438),
.Y(n_3586)
);

INVx8_ASAP7_75t_L g3587 ( 
.A(n_3487),
.Y(n_3587)
);

OR2x6_ASAP7_75t_L g3588 ( 
.A(n_3479),
.B(n_3411),
.Y(n_3588)
);

NOR2xp33_ASAP7_75t_R g3589 ( 
.A(n_3444),
.B(n_3072),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_3440),
.Y(n_3590)
);

INVx2_ASAP7_75t_L g3591 ( 
.A(n_3439),
.Y(n_3591)
);

INVx3_ASAP7_75t_L g3592 ( 
.A(n_3462),
.Y(n_3592)
);

OR2x6_ASAP7_75t_L g3593 ( 
.A(n_3451),
.B(n_3110),
.Y(n_3593)
);

NOR2xp33_ASAP7_75t_L g3594 ( 
.A(n_3516),
.B(n_3266),
.Y(n_3594)
);

AND2x2_ASAP7_75t_L g3595 ( 
.A(n_3534),
.B(n_3580),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_L g3596 ( 
.A(n_3515),
.B(n_3478),
.Y(n_3596)
);

INVx1_ASAP7_75t_L g3597 ( 
.A(n_3575),
.Y(n_3597)
);

BUFx3_ASAP7_75t_L g3598 ( 
.A(n_3533),
.Y(n_3598)
);

BUFx2_ASAP7_75t_L g3599 ( 
.A(n_3587),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_3517),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_L g3601 ( 
.A(n_3547),
.B(n_3486),
.Y(n_3601)
);

OR2x2_ASAP7_75t_L g3602 ( 
.A(n_3519),
.B(n_3457),
.Y(n_3602)
);

OR2x2_ASAP7_75t_L g3603 ( 
.A(n_3520),
.B(n_3458),
.Y(n_3603)
);

AND2x2_ASAP7_75t_L g3604 ( 
.A(n_3565),
.B(n_3506),
.Y(n_3604)
);

INVx2_ASAP7_75t_L g3605 ( 
.A(n_3584),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_3522),
.Y(n_3606)
);

INVx3_ASAP7_75t_L g3607 ( 
.A(n_3587),
.Y(n_3607)
);

BUFx3_ASAP7_75t_L g3608 ( 
.A(n_3536),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3525),
.Y(n_3609)
);

BUFx3_ASAP7_75t_L g3610 ( 
.A(n_3566),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_3532),
.Y(n_3611)
);

INVx5_ASAP7_75t_L g3612 ( 
.A(n_3537),
.Y(n_3612)
);

BUFx2_ASAP7_75t_L g3613 ( 
.A(n_3552),
.Y(n_3613)
);

HB1xp67_ASAP7_75t_L g3614 ( 
.A(n_3526),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3543),
.Y(n_3615)
);

BUFx2_ASAP7_75t_L g3616 ( 
.A(n_3527),
.Y(n_3616)
);

AND2x4_ASAP7_75t_SL g3617 ( 
.A(n_3537),
.B(n_3052),
.Y(n_3617)
);

BUFx2_ASAP7_75t_L g3618 ( 
.A(n_3564),
.Y(n_3618)
);

OR2x2_ASAP7_75t_L g3619 ( 
.A(n_3523),
.B(n_3463),
.Y(n_3619)
);

AND2x2_ASAP7_75t_L g3620 ( 
.A(n_3544),
.B(n_3489),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_3576),
.B(n_3592),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3555),
.Y(n_3622)
);

BUFx3_ASAP7_75t_L g3623 ( 
.A(n_3529),
.Y(n_3623)
);

OR2x2_ASAP7_75t_L g3624 ( 
.A(n_3562),
.B(n_3465),
.Y(n_3624)
);

INVx2_ASAP7_75t_L g3625 ( 
.A(n_3549),
.Y(n_3625)
);

INVx1_ASAP7_75t_L g3626 ( 
.A(n_3563),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_3586),
.Y(n_3627)
);

INVxp67_ASAP7_75t_SL g3628 ( 
.A(n_3572),
.Y(n_3628)
);

HB1xp67_ASAP7_75t_L g3629 ( 
.A(n_3548),
.Y(n_3629)
);

INVx2_ASAP7_75t_L g3630 ( 
.A(n_3550),
.Y(n_3630)
);

NAND2xp33_ASAP7_75t_SL g3631 ( 
.A(n_3556),
.B(n_3496),
.Y(n_3631)
);

AND2x2_ASAP7_75t_L g3632 ( 
.A(n_3570),
.B(n_3491),
.Y(n_3632)
);

BUFx2_ASAP7_75t_L g3633 ( 
.A(n_3546),
.Y(n_3633)
);

AND2x2_ASAP7_75t_L g3634 ( 
.A(n_3554),
.B(n_3483),
.Y(n_3634)
);

OR2x2_ASAP7_75t_L g3635 ( 
.A(n_3551),
.B(n_3472),
.Y(n_3635)
);

INVx3_ASAP7_75t_L g3636 ( 
.A(n_3559),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3590),
.Y(n_3637)
);

INVx3_ASAP7_75t_L g3638 ( 
.A(n_3559),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3561),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_3583),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3591),
.Y(n_3641)
);

BUFx3_ASAP7_75t_L g3642 ( 
.A(n_3518),
.Y(n_3642)
);

NAND2xp5_ASAP7_75t_L g3643 ( 
.A(n_3521),
.B(n_3468),
.Y(n_3643)
);

HB1xp67_ASAP7_75t_L g3644 ( 
.A(n_3560),
.Y(n_3644)
);

OR2x2_ASAP7_75t_L g3645 ( 
.A(n_3579),
.B(n_3441),
.Y(n_3645)
);

INVx2_ASAP7_75t_L g3646 ( 
.A(n_3585),
.Y(n_3646)
);

INVx1_ASAP7_75t_L g3647 ( 
.A(n_3541),
.Y(n_3647)
);

AND2x4_ASAP7_75t_L g3648 ( 
.A(n_3535),
.B(n_3497),
.Y(n_3648)
);

AND2x2_ASAP7_75t_L g3649 ( 
.A(n_3567),
.B(n_3493),
.Y(n_3649)
);

AND2x2_ASAP7_75t_L g3650 ( 
.A(n_3558),
.B(n_3469),
.Y(n_3650)
);

AND2x2_ASAP7_75t_L g3651 ( 
.A(n_3553),
.B(n_3470),
.Y(n_3651)
);

AND2x2_ASAP7_75t_L g3652 ( 
.A(n_3573),
.B(n_3473),
.Y(n_3652)
);

AND2x4_ASAP7_75t_L g3653 ( 
.A(n_3593),
.B(n_3499),
.Y(n_3653)
);

INVx1_ASAP7_75t_L g3654 ( 
.A(n_3521),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3538),
.Y(n_3655)
);

AND2x2_ASAP7_75t_L g3656 ( 
.A(n_3581),
.B(n_3474),
.Y(n_3656)
);

INVx3_ASAP7_75t_L g3657 ( 
.A(n_3574),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_L g3658 ( 
.A(n_3545),
.B(n_3508),
.Y(n_3658)
);

NOR4xp25_ASAP7_75t_SL g3659 ( 
.A(n_3540),
.B(n_3487),
.C(n_3459),
.D(n_3461),
.Y(n_3659)
);

BUFx10_ASAP7_75t_L g3660 ( 
.A(n_3531),
.Y(n_3660)
);

INVx1_ASAP7_75t_L g3661 ( 
.A(n_3601),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_SL g3662 ( 
.A(n_3631),
.B(n_3530),
.Y(n_3662)
);

NAND2x1_ASAP7_75t_L g3663 ( 
.A(n_3613),
.B(n_3593),
.Y(n_3663)
);

AND2x2_ASAP7_75t_L g3664 ( 
.A(n_3633),
.B(n_3542),
.Y(n_3664)
);

INVx2_ASAP7_75t_L g3665 ( 
.A(n_3616),
.Y(n_3665)
);

BUFx12f_ASAP7_75t_L g3666 ( 
.A(n_3618),
.Y(n_3666)
);

BUFx2_ASAP7_75t_L g3667 ( 
.A(n_3599),
.Y(n_3667)
);

AOI21xp5_ASAP7_75t_L g3668 ( 
.A1(n_3628),
.A2(n_3524),
.B(n_3571),
.Y(n_3668)
);

INVx2_ASAP7_75t_SL g3669 ( 
.A(n_3660),
.Y(n_3669)
);

A2O1A1Ixp33_ASAP7_75t_L g3670 ( 
.A1(n_3612),
.A2(n_3578),
.B(n_3582),
.C(n_3557),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3614),
.Y(n_3671)
);

AND2x2_ASAP7_75t_L g3672 ( 
.A(n_3636),
.B(n_3638),
.Y(n_3672)
);

INVx2_ASAP7_75t_L g3673 ( 
.A(n_3629),
.Y(n_3673)
);

INVx2_ASAP7_75t_L g3674 ( 
.A(n_3644),
.Y(n_3674)
);

NAND3xp33_ASAP7_75t_SL g3675 ( 
.A(n_3659),
.B(n_3589),
.C(n_3577),
.Y(n_3675)
);

AO31x2_ASAP7_75t_L g3676 ( 
.A1(n_3654),
.A2(n_3568),
.A3(n_3513),
.B(n_3512),
.Y(n_3676)
);

A2O1A1Ixp33_ASAP7_75t_L g3677 ( 
.A1(n_3612),
.A2(n_3607),
.B(n_3617),
.C(n_3594),
.Y(n_3677)
);

AND2x2_ASAP7_75t_L g3678 ( 
.A(n_3595),
.B(n_3569),
.Y(n_3678)
);

INVx2_ASAP7_75t_L g3679 ( 
.A(n_3635),
.Y(n_3679)
);

INVxp67_ASAP7_75t_SL g3680 ( 
.A(n_3643),
.Y(n_3680)
);

INVx1_ASAP7_75t_L g3681 ( 
.A(n_3596),
.Y(n_3681)
);

OAI21xp33_ASAP7_75t_SL g3682 ( 
.A1(n_3607),
.A2(n_3539),
.B(n_3588),
.Y(n_3682)
);

NAND4xp25_ASAP7_75t_L g3683 ( 
.A(n_3642),
.B(n_3360),
.C(n_3252),
.D(n_3286),
.Y(n_3683)
);

INVx1_ASAP7_75t_L g3684 ( 
.A(n_3597),
.Y(n_3684)
);

INVx2_ASAP7_75t_SL g3685 ( 
.A(n_3660),
.Y(n_3685)
);

AND2x2_ASAP7_75t_L g3686 ( 
.A(n_3648),
.B(n_3528),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_3600),
.Y(n_3687)
);

OR2x6_ASAP7_75t_L g3688 ( 
.A(n_3598),
.B(n_3032),
.Y(n_3688)
);

AOI22xp33_ASAP7_75t_L g3689 ( 
.A1(n_3647),
.A2(n_3012),
.B1(n_3034),
.B2(n_3221),
.Y(n_3689)
);

INVx3_ASAP7_75t_L g3690 ( 
.A(n_3610),
.Y(n_3690)
);

NOR2xp33_ASAP7_75t_SL g3691 ( 
.A(n_3608),
.B(n_3102),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_3606),
.Y(n_3692)
);

A2O1A1Ixp33_ASAP7_75t_L g3693 ( 
.A1(n_3623),
.A2(n_3657),
.B(n_3632),
.C(n_3645),
.Y(n_3693)
);

INVx2_ASAP7_75t_SL g3694 ( 
.A(n_3605),
.Y(n_3694)
);

INVx5_ASAP7_75t_L g3695 ( 
.A(n_3657),
.Y(n_3695)
);

INVx4_ASAP7_75t_R g3696 ( 
.A(n_3634),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3609),
.Y(n_3697)
);

OR2x2_ASAP7_75t_L g3698 ( 
.A(n_3624),
.B(n_3414),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_3611),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3615),
.Y(n_3700)
);

AO21x2_ASAP7_75t_L g3701 ( 
.A1(n_3655),
.A2(n_3452),
.B(n_3484),
.Y(n_3701)
);

NAND2xp5_ASAP7_75t_L g3702 ( 
.A(n_3658),
.B(n_3621),
.Y(n_3702)
);

INVx2_ASAP7_75t_L g3703 ( 
.A(n_3625),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3622),
.Y(n_3704)
);

AND2x2_ASAP7_75t_L g3705 ( 
.A(n_3649),
.B(n_3281),
.Y(n_3705)
);

AND2x2_ASAP7_75t_L g3706 ( 
.A(n_3652),
.B(n_3125),
.Y(n_3706)
);

OAI22xp33_ASAP7_75t_L g3707 ( 
.A1(n_3653),
.A2(n_3146),
.B1(n_3180),
.B2(n_3158),
.Y(n_3707)
);

INVx2_ASAP7_75t_L g3708 ( 
.A(n_3630),
.Y(n_3708)
);

AND4x1_ASAP7_75t_L g3709 ( 
.A(n_3656),
.B(n_3316),
.C(n_3363),
.D(n_3327),
.Y(n_3709)
);

INVx2_ASAP7_75t_L g3710 ( 
.A(n_3667),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3681),
.Y(n_3711)
);

INVx1_ASAP7_75t_L g3712 ( 
.A(n_3671),
.Y(n_3712)
);

HB1xp67_ASAP7_75t_L g3713 ( 
.A(n_3673),
.Y(n_3713)
);

INVx2_ASAP7_75t_L g3714 ( 
.A(n_3674),
.Y(n_3714)
);

AND2x2_ASAP7_75t_L g3715 ( 
.A(n_3672),
.B(n_3620),
.Y(n_3715)
);

OR2x2_ASAP7_75t_L g3716 ( 
.A(n_3661),
.B(n_3619),
.Y(n_3716)
);

NAND2xp5_ASAP7_75t_L g3717 ( 
.A(n_3684),
.B(n_3626),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3687),
.Y(n_3718)
);

AND2x2_ASAP7_75t_L g3719 ( 
.A(n_3664),
.B(n_3669),
.Y(n_3719)
);

INVx1_ASAP7_75t_SL g3720 ( 
.A(n_3666),
.Y(n_3720)
);

INVx1_ASAP7_75t_L g3721 ( 
.A(n_3692),
.Y(n_3721)
);

AND2x2_ASAP7_75t_L g3722 ( 
.A(n_3685),
.B(n_3604),
.Y(n_3722)
);

AND2x4_ASAP7_75t_SL g3723 ( 
.A(n_3688),
.B(n_3651),
.Y(n_3723)
);

OR2x2_ASAP7_75t_L g3724 ( 
.A(n_3702),
.B(n_3602),
.Y(n_3724)
);

INVxp67_ASAP7_75t_L g3725 ( 
.A(n_3690),
.Y(n_3725)
);

AND2x4_ASAP7_75t_SL g3726 ( 
.A(n_3688),
.B(n_3650),
.Y(n_3726)
);

AND2x4_ASAP7_75t_L g3727 ( 
.A(n_3677),
.B(n_3627),
.Y(n_3727)
);

INVx3_ASAP7_75t_L g3728 ( 
.A(n_3663),
.Y(n_3728)
);

HB1xp67_ASAP7_75t_L g3729 ( 
.A(n_3665),
.Y(n_3729)
);

INVx1_ASAP7_75t_L g3730 ( 
.A(n_3697),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3699),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_3700),
.Y(n_3732)
);

OR2x2_ASAP7_75t_L g3733 ( 
.A(n_3679),
.B(n_3603),
.Y(n_3733)
);

AND2x2_ASAP7_75t_L g3734 ( 
.A(n_3686),
.B(n_3646),
.Y(n_3734)
);

INVx2_ASAP7_75t_SL g3735 ( 
.A(n_3696),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3704),
.Y(n_3736)
);

AND2x4_ASAP7_75t_L g3737 ( 
.A(n_3693),
.B(n_3662),
.Y(n_3737)
);

OR2x2_ASAP7_75t_L g3738 ( 
.A(n_3680),
.B(n_3639),
.Y(n_3738)
);

INVx5_ASAP7_75t_SL g3739 ( 
.A(n_3691),
.Y(n_3739)
);

AND2x2_ASAP7_75t_L g3740 ( 
.A(n_3695),
.B(n_3705),
.Y(n_3740)
);

OAI222xp33_ASAP7_75t_L g3741 ( 
.A1(n_3668),
.A2(n_3637),
.B1(n_3641),
.B2(n_3640),
.C1(n_3240),
.C2(n_3267),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3703),
.Y(n_3742)
);

INVx2_ASAP7_75t_L g3743 ( 
.A(n_3708),
.Y(n_3743)
);

AOI22xp5_ASAP7_75t_L g3744 ( 
.A1(n_3683),
.A2(n_3025),
.B1(n_3234),
.B2(n_3152),
.Y(n_3744)
);

INVx1_ASAP7_75t_SL g3745 ( 
.A(n_3678),
.Y(n_3745)
);

AOI222xp33_ASAP7_75t_L g3746 ( 
.A1(n_3682),
.A2(n_3097),
.B1(n_3212),
.B2(n_3402),
.C1(n_3183),
.C2(n_3194),
.Y(n_3746)
);

AO221x2_ASAP7_75t_L g3747 ( 
.A1(n_3707),
.A2(n_3185),
.B1(n_3044),
.B2(n_3020),
.C(n_3291),
.Y(n_3747)
);

AND4x1_ASAP7_75t_L g3748 ( 
.A(n_3670),
.B(n_3396),
.C(n_3248),
.D(n_3249),
.Y(n_3748)
);

OR2x6_ASAP7_75t_SL g3749 ( 
.A(n_3675),
.B(n_3283),
.Y(n_3749)
);

AND2x2_ASAP7_75t_L g3750 ( 
.A(n_3695),
.B(n_3694),
.Y(n_3750)
);

OAI21xp33_ASAP7_75t_SL g3751 ( 
.A1(n_3698),
.A2(n_3345),
.B(n_3341),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3676),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_3676),
.Y(n_3753)
);

INVx1_ASAP7_75t_L g3754 ( 
.A(n_3701),
.Y(n_3754)
);

BUFx3_ASAP7_75t_L g3755 ( 
.A(n_3720),
.Y(n_3755)
);

INVx2_ASAP7_75t_L g3756 ( 
.A(n_3710),
.Y(n_3756)
);

OR2x2_ASAP7_75t_L g3757 ( 
.A(n_3738),
.B(n_3706),
.Y(n_3757)
);

AND2x2_ASAP7_75t_L g3758 ( 
.A(n_3739),
.B(n_3689),
.Y(n_3758)
);

BUFx2_ASAP7_75t_L g3759 ( 
.A(n_3719),
.Y(n_3759)
);

INVx1_ASAP7_75t_L g3760 ( 
.A(n_3729),
.Y(n_3760)
);

BUFx2_ASAP7_75t_L g3761 ( 
.A(n_3735),
.Y(n_3761)
);

NAND3xp33_ASAP7_75t_L g3762 ( 
.A(n_3748),
.B(n_3709),
.C(n_3207),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_L g3763 ( 
.A(n_3711),
.B(n_3712),
.Y(n_3763)
);

NAND2xp67_ASAP7_75t_L g3764 ( 
.A(n_3723),
.B(n_3726),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_3717),
.Y(n_3765)
);

AND2x2_ASAP7_75t_L g3766 ( 
.A(n_3750),
.B(n_3728),
.Y(n_3766)
);

NOR2x1_ASAP7_75t_L g3767 ( 
.A(n_3737),
.B(n_3204),
.Y(n_3767)
);

OR2x2_ASAP7_75t_L g3768 ( 
.A(n_3714),
.B(n_3308),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_3713),
.Y(n_3769)
);

INVx2_ASAP7_75t_L g3770 ( 
.A(n_3716),
.Y(n_3770)
);

AND2x2_ASAP7_75t_L g3771 ( 
.A(n_3725),
.B(n_3291),
.Y(n_3771)
);

INVx2_ASAP7_75t_L g3772 ( 
.A(n_3733),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_3718),
.Y(n_3773)
);

INVx1_ASAP7_75t_L g3774 ( 
.A(n_3721),
.Y(n_3774)
);

INVx1_ASAP7_75t_L g3775 ( 
.A(n_3730),
.Y(n_3775)
);

AND2x4_ASAP7_75t_L g3776 ( 
.A(n_3722),
.B(n_3225),
.Y(n_3776)
);

NAND2x1p5_ASAP7_75t_L g3777 ( 
.A(n_3744),
.B(n_3004),
.Y(n_3777)
);

INVx1_ASAP7_75t_L g3778 ( 
.A(n_3731),
.Y(n_3778)
);

AND2x2_ASAP7_75t_L g3779 ( 
.A(n_3745),
.B(n_3291),
.Y(n_3779)
);

AND2x2_ASAP7_75t_L g3780 ( 
.A(n_3715),
.B(n_3297),
.Y(n_3780)
);

INVx2_ASAP7_75t_L g3781 ( 
.A(n_3743),
.Y(n_3781)
);

INVx1_ASAP7_75t_L g3782 ( 
.A(n_3732),
.Y(n_3782)
);

AND2x2_ASAP7_75t_L g3783 ( 
.A(n_3761),
.B(n_3749),
.Y(n_3783)
);

INVx1_ASAP7_75t_L g3784 ( 
.A(n_3769),
.Y(n_3784)
);

INVx4_ASAP7_75t_L g3785 ( 
.A(n_3755),
.Y(n_3785)
);

AND2x2_ASAP7_75t_L g3786 ( 
.A(n_3758),
.B(n_3727),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3769),
.Y(n_3787)
);

AND2x2_ASAP7_75t_L g3788 ( 
.A(n_3766),
.B(n_3727),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3756),
.Y(n_3789)
);

INVx2_ASAP7_75t_L g3790 ( 
.A(n_3772),
.Y(n_3790)
);

AND2x2_ASAP7_75t_L g3791 ( 
.A(n_3759),
.B(n_3747),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_L g3792 ( 
.A(n_3760),
.B(n_3746),
.Y(n_3792)
);

INVx2_ASAP7_75t_L g3793 ( 
.A(n_3770),
.Y(n_3793)
);

NAND2x1p5_ASAP7_75t_L g3794 ( 
.A(n_3767),
.B(n_3358),
.Y(n_3794)
);

INVx2_ASAP7_75t_L g3795 ( 
.A(n_3757),
.Y(n_3795)
);

AND2x4_ASAP7_75t_L g3796 ( 
.A(n_3771),
.B(n_3740),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_L g3797 ( 
.A(n_3765),
.B(n_3736),
.Y(n_3797)
);

INVxp67_ASAP7_75t_L g3798 ( 
.A(n_3779),
.Y(n_3798)
);

OAI21xp33_ASAP7_75t_L g3799 ( 
.A1(n_3764),
.A2(n_3754),
.B(n_3753),
.Y(n_3799)
);

INVx1_ASAP7_75t_L g3800 ( 
.A(n_3763),
.Y(n_3800)
);

AND2x2_ASAP7_75t_L g3801 ( 
.A(n_3780),
.B(n_3734),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3773),
.Y(n_3802)
);

INVx2_ASAP7_75t_L g3803 ( 
.A(n_3781),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_L g3804 ( 
.A(n_3762),
.B(n_3751),
.Y(n_3804)
);

AND2x2_ASAP7_75t_L g3805 ( 
.A(n_3776),
.B(n_3724),
.Y(n_3805)
);

AND2x2_ASAP7_75t_L g3806 ( 
.A(n_3776),
.B(n_3742),
.Y(n_3806)
);

INVx2_ASAP7_75t_L g3807 ( 
.A(n_3785),
.Y(n_3807)
);

INVx1_ASAP7_75t_L g3808 ( 
.A(n_3790),
.Y(n_3808)
);

INVx2_ASAP7_75t_SL g3809 ( 
.A(n_3796),
.Y(n_3809)
);

INVx1_ASAP7_75t_SL g3810 ( 
.A(n_3783),
.Y(n_3810)
);

INVx2_ASAP7_75t_SL g3811 ( 
.A(n_3796),
.Y(n_3811)
);

INVx2_ASAP7_75t_L g3812 ( 
.A(n_3795),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3789),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3789),
.Y(n_3814)
);

INVx1_ASAP7_75t_L g3815 ( 
.A(n_3793),
.Y(n_3815)
);

INVx1_ASAP7_75t_SL g3816 ( 
.A(n_3791),
.Y(n_3816)
);

INVx1_ASAP7_75t_L g3817 ( 
.A(n_3784),
.Y(n_3817)
);

NAND2xp5_ASAP7_75t_L g3818 ( 
.A(n_3800),
.B(n_3774),
.Y(n_3818)
);

OAI31xp33_ASAP7_75t_SL g3819 ( 
.A1(n_3799),
.A2(n_3752),
.A3(n_3778),
.B(n_3775),
.Y(n_3819)
);

AND2x2_ASAP7_75t_L g3820 ( 
.A(n_3788),
.B(n_3777),
.Y(n_3820)
);

INVx4_ASAP7_75t_L g3821 ( 
.A(n_3803),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_3787),
.Y(n_3822)
);

INVx3_ASAP7_75t_L g3823 ( 
.A(n_3806),
.Y(n_3823)
);

NOR2xp33_ASAP7_75t_L g3824 ( 
.A(n_3792),
.B(n_3741),
.Y(n_3824)
);

OR2x2_ASAP7_75t_L g3825 ( 
.A(n_3797),
.B(n_3768),
.Y(n_3825)
);

INVxp67_ASAP7_75t_L g3826 ( 
.A(n_3786),
.Y(n_3826)
);

NOR2xp33_ASAP7_75t_L g3827 ( 
.A(n_3798),
.B(n_3775),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_3802),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_L g3829 ( 
.A(n_3805),
.B(n_3782),
.Y(n_3829)
);

INVx2_ASAP7_75t_L g3830 ( 
.A(n_3794),
.Y(n_3830)
);

INVx1_ASAP7_75t_L g3831 ( 
.A(n_3801),
.Y(n_3831)
);

NAND2xp5_ASAP7_75t_L g3832 ( 
.A(n_3807),
.B(n_3782),
.Y(n_3832)
);

AND2x4_ASAP7_75t_L g3833 ( 
.A(n_3809),
.B(n_3804),
.Y(n_3833)
);

AND2x4_ASAP7_75t_L g3834 ( 
.A(n_3811),
.B(n_3184),
.Y(n_3834)
);

NAND2xp5_ASAP7_75t_L g3835 ( 
.A(n_3816),
.B(n_3397),
.Y(n_3835)
);

AND2x2_ASAP7_75t_L g3836 ( 
.A(n_3810),
.B(n_3181),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_3821),
.B(n_3397),
.Y(n_3837)
);

AND2x2_ASAP7_75t_L g3838 ( 
.A(n_3820),
.B(n_3117),
.Y(n_3838)
);

NAND2xp5_ASAP7_75t_L g3839 ( 
.A(n_3821),
.B(n_581),
.Y(n_3839)
);

INVx2_ASAP7_75t_L g3840 ( 
.A(n_3812),
.Y(n_3840)
);

OR2x2_ASAP7_75t_L g3841 ( 
.A(n_3808),
.B(n_581),
.Y(n_3841)
);

HB1xp67_ASAP7_75t_L g3842 ( 
.A(n_3815),
.Y(n_3842)
);

AND2x2_ASAP7_75t_L g3843 ( 
.A(n_3823),
.B(n_3230),
.Y(n_3843)
);

OR2x2_ASAP7_75t_L g3844 ( 
.A(n_3829),
.B(n_582),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_3813),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_3814),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_L g3847 ( 
.A(n_3826),
.B(n_582),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_L g3848 ( 
.A(n_3824),
.B(n_583),
.Y(n_3848)
);

INVx2_ASAP7_75t_L g3849 ( 
.A(n_3831),
.Y(n_3849)
);

NAND2xp5_ASAP7_75t_L g3850 ( 
.A(n_3827),
.B(n_583),
.Y(n_3850)
);

AND2x2_ASAP7_75t_L g3851 ( 
.A(n_3830),
.B(n_3386),
.Y(n_3851)
);

INVx2_ASAP7_75t_L g3852 ( 
.A(n_3825),
.Y(n_3852)
);

INVx2_ASAP7_75t_L g3853 ( 
.A(n_3828),
.Y(n_3853)
);

AND2x2_ASAP7_75t_L g3854 ( 
.A(n_3819),
.B(n_3365),
.Y(n_3854)
);

OR2x2_ASAP7_75t_L g3855 ( 
.A(n_3818),
.B(n_584),
.Y(n_3855)
);

OAI21xp33_ASAP7_75t_L g3856 ( 
.A1(n_3833),
.A2(n_3822),
.B(n_3817),
.Y(n_3856)
);

INVx1_ASAP7_75t_SL g3857 ( 
.A(n_3838),
.Y(n_3857)
);

AND2x4_ASAP7_75t_L g3858 ( 
.A(n_3834),
.B(n_3362),
.Y(n_3858)
);

INVx1_ASAP7_75t_L g3859 ( 
.A(n_3842),
.Y(n_3859)
);

NAND5xp2_ASAP7_75t_SL g3860 ( 
.A(n_3854),
.B(n_587),
.C(n_585),
.D(n_586),
.E(n_588),
.Y(n_3860)
);

AOI322xp5_ASAP7_75t_L g3861 ( 
.A1(n_3849),
.A2(n_3228),
.A3(n_3155),
.B1(n_3359),
.B2(n_3370),
.C1(n_3366),
.C2(n_3071),
.Y(n_3861)
);

AND2x2_ASAP7_75t_L g3862 ( 
.A(n_3836),
.B(n_588),
.Y(n_3862)
);

AND2x2_ASAP7_75t_SL g3863 ( 
.A(n_3841),
.B(n_3270),
.Y(n_3863)
);

OAI21xp33_ASAP7_75t_SL g3864 ( 
.A1(n_3832),
.A2(n_3395),
.B(n_3394),
.Y(n_3864)
);

INVx1_ASAP7_75t_L g3865 ( 
.A(n_3847),
.Y(n_3865)
);

AOI22xp33_ASAP7_75t_L g3866 ( 
.A1(n_3852),
.A2(n_3019),
.B1(n_3255),
.B2(n_3270),
.Y(n_3866)
);

NAND2xp5_ASAP7_75t_L g3867 ( 
.A(n_3834),
.B(n_589),
.Y(n_3867)
);

OAI21xp5_ASAP7_75t_SL g3868 ( 
.A1(n_3835),
.A2(n_589),
.B(n_591),
.Y(n_3868)
);

INVx1_ASAP7_75t_L g3869 ( 
.A(n_3844),
.Y(n_3869)
);

NAND2x1_ASAP7_75t_SL g3870 ( 
.A(n_3853),
.B(n_591),
.Y(n_3870)
);

AOI22xp33_ASAP7_75t_L g3871 ( 
.A1(n_3851),
.A2(n_3019),
.B1(n_3010),
.B2(n_3051),
.Y(n_3871)
);

NAND2xp33_ASAP7_75t_SL g3872 ( 
.A(n_3855),
.B(n_3055),
.Y(n_3872)
);

INVx3_ASAP7_75t_L g3873 ( 
.A(n_3843),
.Y(n_3873)
);

INVxp33_ASAP7_75t_L g3874 ( 
.A(n_3850),
.Y(n_3874)
);

INVx1_ASAP7_75t_L g3875 ( 
.A(n_3837),
.Y(n_3875)
);

NAND2xp5_ASAP7_75t_SL g3876 ( 
.A(n_3846),
.B(n_3017),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3845),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3845),
.Y(n_3878)
);

AND2x2_ASAP7_75t_L g3879 ( 
.A(n_3838),
.B(n_593),
.Y(n_3879)
);

OR2x2_ASAP7_75t_L g3880 ( 
.A(n_3839),
.B(n_593),
.Y(n_3880)
);

NAND2xp5_ASAP7_75t_L g3881 ( 
.A(n_3833),
.B(n_594),
.Y(n_3881)
);

OAI21xp5_ASAP7_75t_L g3882 ( 
.A1(n_3848),
.A2(n_3384),
.B(n_3357),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_L g3883 ( 
.A(n_3833),
.B(n_594),
.Y(n_3883)
);

O2A1O1Ixp33_ASAP7_75t_L g3884 ( 
.A1(n_3848),
.A2(n_597),
.B(n_595),
.C(n_596),
.Y(n_3884)
);

INVx2_ASAP7_75t_L g3885 ( 
.A(n_3840),
.Y(n_3885)
);

NAND2xp5_ASAP7_75t_L g3886 ( 
.A(n_3833),
.B(n_596),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3881),
.Y(n_3887)
);

INVxp67_ASAP7_75t_L g3888 ( 
.A(n_3879),
.Y(n_3888)
);

AOI21xp5_ASAP7_75t_L g3889 ( 
.A1(n_3883),
.A2(n_3314),
.B(n_3339),
.Y(n_3889)
);

AND2x2_ASAP7_75t_L g3890 ( 
.A(n_3857),
.B(n_596),
.Y(n_3890)
);

AND2x2_ASAP7_75t_L g3891 ( 
.A(n_3862),
.B(n_598),
.Y(n_3891)
);

INVx1_ASAP7_75t_SL g3892 ( 
.A(n_3867),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_SL g3893 ( 
.A(n_3885),
.B(n_2950),
.Y(n_3893)
);

AND2x2_ASAP7_75t_L g3894 ( 
.A(n_3873),
.B(n_599),
.Y(n_3894)
);

INVx1_ASAP7_75t_L g3895 ( 
.A(n_3886),
.Y(n_3895)
);

NAND2xp5_ASAP7_75t_L g3896 ( 
.A(n_3859),
.B(n_599),
.Y(n_3896)
);

INVx1_ASAP7_75t_L g3897 ( 
.A(n_3880),
.Y(n_3897)
);

INVx1_ASAP7_75t_L g3898 ( 
.A(n_3870),
.Y(n_3898)
);

AND2x4_ASAP7_75t_L g3899 ( 
.A(n_3869),
.B(n_600),
.Y(n_3899)
);

NOR2xp33_ASAP7_75t_L g3900 ( 
.A(n_3856),
.B(n_601),
.Y(n_3900)
);

OR2x2_ASAP7_75t_L g3901 ( 
.A(n_3875),
.B(n_601),
.Y(n_3901)
);

INVx2_ASAP7_75t_L g3902 ( 
.A(n_3858),
.Y(n_3902)
);

INVx1_ASAP7_75t_L g3903 ( 
.A(n_3877),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_L g3904 ( 
.A(n_3864),
.B(n_602),
.Y(n_3904)
);

NAND2xp5_ASAP7_75t_L g3905 ( 
.A(n_3868),
.B(n_602),
.Y(n_3905)
);

INVx1_ASAP7_75t_L g3906 ( 
.A(n_3878),
.Y(n_3906)
);

OR2x6_ASAP7_75t_L g3907 ( 
.A(n_3884),
.B(n_3101),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_3863),
.Y(n_3908)
);

NOR2xp33_ASAP7_75t_L g3909 ( 
.A(n_3874),
.B(n_3876),
.Y(n_3909)
);

INVx1_ASAP7_75t_SL g3910 ( 
.A(n_3872),
.Y(n_3910)
);

INVxp33_ASAP7_75t_L g3911 ( 
.A(n_3865),
.Y(n_3911)
);

INVx1_ASAP7_75t_L g3912 ( 
.A(n_3894),
.Y(n_3912)
);

NOR2xp33_ASAP7_75t_L g3913 ( 
.A(n_3898),
.B(n_3871),
.Y(n_3913)
);

NOR2xp33_ASAP7_75t_L g3914 ( 
.A(n_3910),
.B(n_3882),
.Y(n_3914)
);

NAND2xp5_ASAP7_75t_SL g3915 ( 
.A(n_3904),
.B(n_3866),
.Y(n_3915)
);

AND2x2_ASAP7_75t_L g3916 ( 
.A(n_3891),
.B(n_3860),
.Y(n_3916)
);

NAND2xp5_ASAP7_75t_L g3917 ( 
.A(n_3899),
.B(n_3861),
.Y(n_3917)
);

AOI211xp5_ASAP7_75t_L g3918 ( 
.A1(n_3900),
.A2(n_604),
.B(n_602),
.C(n_603),
.Y(n_3918)
);

HB1xp67_ASAP7_75t_L g3919 ( 
.A(n_3902),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_3901),
.Y(n_3920)
);

HB1xp67_ASAP7_75t_L g3921 ( 
.A(n_3897),
.Y(n_3921)
);

INVx2_ASAP7_75t_L g3922 ( 
.A(n_3907),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_3896),
.Y(n_3923)
);

NOR2xp33_ASAP7_75t_L g3924 ( 
.A(n_3888),
.B(n_603),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3905),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3908),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3903),
.Y(n_3927)
);

INVx1_ASAP7_75t_SL g3928 ( 
.A(n_3893),
.Y(n_3928)
);

OAI22xp5_ASAP7_75t_L g3929 ( 
.A1(n_3911),
.A2(n_3083),
.B1(n_3096),
.B2(n_3067),
.Y(n_3929)
);

INVx1_ASAP7_75t_L g3930 ( 
.A(n_3906),
.Y(n_3930)
);

AND2x4_ASAP7_75t_L g3931 ( 
.A(n_3907),
.B(n_3098),
.Y(n_3931)
);

AND2x2_ASAP7_75t_L g3932 ( 
.A(n_3892),
.B(n_605),
.Y(n_3932)
);

NAND2xp5_ASAP7_75t_L g3933 ( 
.A(n_3889),
.B(n_605),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_L g3934 ( 
.A(n_3887),
.B(n_606),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3895),
.Y(n_3935)
);

CKINVDCx16_ASAP7_75t_R g3936 ( 
.A(n_3909),
.Y(n_3936)
);

NAND2xp5_ASAP7_75t_L g3937 ( 
.A(n_3890),
.B(n_607),
.Y(n_3937)
);

NAND4xp25_ASAP7_75t_L g3938 ( 
.A(n_3913),
.B(n_610),
.C(n_608),
.D(n_609),
.Y(n_3938)
);

NAND3xp33_ASAP7_75t_L g3939 ( 
.A(n_3919),
.B(n_609),
.C(n_610),
.Y(n_3939)
);

NAND2xp5_ASAP7_75t_L g3940 ( 
.A(n_3936),
.B(n_610),
.Y(n_3940)
);

XOR2x2_ASAP7_75t_L g3941 ( 
.A(n_3916),
.B(n_611),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3932),
.Y(n_3942)
);

NAND4xp75_ASAP7_75t_L g3943 ( 
.A(n_3924),
.B(n_614),
.C(n_612),
.D(n_613),
.Y(n_3943)
);

NAND5xp2_ASAP7_75t_L g3944 ( 
.A(n_3914),
.B(n_616),
.C(n_614),
.D(n_615),
.E(n_617),
.Y(n_3944)
);

AND2x4_ASAP7_75t_L g3945 ( 
.A(n_3922),
.B(n_3100),
.Y(n_3945)
);

HB1xp67_ASAP7_75t_L g3946 ( 
.A(n_3921),
.Y(n_3946)
);

OAI22xp33_ASAP7_75t_L g3947 ( 
.A1(n_3933),
.A2(n_3103),
.B1(n_2978),
.B2(n_2980),
.Y(n_3947)
);

OAI211xp5_ASAP7_75t_L g3948 ( 
.A1(n_3918),
.A2(n_618),
.B(n_616),
.C(n_617),
.Y(n_3948)
);

NOR2xp33_ASAP7_75t_L g3949 ( 
.A(n_3937),
.B(n_619),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3934),
.Y(n_3950)
);

NOR3xp33_ASAP7_75t_L g3951 ( 
.A(n_3926),
.B(n_619),
.C(n_620),
.Y(n_3951)
);

AND2x2_ASAP7_75t_L g3952 ( 
.A(n_3912),
.B(n_620),
.Y(n_3952)
);

NOR3xp33_ASAP7_75t_L g3953 ( 
.A(n_3935),
.B(n_620),
.C(n_621),
.Y(n_3953)
);

NAND3x1_ASAP7_75t_L g3954 ( 
.A(n_3917),
.B(n_621),
.C(n_622),
.Y(n_3954)
);

OAI22xp5_ASAP7_75t_L g3955 ( 
.A1(n_3928),
.A2(n_3114),
.B1(n_3132),
.B2(n_3128),
.Y(n_3955)
);

AOI22xp33_ASAP7_75t_L g3956 ( 
.A1(n_3931),
.A2(n_3114),
.B1(n_3128),
.B2(n_3275),
.Y(n_3956)
);

AOI21xp33_ASAP7_75t_L g3957 ( 
.A1(n_3927),
.A2(n_623),
.B(n_624),
.Y(n_3957)
);

NAND3xp33_ASAP7_75t_L g3958 ( 
.A(n_3930),
.B(n_623),
.C(n_624),
.Y(n_3958)
);

NOR4xp25_ASAP7_75t_L g3959 ( 
.A(n_3925),
.B(n_626),
.C(n_624),
.D(n_625),
.Y(n_3959)
);

NOR3x1_ASAP7_75t_L g3960 ( 
.A(n_3915),
.B(n_625),
.C(n_626),
.Y(n_3960)
);

NAND4xp25_ASAP7_75t_L g3961 ( 
.A(n_3920),
.B(n_628),
.C(n_625),
.D(n_627),
.Y(n_3961)
);

OR3x1_ASAP7_75t_L g3962 ( 
.A(n_3944),
.B(n_3923),
.C(n_3929),
.Y(n_3962)
);

AND2x4_ASAP7_75t_L g3963 ( 
.A(n_3945),
.B(n_629),
.Y(n_3963)
);

OAI22xp5_ASAP7_75t_L g3964 ( 
.A1(n_3940),
.A2(n_3015),
.B1(n_3040),
.B2(n_2983),
.Y(n_3964)
);

CKINVDCx20_ASAP7_75t_R g3965 ( 
.A(n_3941),
.Y(n_3965)
);

OAI221xp5_ASAP7_75t_L g3966 ( 
.A1(n_3959),
.A2(n_632),
.B1(n_630),
.B2(n_631),
.C(n_633),
.Y(n_3966)
);

A2O1A1Ixp33_ASAP7_75t_L g3967 ( 
.A1(n_3949),
.A2(n_3280),
.B(n_632),
.C(n_630),
.Y(n_3967)
);

NOR2xp33_ASAP7_75t_L g3968 ( 
.A(n_3939),
.B(n_630),
.Y(n_3968)
);

INVx1_ASAP7_75t_L g3969 ( 
.A(n_3946),
.Y(n_3969)
);

OAI211xp5_ASAP7_75t_L g3970 ( 
.A1(n_3938),
.A2(n_634),
.B(n_631),
.C(n_633),
.Y(n_3970)
);

AOI21xp33_ASAP7_75t_L g3971 ( 
.A1(n_3948),
.A2(n_3958),
.B(n_3952),
.Y(n_3971)
);

OAI21xp5_ASAP7_75t_L g3972 ( 
.A1(n_3954),
.A2(n_631),
.B(n_634),
.Y(n_3972)
);

OAI221xp5_ASAP7_75t_L g3973 ( 
.A1(n_3961),
.A2(n_635),
.B1(n_636),
.B2(n_3015),
.C(n_2983),
.Y(n_3973)
);

AOI211xp5_ASAP7_75t_SL g3974 ( 
.A1(n_3957),
.A2(n_635),
.B(n_636),
.C(n_692),
.Y(n_3974)
);

OAI221xp5_ASAP7_75t_L g3975 ( 
.A1(n_3951),
.A2(n_3059),
.B1(n_3040),
.B2(n_3093),
.C(n_3092),
.Y(n_3975)
);

O2A1O1Ixp33_ASAP7_75t_L g3976 ( 
.A1(n_3953),
.A2(n_695),
.B(n_693),
.C(n_694),
.Y(n_3976)
);

AOI211xp5_ASAP7_75t_SL g3977 ( 
.A1(n_3942),
.A2(n_700),
.B(n_698),
.C(n_699),
.Y(n_3977)
);

NOR2xp33_ASAP7_75t_L g3978 ( 
.A(n_3943),
.B(n_701),
.Y(n_3978)
);

OAI31xp33_ASAP7_75t_L g3979 ( 
.A1(n_3947),
.A2(n_704),
.A3(n_702),
.B(n_703),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_SL g3980 ( 
.A(n_3950),
.B(n_3059),
.Y(n_3980)
);

O2A1O1Ixp33_ASAP7_75t_L g3981 ( 
.A1(n_3960),
.A2(n_705),
.B(n_703),
.C(n_704),
.Y(n_3981)
);

OAI21xp33_ASAP7_75t_SL g3982 ( 
.A1(n_3956),
.A2(n_705),
.B(n_706),
.Y(n_3982)
);

NAND3xp33_ASAP7_75t_L g3983 ( 
.A(n_3955),
.B(n_706),
.C(n_708),
.Y(n_3983)
);

OAI211xp5_ASAP7_75t_SL g3984 ( 
.A1(n_3974),
.A2(n_712),
.B(n_709),
.C(n_711),
.Y(n_3984)
);

CKINVDCx20_ASAP7_75t_R g3985 ( 
.A(n_3965),
.Y(n_3985)
);

AOI211xp5_ASAP7_75t_SL g3986 ( 
.A1(n_3970),
.A2(n_3971),
.B(n_3978),
.C(n_3966),
.Y(n_3986)
);

INVxp67_ASAP7_75t_SL g3987 ( 
.A(n_3981),
.Y(n_3987)
);

AOI211xp5_ASAP7_75t_SL g3988 ( 
.A1(n_3968),
.A2(n_713),
.B(n_709),
.C(n_711),
.Y(n_3988)
);

AOI221xp5_ASAP7_75t_SL g3989 ( 
.A1(n_3973),
.A2(n_3104),
.B1(n_3108),
.B2(n_3093),
.C(n_3092),
.Y(n_3989)
);

AOI221xp5_ASAP7_75t_L g3990 ( 
.A1(n_3976),
.A2(n_716),
.B1(n_714),
.B2(n_715),
.C(n_717),
.Y(n_3990)
);

OAI32xp33_ASAP7_75t_L g3991 ( 
.A1(n_3969),
.A2(n_718),
.A3(n_714),
.B1(n_717),
.B2(n_719),
.Y(n_3991)
);

AOI22xp5_ASAP7_75t_L g3992 ( 
.A1(n_3962),
.A2(n_3166),
.B1(n_3165),
.B2(n_3075),
.Y(n_3992)
);

AOI221xp5_ASAP7_75t_L g3993 ( 
.A1(n_3972),
.A2(n_721),
.B1(n_719),
.B2(n_720),
.C(n_722),
.Y(n_3993)
);

AOI22xp33_ASAP7_75t_SL g3994 ( 
.A1(n_3963),
.A2(n_3075),
.B1(n_3050),
.B2(n_723),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_L g3995 ( 
.A(n_3963),
.B(n_724),
.Y(n_3995)
);

OAI211xp5_ASAP7_75t_L g3996 ( 
.A1(n_3979),
.A2(n_727),
.B(n_725),
.C(n_726),
.Y(n_3996)
);

NAND5xp2_ASAP7_75t_L g3997 ( 
.A(n_3977),
.B(n_730),
.C(n_728),
.D(n_729),
.E(n_731),
.Y(n_3997)
);

OAI21xp5_ASAP7_75t_L g3998 ( 
.A1(n_3982),
.A2(n_728),
.B(n_730),
.Y(n_3998)
);

OAI211xp5_ASAP7_75t_L g3999 ( 
.A1(n_3983),
.A2(n_734),
.B(n_731),
.C(n_733),
.Y(n_3999)
);

NAND3x1_ASAP7_75t_L g4000 ( 
.A(n_3995),
.B(n_3980),
.C(n_3967),
.Y(n_4000)
);

NAND3xp33_ASAP7_75t_L g4001 ( 
.A(n_3986),
.B(n_3964),
.C(n_3975),
.Y(n_4001)
);

AOI22xp33_ASAP7_75t_L g4002 ( 
.A1(n_3987),
.A2(n_3075),
.B1(n_3050),
.B2(n_736),
.Y(n_4002)
);

AND2x2_ASAP7_75t_SL g4003 ( 
.A(n_3990),
.B(n_737),
.Y(n_4003)
);

AOI321xp33_ASAP7_75t_L g4004 ( 
.A1(n_3996),
.A2(n_739),
.A3(n_741),
.B1(n_737),
.B2(n_738),
.C(n_740),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_L g4005 ( 
.A(n_3989),
.B(n_739),
.Y(n_4005)
);

NAND3xp33_ASAP7_75t_L g4006 ( 
.A(n_3993),
.B(n_741),
.C(n_742),
.Y(n_4006)
);

OAI22xp33_ASAP7_75t_L g4007 ( 
.A1(n_3988),
.A2(n_744),
.B1(n_742),
.B2(n_743),
.Y(n_4007)
);

NOR3xp33_ASAP7_75t_L g4008 ( 
.A(n_3984),
.B(n_3999),
.C(n_3991),
.Y(n_4008)
);

AND2x2_ASAP7_75t_L g4009 ( 
.A(n_3998),
.B(n_744),
.Y(n_4009)
);

AOI21xp5_ASAP7_75t_L g4010 ( 
.A1(n_3997),
.A2(n_745),
.B(n_746),
.Y(n_4010)
);

NOR2x1p5_ASAP7_75t_L g4011 ( 
.A(n_3994),
.B(n_747),
.Y(n_4011)
);

NAND2x1p5_ASAP7_75t_L g4012 ( 
.A(n_3992),
.B(n_748),
.Y(n_4012)
);

AOI22xp5_ASAP7_75t_L g4013 ( 
.A1(n_3985),
.A2(n_3075),
.B1(n_3050),
.B2(n_751),
.Y(n_4013)
);

AOI21xp33_ASAP7_75t_SL g4014 ( 
.A1(n_3995),
.A2(n_749),
.B(n_750),
.Y(n_4014)
);

NOR4xp25_ASAP7_75t_L g4015 ( 
.A(n_4001),
.B(n_754),
.C(n_752),
.D(n_753),
.Y(n_4015)
);

NAND2xp5_ASAP7_75t_L g4016 ( 
.A(n_4010),
.B(n_757),
.Y(n_4016)
);

NOR2xp33_ASAP7_75t_SL g4017 ( 
.A(n_4005),
.B(n_757),
.Y(n_4017)
);

AOI322xp5_ASAP7_75t_L g4018 ( 
.A1(n_4007),
.A2(n_758),
.A3(n_759),
.B1(n_760),
.B2(n_761),
.C1(n_762),
.C2(n_763),
.Y(n_4018)
);

NAND5xp2_ASAP7_75t_L g4019 ( 
.A(n_4004),
.B(n_760),
.C(n_758),
.D(n_759),
.E(n_763),
.Y(n_4019)
);

INVx2_ASAP7_75t_L g4020 ( 
.A(n_4012),
.Y(n_4020)
);

NAND4xp25_ASAP7_75t_L g4021 ( 
.A(n_4008),
.B(n_766),
.C(n_764),
.D(n_765),
.Y(n_4021)
);

AND2x2_ASAP7_75t_L g4022 ( 
.A(n_4009),
.B(n_766),
.Y(n_4022)
);

AOI221xp5_ASAP7_75t_L g4023 ( 
.A1(n_4014),
.A2(n_4006),
.B1(n_4002),
.B2(n_4013),
.C(n_4000),
.Y(n_4023)
);

AOI22xp33_ASAP7_75t_L g4024 ( 
.A1(n_4003),
.A2(n_4011),
.B1(n_3050),
.B2(n_768),
.Y(n_4024)
);

NAND2xp5_ASAP7_75t_SL g4025 ( 
.A(n_4005),
.B(n_767),
.Y(n_4025)
);

BUFx6f_ASAP7_75t_L g4026 ( 
.A(n_4020),
.Y(n_4026)
);

NOR2xp33_ASAP7_75t_L g4027 ( 
.A(n_4016),
.B(n_768),
.Y(n_4027)
);

AOI211xp5_ASAP7_75t_L g4028 ( 
.A1(n_4021),
.A2(n_772),
.B(n_770),
.C(n_771),
.Y(n_4028)
);

AOI221xp5_ASAP7_75t_L g4029 ( 
.A1(n_4015),
.A2(n_773),
.B1(n_770),
.B2(n_771),
.C(n_774),
.Y(n_4029)
);

CKINVDCx20_ASAP7_75t_R g4030 ( 
.A(n_4022),
.Y(n_4030)
);

OR2x2_ASAP7_75t_L g4031 ( 
.A(n_4019),
.B(n_773),
.Y(n_4031)
);

XNOR2x1_ASAP7_75t_L g4032 ( 
.A(n_4031),
.B(n_4018),
.Y(n_4032)
);

NAND2xp5_ASAP7_75t_L g4033 ( 
.A(n_4029),
.B(n_4017),
.Y(n_4033)
);

OAI22xp5_ASAP7_75t_L g4034 ( 
.A1(n_4030),
.A2(n_4024),
.B1(n_4025),
.B2(n_4023),
.Y(n_4034)
);

XOR2xp5_ASAP7_75t_L g4035 ( 
.A(n_4026),
.B(n_878),
.Y(n_4035)
);

XNOR2xp5_ASAP7_75t_L g4036 ( 
.A(n_4028),
.B(n_778),
.Y(n_4036)
);

NAND2xp5_ASAP7_75t_L g4037 ( 
.A(n_4036),
.B(n_4027),
.Y(n_4037)
);

INVxp67_ASAP7_75t_SL g4038 ( 
.A(n_4032),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_4038),
.Y(n_4039)
);

OAI22xp33_ASAP7_75t_SL g4040 ( 
.A1(n_4039),
.A2(n_4033),
.B1(n_4037),
.B2(n_4034),
.Y(n_4040)
);

INVx1_ASAP7_75t_L g4041 ( 
.A(n_4040),
.Y(n_4041)
);

XNOR2xp5_ASAP7_75t_L g4042 ( 
.A(n_4041),
.B(n_4035),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_4042),
.Y(n_4043)
);

AOI22xp5_ASAP7_75t_SL g4044 ( 
.A1(n_4043),
.A2(n_782),
.B1(n_780),
.B2(n_781),
.Y(n_4044)
);

AO21x2_ASAP7_75t_L g4045 ( 
.A1(n_4044),
.A2(n_784),
.B(n_785),
.Y(n_4045)
);

AOI22xp5_ASAP7_75t_L g4046 ( 
.A1(n_4045),
.A2(n_788),
.B1(n_786),
.B2(n_787),
.Y(n_4046)
);

AOI211xp5_ASAP7_75t_L g4047 ( 
.A1(n_4046),
.A2(n_791),
.B(n_789),
.C(n_790),
.Y(n_4047)
);


endmodule