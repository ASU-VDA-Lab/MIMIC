module fake_jpeg_21146_n_101 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_101);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_101;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

HB1xp67_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_7),
.B(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_28),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_26),
.A2(n_27),
.B1(n_32),
.B2(n_22),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_20),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_21),
.B(n_3),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_31),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_4),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_13),
.B(n_19),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_13),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_29),
.A2(n_19),
.B1(n_12),
.B2(n_22),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_12),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_17),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_17),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_32),
.B1(n_25),
.B2(n_18),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_43),
.B(n_25),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_46),
.B(n_10),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_27),
.B1(n_26),
.B2(n_29),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_50),
.Y(n_62)
);

INVxp33_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_8),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_52),
.B(n_57),
.Y(n_69)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_24),
.B1(n_23),
.B2(n_16),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_56),
.Y(n_64)
);

OAI32xp33_ASAP7_75t_L g56 ( 
.A1(n_33),
.A2(n_15),
.A3(n_24),
.B1(n_14),
.B2(n_5),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_33),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_60),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_24),
.Y(n_60)
);

NOR3xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_15),
.C(n_14),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_11),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_8),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_68),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_72),
.C(n_49),
.Y(n_78)
);

XOR2x2_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_10),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_46),
.C(n_59),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_56),
.B1(n_47),
.B2(n_44),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_79),
.B1(n_44),
.B2(n_66),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_77),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_50),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_59),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_70),
.C(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_60),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_78),
.A2(n_65),
.B1(n_49),
.B2(n_69),
.Y(n_82)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_84),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_75),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_83),
.A2(n_65),
.B1(n_64),
.B2(n_71),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_64),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_77),
.C(n_63),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_90),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_89),
.Y(n_94)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

NAND3xp33_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_74),
.C(n_71),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_92),
.B(n_93),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_86),
.A2(n_80),
.B1(n_79),
.B2(n_85),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_54),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_45),
.C(n_55),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_92),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_63),
.B(n_67),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_98),
.A2(n_99),
.B1(n_97),
.B2(n_60),
.Y(n_100)
);

AOI221xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_95),
.B1(n_84),
.B2(n_86),
.C(n_91),
.Y(n_101)
);


endmodule