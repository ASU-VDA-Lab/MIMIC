module fake_netlist_1_12160_n_42 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_42);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_42;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_30;
wire n_33;
wire n_26;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
HB1xp67_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_4), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_12), .Y(n_18) );
OAI22xp5_ASAP7_75t_SL g19 ( .A1(n_14), .A2(n_13), .B1(n_3), .B2(n_11), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_0), .Y(n_20) );
CKINVDCx20_ASAP7_75t_R g21 ( .A(n_8), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_10), .B(n_1), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_4), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
AOI21xp5_ASAP7_75t_L g25 ( .A1(n_16), .A2(n_9), .B(n_1), .Y(n_25) );
INVx2_ASAP7_75t_SL g26 ( .A(n_18), .Y(n_26) );
BUFx2_ASAP7_75t_L g27 ( .A(n_17), .Y(n_27) );
OR2x2_ASAP7_75t_L g28 ( .A(n_27), .B(n_20), .Y(n_28) );
AOI21x1_ASAP7_75t_L g29 ( .A1(n_25), .A2(n_18), .B(n_22), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_29), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
AO221x2_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_19), .B1(n_23), .B2(n_24), .C(n_5), .Y(n_32) );
AND2x2_ASAP7_75t_L g33 ( .A(n_30), .B(n_27), .Y(n_33) );
AND2x2_ASAP7_75t_L g34 ( .A(n_33), .B(n_32), .Y(n_34) );
NOR3xp33_ASAP7_75t_L g35 ( .A(n_32), .B(n_26), .C(n_24), .Y(n_35) );
NAND4xp25_ASAP7_75t_L g36 ( .A(n_35), .B(n_30), .C(n_2), .D(n_3), .Y(n_36) );
NOR2xp67_ASAP7_75t_L g37 ( .A(n_34), .B(n_0), .Y(n_37) );
O2A1O1Ixp33_ASAP7_75t_L g38 ( .A1(n_36), .A2(n_26), .B(n_21), .C(n_7), .Y(n_38) );
OAI211xp5_ASAP7_75t_L g39 ( .A1(n_37), .A2(n_5), .B(n_6), .C(n_7), .Y(n_39) );
INVx2_ASAP7_75t_L g40 ( .A(n_39), .Y(n_40) );
OAI21xp5_ASAP7_75t_L g41 ( .A1(n_40), .A2(n_38), .B(n_6), .Y(n_41) );
INVx1_ASAP7_75t_L g42 ( .A(n_41), .Y(n_42) );
endmodule