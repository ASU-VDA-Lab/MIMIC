module fake_jpeg_16831_n_333 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_40),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_41),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_22),
.B(n_10),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_43),
.B(n_45),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_22),
.B(n_9),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_47),
.B(n_58),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_15),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_64),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_20),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_59),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_24),
.B(n_29),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_28),
.B(n_7),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_15),
.B(n_0),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_30),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_67),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_24),
.B(n_7),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_70),
.A2(n_26),
.B1(n_38),
.B2(n_30),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_71),
.A2(n_75),
.B(n_119),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_72),
.B(n_114),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_26),
.B1(n_38),
.B2(n_64),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_74),
.A2(n_5),
.B1(n_75),
.B2(n_108),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_39),
.A2(n_26),
.B1(n_38),
.B2(n_35),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_47),
.A2(n_29),
.B(n_34),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_78),
.B(n_102),
.Y(n_149)
);

AOI21xp33_ASAP7_75t_SL g80 ( 
.A1(n_56),
.A2(n_35),
.B(n_17),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_L g136 ( 
.A1(n_80),
.A2(n_0),
.B(n_1),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_55),
.A2(n_21),
.B1(n_33),
.B2(n_31),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_88),
.A2(n_103),
.B1(n_121),
.B2(n_16),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_61),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_92),
.B(n_100),
.Y(n_152)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_45),
.B(n_37),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_52),
.B(n_37),
.Y(n_102)
);

OA22x2_ASAP7_75t_L g103 ( 
.A1(n_63),
.A2(n_21),
.B1(n_31),
.B2(n_33),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_54),
.B(n_17),
.C(n_33),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_111),
.Y(n_122)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_54),
.B(n_17),
.C(n_31),
.Y(n_111)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_48),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_62),
.B(n_34),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_116),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_44),
.B(n_27),
.C(n_18),
.Y(n_116)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_118),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_40),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_65),
.A2(n_27),
.B1(n_18),
.B2(n_16),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_119),
.Y(n_123)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_125),
.A2(n_140),
.B1(n_150),
.B2(n_161),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_86),
.A2(n_32),
.B1(n_6),
.B2(n_7),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_126),
.A2(n_132),
.B1(n_141),
.B2(n_160),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_127),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_120),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_130),
.B(n_145),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_81),
.B(n_50),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_142),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_83),
.A2(n_32),
.B1(n_6),
.B2(n_2),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_133),
.Y(n_175)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_136),
.B(n_151),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_73),
.A2(n_41),
.B1(n_42),
.B2(n_4),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_137),
.A2(n_154),
.B1(n_142),
.B2(n_130),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_79),
.B(n_1),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_139),
.B(n_153),
.Y(n_183)
);

OA21x2_ASAP7_75t_L g140 ( 
.A1(n_103),
.A2(n_1),
.B(n_3),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_98),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_87),
.B(n_3),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_99),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_144),
.B(n_147),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_85),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_147),
.B(n_159),
.Y(n_189)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

OR2x2_ASAP7_75t_SL g151 ( 
.A(n_82),
.B(n_5),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_91),
.B(n_5),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_103),
.A2(n_106),
.B1(n_90),
.B2(n_89),
.Y(n_154)
);

AO22x1_ASAP7_75t_L g156 ( 
.A1(n_88),
.A2(n_121),
.B1(n_114),
.B2(n_71),
.Y(n_156)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_76),
.A2(n_105),
.B1(n_113),
.B2(n_97),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_95),
.B(n_112),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_158),
.B(n_166),
.Y(n_184)
);

AOI32xp33_ASAP7_75t_L g159 ( 
.A1(n_76),
.A2(n_118),
.A3(n_99),
.B1(n_101),
.B2(n_110),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_85),
.A2(n_84),
.B1(n_101),
.B2(n_119),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_112),
.B(n_110),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_167),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_71),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_157),
.Y(n_190)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_102),
.Y(n_164)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_93),
.Y(n_165)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_165),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_79),
.B(n_100),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_81),
.B(n_74),
.Y(n_167)
);

AO21x2_ASAP7_75t_L g168 ( 
.A1(n_140),
.A2(n_156),
.B(n_161),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_168),
.A2(n_194),
.B1(n_202),
.B2(n_176),
.Y(n_225)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_169),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_163),
.A2(n_122),
.B1(n_140),
.B2(n_156),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_172),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_149),
.B(n_164),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_179),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_131),
.C(n_129),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_174),
.B(n_170),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_181),
.B(n_188),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_122),
.B(n_149),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_191),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_152),
.B(n_151),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_190),
.A2(n_168),
.B(n_188),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_122),
.B(n_162),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_138),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_197),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_125),
.A2(n_165),
.B1(n_135),
.B2(n_143),
.Y(n_194)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_124),
.Y(n_196)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_128),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_124),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_204),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_144),
.B(n_148),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_203),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_143),
.B(n_155),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_134),
.B(n_155),
.Y(n_204)
);

INVx13_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_175),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_191),
.B(n_145),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_206),
.B(n_215),
.C(n_219),
.Y(n_242)
);

AND2x6_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_123),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_210),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_199),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_222),
.Y(n_246)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_201),
.Y(n_213)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_203),
.Y(n_214)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_214),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_186),
.B(n_133),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_187),
.A2(n_146),
.B(n_123),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_217),
.A2(n_223),
.B(n_224),
.Y(n_247)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_218),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_174),
.B(n_146),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_172),
.B(n_127),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_182),
.B(n_187),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_225),
.B(n_198),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_168),
.A2(n_176),
.B(n_189),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_226),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_168),
.A2(n_200),
.B(n_182),
.Y(n_227)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_227),
.B(n_231),
.CI(n_225),
.CON(n_258),
.SN(n_258)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_194),
.A2(n_193),
.B1(n_170),
.B2(n_173),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_231),
.A2(n_214),
.B1(n_207),
.B2(n_216),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_171),
.C(n_185),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_184),
.B(n_192),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_171),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_200),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_181),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_200),
.A2(n_178),
.B(n_180),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_196),
.Y(n_253)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_238),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_239),
.A2(n_250),
.B(n_254),
.Y(n_280)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_241),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_183),
.Y(n_243)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_243),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_209),
.B(n_185),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_245),
.B(n_248),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_253),
.C(n_259),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_252),
.A2(n_223),
.B1(n_211),
.B2(n_208),
.Y(n_268)
);

AOI211xp5_ASAP7_75t_SL g254 ( 
.A1(n_210),
.A2(n_175),
.B(n_195),
.C(n_216),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_195),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_256),
.B(n_260),
.Y(n_277)
);

NOR4xp25_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_207),
.C(n_234),
.D(n_220),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_257),
.B(n_261),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_258),
.A2(n_223),
.B(n_224),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_219),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_230),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_206),
.B(n_215),
.C(n_227),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_255),
.A2(n_217),
.B1(n_226),
.B2(n_213),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_264),
.A2(n_266),
.B1(n_268),
.B2(n_281),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_246),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_265),
.B(n_279),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_255),
.A2(n_250),
.B1(n_239),
.B2(n_244),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_267),
.A2(n_247),
.B(n_245),
.Y(n_288)
);

AOI322xp5_ASAP7_75t_L g270 ( 
.A1(n_252),
.A2(n_235),
.A3(n_211),
.B1(n_229),
.B2(n_218),
.C1(n_205),
.C2(n_212),
.Y(n_270)
);

OAI21x1_ASAP7_75t_L g291 ( 
.A1(n_270),
.A2(n_237),
.B(n_259),
.Y(n_291)
);

AOI321xp33_ASAP7_75t_L g272 ( 
.A1(n_257),
.A2(n_205),
.A3(n_221),
.B1(n_222),
.B2(n_261),
.C(n_242),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_272),
.A2(n_273),
.B(n_278),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_246),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_241),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_253),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_237),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_240),
.A2(n_254),
.B1(n_258),
.B2(n_236),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_242),
.B(n_249),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_271),
.C(n_263),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_262),
.B(n_243),
.Y(n_285)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_285),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_274),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_291),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_280),
.A2(n_247),
.B(n_258),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_287),
.A2(n_288),
.B(n_278),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_236),
.Y(n_290)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_290),
.Y(n_300)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_269),
.Y(n_292)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_292),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_278),
.A2(n_251),
.B1(n_273),
.B2(n_280),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_293),
.A2(n_268),
.B1(n_277),
.B2(n_266),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_264),
.Y(n_307)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_269),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_251),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_262),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_296),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_283),
.A2(n_281),
.B(n_267),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_287),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_307),
.Y(n_316)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_299),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_271),
.C(n_282),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_301),
.B(n_306),
.Y(n_312)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_303),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_263),
.C(n_272),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_276),
.Y(n_309)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_309),
.Y(n_319)
);

AO21x1_ASAP7_75t_L g323 ( 
.A1(n_310),
.A2(n_314),
.B(n_309),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_299),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_305),
.Y(n_322)
);

AOI31xp33_ASAP7_75t_L g314 ( 
.A1(n_302),
.A2(n_276),
.A3(n_288),
.B(n_289),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_303),
.B(n_284),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_304),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_300),
.A2(n_293),
.B1(n_292),
.B2(n_295),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_318),
.B(n_298),
.C(n_297),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_320),
.A2(n_317),
.B(n_306),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_321),
.A2(n_324),
.B1(n_325),
.B2(n_313),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_323),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_300),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_308),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_326),
.B(n_328),
.C(n_316),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_329),
.B(n_330),
.Y(n_331)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_327),
.B(n_296),
.Y(n_330)
);

NAND2x1_ASAP7_75t_SL g332 ( 
.A(n_331),
.B(n_316),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_312),
.Y(n_333)
);


endmodule