module fake_jpeg_17999_n_296 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_296);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_296;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_181;
wire n_38;
wire n_26;
wire n_28;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_265;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_SL g19 ( 
.A(n_11),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g43 ( 
.A(n_33),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_21),
.Y(n_34)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_33),
.A2(n_24),
.B1(n_17),
.B2(n_16),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_44),
.A2(n_47),
.B1(n_52),
.B2(n_20),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_24),
.B1(n_17),
.B2(n_16),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_32),
.A2(n_27),
.B(n_29),
.C(n_22),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_48),
.A2(n_59),
.B(n_27),
.C(n_29),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_15),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_49),
.B(n_53),
.Y(n_86)
);

CKINVDCx11_ASAP7_75t_R g50 ( 
.A(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_58),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_24),
.B1(n_17),
.B2(n_16),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_15),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_15),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_22),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_56),
.B(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_80),
.Y(n_92)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_48),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_67),
.B(n_71),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_68),
.B(n_26),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_78),
.Y(n_90)
);

FAx1_ASAP7_75t_SL g71 ( 
.A(n_49),
.B(n_34),
.CI(n_35),
.CON(n_71),
.SN(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_50),
.A2(n_17),
.B1(n_24),
.B2(n_25),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_76),
.A2(n_83),
.B1(n_51),
.B2(n_43),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_47),
.A2(n_20),
.B1(n_16),
.B2(n_29),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_77),
.A2(n_84),
.B(n_25),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_60),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_40),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_60),
.B(n_36),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_26),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_61),
.A2(n_20),
.B1(n_26),
.B2(n_25),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_62),
.A2(n_20),
.B1(n_36),
.B2(n_35),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_34),
.B1(n_36),
.B2(n_61),
.Y(n_91)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

CKINVDCx6p67_ASAP7_75t_R g88 ( 
.A(n_45),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_91),
.A2(n_109),
.B1(n_113),
.B2(n_89),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_103),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_86),
.B(n_52),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_98),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_44),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_96),
.B(n_97),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_63),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_63),
.Y(n_99)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_34),
.C(n_43),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_100),
.B(n_101),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_40),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_27),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_67),
.A2(n_51),
.B1(n_42),
.B2(n_38),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_68),
.Y(n_118)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_118),
.A2(n_127),
.B(n_95),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_134),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_64),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_126),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_112),
.A2(n_77),
.B1(n_83),
.B2(n_80),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_123),
.A2(n_125),
.B1(n_131),
.B2(n_116),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_102),
.A2(n_78),
.B1(n_84),
.B2(n_65),
.Y(n_125)
);

OAI32xp33_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_82),
.A3(n_75),
.B1(n_65),
.B2(n_85),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_102),
.A2(n_74),
.B1(n_87),
.B2(n_75),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_133),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_31),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_137),
.Y(n_151)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_92),
.B(n_46),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_106),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_107),
.A2(n_89),
.B1(n_76),
.B2(n_88),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_139),
.A2(n_108),
.B1(n_115),
.B2(n_111),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_105),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_140),
.Y(n_146)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_105),
.Y(n_141)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_98),
.B(n_30),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_142),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_144),
.A2(n_152),
.B(n_160),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_128),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_148),
.B(n_150),
.Y(n_170)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

AND2x6_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_100),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_154),
.A2(n_147),
.B(n_149),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_118),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_130),
.A2(n_92),
.B1(n_109),
.B2(n_106),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_159),
.A2(n_162),
.B1(n_163),
.B2(n_165),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_130),
.A2(n_97),
.B(n_110),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_128),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_161),
.B(n_120),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_127),
.A2(n_91),
.B1(n_115),
.B2(n_108),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_117),
.A2(n_110),
.B1(n_111),
.B2(n_42),
.Y(n_163)
);

INVx13_ASAP7_75t_L g164 ( 
.A(n_119),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_135),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_38),
.Y(n_165)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_165),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_126),
.B(n_38),
.Y(n_166)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_43),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_129),
.C(n_21),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_181),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_166),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_171),
.A2(n_188),
.B1(n_190),
.B2(n_88),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_121),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_183),
.C(n_187),
.Y(n_211)
);

XNOR2x1_ASAP7_75t_SL g173 ( 
.A(n_157),
.B(n_124),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_173),
.A2(n_178),
.B(n_182),
.Y(n_199)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_174),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_145),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_145),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_176),
.A2(n_154),
.B1(n_158),
.B2(n_88),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_155),
.A2(n_131),
.B1(n_133),
.B2(n_137),
.Y(n_178)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_122),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_43),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_144),
.A2(n_132),
.B(n_129),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_185),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_159),
.A2(n_30),
.B1(n_18),
.B2(n_31),
.Y(n_188)
);

OAI21x1_ASAP7_75t_L g189 ( 
.A1(n_150),
.A2(n_18),
.B(n_30),
.Y(n_189)
);

NOR3xp33_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_143),
.C(n_151),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_153),
.A2(n_88),
.B1(n_42),
.B2(n_46),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_23),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_192),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_147),
.B(n_23),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_146),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_194),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_185),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_203),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_152),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_200),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_160),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_204),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_164),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_207),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_163),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_206),
.B(n_31),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_158),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_162),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_210),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_209),
.A2(n_31),
.B1(n_30),
.B2(n_18),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_190),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_169),
.B(n_18),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_212),
.B(n_46),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_214),
.A2(n_210),
.B1(n_194),
.B2(n_168),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_197),
.A2(n_186),
.B1(n_182),
.B2(n_171),
.Y(n_216)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

A2O1A1Ixp33_ASAP7_75t_SL g218 ( 
.A1(n_208),
.A2(n_177),
.B(n_186),
.C(n_168),
.Y(n_218)
);

AOI22x1_ASAP7_75t_L g243 ( 
.A1(n_218),
.A2(n_28),
.B1(n_23),
.B2(n_31),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_213),
.A2(n_175),
.B(n_177),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_219),
.A2(n_231),
.B(n_1),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_209),
.A2(n_184),
.B1(n_192),
.B2(n_187),
.Y(n_221)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_221),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_206),
.A2(n_173),
.B1(n_183),
.B2(n_2),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_222),
.A2(n_225),
.B1(n_232),
.B2(n_0),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_200),
.A2(n_199),
.B1(n_196),
.B2(n_195),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_228),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_196),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_211),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_199),
.A2(n_9),
.B(n_13),
.Y(n_231)
);

XNOR2x1_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_229),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_235),
.A2(n_239),
.B1(n_243),
.B2(n_244),
.Y(n_249)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_236),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_198),
.C(n_211),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_240),
.C(n_247),
.Y(n_252)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_219),
.A2(n_202),
.B(n_201),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_202),
.Y(n_242)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_242),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_227),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_30),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_224),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_28),
.C(n_18),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_234),
.Y(n_251)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_251),
.Y(n_265)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_220),
.C(n_215),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_237),
.C(n_233),
.Y(n_262)
);

AOI322xp5_ASAP7_75t_SL g255 ( 
.A1(n_235),
.A2(n_217),
.A3(n_231),
.B1(n_222),
.B2(n_216),
.C1(n_218),
.C2(n_6),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_259),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_241),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_239),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_246),
.A2(n_218),
.B(n_7),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_258),
.A2(n_6),
.B(n_12),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_218),
.Y(n_259)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_261),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_264),
.C(n_266),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_256),
.A2(n_243),
.B(n_244),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_267),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_247),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_28),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_258),
.A2(n_7),
.B(n_12),
.Y(n_267)
);

XOR2x1_ASAP7_75t_SL g268 ( 
.A(n_249),
.B(n_7),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_250),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_269),
.A2(n_260),
.B(n_268),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_273),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_270),
.B(n_248),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_249),
.Y(n_274)
);

AO21x1_ASAP7_75t_L g280 ( 
.A1(n_274),
.A2(n_264),
.B(n_266),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_276),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_252),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_5),
.Y(n_278)
);

NAND3xp33_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_8),
.C(n_10),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_283),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_274),
.A2(n_5),
.B(n_11),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_282),
.A2(n_271),
.B(n_286),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_279),
.A2(n_4),
.B(n_8),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_28),
.C(n_4),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_284),
.B(n_1),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_8),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_286),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_288),
.Y(n_292)
);

AOI21x1_ASAP7_75t_L g293 ( 
.A1(n_290),
.A2(n_291),
.B(n_10),
.Y(n_293)
);

OAI221xp5_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_289),
.B1(n_281),
.B2(n_10),
.C(n_3),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_294),
.A2(n_292),
.B(n_2),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_28),
.Y(n_296)
);


endmodule