module real_jpeg_26988_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_249;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_244;
wire n_213;
wire n_128;
wire n_179;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_0),
.A2(n_59),
.B1(n_65),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_0),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_0),
.A2(n_49),
.B1(n_50),
.B2(n_68),
.Y(n_109)
);

INVx11_ASAP7_75t_SL g60 ( 
.A(n_1),
.Y(n_60)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_5),
.Y(n_137)
);

AOI21xp33_ASAP7_75t_SL g138 ( 
.A1(n_5),
.A2(n_29),
.B(n_33),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_137),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_5),
.B(n_31),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_5),
.A2(n_49),
.B(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_5),
.B(n_49),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_5),
.B(n_54),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_5),
.A2(n_57),
.B1(n_66),
.B2(n_225),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_5),
.A2(n_32),
.B(n_240),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_6),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_144),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_6),
.A2(n_49),
.B1(n_50),
.B2(n_144),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_6),
.A2(n_59),
.B1(n_65),
.B2(n_144),
.Y(n_225)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_8),
.A2(n_25),
.B1(n_32),
.B2(n_33),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_8),
.A2(n_25),
.B1(n_59),
.B2(n_65),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_8),
.A2(n_25),
.B1(n_49),
.B2(n_50),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_9),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g161 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_98),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_9),
.A2(n_49),
.B1(n_50),
.B2(n_98),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_9),
.A2(n_59),
.B1(n_65),
.B2(n_98),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_10),
.A2(n_49),
.B1(n_50),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_10),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_10),
.A2(n_59),
.B1(n_65),
.B2(n_77),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_77),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_11),
.A2(n_37),
.B1(n_49),
.B2(n_50),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_11),
.A2(n_37),
.B1(n_59),
.B2(n_65),
.Y(n_214)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_12),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_13),
.A2(n_59),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_13),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_13),
.A2(n_49),
.B1(n_50),
.B2(n_64),
.Y(n_84)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_15),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_16),
.A2(n_32),
.B1(n_33),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_16),
.A2(n_40),
.B1(n_49),
.B2(n_50),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_16),
.A2(n_26),
.B1(n_27),
.B2(n_40),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_16),
.A2(n_40),
.B1(n_59),
.B2(n_65),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_17),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_17),
.A2(n_49),
.B1(n_50),
.B2(n_53),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_17),
.A2(n_53),
.B1(n_59),
.B2(n_65),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_126),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_124),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_101),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_21),
.B(n_101),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_78),
.C(n_88),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_22),
.B(n_78),
.Y(n_148)
);

BUFx24_ASAP7_75t_SL g276 ( 
.A(n_22),
.Y(n_276)
);

FAx1_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_38),
.CI(n_55),
.CON(n_22),
.SN(n_22)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_23),
.B(n_38),
.C(n_55),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B1(n_31),
.B2(n_36),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_24),
.A2(n_28),
.B1(n_31),
.B2(n_97),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_26),
.A2(n_35),
.B(n_137),
.C(n_138),
.Y(n_136)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_27),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g30 ( 
.A(n_27),
.B(n_29),
.Y(n_30)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_28),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_28),
.A2(n_31),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

AO22x1_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_31),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_43),
.B(n_45),
.C(n_48),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_46),
.Y(n_45)
);

OAI32xp33_ASAP7_75t_L g248 ( 
.A1(n_32),
.A2(n_43),
.A3(n_50),
.B1(n_241),
.B2(n_249),
.Y(n_248)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_33),
.B(n_137),
.Y(n_241)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_36),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_41),
.B1(n_52),
.B2(n_54),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_39),
.A2(n_41),
.B1(n_54),
.B2(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_41),
.A2(n_54),
.B1(n_161),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_42),
.A2(n_48),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_42),
.A2(n_48),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_42),
.A2(n_48),
.B1(n_133),
.B2(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_42),
.A2(n_48),
.B1(n_182),
.B2(n_239),
.Y(n_238)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_49),
.A2(n_50),
.B1(n_73),
.B2(n_74),
.Y(n_75)
);

OAI32xp33_ASAP7_75t_L g202 ( 
.A1(n_49),
.A2(n_65),
.A3(n_73),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_49),
.B(n_51),
.Y(n_249)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_52),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_69),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_56),
.B(n_69),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_63),
.B1(n_66),
.B2(n_67),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_57),
.A2(n_66),
.B(n_67),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_57),
.A2(n_63),
.B1(n_66),
.B2(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_57),
.A2(n_66),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_57),
.A2(n_66),
.B1(n_219),
.B2(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_57),
.A2(n_66),
.B1(n_214),
.B2(n_251),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_58),
.A2(n_92),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_58),
.A2(n_61),
.B1(n_140),
.B2(n_184),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_58),
.A2(n_141),
.B1(n_218),
.B2(n_220),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_61),
.Y(n_58)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_65),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_59),
.B(n_74),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_59),
.B(n_230),
.Y(n_229)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_66),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_66),
.B(n_137),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_76),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_71),
.A2(n_72),
.B1(n_84),
.B2(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_71),
.A2(n_72),
.B1(n_198),
.B2(n_200),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_71),
.A2(n_72),
.B1(n_200),
.B2(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_71),
.A2(n_72),
.B1(n_167),
.B2(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_72),
.B(n_137),
.Y(n_226)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_76),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_86),
.B2(n_87),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_79),
.B(n_87),
.Y(n_120)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_82),
.A2(n_85),
.B1(n_95),
.B2(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_82),
.A2(n_85),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_86),
.A2(n_87),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_88),
.B(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_96),
.C(n_99),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_89),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_90),
.B(n_93),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_99),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_97),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_100),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_122),
.B2(n_123),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_111),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_108),
.B(n_110),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_108),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_111)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_116),
.A2(n_118),
.B1(n_143),
.B2(n_145),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_122),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_149),
.B(n_275),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_147),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_128),
.B(n_147),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.C(n_146),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_129),
.B(n_146),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.C(n_142),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_142),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_135),
.B(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_139),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_143),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_187),
.Y(n_149)
);

INVxp33_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI21xp33_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_170),
.B(n_186),
.Y(n_151)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_168),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_153),
.B(n_168),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.C(n_157),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_157),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_162),
.C(n_165),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_158),
.A2(n_159),
.B1(n_165),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_173),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.C(n_178),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_174),
.B(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_273),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_177),
.Y(n_273)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.C(n_185),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_180),
.B(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_183),
.B(n_185),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_184),
.Y(n_251)
);

NOR3xp33_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_189),
.C(n_190),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_269),
.B(n_274),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_255),
.B(n_268),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_234),
.B(n_254),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_215),
.B(n_233),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_205),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_195),
.B(n_205),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_201),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_196),
.A2(n_197),
.B1(n_201),
.B2(n_202),
.Y(n_221)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_199),
.Y(n_203)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_212),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_210),
.C(n_212),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_211),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_213),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_222),
.B(n_232),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_221),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_217),
.B(n_221),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_227),
.B(n_231),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_224),
.B(n_226),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_235),
.B(n_236),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_247),
.B1(n_252),
.B2(n_253),
.Y(n_236)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_237),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_242),
.B1(n_245),
.B2(n_246),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_238),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_242),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_246),
.C(n_253),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_244),
.Y(n_265)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_247),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_250),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_250),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_256),
.B(n_257),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_261),
.B2(n_262),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_264),
.C(n_266),
.Y(n_270)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_266),
.B2(n_267),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_263),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_264),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_270),
.B(n_271),
.Y(n_274)
);


endmodule