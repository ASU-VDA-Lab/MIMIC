module fake_aes_2496_n_1166 (n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_292, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_297, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_291, n_170, n_294, n_40, n_111, n_157, n_296, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_295, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_283, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_293, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_290, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1166);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_292;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_297;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_291;
input n_170;
input n_294;
input n_40;
input n_111;
input n_157;
input n_296;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_295;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_283;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_293;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1166;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1092;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_667;
wire n_496;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_1158;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_1122;
wire n_528;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_1128;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_1161;
wire n_987;
wire n_1030;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_1163;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_384;
wire n_617;
wire n_434;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_1090;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1024;
wire n_1016;
wire n_1078;
wire n_572;
wire n_1017;
wire n_324;
wire n_1097;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_303;
wire n_975;
wire n_1042;
wire n_437;
wire n_512;
wire n_326;
wire n_333;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_945;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_1025;
wire n_1011;
wire n_1132;
wire n_880;
wire n_1101;
wire n_1159;
wire n_630;
wire n_1155;
wire n_511;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_624;
wire n_426;
wire n_769;
wire n_725;
wire n_844;
wire n_818;
wire n_1160;
wire n_1018;
wire n_738;
wire n_979;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_1138;
wire n_506;
wire n_533;
wire n_490;
wire n_393;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_1154;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_1091;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_935;
wire n_427;
wire n_950;
wire n_910;
wire n_460;
wire n_1046;
wire n_478;
wire n_482;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_1145;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_1140;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_1147;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_685;
wire n_362;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_601;
wire n_439;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_446;
wire n_420;
wire n_621;
wire n_423;
wire n_342;
wire n_666;
wire n_799;
wire n_1089;
wire n_1058;
wire n_370;
wire n_1050;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_806;
wire n_1066;
wire n_539;
wire n_1055;
wire n_1157;
wire n_974;
wire n_1153;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_1135;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_363;
wire n_315;
wire n_409;
wire n_733;
wire n_861;
wire n_899;
wire n_654;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_1144;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_756;
wire n_520;
wire n_1057;
wire n_1152;
wire n_681;
wire n_1139;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_1149;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_419;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_1125;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_1133;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_553;
wire n_440;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_1110;
wire n_325;
wire n_1131;
wire n_1102;
wire n_498;
wire n_597;
wire n_349;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1123;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_1156;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_924;
wire n_912;
wire n_947;
wire n_1043;
wire n_582;
wire n_378;
wire n_1141;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_1096;
wire n_335;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_1136;
wire n_397;
wire n_1142;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1027;
wire n_1007;
wire n_859;
wire n_1117;
wire n_1040;
wire n_1165;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_1143;
wire n_629;
wire n_569;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_1112;
wire n_675;
wire n_967;
wire n_504;
wire n_581;
wire n_458;
wire n_493;
wire n_418;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_1164;
wire n_1038;
wire n_341;
wire n_1162;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_1150;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_695;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_1104;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_1134;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_1146;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_1137;
wire n_781;
wire n_916;
wire n_421;
wire n_1148;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_819;
wire n_405;
wire n_772;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_992;
wire n_1127;
INVx1_ASAP7_75t_L g298 ( .A(n_27), .Y(n_298) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_146), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_109), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_179), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_124), .Y(n_302) );
BUFx10_ASAP7_75t_L g303 ( .A(n_32), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_186), .Y(n_304) );
NOR2xp67_ASAP7_75t_L g305 ( .A(n_6), .B(n_130), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_71), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_201), .Y(n_307) );
INVxp67_ASAP7_75t_SL g308 ( .A(n_229), .Y(n_308) );
BUFx3_ASAP7_75t_L g309 ( .A(n_122), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_249), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_172), .Y(n_311) );
INVxp67_ASAP7_75t_L g312 ( .A(n_94), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_268), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_214), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_151), .Y(n_315) );
BUFx3_ASAP7_75t_L g316 ( .A(n_296), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_241), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_28), .Y(n_318) );
CKINVDCx20_ASAP7_75t_R g319 ( .A(n_67), .Y(n_319) );
BUFx2_ASAP7_75t_L g320 ( .A(n_219), .Y(n_320) );
INVx1_ASAP7_75t_SL g321 ( .A(n_171), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_254), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_173), .Y(n_323) );
INVxp67_ASAP7_75t_SL g324 ( .A(n_142), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_128), .Y(n_325) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_50), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_162), .Y(n_327) );
BUFx10_ASAP7_75t_L g328 ( .A(n_231), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_200), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_15), .Y(n_330) );
INVxp33_ASAP7_75t_SL g331 ( .A(n_239), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_13), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_287), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_259), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_56), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_152), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_150), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_267), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_208), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_58), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_78), .Y(n_341) );
CKINVDCx20_ASAP7_75t_R g342 ( .A(n_188), .Y(n_342) );
INVxp67_ASAP7_75t_L g343 ( .A(n_66), .Y(n_343) );
INVxp67_ASAP7_75t_SL g344 ( .A(n_163), .Y(n_344) );
INVx1_ASAP7_75t_SL g345 ( .A(n_70), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_111), .Y(n_346) );
BUFx2_ASAP7_75t_L g347 ( .A(n_297), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_66), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_79), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_72), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_193), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_61), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_192), .Y(n_353) );
INVxp67_ASAP7_75t_SL g354 ( .A(n_82), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_243), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_251), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_140), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_50), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_6), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_294), .Y(n_360) );
BUFx2_ASAP7_75t_L g361 ( .A(n_256), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_271), .Y(n_362) );
CKINVDCx20_ASAP7_75t_R g363 ( .A(n_16), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_7), .Y(n_364) );
BUFx3_ASAP7_75t_L g365 ( .A(n_120), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_196), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_22), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_123), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_199), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_9), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_289), .Y(n_371) );
INVxp67_ASAP7_75t_SL g372 ( .A(n_36), .Y(n_372) );
CKINVDCx20_ASAP7_75t_R g373 ( .A(n_77), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_57), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_278), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_255), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_264), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_92), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_250), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_265), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_207), .Y(n_381) );
CKINVDCx20_ASAP7_75t_R g382 ( .A(n_285), .Y(n_382) );
INVxp67_ASAP7_75t_SL g383 ( .A(n_292), .Y(n_383) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_215), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_0), .Y(n_385) );
BUFx3_ASAP7_75t_L g386 ( .A(n_141), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_204), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_242), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_119), .Y(n_389) );
INVxp67_ASAP7_75t_SL g390 ( .A(n_222), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_258), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_252), .Y(n_392) );
CKINVDCx20_ASAP7_75t_R g393 ( .A(n_43), .Y(n_393) );
INVxp67_ASAP7_75t_L g394 ( .A(n_45), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g395 ( .A(n_167), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_101), .Y(n_396) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_15), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_270), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_68), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_24), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_183), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_10), .Y(n_402) );
BUFx3_ASAP7_75t_L g403 ( .A(n_180), .Y(n_403) );
INVx1_ASAP7_75t_SL g404 ( .A(n_85), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_263), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_23), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_135), .Y(n_407) );
INVxp67_ASAP7_75t_L g408 ( .A(n_181), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_205), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_88), .Y(n_410) );
CKINVDCx20_ASAP7_75t_R g411 ( .A(n_18), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_20), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_190), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_266), .Y(n_414) );
CKINVDCx5p33_ASAP7_75t_R g415 ( .A(n_281), .Y(n_415) );
INVxp33_ASAP7_75t_SL g416 ( .A(n_42), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_211), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_154), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_238), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_113), .Y(n_420) );
INVxp67_ASAP7_75t_SL g421 ( .A(n_10), .Y(n_421) );
BUFx3_ASAP7_75t_L g422 ( .A(n_121), .Y(n_422) );
CKINVDCx14_ASAP7_75t_R g423 ( .A(n_178), .Y(n_423) );
CKINVDCx5p33_ASAP7_75t_R g424 ( .A(n_76), .Y(n_424) );
INVxp33_ASAP7_75t_L g425 ( .A(n_24), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_160), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_286), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_65), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_39), .Y(n_429) );
CKINVDCx16_ASAP7_75t_R g430 ( .A(n_64), .Y(n_430) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_145), .Y(n_431) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_197), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_29), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_276), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_7), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_237), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_275), .Y(n_437) );
INVx3_ASAP7_75t_L g438 ( .A(n_14), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_104), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_272), .Y(n_440) );
CKINVDCx16_ASAP7_75t_R g441 ( .A(n_37), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_44), .Y(n_442) );
INVxp67_ASAP7_75t_SL g443 ( .A(n_90), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_218), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_102), .Y(n_445) );
CKINVDCx5p33_ASAP7_75t_R g446 ( .A(n_36), .Y(n_446) );
CKINVDCx5p33_ASAP7_75t_R g447 ( .A(n_98), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_93), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_5), .Y(n_449) );
CKINVDCx5p33_ASAP7_75t_R g450 ( .A(n_158), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_22), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_117), .Y(n_452) );
BUFx5_ASAP7_75t_L g453 ( .A(n_138), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_438), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_453), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_438), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_340), .Y(n_457) );
CKINVDCx5p33_ASAP7_75t_R g458 ( .A(n_342), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_453), .Y(n_459) );
OAI22xp5_ASAP7_75t_SL g460 ( .A1(n_319), .A2(n_2), .B1(n_0), .B2(n_1), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_377), .B(n_1), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_340), .Y(n_462) );
OA21x2_ASAP7_75t_L g463 ( .A1(n_337), .A2(n_73), .B(n_69), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_428), .Y(n_464) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_299), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_320), .B(n_2), .Y(n_466) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_299), .Y(n_467) );
OA21x2_ASAP7_75t_L g468 ( .A1(n_337), .A2(n_75), .B(n_74), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_326), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_453), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_428), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_412), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_433), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_433), .Y(n_474) );
NOR2xp33_ASAP7_75t_R g475 ( .A(n_423), .B(n_80), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_453), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_347), .B(n_3), .Y(n_477) );
AOI22x1_ASAP7_75t_SL g478 ( .A1(n_319), .A2(n_5), .B1(n_3), .B2(n_4), .Y(n_478) );
XOR2xp5_ASAP7_75t_L g479 ( .A(n_363), .B(n_8), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_361), .B(n_8), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_300), .Y(n_481) );
BUFx8_ASAP7_75t_L g482 ( .A(n_453), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_301), .Y(n_483) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_299), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_380), .B(n_9), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_453), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_302), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_425), .B(n_11), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_304), .Y(n_489) );
NOR2xp33_ASAP7_75t_R g490 ( .A(n_423), .B(n_81), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_488), .B(n_425), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_488), .B(n_303), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_469), .B(n_303), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_455), .Y(n_494) );
INVx4_ASAP7_75t_L g495 ( .A(n_477), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_481), .B(n_446), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_455), .Y(n_497) );
AND2x6_ASAP7_75t_L g498 ( .A(n_477), .B(n_309), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_455), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_482), .B(n_328), .Y(n_500) );
INVx4_ASAP7_75t_L g501 ( .A(n_477), .Y(n_501) );
INVx1_ASAP7_75t_SL g502 ( .A(n_472), .Y(n_502) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_465), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_481), .B(n_446), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_459), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_459), .Y(n_506) );
NAND2xp33_ASAP7_75t_L g507 ( .A(n_475), .B(n_453), .Y(n_507) );
BUFx3_ASAP7_75t_L g508 ( .A(n_482), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_477), .B(n_298), .Y(n_509) );
CKINVDCx5p33_ASAP7_75t_R g510 ( .A(n_458), .Y(n_510) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_465), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_459), .Y(n_512) );
INVxp67_ASAP7_75t_L g513 ( .A(n_480), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_482), .B(n_328), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_470), .Y(n_515) );
INVx4_ASAP7_75t_L g516 ( .A(n_463), .Y(n_516) );
INVx4_ASAP7_75t_L g517 ( .A(n_463), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_454), .B(n_312), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_483), .B(n_334), .Y(n_519) );
NOR2x1p5_ASAP7_75t_L g520 ( .A(n_485), .B(n_334), .Y(n_520) );
OR2x6_ASAP7_75t_L g521 ( .A(n_460), .B(n_318), .Y(n_521) );
INVx4_ASAP7_75t_L g522 ( .A(n_463), .Y(n_522) );
BUFx2_ASAP7_75t_L g523 ( .A(n_482), .Y(n_523) );
BUFx4f_ASAP7_75t_L g524 ( .A(n_463), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_470), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_470), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_476), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_476), .Y(n_528) );
AND2x2_ASAP7_75t_SL g529 ( .A(n_468), .B(n_397), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_490), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_476), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_483), .B(n_328), .Y(n_532) );
AND2x4_ASAP7_75t_L g533 ( .A(n_509), .B(n_466), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_513), .B(n_487), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_519), .B(n_487), .Y(n_535) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_508), .Y(n_536) );
INVx2_ASAP7_75t_SL g537 ( .A(n_502), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_491), .B(n_489), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_505), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_505), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_491), .B(n_489), .Y(n_541) );
BUFx2_ASAP7_75t_L g542 ( .A(n_493), .Y(n_542) );
AND2x4_ASAP7_75t_SL g543 ( .A(n_493), .B(n_342), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_492), .Y(n_544) );
INVx3_ASAP7_75t_L g545 ( .A(n_495), .Y(n_545) );
BUFx6f_ASAP7_75t_L g546 ( .A(n_508), .Y(n_546) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_510), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_492), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_509), .Y(n_549) );
BUFx2_ASAP7_75t_L g550 ( .A(n_510), .Y(n_550) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_523), .Y(n_551) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_529), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_495), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_495), .B(n_486), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_501), .B(n_486), .Y(n_555) );
INVx2_ASAP7_75t_SL g556 ( .A(n_520), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_528), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_501), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_496), .B(n_454), .Y(n_559) );
BUFx8_ASAP7_75t_SL g560 ( .A(n_521), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_504), .B(n_456), .Y(n_561) );
BUFx3_ASAP7_75t_L g562 ( .A(n_498), .Y(n_562) );
CKINVDCx8_ASAP7_75t_R g563 ( .A(n_521), .Y(n_563) );
NAND2x1p5_ASAP7_75t_L g564 ( .A(n_500), .B(n_330), .Y(n_564) );
AND2x6_ASAP7_75t_SL g565 ( .A(n_521), .B(n_479), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_532), .B(n_456), .Y(n_566) );
NAND3xp33_ASAP7_75t_SL g567 ( .A(n_530), .B(n_373), .C(n_369), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_528), .Y(n_568) );
XOR2xp5_ASAP7_75t_L g569 ( .A(n_530), .B(n_479), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_498), .B(n_461), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_518), .Y(n_571) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_529), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_514), .B(n_331), .Y(n_573) );
INVx5_ASAP7_75t_L g574 ( .A(n_498), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_494), .Y(n_575) );
INVx3_ASAP7_75t_L g576 ( .A(n_498), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_494), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_498), .B(n_392), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_497), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_497), .Y(n_580) );
NAND2x1p5_ASAP7_75t_L g581 ( .A(n_524), .B(n_332), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_524), .B(n_486), .Y(n_582) );
O2A1O1Ixp5_ASAP7_75t_L g583 ( .A1(n_516), .A2(n_308), .B(n_344), .C(n_324), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_499), .B(n_395), .Y(n_584) );
NAND3xp33_ASAP7_75t_SL g585 ( .A(n_499), .B(n_373), .C(n_369), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_506), .Y(n_586) );
AND2x4_ASAP7_75t_SL g587 ( .A(n_521), .B(n_382), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_506), .B(n_395), .Y(n_588) );
NOR2x2_ASAP7_75t_L g589 ( .A(n_507), .B(n_478), .Y(n_589) );
OAI21xp5_ASAP7_75t_L g590 ( .A1(n_516), .A2(n_468), .B(n_310), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_512), .B(n_415), .Y(n_591) );
INVx2_ASAP7_75t_SL g592 ( .A(n_516), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_515), .Y(n_593) );
AND2x4_ASAP7_75t_L g594 ( .A(n_517), .B(n_382), .Y(n_594) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_515), .Y(n_595) );
BUFx2_ASAP7_75t_L g596 ( .A(n_525), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_525), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_517), .A2(n_416), .B1(n_462), .B2(n_457), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_517), .A2(n_416), .B1(n_462), .B2(n_457), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_526), .B(n_450), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_522), .A2(n_471), .B1(n_473), .B2(n_464), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_534), .B(n_526), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_544), .A2(n_522), .B1(n_531), .B2(n_527), .Y(n_603) );
AOI22x1_ASAP7_75t_L g604 ( .A1(n_590), .A2(n_522), .B1(n_531), .B2(n_527), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_595), .Y(n_605) );
INVx5_ASAP7_75t_L g606 ( .A(n_536), .Y(n_606) );
INVx4_ASAP7_75t_L g607 ( .A(n_574), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_538), .B(n_430), .Y(n_608) );
BUFx3_ASAP7_75t_L g609 ( .A(n_537), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_596), .Y(n_610) );
BUFx12f_ASAP7_75t_L g611 ( .A(n_547), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_553), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_595), .Y(n_613) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_536), .Y(n_614) );
AOI21x1_ASAP7_75t_L g615 ( .A1(n_582), .A2(n_468), .B(n_311), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_579), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g617 ( .A1(n_583), .A2(n_468), .B(n_383), .Y(n_617) );
A2O1A1Ixp33_ASAP7_75t_L g618 ( .A1(n_535), .A2(n_348), .B(n_352), .C(n_335), .Y(n_618) );
BUFx6f_ASAP7_75t_L g619 ( .A(n_536), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_594), .A2(n_431), .B1(n_432), .B2(n_384), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_558), .Y(n_621) );
AND2x4_ASAP7_75t_L g622 ( .A(n_548), .B(n_372), .Y(n_622) );
A2O1A1Ixp33_ASAP7_75t_SL g623 ( .A1(n_573), .A2(n_471), .B(n_473), .C(n_464), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_549), .Y(n_624) );
AND2x4_ASAP7_75t_L g625 ( .A(n_551), .B(n_533), .Y(n_625) );
A2O1A1Ixp33_ASAP7_75t_L g626 ( .A1(n_571), .A2(n_358), .B(n_364), .C(n_359), .Y(n_626) );
INVx1_ASAP7_75t_SL g627 ( .A(n_543), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_541), .B(n_441), .Y(n_628) );
NAND2xp5_ASAP7_75t_SL g629 ( .A(n_546), .B(n_331), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_579), .Y(n_630) );
OAI22xp5_ASAP7_75t_SL g631 ( .A1(n_563), .A2(n_569), .B1(n_393), .B2(n_411), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_580), .Y(n_632) );
OAI21x1_ASAP7_75t_L g633 ( .A1(n_582), .A2(n_353), .B(n_339), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g634 ( .A(n_546), .B(n_306), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_542), .B(n_363), .Y(n_635) );
INVx3_ASAP7_75t_L g636 ( .A(n_546), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_580), .Y(n_637) );
A2O1A1Ixp33_ASAP7_75t_L g638 ( .A1(n_575), .A2(n_367), .B(n_374), .C(n_370), .Y(n_638) );
A2O1A1Ixp33_ASAP7_75t_L g639 ( .A1(n_577), .A2(n_385), .B(n_400), .C(n_399), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_593), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_593), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_597), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_533), .B(n_343), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_597), .Y(n_644) );
BUFx3_ASAP7_75t_L g645 ( .A(n_550), .Y(n_645) );
AO22x1_ASAP7_75t_L g646 ( .A1(n_574), .A2(n_478), .B1(n_449), .B2(n_421), .Y(n_646) );
O2A1O1Ixp33_ASAP7_75t_L g647 ( .A1(n_559), .A2(n_394), .B(n_406), .C(n_402), .Y(n_647) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_546), .Y(n_648) );
AOI21xp5_ASAP7_75t_L g649 ( .A1(n_592), .A2(n_390), .B(n_354), .Y(n_649) );
INVx5_ASAP7_75t_L g650 ( .A(n_574), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_586), .Y(n_651) );
OAI221xp5_ASAP7_75t_L g652 ( .A1(n_598), .A2(n_442), .B1(n_451), .B2(n_435), .C(n_429), .Y(n_652) );
A2O1A1Ixp33_ASAP7_75t_L g653 ( .A1(n_561), .A2(n_305), .B(n_474), .C(n_313), .Y(n_653) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_562), .Y(n_654) );
OAI321xp33_ASAP7_75t_L g655 ( .A1(n_599), .A2(n_397), .A3(n_307), .B1(n_389), .B2(n_323), .C(n_325), .Y(n_655) );
BUFx6f_ASAP7_75t_L g656 ( .A(n_562), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_599), .A2(n_397), .B1(n_315), .B2(n_317), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_545), .Y(n_658) );
A2O1A1Ixp33_ASAP7_75t_L g659 ( .A1(n_566), .A2(n_322), .B(n_327), .C(n_314), .Y(n_659) );
AND2x4_ASAP7_75t_L g660 ( .A(n_556), .B(n_443), .Y(n_660) );
INVx1_ASAP7_75t_SL g661 ( .A(n_587), .Y(n_661) );
BUFx2_ASAP7_75t_L g662 ( .A(n_581), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_539), .Y(n_663) );
OAI22xp33_ASAP7_75t_L g664 ( .A1(n_585), .A2(n_397), .B1(n_408), .B2(n_338), .Y(n_664) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_574), .Y(n_665) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_581), .Y(n_666) );
INVx3_ASAP7_75t_L g667 ( .A(n_545), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_539), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_540), .Y(n_669) );
INVxp67_ASAP7_75t_L g670 ( .A(n_584), .Y(n_670) );
INVx2_ASAP7_75t_SL g671 ( .A(n_564), .Y(n_671) );
AOI21xp5_ASAP7_75t_L g672 ( .A1(n_554), .A2(n_333), .B(n_329), .Y(n_672) );
INVxp67_ASAP7_75t_SL g673 ( .A(n_552), .Y(n_673) );
BUFx6f_ASAP7_75t_L g674 ( .A(n_552), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_540), .Y(n_675) );
INVx2_ASAP7_75t_SL g676 ( .A(n_564), .Y(n_676) );
BUFx3_ASAP7_75t_L g677 ( .A(n_560), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_557), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_568), .Y(n_679) );
CKINVDCx6p67_ASAP7_75t_R g680 ( .A(n_588), .Y(n_680) );
NAND2xp5_ASAP7_75t_SL g681 ( .A(n_576), .B(n_336), .Y(n_681) );
BUFx12f_ASAP7_75t_L g682 ( .A(n_565), .Y(n_682) );
INVx2_ASAP7_75t_SL g683 ( .A(n_591), .Y(n_683) );
CKINVDCx20_ASAP7_75t_R g684 ( .A(n_560), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_554), .A2(n_346), .B(n_341), .Y(n_685) );
OR2x6_ASAP7_75t_L g686 ( .A(n_573), .B(n_351), .Y(n_686) );
CKINVDCx20_ASAP7_75t_R g687 ( .A(n_567), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_566), .A2(n_356), .B1(n_357), .B2(n_355), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_601), .A2(n_362), .B1(n_366), .B2(n_360), .Y(n_689) );
A2O1A1Ixp33_ASAP7_75t_L g690 ( .A1(n_601), .A2(n_375), .B(n_376), .C(n_371), .Y(n_690) );
BUFx2_ASAP7_75t_L g691 ( .A(n_600), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_568), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_570), .A2(n_379), .B1(n_381), .B2(n_378), .Y(n_693) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_552), .A2(n_410), .B1(n_387), .B2(n_388), .C(n_391), .Y(n_694) );
NOR2xp33_ASAP7_75t_SL g695 ( .A(n_576), .B(n_349), .Y(n_695) );
OA21x2_ASAP7_75t_L g696 ( .A1(n_604), .A2(n_353), .B(n_339), .Y(n_696) );
OAI21x1_ASAP7_75t_L g697 ( .A1(n_615), .A2(n_555), .B(n_407), .Y(n_697) );
CKINVDCx11_ASAP7_75t_R g698 ( .A(n_611), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_610), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_605), .B(n_552), .Y(n_700) );
OA21x2_ASAP7_75t_L g701 ( .A1(n_633), .A2(n_407), .B(n_368), .Y(n_701) );
NAND2x1p5_ASAP7_75t_L g702 ( .A(n_662), .B(n_572), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_605), .B(n_572), .Y(n_703) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_647), .A2(n_405), .B1(n_418), .B2(n_414), .C(n_420), .Y(n_704) );
OAI21x1_ASAP7_75t_L g705 ( .A1(n_617), .A2(n_555), .B(n_409), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_651), .B(n_572), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_651), .Y(n_707) );
AND2x4_ASAP7_75t_L g708 ( .A(n_609), .B(n_572), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_616), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_616), .Y(n_710) );
O2A1O1Ixp33_ASAP7_75t_L g711 ( .A1(n_618), .A2(n_578), .B(n_409), .C(n_440), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_613), .B(n_396), .Y(n_712) );
OAI21x1_ASAP7_75t_L g713 ( .A1(n_636), .A2(n_440), .B(n_368), .Y(n_713) );
A2O1A1Ixp33_ASAP7_75t_L g714 ( .A1(n_670), .A2(n_401), .B(n_413), .C(n_398), .Y(n_714) );
OAI21x1_ASAP7_75t_L g715 ( .A1(n_636), .A2(n_426), .B(n_417), .Y(n_715) );
INVx2_ASAP7_75t_L g716 ( .A(n_640), .Y(n_716) );
AOI22xp33_ASAP7_75t_SL g717 ( .A1(n_631), .A2(n_589), .B1(n_309), .B2(n_365), .Y(n_717) );
OAI21x1_ASAP7_75t_L g718 ( .A1(n_640), .A2(n_434), .B(n_427), .Y(n_718) );
OAI21xp5_ASAP7_75t_L g719 ( .A1(n_603), .A2(n_437), .B(n_436), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_641), .B(n_439), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_624), .Y(n_721) );
OR3x4_ASAP7_75t_SL g722 ( .A(n_682), .B(n_12), .C(n_13), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_612), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_652), .A2(n_452), .B1(n_445), .B2(n_316), .Y(n_724) );
AOI22xp33_ASAP7_75t_SL g725 ( .A1(n_661), .A2(n_316), .B1(n_386), .B2(n_365), .Y(n_725) );
NOR2xp67_ASAP7_75t_L g726 ( .A(n_620), .B(n_12), .Y(n_726) );
OAI21x1_ASAP7_75t_L g727 ( .A1(n_641), .A2(n_299), .B(n_386), .Y(n_727) );
OA21x2_ASAP7_75t_L g728 ( .A1(n_653), .A2(n_345), .B(n_321), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_621), .Y(n_729) );
OA21x2_ASAP7_75t_L g730 ( .A1(n_655), .A2(n_404), .B(n_350), .Y(n_730) );
AO21x2_ASAP7_75t_L g731 ( .A1(n_623), .A2(n_467), .B(n_465), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_635), .A2(n_419), .B1(n_444), .B2(n_424), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_644), .Y(n_733) );
AND2x4_ASAP7_75t_L g734 ( .A(n_625), .B(n_403), .Y(n_734) );
OA21x2_ASAP7_75t_L g735 ( .A1(n_690), .A2(n_448), .B(n_447), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_622), .Y(n_736) );
CKINVDCx5p33_ASAP7_75t_R g737 ( .A(n_684), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_602), .Y(n_738) );
AO21x2_ASAP7_75t_L g739 ( .A1(n_659), .A2(n_467), .B(n_465), .Y(n_739) );
OAI21x1_ASAP7_75t_L g740 ( .A1(n_644), .A2(n_422), .B(n_403), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_663), .B(n_16), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_663), .Y(n_742) );
OA21x2_ASAP7_75t_L g743 ( .A1(n_669), .A2(n_422), .B(n_465), .Y(n_743) );
AOI22x1_ASAP7_75t_L g744 ( .A1(n_672), .A2(n_467), .B1(n_484), .B2(n_465), .Y(n_744) );
OAI21xp5_ASAP7_75t_L g745 ( .A1(n_669), .A2(n_484), .B(n_467), .Y(n_745) );
BUFx10_ASAP7_75t_L g746 ( .A(n_625), .Y(n_746) );
OAI21xp5_ASAP7_75t_L g747 ( .A1(n_678), .A2(n_484), .B(n_467), .Y(n_747) );
CKINVDCx5p33_ASAP7_75t_R g748 ( .A(n_677), .Y(n_748) );
AO21x2_ASAP7_75t_L g749 ( .A1(n_685), .A2(n_484), .B(n_467), .Y(n_749) );
OAI21x1_ASAP7_75t_SL g750 ( .A1(n_671), .A2(n_17), .B(n_18), .Y(n_750) );
O2A1O1Ixp33_ASAP7_75t_SL g751 ( .A1(n_678), .A2(n_84), .B(n_86), .C(n_83), .Y(n_751) );
AOI21xp5_ASAP7_75t_L g752 ( .A1(n_668), .A2(n_511), .B(n_503), .Y(n_752) );
OAI22xp5_ASAP7_75t_L g753 ( .A1(n_632), .A2(n_484), .B1(n_511), .B2(n_503), .Y(n_753) );
OAI21x1_ASAP7_75t_L g754 ( .A1(n_630), .A2(n_484), .B(n_89), .Y(n_754) );
OAI21x1_ASAP7_75t_L g755 ( .A1(n_637), .A2(n_91), .B(n_87), .Y(n_755) );
OAI21x1_ASAP7_75t_L g756 ( .A1(n_642), .A2(n_96), .B(n_95), .Y(n_756) );
OAI22xp33_ASAP7_75t_L g757 ( .A1(n_686), .A2(n_19), .B1(n_20), .B2(n_21), .Y(n_757) );
AOI221xp5_ASAP7_75t_L g758 ( .A1(n_626), .A2(n_511), .B1(n_503), .B2(n_25), .C(n_26), .Y(n_758) );
OAI21xp5_ASAP7_75t_L g759 ( .A1(n_675), .A2(n_511), .B(n_503), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_643), .Y(n_760) );
OA21x2_ASAP7_75t_L g761 ( .A1(n_694), .A2(n_99), .B(n_97), .Y(n_761) );
INVx6_ASAP7_75t_L g762 ( .A(n_606), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_683), .B(n_21), .Y(n_763) );
AND2x2_ASAP7_75t_L g764 ( .A(n_608), .B(n_628), .Y(n_764) );
AND2x4_ASAP7_75t_L g765 ( .A(n_666), .B(n_23), .Y(n_765) );
HB1xp67_ASAP7_75t_L g766 ( .A(n_645), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_691), .B(n_28), .Y(n_767) );
AND2x4_ASAP7_75t_L g768 ( .A(n_676), .B(n_29), .Y(n_768) );
O2A1O1Ixp33_ASAP7_75t_L g769 ( .A1(n_638), .A2(n_30), .B(n_31), .C(n_32), .Y(n_769) );
INVx2_ASAP7_75t_L g770 ( .A(n_679), .Y(n_770) );
BUFx3_ASAP7_75t_L g771 ( .A(n_606), .Y(n_771) );
OAI21x1_ASAP7_75t_L g772 ( .A1(n_692), .A2(n_103), .B(n_100), .Y(n_772) );
BUFx6f_ASAP7_75t_L g773 ( .A(n_614), .Y(n_773) );
BUFx3_ASAP7_75t_L g774 ( .A(n_687), .Y(n_774) );
BUFx2_ASAP7_75t_L g775 ( .A(n_627), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_693), .B(n_30), .Y(n_776) );
BUFx6f_ASAP7_75t_L g777 ( .A(n_614), .Y(n_777) );
AOI21xp5_ASAP7_75t_L g778 ( .A1(n_649), .A2(n_106), .B(n_105), .Y(n_778) );
CKINVDCx11_ASAP7_75t_R g779 ( .A(n_680), .Y(n_779) );
INVx1_ASAP7_75t_SL g780 ( .A(n_674), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_657), .B(n_31), .Y(n_781) );
AO21x2_ASAP7_75t_L g782 ( .A1(n_639), .A2(n_108), .B(n_107), .Y(n_782) );
OAI21x1_ASAP7_75t_L g783 ( .A1(n_634), .A2(n_112), .B(n_110), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_686), .B(n_33), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_689), .B(n_34), .Y(n_785) );
OAI21x1_ASAP7_75t_L g786 ( .A1(n_681), .A2(n_115), .B(n_114), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_629), .Y(n_787) );
OR2x6_ASAP7_75t_L g788 ( .A(n_646), .B(n_35), .Y(n_788) );
OA21x2_ASAP7_75t_L g789 ( .A1(n_688), .A2(n_118), .B(n_116), .Y(n_789) );
OAI21x1_ASAP7_75t_L g790 ( .A1(n_667), .A2(n_126), .B(n_125), .Y(n_790) );
OAI21x1_ASAP7_75t_L g791 ( .A1(n_673), .A2(n_129), .B(n_127), .Y(n_791) );
OAI21x1_ASAP7_75t_L g792 ( .A1(n_658), .A2(n_132), .B(n_131), .Y(n_792) );
AO21x2_ASAP7_75t_L g793 ( .A1(n_664), .A2(n_134), .B(n_133), .Y(n_793) );
NAND2x1_ASAP7_75t_L g794 ( .A(n_607), .B(n_136), .Y(n_794) );
OAI21x1_ASAP7_75t_L g795 ( .A1(n_619), .A2(n_139), .B(n_137), .Y(n_795) );
OAI21xp5_ASAP7_75t_L g796 ( .A1(n_705), .A2(n_660), .B(n_695), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_699), .Y(n_797) );
AND2x2_ASAP7_75t_L g798 ( .A(n_764), .B(n_765), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_738), .B(n_760), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_707), .B(n_674), .Y(n_800) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_785), .A2(n_619), .B1(n_648), .B2(n_656), .Y(n_801) );
AO31x2_ASAP7_75t_L g802 ( .A1(n_741), .A2(n_607), .A3(n_648), .B(n_619), .Y(n_802) );
INVx2_ASAP7_75t_L g803 ( .A(n_742), .Y(n_803) );
AOI222xp33_ASAP7_75t_L g804 ( .A1(n_726), .A2(n_654), .B1(n_650), .B2(n_648), .C1(n_665), .C2(n_40), .Y(n_804) );
AOI222xp33_ASAP7_75t_L g805 ( .A1(n_757), .A2(n_650), .B1(n_665), .B2(n_38), .C1(n_39), .C2(n_41), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_717), .A2(n_665), .B1(n_650), .B2(n_41), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_736), .Y(n_807) );
AOI221xp5_ASAP7_75t_L g808 ( .A1(n_704), .A2(n_43), .B1(n_44), .B2(n_46), .C(n_47), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_717), .B(n_46), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_721), .Y(n_810) );
AOI21xp5_ASAP7_75t_L g811 ( .A1(n_752), .A2(n_195), .B(n_295), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_788), .A2(n_48), .B1(n_49), .B2(n_51), .Y(n_812) );
A2O1A1Ixp33_ASAP7_75t_L g813 ( .A1(n_711), .A2(n_48), .B(n_49), .C(n_51), .Y(n_813) );
AOI21xp33_ASAP7_75t_L g814 ( .A1(n_711), .A2(n_52), .B(n_53), .Y(n_814) );
AOI21xp5_ASAP7_75t_L g815 ( .A1(n_752), .A2(n_202), .B(n_293), .Y(n_815) );
AOI322xp5_ASAP7_75t_L g816 ( .A1(n_757), .A2(n_54), .A3(n_55), .B1(n_56), .B2(n_58), .C1(n_59), .C2(n_60), .Y(n_816) );
OAI221xp5_ASAP7_75t_L g817 ( .A1(n_704), .A2(n_54), .B1(n_55), .B2(n_59), .C(n_60), .Y(n_817) );
AOI21xp5_ASAP7_75t_L g818 ( .A1(n_759), .A2(n_210), .B(n_291), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_768), .Y(n_819) );
BUFx12f_ASAP7_75t_L g820 ( .A(n_698), .Y(n_820) );
HB1xp67_ASAP7_75t_L g821 ( .A(n_766), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_741), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_763), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_763), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_723), .Y(n_825) );
BUFx6f_ASAP7_75t_L g826 ( .A(n_773), .Y(n_826) );
OAI21x1_ASAP7_75t_L g827 ( .A1(n_697), .A2(n_213), .B(n_290), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_729), .Y(n_828) );
HB1xp67_ASAP7_75t_L g829 ( .A(n_775), .Y(n_829) );
BUFx8_ASAP7_75t_L g830 ( .A(n_779), .Y(n_830) );
OAI22xp5_ASAP7_75t_L g831 ( .A1(n_724), .A2(n_62), .B1(n_63), .B2(n_64), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_767), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_767), .Y(n_833) );
AO21x2_ASAP7_75t_L g834 ( .A1(n_745), .A2(n_143), .B(n_144), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_776), .A2(n_147), .B1(n_148), .B2(n_149), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_776), .A2(n_153), .B1(n_155), .B2(n_156), .Y(n_836) );
INVx2_ASAP7_75t_L g837 ( .A(n_709), .Y(n_837) );
BUFx12f_ASAP7_75t_L g838 ( .A(n_737), .Y(n_838) );
A2O1A1Ixp33_ASAP7_75t_L g839 ( .A1(n_769), .A2(n_157), .B(n_159), .C(n_161), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_784), .A2(n_164), .B1(n_165), .B2(n_166), .Y(n_840) );
AOI21xp5_ASAP7_75t_L g841 ( .A1(n_759), .A2(n_168), .B(n_169), .Y(n_841) );
AND2x2_ASAP7_75t_L g842 ( .A(n_746), .B(n_170), .Y(n_842) );
O2A1O1Ixp33_ASAP7_75t_L g843 ( .A1(n_714), .A2(n_174), .B(n_175), .C(n_176), .Y(n_843) );
AND2x4_ASAP7_75t_L g844 ( .A(n_708), .B(n_177), .Y(n_844) );
OR2x6_ASAP7_75t_L g845 ( .A(n_702), .B(n_182), .Y(n_845) );
OR2x6_ASAP7_75t_L g846 ( .A(n_702), .B(n_184), .Y(n_846) );
OA21x2_ASAP7_75t_L g847 ( .A1(n_740), .A2(n_185), .B(n_187), .Y(n_847) );
AOI21xp5_ASAP7_75t_L g848 ( .A1(n_696), .A2(n_189), .B(n_191), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_785), .A2(n_194), .B1(n_198), .B2(n_203), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_724), .B(n_712), .Y(n_850) );
AOI21xp33_ASAP7_75t_L g851 ( .A1(n_735), .A2(n_206), .B(n_209), .Y(n_851) );
OAI22xp5_ASAP7_75t_L g852 ( .A1(n_710), .A2(n_212), .B1(n_216), .B2(n_217), .Y(n_852) );
AOI21xp5_ASAP7_75t_L g853 ( .A1(n_701), .A2(n_220), .B(n_221), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_720), .A2(n_223), .B1(n_224), .B2(n_225), .Y(n_854) );
AND2x2_ASAP7_75t_L g855 ( .A(n_746), .B(n_226), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_716), .Y(n_856) );
OAI21xp5_ASAP7_75t_L g857 ( .A1(n_706), .A2(n_227), .B(n_228), .Y(n_857) );
A2O1A1Ixp33_ASAP7_75t_L g858 ( .A1(n_769), .A2(n_230), .B(n_232), .C(n_233), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_734), .A2(n_234), .B1(n_235), .B2(n_236), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_774), .A2(n_240), .B1(n_244), .B2(n_245), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_728), .A2(n_246), .B1(n_247), .B2(n_248), .Y(n_861) );
BUFx6f_ASAP7_75t_L g862 ( .A(n_773), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_733), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_728), .A2(n_253), .B1(n_257), .B2(n_260), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_720), .Y(n_865) );
AND2x2_ASAP7_75t_L g866 ( .A(n_732), .B(n_261), .Y(n_866) );
AND2x2_ASAP7_75t_L g867 ( .A(n_787), .B(n_262), .Y(n_867) );
AO21x2_ASAP7_75t_L g868 ( .A1(n_747), .A2(n_269), .B(n_273), .Y(n_868) );
OAI22xp5_ASAP7_75t_L g869 ( .A1(n_706), .A2(n_274), .B1(n_277), .B2(n_279), .Y(n_869) );
AND2x2_ASAP7_75t_L g870 ( .A(n_725), .B(n_280), .Y(n_870) );
NAND3xp33_ASAP7_75t_L g871 ( .A(n_758), .B(n_282), .C(n_283), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_750), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g873 ( .A1(n_700), .A2(n_284), .B1(n_288), .B2(n_703), .Y(n_873) );
OR2x2_ASAP7_75t_L g874 ( .A(n_700), .B(n_703), .Y(n_874) );
AND2x2_ASAP7_75t_L g875 ( .A(n_708), .B(n_771), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_770), .Y(n_876) );
AOI21xp5_ASAP7_75t_L g877 ( .A1(n_701), .A2(n_747), .B(n_731), .Y(n_877) );
NOR2xp33_ASAP7_75t_L g878 ( .A(n_748), .B(n_781), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_719), .B(n_762), .Y(n_879) );
O2A1O1Ixp33_ASAP7_75t_L g880 ( .A1(n_778), .A2(n_751), .B(n_739), .C(n_782), .Y(n_880) );
AOI221xp5_ASAP7_75t_L g881 ( .A1(n_778), .A2(n_753), .B1(n_739), .B2(n_782), .C(n_793), .Y(n_881) );
AND2x2_ASAP7_75t_L g882 ( .A(n_762), .B(n_718), .Y(n_882) );
BUFx10_ASAP7_75t_L g883 ( .A(n_773), .Y(n_883) );
AO221x2_ASAP7_75t_L g884 ( .A1(n_722), .A2(n_753), .B1(n_789), .B2(n_793), .C(n_730), .Y(n_884) );
INVx1_ASAP7_75t_SL g885 ( .A(n_780), .Y(n_885) );
OAI22xp5_ASAP7_75t_L g886 ( .A1(n_761), .A2(n_789), .B1(n_780), .B2(n_777), .Y(n_886) );
INVx1_ASAP7_75t_SL g887 ( .A(n_777), .Y(n_887) );
INVx2_ASAP7_75t_L g888 ( .A(n_803), .Y(n_888) );
AND2x2_ASAP7_75t_L g889 ( .A(n_837), .B(n_743), .Y(n_889) );
OA21x2_ASAP7_75t_L g890 ( .A1(n_877), .A2(n_727), .B(n_754), .Y(n_890) );
HB1xp67_ASAP7_75t_L g891 ( .A(n_821), .Y(n_891) );
INVx2_ASAP7_75t_L g892 ( .A(n_874), .Y(n_892) );
BUFx3_ASAP7_75t_L g893 ( .A(n_883), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_799), .B(n_715), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_797), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_810), .Y(n_896) );
OR2x2_ASAP7_75t_L g897 ( .A(n_832), .B(n_743), .Y(n_897) );
INVx2_ASAP7_75t_L g898 ( .A(n_856), .Y(n_898) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_798), .B(n_731), .Y(n_899) );
INVx4_ASAP7_75t_R g900 ( .A(n_830), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_822), .Y(n_901) );
AND2x2_ASAP7_75t_L g902 ( .A(n_863), .B(n_777), .Y(n_902) );
INVx2_ASAP7_75t_L g903 ( .A(n_802), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_825), .Y(n_904) );
BUFx6f_ASAP7_75t_L g905 ( .A(n_826), .Y(n_905) );
INVx2_ASAP7_75t_L g906 ( .A(n_802), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_828), .Y(n_907) );
AND2x2_ASAP7_75t_L g908 ( .A(n_876), .B(n_713), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_833), .B(n_783), .Y(n_909) );
AND2x4_ASAP7_75t_L g910 ( .A(n_845), .B(n_791), .Y(n_910) );
INVx2_ASAP7_75t_L g911 ( .A(n_802), .Y(n_911) );
NOR2xp33_ASAP7_75t_L g912 ( .A(n_878), .B(n_794), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_807), .Y(n_913) );
INVx2_ASAP7_75t_L g914 ( .A(n_826), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_823), .Y(n_915) );
AND2x2_ASAP7_75t_L g916 ( .A(n_865), .B(n_790), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_824), .Y(n_917) );
BUFx6f_ASAP7_75t_L g918 ( .A(n_826), .Y(n_918) );
INVx2_ASAP7_75t_L g919 ( .A(n_862), .Y(n_919) );
AOI221xp5_ASAP7_75t_L g920 ( .A1(n_817), .A2(n_749), .B1(n_786), .B2(n_744), .C(n_792), .Y(n_920) );
INVx2_ASAP7_75t_L g921 ( .A(n_862), .Y(n_921) );
INVx6_ASAP7_75t_L g922 ( .A(n_875), .Y(n_922) );
HB1xp67_ASAP7_75t_L g923 ( .A(n_829), .Y(n_923) );
BUFx2_ASAP7_75t_L g924 ( .A(n_845), .Y(n_924) );
OR2x2_ASAP7_75t_L g925 ( .A(n_879), .B(n_755), .Y(n_925) );
BUFx6f_ASAP7_75t_L g926 ( .A(n_862), .Y(n_926) );
INVx2_ASAP7_75t_L g927 ( .A(n_827), .Y(n_927) );
BUFx6f_ASAP7_75t_L g928 ( .A(n_845), .Y(n_928) );
AND2x2_ASAP7_75t_L g929 ( .A(n_805), .B(n_795), .Y(n_929) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_819), .B(n_756), .Y(n_930) );
AND2x2_ASAP7_75t_L g931 ( .A(n_805), .B(n_772), .Y(n_931) );
INVx3_ASAP7_75t_L g932 ( .A(n_846), .Y(n_932) );
INVx2_ASAP7_75t_L g933 ( .A(n_847), .Y(n_933) );
OAI22xp5_ASAP7_75t_L g934 ( .A1(n_850), .A2(n_846), .B1(n_806), .B2(n_812), .Y(n_934) );
AND2x2_ASAP7_75t_L g935 ( .A(n_816), .B(n_809), .Y(n_935) );
INVx2_ASAP7_75t_L g936 ( .A(n_800), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_831), .Y(n_937) );
AND2x2_ASAP7_75t_L g938 ( .A(n_882), .B(n_870), .Y(n_938) );
OR2x2_ASAP7_75t_SL g939 ( .A(n_871), .B(n_872), .Y(n_939) );
INVx2_ASAP7_75t_SL g940 ( .A(n_844), .Y(n_940) );
INVx1_ASAP7_75t_L g941 ( .A(n_801), .Y(n_941) );
INVx2_ASAP7_75t_L g942 ( .A(n_834), .Y(n_942) );
AND2x2_ASAP7_75t_L g943 ( .A(n_844), .B(n_804), .Y(n_943) );
INVx2_ASAP7_75t_L g944 ( .A(n_834), .Y(n_944) );
BUFx2_ASAP7_75t_L g945 ( .A(n_801), .Y(n_945) );
BUFx3_ASAP7_75t_L g946 ( .A(n_830), .Y(n_946) );
AO21x2_ASAP7_75t_L g947 ( .A1(n_886), .A2(n_880), .B(n_796), .Y(n_947) );
AND2x2_ASAP7_75t_L g948 ( .A(n_804), .B(n_885), .Y(n_948) );
HB1xp67_ASAP7_75t_L g949 ( .A(n_842), .Y(n_949) );
BUFx3_ASAP7_75t_L g950 ( .A(n_887), .Y(n_950) );
AND2x2_ASAP7_75t_L g951 ( .A(n_867), .B(n_866), .Y(n_951) );
INVx2_ASAP7_75t_L g952 ( .A(n_868), .Y(n_952) );
AND2x2_ASAP7_75t_L g953 ( .A(n_808), .B(n_887), .Y(n_953) );
AND2x4_ASAP7_75t_L g954 ( .A(n_857), .B(n_855), .Y(n_954) );
INVx2_ASAP7_75t_L g955 ( .A(n_868), .Y(n_955) );
INVx3_ASAP7_75t_L g956 ( .A(n_884), .Y(n_956) );
INVxp67_ASAP7_75t_SL g957 ( .A(n_854), .Y(n_957) );
OAI22xp33_ASAP7_75t_L g958 ( .A1(n_854), .A2(n_820), .B1(n_857), .B2(n_873), .Y(n_958) );
AND2x2_ASAP7_75t_L g959 ( .A(n_813), .B(n_861), .Y(n_959) );
INVx2_ASAP7_75t_L g960 ( .A(n_886), .Y(n_960) );
NOR2xp33_ASAP7_75t_L g961 ( .A(n_838), .B(n_814), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_851), .A2(n_796), .B1(n_864), .B2(n_881), .Y(n_962) );
OR2x2_ASAP7_75t_L g963 ( .A(n_839), .B(n_858), .Y(n_963) );
BUFx6f_ASAP7_75t_L g964 ( .A(n_818), .Y(n_964) );
AND2x4_ASAP7_75t_L g965 ( .A(n_811), .B(n_815), .Y(n_965) );
AND2x2_ASAP7_75t_L g966 ( .A(n_849), .B(n_835), .Y(n_966) );
INVx2_ASAP7_75t_L g967 ( .A(n_869), .Y(n_967) );
BUFx2_ASAP7_75t_L g968 ( .A(n_852), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g969 ( .A(n_892), .B(n_840), .Y(n_969) );
AND2x4_ASAP7_75t_L g970 ( .A(n_932), .B(n_853), .Y(n_970) );
OAI221xp5_ASAP7_75t_SL g971 ( .A1(n_943), .A2(n_859), .B1(n_860), .B2(n_836), .C(n_843), .Y(n_971) );
NOR2xp33_ASAP7_75t_R g972 ( .A(n_946), .B(n_841), .Y(n_972) );
AND2x2_ASAP7_75t_L g973 ( .A(n_938), .B(n_848), .Y(n_973) );
HB1xp67_ASAP7_75t_L g974 ( .A(n_891), .Y(n_974) );
AND2x2_ASAP7_75t_L g975 ( .A(n_938), .B(n_898), .Y(n_975) );
AND4x1_ASAP7_75t_L g976 ( .A(n_900), .B(n_961), .C(n_946), .D(n_943), .Y(n_976) );
HB1xp67_ASAP7_75t_L g977 ( .A(n_923), .Y(n_977) );
AND2x2_ASAP7_75t_L g978 ( .A(n_898), .B(n_888), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_895), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g980 ( .A(n_935), .B(n_901), .Y(n_980) );
INVx1_ASAP7_75t_L g981 ( .A(n_896), .Y(n_981) );
AND2x2_ASAP7_75t_L g982 ( .A(n_888), .B(n_901), .Y(n_982) );
INVx2_ASAP7_75t_L g983 ( .A(n_903), .Y(n_983) );
AND2x4_ASAP7_75t_L g984 ( .A(n_932), .B(n_924), .Y(n_984) );
INVx2_ASAP7_75t_L g985 ( .A(n_903), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_904), .Y(n_986) );
AND2x2_ASAP7_75t_L g987 ( .A(n_915), .B(n_917), .Y(n_987) );
INVx2_ASAP7_75t_L g988 ( .A(n_906), .Y(n_988) );
O2A1O1Ixp33_ASAP7_75t_SL g989 ( .A1(n_958), .A2(n_932), .B(n_940), .C(n_957), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_907), .Y(n_990) );
BUFx3_ASAP7_75t_L g991 ( .A(n_893), .Y(n_991) );
AND2x2_ASAP7_75t_L g992 ( .A(n_936), .B(n_956), .Y(n_992) );
OR2x2_ASAP7_75t_L g993 ( .A(n_956), .B(n_936), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_913), .Y(n_994) );
INVx2_ASAP7_75t_L g995 ( .A(n_911), .Y(n_995) );
AND2x2_ASAP7_75t_L g996 ( .A(n_956), .B(n_889), .Y(n_996) );
NAND4xp25_ASAP7_75t_L g997 ( .A(n_912), .B(n_948), .C(n_934), .D(n_951), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_897), .Y(n_998) );
AND2x2_ASAP7_75t_L g999 ( .A(n_889), .B(n_902), .Y(n_999) );
AND2x2_ASAP7_75t_L g1000 ( .A(n_902), .B(n_941), .Y(n_1000) );
OAI221xp5_ASAP7_75t_SL g1001 ( .A1(n_929), .A2(n_940), .B1(n_931), .B2(n_962), .C(n_945), .Y(n_1001) );
BUFx6f_ASAP7_75t_L g1002 ( .A(n_905), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_897), .Y(n_1003) );
INVx2_ASAP7_75t_L g1004 ( .A(n_911), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_922), .Y(n_1005) );
OAI22xp5_ASAP7_75t_SL g1006 ( .A1(n_928), .A2(n_922), .B1(n_939), .B2(n_949), .Y(n_1006) );
INVx2_ASAP7_75t_L g1007 ( .A(n_960), .Y(n_1007) );
HB1xp67_ASAP7_75t_L g1008 ( .A(n_950), .Y(n_1008) );
INVx3_ASAP7_75t_L g1009 ( .A(n_928), .Y(n_1009) );
AND2x2_ASAP7_75t_L g1010 ( .A(n_941), .B(n_899), .Y(n_1010) );
INVx1_ASAP7_75t_L g1011 ( .A(n_922), .Y(n_1011) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_916), .B(n_908), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_916), .B(n_908), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_894), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_937), .B(n_953), .Y(n_1015) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_954), .B(n_928), .Y(n_1016) );
BUFx3_ASAP7_75t_L g1017 ( .A(n_893), .Y(n_1017) );
INVxp67_ASAP7_75t_SL g1018 ( .A(n_928), .Y(n_1018) );
INVx2_ASAP7_75t_L g1019 ( .A(n_960), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_954), .B(n_914), .Y(n_1020) );
INVx2_ASAP7_75t_L g1021 ( .A(n_933), .Y(n_1021) );
BUFx2_ASAP7_75t_L g1022 ( .A(n_910), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_919), .B(n_921), .Y(n_1023) );
INVx4_ASAP7_75t_SL g1024 ( .A(n_910), .Y(n_1024) );
OR2x2_ASAP7_75t_L g1025 ( .A(n_925), .B(n_909), .Y(n_1025) );
AOI22xp5_ASAP7_75t_L g1026 ( .A1(n_966), .A2(n_959), .B1(n_968), .B2(n_967), .Y(n_1026) );
AND2x4_ASAP7_75t_L g1027 ( .A(n_910), .B(n_905), .Y(n_1027) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_947), .B(n_925), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_959), .B(n_966), .Y(n_1029) );
OR2x2_ASAP7_75t_L g1030 ( .A(n_939), .B(n_947), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_930), .B(n_905), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_918), .B(n_926), .Y(n_1032) );
NAND4xp25_ASAP7_75t_L g1033 ( .A(n_963), .B(n_920), .C(n_967), .D(n_965), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_918), .B(n_926), .Y(n_1034) );
AOI31xp33_ASAP7_75t_L g1035 ( .A1(n_963), .A2(n_965), .A3(n_942), .B(n_944), .Y(n_1035) );
OAI21xp5_ASAP7_75t_L g1036 ( .A1(n_969), .A2(n_965), .B(n_944), .Y(n_1036) );
OR2x2_ASAP7_75t_L g1037 ( .A(n_975), .B(n_918), .Y(n_1037) );
INVx3_ASAP7_75t_L g1038 ( .A(n_991), .Y(n_1038) );
OR2x2_ASAP7_75t_L g1039 ( .A(n_975), .B(n_926), .Y(n_1039) );
INVx1_ASAP7_75t_L g1040 ( .A(n_979), .Y(n_1040) );
INVx2_ASAP7_75t_L g1041 ( .A(n_978), .Y(n_1041) );
AND2x4_ASAP7_75t_L g1042 ( .A(n_1024), .B(n_926), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_999), .B(n_952), .Y(n_1043) );
INVx3_ASAP7_75t_L g1044 ( .A(n_991), .Y(n_1044) );
INVx1_ASAP7_75t_L g1045 ( .A(n_981), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_986), .Y(n_1046) );
NAND2x1p5_ASAP7_75t_L g1047 ( .A(n_1017), .B(n_927), .Y(n_1047) );
NAND2xp5_ASAP7_75t_L g1048 ( .A(n_1015), .B(n_955), .Y(n_1048) );
INVx2_ASAP7_75t_L g1049 ( .A(n_1021), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g1050 ( .A(n_998), .B(n_955), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_990), .Y(n_1051) );
AND2x2_ASAP7_75t_L g1052 ( .A(n_992), .B(n_890), .Y(n_1052) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_1003), .B(n_964), .Y(n_1053) );
OR2x2_ASAP7_75t_L g1054 ( .A(n_974), .B(n_890), .Y(n_1054) );
OR2x2_ASAP7_75t_L g1055 ( .A(n_977), .B(n_890), .Y(n_1055) );
NAND2xp33_ASAP7_75t_SL g1056 ( .A(n_1006), .B(n_964), .Y(n_1056) );
NAND2x1_ASAP7_75t_L g1057 ( .A(n_984), .B(n_964), .Y(n_1057) );
INVx2_ASAP7_75t_L g1058 ( .A(n_982), .Y(n_1058) );
INVxp67_ASAP7_75t_SL g1059 ( .A(n_983), .Y(n_1059) );
INVx1_ASAP7_75t_L g1060 ( .A(n_994), .Y(n_1060) );
NOR2xp33_ASAP7_75t_L g1061 ( .A(n_1029), .B(n_997), .Y(n_1061) );
AND2x4_ASAP7_75t_L g1062 ( .A(n_1024), .B(n_984), .Y(n_1062) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_996), .B(n_987), .Y(n_1063) );
NAND2x1_ASAP7_75t_L g1064 ( .A(n_984), .B(n_1022), .Y(n_1064) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_1026), .B(n_1014), .Y(n_1065) );
NAND2xp5_ASAP7_75t_L g1066 ( .A(n_1010), .B(n_1000), .Y(n_1066) );
INVxp67_ASAP7_75t_L g1067 ( .A(n_1008), .Y(n_1067) );
INVx4_ASAP7_75t_L g1068 ( .A(n_1009), .Y(n_1068) );
INVx1_ASAP7_75t_L g1069 ( .A(n_980), .Y(n_1069) );
CKINVDCx16_ASAP7_75t_R g1070 ( .A(n_972), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_993), .Y(n_1071) );
INVx2_ASAP7_75t_L g1072 ( .A(n_1021), .Y(n_1072) );
INVx2_ASAP7_75t_L g1073 ( .A(n_983), .Y(n_1073) );
AND2x4_ASAP7_75t_L g1074 ( .A(n_1024), .B(n_1016), .Y(n_1074) );
AND2x4_ASAP7_75t_L g1075 ( .A(n_1024), .B(n_1016), .Y(n_1075) );
OR2x2_ASAP7_75t_L g1076 ( .A(n_1012), .B(n_1013), .Y(n_1076) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_1028), .B(n_1025), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g1078 ( .A(n_1028), .B(n_1025), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1023), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_1005), .B(n_1011), .Y(n_1080) );
OR2x2_ASAP7_75t_L g1081 ( .A(n_1020), .B(n_1018), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_985), .Y(n_1082) );
HB1xp67_ASAP7_75t_L g1083 ( .A(n_1067), .Y(n_1083) );
NAND2xp5_ASAP7_75t_L g1084 ( .A(n_1069), .B(n_973), .Y(n_1084) );
OR2x6_ASAP7_75t_L g1085 ( .A(n_1064), .B(n_1030), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_1063), .B(n_1031), .Y(n_1086) );
INVx2_ASAP7_75t_L g1087 ( .A(n_1049), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1040), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1089 ( .A(n_1076), .B(n_1031), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1045), .Y(n_1090) );
OR2x2_ASAP7_75t_L g1091 ( .A(n_1077), .B(n_1033), .Y(n_1091) );
AOI21xp5_ASAP7_75t_L g1092 ( .A1(n_1056), .A2(n_989), .B(n_1035), .Y(n_1092) );
AOI211xp5_ASAP7_75t_L g1093 ( .A1(n_1061), .A2(n_989), .B(n_1001), .C(n_971), .Y(n_1093) );
AOI21xp33_ASAP7_75t_SL g1094 ( .A1(n_1070), .A2(n_976), .B(n_1030), .Y(n_1094) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_1043), .B(n_1027), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1046), .Y(n_1096) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_1066), .B(n_1027), .Y(n_1097) );
HB1xp67_ASAP7_75t_L g1098 ( .A(n_1067), .Y(n_1098) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1058), .Y(n_1099) );
OAI221xp5_ASAP7_75t_SL g1100 ( .A1(n_1061), .A2(n_995), .B1(n_1004), .B2(n_985), .C(n_988), .Y(n_1100) );
INVx2_ASAP7_75t_SL g1101 ( .A(n_1038), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1051), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_1052), .B(n_1004), .Y(n_1103) );
INVx2_ASAP7_75t_L g1104 ( .A(n_1049), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1060), .Y(n_1105) );
INVx2_ASAP7_75t_L g1106 ( .A(n_1072), .Y(n_1106) );
OR2x6_ASAP7_75t_L g1107 ( .A(n_1062), .B(n_970), .Y(n_1107) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1041), .Y(n_1108) );
AND2x2_ASAP7_75t_SL g1109 ( .A(n_1062), .B(n_970), .Y(n_1109) );
AOI221x1_ASAP7_75t_L g1110 ( .A1(n_1056), .A2(n_1034), .B1(n_1032), .B2(n_1002), .C(n_1019), .Y(n_1110) );
INVx2_ASAP7_75t_SL g1111 ( .A(n_1044), .Y(n_1111) );
OR2x2_ASAP7_75t_L g1112 ( .A(n_1077), .B(n_1007), .Y(n_1112) );
OR2x2_ASAP7_75t_L g1113 ( .A(n_1078), .B(n_1019), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1088), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1090), .Y(n_1115) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_1091), .B(n_1065), .Y(n_1116) );
NAND2xp5_ASAP7_75t_L g1117 ( .A(n_1091), .B(n_1079), .Y(n_1117) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1096), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1102), .Y(n_1119) );
AOI22xp33_ASAP7_75t_SL g1120 ( .A1(n_1109), .A2(n_1074), .B1(n_1075), .B2(n_1071), .Y(n_1120) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1105), .Y(n_1121) );
OAI22xp5_ASAP7_75t_L g1122 ( .A1(n_1093), .A2(n_1075), .B1(n_1037), .B2(n_1039), .Y(n_1122) );
NAND3xp33_ASAP7_75t_L g1123 ( .A(n_1083), .B(n_1055), .C(n_1054), .Y(n_1123) );
NOR2xp33_ASAP7_75t_L g1124 ( .A(n_1098), .B(n_1048), .Y(n_1124) );
XNOR2xp5_ASAP7_75t_L g1125 ( .A(n_1089), .B(n_1080), .Y(n_1125) );
A2O1A1Ixp33_ASAP7_75t_L g1126 ( .A1(n_1094), .A2(n_1042), .B(n_1081), .C(n_1057), .Y(n_1126) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1097), .Y(n_1127) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1099), .Y(n_1128) );
OAI22xp5_ASAP7_75t_L g1129 ( .A1(n_1092), .A2(n_1047), .B1(n_1068), .B2(n_1059), .Y(n_1129) );
NAND2xp5_ASAP7_75t_L g1130 ( .A(n_1099), .B(n_1053), .Y(n_1130) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1128), .Y(n_1131) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1114), .Y(n_1132) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1115), .Y(n_1133) );
XNOR2x1_ASAP7_75t_L g1134 ( .A(n_1122), .B(n_1086), .Y(n_1134) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1118), .Y(n_1135) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1119), .Y(n_1136) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1121), .Y(n_1137) );
XNOR2x1_ASAP7_75t_L g1138 ( .A(n_1125), .B(n_1095), .Y(n_1138) );
OAI21xp5_ASAP7_75t_L g1139 ( .A1(n_1129), .A2(n_1101), .B(n_1111), .Y(n_1139) );
NOR2xp33_ASAP7_75t_L g1140 ( .A(n_1116), .B(n_1084), .Y(n_1140) );
NAND2xp5_ASAP7_75t_L g1141 ( .A(n_1124), .B(n_1108), .Y(n_1141) );
NAND4xp25_ASAP7_75t_L g1142 ( .A(n_1126), .B(n_1110), .C(n_1100), .D(n_1036), .Y(n_1142) );
OAI21xp33_ASAP7_75t_L g1143 ( .A1(n_1134), .A2(n_1120), .B(n_1117), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1131), .Y(n_1144) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1132), .Y(n_1145) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1133), .Y(n_1146) );
NAND2xp5_ASAP7_75t_L g1147 ( .A(n_1140), .B(n_1127), .Y(n_1147) );
NAND2xp5_ASAP7_75t_L g1148 ( .A(n_1140), .B(n_1123), .Y(n_1148) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1135), .Y(n_1149) );
AOI21xp33_ASAP7_75t_L g1150 ( .A1(n_1139), .A2(n_1085), .B(n_1130), .Y(n_1150) );
AOI221xp5_ASAP7_75t_L g1151 ( .A1(n_1143), .A2(n_1142), .B1(n_1136), .B2(n_1137), .C(n_1141), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1145), .Y(n_1152) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1146), .Y(n_1153) );
AO22x2_ASAP7_75t_L g1154 ( .A1(n_1148), .A2(n_1138), .B1(n_1112), .B2(n_1113), .Y(n_1154) );
OR2x2_ASAP7_75t_L g1155 ( .A(n_1152), .B(n_1147), .Y(n_1155) );
HB1xp67_ASAP7_75t_L g1156 ( .A(n_1153), .Y(n_1156) );
AND2x2_ASAP7_75t_SL g1157 ( .A(n_1151), .B(n_1149), .Y(n_1157) );
NAND3xp33_ASAP7_75t_L g1158 ( .A(n_1154), .B(n_1150), .C(n_1144), .Y(n_1158) );
AOI22xp5_ASAP7_75t_L g1159 ( .A1(n_1157), .A2(n_1107), .B1(n_1103), .B2(n_1106), .Y(n_1159) );
AND4x1_ASAP7_75t_L g1160 ( .A(n_1158), .B(n_1032), .C(n_1034), .D(n_1107), .Y(n_1160) );
CKINVDCx20_ASAP7_75t_R g1161 ( .A(n_1159), .Y(n_1161) );
AOI22xp5_ASAP7_75t_L g1162 ( .A1(n_1161), .A2(n_1156), .B1(n_1155), .B2(n_1160), .Y(n_1162) );
OAI22xp5_ASAP7_75t_L g1163 ( .A1(n_1162), .A2(n_1106), .B1(n_1087), .B2(n_1104), .Y(n_1163) );
AOI22xp33_ASAP7_75t_SL g1164 ( .A1(n_1163), .A2(n_1002), .B1(n_1050), .B2(n_1082), .Y(n_1164) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1164), .Y(n_1165) );
AOI21xp5_ASAP7_75t_L g1166 ( .A1(n_1165), .A2(n_1073), .B(n_1002), .Y(n_1166) );
endmodule