module fake_jpeg_2414_n_358 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_358);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_358;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_15),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_52),
.Y(n_83)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx5_ASAP7_75t_SL g111 ( 
.A(n_47),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_17),
.B(n_14),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_17),
.B(n_15),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_54),
.B(n_57),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_19),
.B(n_14),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_42),
.Y(n_60)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_42),
.Y(n_64)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g117 ( 
.A(n_65),
.Y(n_117)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_19),
.B(n_13),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_68),
.B(n_73),
.Y(n_118)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

BUFx4f_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_25),
.B(n_13),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_25),
.B(n_10),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_74),
.B(n_26),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_28),
.B(n_13),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_32),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_18),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_76),
.B(n_80),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_75),
.A2(n_22),
.B1(n_24),
.B2(n_37),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_78),
.A2(n_79),
.B1(n_113),
.B2(n_29),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_55),
.A2(n_38),
.B1(n_21),
.B2(n_41),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_47),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_84),
.B(n_86),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_47),
.Y(n_86)
);

BUFx6f_ASAP7_75t_SL g89 ( 
.A(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_26),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_58),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_95),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_56),
.A2(n_27),
.B1(n_36),
.B2(n_24),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g135 ( 
.A1(n_97),
.A2(n_116),
.B1(n_42),
.B2(n_39),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_51),
.B(n_32),
.Y(n_98)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_98),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_45),
.B(n_37),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_22),
.Y(n_126)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_106),
.Y(n_140)
);

BUFx10_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_72),
.A2(n_28),
.B1(n_24),
.B2(n_41),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_65),
.A2(n_27),
.B1(n_36),
.B2(n_18),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_67),
.B(n_21),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_16),
.C(n_31),
.Y(n_134)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_50),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_61),
.B(n_35),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_124),
.A2(n_35),
.B1(n_31),
.B2(n_33),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_126),
.B(n_164),
.Y(n_179)
);

OR2x4_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_83),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_128),
.B(n_137),
.Y(n_181)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_131),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_132),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_134),
.B(n_7),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_135),
.A2(n_141),
.B1(n_157),
.B2(n_159),
.Y(n_171)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_136),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_119),
.A2(n_16),
.B1(n_33),
.B2(n_71),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_139),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_92),
.A2(n_27),
.B1(n_70),
.B2(n_42),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_79),
.A2(n_63),
.B1(n_62),
.B2(n_42),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g172 ( 
.A1(n_142),
.A2(n_147),
.B1(n_103),
.B2(n_123),
.Y(n_172)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_143),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_97),
.A2(n_116),
.B1(n_115),
.B2(n_96),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_144),
.A2(n_123),
.B1(n_101),
.B2(n_102),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_76),
.A2(n_22),
.B1(n_29),
.B2(n_39),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_145),
.A2(n_151),
.B1(n_152),
.B2(n_143),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

INVxp33_ASAP7_75t_L g203 ( 
.A(n_146),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_29),
.B1(n_39),
.B2(n_2),
.Y(n_147)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_82),
.B(n_0),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_156),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_77),
.B(n_99),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_121),
.A2(n_29),
.B1(n_1),
.B2(n_2),
.Y(n_157)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_93),
.Y(n_158)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_121),
.A2(n_29),
.B1(n_1),
.B2(n_4),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_120),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_161),
.A2(n_162),
.B1(n_81),
.B2(n_85),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_120),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_162)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_104),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_91),
.B(n_5),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_7),
.Y(n_189)
);

A2O1A1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_105),
.A2(n_9),
.B(n_10),
.C(n_8),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_166),
.B(n_5),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_125),
.A2(n_81),
.B(n_114),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_167),
.A2(n_176),
.B(n_185),
.Y(n_214)
);

NOR3xp33_ASAP7_75t_L g236 ( 
.A(n_168),
.B(n_175),
.C(n_178),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_109),
.C(n_114),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_169),
.B(n_197),
.C(n_129),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_173),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_133),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_135),
.A2(n_85),
.B1(n_107),
.B2(n_110),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_156),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_166),
.A2(n_111),
.B(n_112),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_182),
.A2(n_200),
.B(n_134),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_160),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_184),
.B(n_187),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_132),
.B(n_111),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_188),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_163),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_107),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_189),
.B(n_168),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_138),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_135),
.A2(n_107),
.B1(n_110),
.B2(n_112),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_191),
.A2(n_149),
.B(n_136),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_193),
.A2(n_140),
.B1(n_164),
.B2(n_139),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_103),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_196),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_138),
.B(n_110),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_128),
.B(n_101),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_135),
.A2(n_7),
.B(n_8),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_140),
.B(n_102),
.Y(n_201)
);

XNOR2x1_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_188),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_126),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_205),
.B(n_223),
.Y(n_264)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_192),
.Y(n_207)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_207),
.Y(n_255)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_201),
.Y(n_208)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_208),
.Y(n_262)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_204),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_209),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_193),
.A2(n_137),
.B1(n_145),
.B2(n_153),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_210),
.A2(n_215),
.B1(n_221),
.B2(n_228),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_211),
.A2(n_222),
.B(n_188),
.Y(n_245)
);

OAI21xp33_ASAP7_75t_L g251 ( 
.A1(n_212),
.A2(n_203),
.B(n_175),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_220),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_131),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_217),
.A2(n_234),
.B(n_196),
.Y(n_248)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_201),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_178),
.A2(n_158),
.B1(n_150),
.B2(n_108),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_180),
.B(n_130),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_233),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_148),
.Y(n_225)
);

INVxp33_ASAP7_75t_L g238 ( 
.A(n_225),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_180),
.B(n_148),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_226),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_184),
.B(n_149),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_231),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_186),
.A2(n_200),
.B1(n_181),
.B2(n_195),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_181),
.A2(n_108),
.B1(n_127),
.B2(n_8),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_229),
.A2(n_215),
.B1(n_170),
.B2(n_194),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_181),
.A2(n_127),
.B1(n_179),
.B2(n_185),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_230),
.A2(n_170),
.B1(n_183),
.B2(n_194),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_202),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_235),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_185),
.A2(n_167),
.B(n_171),
.Y(n_234)
);

NOR2x1_ASAP7_75t_L g235 ( 
.A(n_177),
.B(n_188),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_179),
.B(n_189),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_219),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_240),
.A2(n_249),
.B1(n_251),
.B2(n_253),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_213),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_241),
.Y(n_285)
);

FAx1_ASAP7_75t_SL g243 ( 
.A(n_223),
.B(n_169),
.CI(n_190),
.CON(n_243),
.SN(n_243)
);

AO21x1_ASAP7_75t_L g268 ( 
.A1(n_243),
.A2(n_245),
.B(n_248),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_244),
.B(n_232),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_228),
.A2(n_172),
.B1(n_204),
.B2(n_192),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_217),
.Y(n_252)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

A2O1A1O1Ixp25_ASAP7_75t_L g254 ( 
.A1(n_219),
.A2(n_183),
.B(n_198),
.C(n_174),
.D(n_172),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_254),
.A2(n_234),
.B(n_218),
.Y(n_277)
);

INVx13_ASAP7_75t_L g256 ( 
.A(n_217),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_256),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_198),
.Y(n_258)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_224),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_258),
.Y(n_284)
);

AND2x6_ASAP7_75t_L g260 ( 
.A(n_211),
.B(n_172),
.Y(n_260)
);

AO21x2_ASAP7_75t_L g272 ( 
.A1(n_260),
.A2(n_214),
.B(n_222),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_174),
.Y(n_263)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_263),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_205),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_265),
.B(n_266),
.C(n_270),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_264),
.B(n_226),
.C(n_216),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_263),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_276),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_230),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_272),
.A2(n_280),
.B1(n_277),
.B2(n_248),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_235),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_257),
.Y(n_288)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_277),
.A2(n_247),
.B(n_261),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_259),
.A2(n_206),
.B1(n_214),
.B2(n_218),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_278),
.A2(n_284),
.B1(n_286),
.B2(n_249),
.Y(n_293)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_242),
.Y(n_279)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_279),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_252),
.A2(n_206),
.B1(n_218),
.B2(n_210),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_281),
.B(n_257),
.Y(n_289)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_242),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_238),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_246),
.A2(n_206),
.B1(n_220),
.B2(n_208),
.Y(n_286)
);

MAJx2_ASAP7_75t_L g319 ( 
.A(n_288),
.B(n_289),
.C(n_296),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_290),
.A2(n_272),
.B1(n_283),
.B2(n_267),
.Y(n_306)
);

INVxp33_ASAP7_75t_L g311 ( 
.A(n_291),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_247),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_297),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_293),
.A2(n_294),
.B1(n_295),
.B2(n_288),
.Y(n_316)
);

NOR3xp33_ASAP7_75t_SL g294 ( 
.A(n_285),
.B(n_241),
.C(n_236),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_271),
.A2(n_246),
.B1(n_239),
.B2(n_253),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_268),
.A2(n_245),
.B(n_254),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_266),
.B(n_268),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_298),
.A2(n_262),
.B(n_254),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_273),
.B(n_243),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_301),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_270),
.B(n_243),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_239),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_275),
.C(n_271),
.Y(n_305)
);

AO22x2_ASAP7_75t_L g303 ( 
.A1(n_283),
.A2(n_278),
.B1(n_286),
.B2(n_274),
.Y(n_303)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_303),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_317),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_306),
.A2(n_309),
.B1(n_315),
.B2(n_316),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_262),
.C(n_284),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_307),
.B(n_312),
.C(n_250),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_287),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_301),
.C(n_299),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_298),
.A2(n_272),
.B(n_256),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_272),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_300),
.A2(n_284),
.B1(n_272),
.B2(n_280),
.Y(n_315)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_303),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_318),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g337 ( 
.A(n_321),
.B(n_306),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_311),
.B(n_302),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_324),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_307),
.B(n_289),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_305),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_328),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_310),
.A2(n_303),
.B1(n_260),
.B2(n_297),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_326),
.A2(n_327),
.B1(n_329),
.B2(n_315),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_310),
.A2(n_303),
.B1(n_260),
.B2(n_292),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_318),
.A2(n_240),
.B1(n_256),
.B2(n_276),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_317),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_309),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_334),
.B(n_326),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_335),
.B(n_336),
.Y(n_343)
);

OAI322xp33_ASAP7_75t_L g336 ( 
.A1(n_330),
.A2(n_319),
.A3(n_313),
.B1(n_312),
.B2(n_308),
.C1(n_294),
.C2(n_314),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_337),
.A2(n_329),
.B1(n_320),
.B2(n_327),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_322),
.B(n_331),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_338),
.A2(n_207),
.B1(n_209),
.B2(n_199),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_308),
.C(n_313),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_339),
.B(n_340),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_322),
.B(n_319),
.C(n_255),
.Y(n_340)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_341),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_342),
.B(n_347),
.Y(n_349)
);

O2A1O1Ixp33_ASAP7_75t_SL g344 ( 
.A1(n_337),
.A2(n_229),
.B(n_221),
.C(n_172),
.Y(n_344)
);

OAI31xp33_ASAP7_75t_L g351 ( 
.A1(n_344),
.A2(n_334),
.A3(n_340),
.B(n_339),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_332),
.B(n_333),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_346),
.B(n_338),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_350),
.B(n_351),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_348),
.B(n_345),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_352),
.B(n_343),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_354),
.B(n_353),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_355),
.A2(n_349),
.B(n_342),
.Y(n_356)
);

AO21x1_ASAP7_75t_L g357 ( 
.A1(n_356),
.A2(n_349),
.B(n_344),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_357),
.B(n_199),
.Y(n_358)
);


endmodule