module fake_jpeg_13100_n_114 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_114);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_114;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx11_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_27),
.A2(n_29),
.B1(n_26),
.B2(n_28),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_16),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_28),
.B(n_33),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_35),
.Y(n_47)
);

AOI21xp33_ASAP7_75t_L g33 ( 
.A1(n_12),
.A2(n_0),
.B(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_16),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_36),
.B(n_25),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_20),
.A2(n_24),
.B1(n_19),
.B2(n_14),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_40),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_20),
.A2(n_9),
.B1(n_10),
.B2(n_19),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_14),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_44),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_57),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_21),
.C(n_23),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_62),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_63),
.B(n_64),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_31),
.A2(n_23),
.B1(n_25),
.B2(n_15),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_45),
.B1(n_48),
.B2(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_15),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_15),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_SL g73 ( 
.A(n_59),
.B(n_61),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_15),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_29),
.A2(n_41),
.B1(n_35),
.B2(n_34),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_36),
.B(n_29),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_49),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_30),
.B1(n_38),
.B2(n_50),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_80),
.B1(n_58),
.B2(n_74),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_54),
.A2(n_65),
.B1(n_55),
.B2(n_59),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_SL g83 ( 
.A(n_69),
.B(n_58),
.C(n_66),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_47),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_72),
.C(n_73),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_61),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_48),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_78),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_58),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_46),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_52),
.B(n_60),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_79),
.A2(n_75),
.B(n_70),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_58),
.A2(n_54),
.B1(n_50),
.B2(n_59),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_82),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_84),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_72),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_90),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_73),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_80),
.B1(n_77),
.B2(n_76),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_84),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_96),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_89),
.A2(n_87),
.B1(n_81),
.B2(n_86),
.Y(n_94)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

OAI31xp33_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_83),
.A3(n_88),
.B(n_85),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_97),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_100),
.B(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_103),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_92),
.C(n_96),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_105),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

NOR2x1_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_102),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_108),
.A2(n_99),
.B(n_101),
.Y(n_111)
);

AOI322xp5_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_111),
.A3(n_107),
.B1(n_101),
.B2(n_97),
.C1(n_105),
.C2(n_93),
.Y(n_113)
);

BUFx24_ASAP7_75t_SL g114 ( 
.A(n_113),
.Y(n_114)
);


endmodule