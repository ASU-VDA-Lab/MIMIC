module fake_netlist_6_3857_n_1904 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1904);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1904;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_268;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_811;
wire n_683;
wire n_474;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1851;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g179 ( 
.A(n_72),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_68),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_119),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_32),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_149),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_42),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_105),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_127),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_116),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_68),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_133),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_94),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_65),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_82),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_59),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_16),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g196 ( 
.A(n_29),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_69),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_97),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_12),
.Y(n_199)
);

BUFx8_ASAP7_75t_SL g200 ( 
.A(n_90),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_112),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_86),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_79),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_164),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_67),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_35),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_52),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_135),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_161),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_36),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_31),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_44),
.Y(n_212)
);

BUFx10_ASAP7_75t_L g213 ( 
.A(n_88),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_24),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_89),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_139),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_25),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_42),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_129),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_78),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_177),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_156),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_155),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_172),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_99),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_101),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_0),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_71),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_115),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_70),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_83),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_150),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_59),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_76),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_80),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_14),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_43),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_21),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_159),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_9),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_54),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_69),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_123),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_20),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_117),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_141),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_24),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_8),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_125),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_146),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_19),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_74),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_142),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_136),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_148),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_14),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_126),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_44),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_45),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_137),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_113),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_173),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_170),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_19),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_174),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_41),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_77),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_25),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_106),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_160),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_30),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_17),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_16),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_58),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_71),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_11),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_131),
.Y(n_278)
);

BUFx8_ASAP7_75t_SL g279 ( 
.A(n_165),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_114),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_122),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_30),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_107),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_138),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_53),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_43),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_166),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_47),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_40),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_54),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_38),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_62),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_10),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_98),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_81),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_0),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_41),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_84),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_134),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_104),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_12),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_67),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_162),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_39),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_100),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_26),
.Y(n_306)
);

BUFx2_ASAP7_75t_R g307 ( 
.A(n_167),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_70),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_93),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_176),
.Y(n_310)
);

BUFx5_ASAP7_75t_L g311 ( 
.A(n_56),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_37),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_11),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_36),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_73),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_152),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_75),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_64),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_144),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_53),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_109),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_1),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_2),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_143),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_96),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_22),
.Y(n_326)
);

BUFx10_ASAP7_75t_L g327 ( 
.A(n_9),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_118),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_35),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_85),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_163),
.Y(n_331)
);

BUFx10_ASAP7_75t_L g332 ( 
.A(n_23),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_92),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_22),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_37),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_2),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_52),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_10),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_7),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_111),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_158),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_102),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_40),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_62),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_175),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_18),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_38),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_147),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_49),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_7),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_34),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_48),
.Y(n_352)
);

BUFx10_ASAP7_75t_L g353 ( 
.A(n_56),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_8),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_171),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_168),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_200),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_196),
.Y(n_358)
);

BUFx2_ASAP7_75t_SL g359 ( 
.A(n_202),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_190),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_279),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_254),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_213),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_196),
.Y(n_364)
);

OR2x2_ASAP7_75t_L g365 ( 
.A(n_195),
.B(n_1),
.Y(n_365)
);

OR2x2_ASAP7_75t_L g366 ( 
.A(n_197),
.B(n_3),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_220),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_215),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_204),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_222),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_225),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_226),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_196),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_233),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_196),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_196),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_235),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_263),
.Y(n_378)
);

INVxp33_ASAP7_75t_SL g379 ( 
.A(n_184),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_196),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_196),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_327),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_236),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_240),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_270),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_251),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_266),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_280),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_327),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_230),
.B(n_3),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_196),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_278),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_311),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_311),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_311),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_283),
.Y(n_396)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_261),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_281),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_284),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_311),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_287),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_202),
.B(n_4),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_311),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_311),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_311),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_311),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_180),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_295),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_191),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_180),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_180),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_180),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_298),
.Y(n_413)
);

INVxp33_ASAP7_75t_L g414 ( 
.A(n_207),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_184),
.Y(n_415)
);

NOR2xp67_ASAP7_75t_L g416 ( 
.A(n_253),
.B(n_4),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_327),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_303),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_180),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_319),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_305),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_354),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_354),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_354),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_354),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_340),
.B(n_5),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_354),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_261),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_315),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_199),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_199),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_316),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g433 ( 
.A(n_212),
.B(n_5),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_214),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_317),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_214),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_269),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_269),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_183),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_183),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_217),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_185),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_210),
.B(n_290),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_347),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_228),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_340),
.B(n_6),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_365),
.A2(n_277),
.B1(n_352),
.B2(n_351),
.Y(n_447)
);

AND2x6_ASAP7_75t_L g448 ( 
.A(n_409),
.B(n_253),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_410),
.Y(n_449)
);

AND2x2_ASAP7_75t_SL g450 ( 
.A(n_390),
.B(n_247),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_397),
.B(n_185),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_428),
.B(n_446),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_410),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_359),
.B(n_253),
.Y(n_454)
);

AND3x2_ASAP7_75t_L g455 ( 
.A(n_402),
.B(n_182),
.C(n_247),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_380),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_411),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_411),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_412),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_441),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_380),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_443),
.B(n_299),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_407),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_426),
.B(n_186),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_412),
.B(n_186),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_443),
.B(n_432),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_407),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_419),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_416),
.B(n_316),
.Y(n_469)
);

INVx4_ASAP7_75t_L g470 ( 
.A(n_409),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_427),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_415),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_427),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_419),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_422),
.B(n_423),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_422),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_358),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_423),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_367),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_358),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_416),
.B(n_299),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_364),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_424),
.B(n_189),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_424),
.B(n_299),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_432),
.B(n_210),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_425),
.B(n_364),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_359),
.B(n_181),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_425),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_373),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_373),
.B(n_179),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_375),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_375),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_376),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_376),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_381),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_381),
.Y(n_496)
);

NAND2xp33_ASAP7_75t_L g497 ( 
.A(n_445),
.B(n_192),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_391),
.Y(n_498)
);

AND2x6_ASAP7_75t_L g499 ( 
.A(n_409),
.B(n_218),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_391),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_393),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_393),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_394),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_432),
.B(n_189),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_394),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_395),
.B(n_221),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_395),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_400),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_400),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_403),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_403),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_404),
.B(n_290),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_370),
.B(n_187),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_404),
.B(n_193),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_405),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_405),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_360),
.B(n_368),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_406),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_406),
.B(n_223),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_372),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_369),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_430),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_430),
.B(n_431),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_431),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_454),
.B(n_374),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_466),
.B(n_444),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_456),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_466),
.B(n_444),
.Y(n_528)
);

INVxp33_ASAP7_75t_L g529 ( 
.A(n_466),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_463),
.Y(n_530)
);

OAI21xp33_ASAP7_75t_SL g531 ( 
.A1(n_450),
.A2(n_320),
.B(n_219),
.Y(n_531)
);

AND2x6_ASAP7_75t_L g532 ( 
.A(n_481),
.B(n_218),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_513),
.B(n_377),
.Y(n_533)
);

NAND2xp33_ASAP7_75t_SL g534 ( 
.A(n_464),
.B(n_219),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_470),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_504),
.B(n_362),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_490),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_456),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_463),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_462),
.B(n_434),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_SL g541 ( 
.A(n_479),
.B(n_307),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_521),
.B(n_383),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_454),
.B(n_384),
.Y(n_543)
);

NOR2x1p5_ASAP7_75t_L g544 ( 
.A(n_520),
.B(n_357),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_456),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_472),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_470),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_462),
.B(n_386),
.Y(n_548)
);

INVx8_ASAP7_75t_L g549 ( 
.A(n_469),
.Y(n_549)
);

BUFx8_ASAP7_75t_SL g550 ( 
.A(n_460),
.Y(n_550)
);

INVx4_ASAP7_75t_L g551 ( 
.A(n_480),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_489),
.Y(n_552)
);

OR2x6_ASAP7_75t_L g553 ( 
.A(n_520),
.B(n_365),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_SL g554 ( 
.A1(n_447),
.A2(n_363),
.B1(n_237),
.B2(n_259),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_450),
.A2(n_320),
.B1(n_366),
.B2(n_433),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_450),
.A2(n_366),
.B1(n_433),
.B2(n_347),
.Y(n_556)
);

INVx6_ASAP7_75t_L g557 ( 
.A(n_470),
.Y(n_557)
);

INVx5_ASAP7_75t_L g558 ( 
.A(n_499),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_463),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_462),
.B(n_387),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_487),
.B(n_392),
.Y(n_561)
);

OAI21xp33_ASAP7_75t_SL g562 ( 
.A1(n_452),
.A2(n_464),
.B(n_512),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_452),
.B(n_396),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_470),
.Y(n_564)
);

OR2x6_ASAP7_75t_L g565 ( 
.A(n_520),
.B(n_308),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_489),
.Y(n_566)
);

AND2x6_ASAP7_75t_L g567 ( 
.A(n_481),
.B(n_218),
.Y(n_567)
);

AO22x2_ASAP7_75t_L g568 ( 
.A1(n_447),
.A2(n_249),
.B1(n_344),
.B2(n_306),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_491),
.Y(n_569)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_485),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_517),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_521),
.B(n_399),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_491),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_504),
.B(n_451),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_497),
.A2(n_440),
.B1(n_442),
.B2(n_439),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_512),
.B(n_434),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_492),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_469),
.B(n_401),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_469),
.B(n_408),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_451),
.B(n_362),
.Y(n_580)
);

INVx1_ASAP7_75t_SL g581 ( 
.A(n_517),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_514),
.B(n_418),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_514),
.B(n_363),
.Y(n_583)
);

BUFx10_ASAP7_75t_L g584 ( 
.A(n_469),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_471),
.Y(n_585)
);

BUFx10_ASAP7_75t_L g586 ( 
.A(n_469),
.Y(n_586)
);

INVx4_ASAP7_75t_L g587 ( 
.A(n_480),
.Y(n_587)
);

BUFx8_ASAP7_75t_SL g588 ( 
.A(n_460),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_492),
.Y(n_589)
);

NAND2xp33_ASAP7_75t_L g590 ( 
.A(n_448),
.B(n_218),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_472),
.A2(n_379),
.B1(n_435),
.B2(n_429),
.Y(n_591)
);

INVxp33_ASAP7_75t_L g592 ( 
.A(n_485),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_493),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_490),
.Y(n_594)
);

OAI22xp33_ASAP7_75t_SL g595 ( 
.A1(n_465),
.A2(n_382),
.B1(n_389),
.B2(n_417),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_465),
.B(n_421),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_471),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_471),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_456),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_493),
.B(n_203),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_485),
.B(n_361),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_490),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_473),
.Y(n_603)
);

AND2x6_ASAP7_75t_L g604 ( 
.A(n_481),
.B(n_218),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_496),
.B(n_333),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_SL g606 ( 
.A(n_483),
.B(n_245),
.Y(n_606)
);

NAND2xp33_ASAP7_75t_L g607 ( 
.A(n_448),
.B(n_271),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_496),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_512),
.B(n_436),
.Y(n_609)
);

BUFx4f_ASAP7_75t_L g610 ( 
.A(n_480),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_500),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_483),
.B(n_414),
.Y(n_612)
);

OR2x6_ASAP7_75t_L g613 ( 
.A(n_523),
.B(n_308),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g614 ( 
.A(n_490),
.B(n_188),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_500),
.B(n_371),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_501),
.B(n_378),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_501),
.B(n_385),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_490),
.B(n_213),
.Y(n_618)
);

INVx1_ASAP7_75t_SL g619 ( 
.A(n_455),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_502),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_502),
.B(n_388),
.Y(n_621)
);

NAND3xp33_ASAP7_75t_L g622 ( 
.A(n_506),
.B(n_234),
.C(n_231),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_481),
.A2(n_506),
.B1(n_519),
.B2(n_508),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_456),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_506),
.Y(n_625)
);

OR2x6_ASAP7_75t_L g626 ( 
.A(n_523),
.B(n_343),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_503),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_456),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_503),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_473),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_524),
.B(n_438),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_456),
.Y(n_632)
);

OR2x6_ASAP7_75t_L g633 ( 
.A(n_506),
.B(n_343),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_508),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_473),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_461),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_455),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_506),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_510),
.Y(n_639)
);

AND2x2_ASAP7_75t_SL g640 ( 
.A(n_481),
.B(n_271),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_519),
.B(n_213),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_461),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_461),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_510),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_511),
.Y(n_645)
);

BUFx10_ASAP7_75t_L g646 ( 
.A(n_519),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_511),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_461),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_515),
.Y(n_649)
);

HB1xp67_ASAP7_75t_L g650 ( 
.A(n_524),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_515),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_477),
.Y(n_652)
);

INVxp67_ASAP7_75t_L g653 ( 
.A(n_519),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_486),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_486),
.Y(n_655)
);

OR2x6_ASAP7_75t_L g656 ( 
.A(n_519),
.B(n_242),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_486),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_486),
.Y(n_658)
);

NAND2xp33_ASAP7_75t_L g659 ( 
.A(n_448),
.B(n_271),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_486),
.B(n_193),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_522),
.B(n_438),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_516),
.B(n_229),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_484),
.A2(n_289),
.B1(n_292),
.B2(n_293),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_516),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_484),
.Y(n_665)
);

AND2x2_ASAP7_75t_SL g666 ( 
.A(n_484),
.B(n_271),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_516),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_516),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_477),
.Y(n_669)
);

BUFx4f_ASAP7_75t_L g670 ( 
.A(n_480),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_477),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_482),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_482),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_482),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_494),
.B(n_224),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_484),
.A2(n_243),
.B1(n_334),
.B2(n_260),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_522),
.B(n_436),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_563),
.B(n_398),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_526),
.Y(n_679)
);

NAND3xp33_ASAP7_75t_L g680 ( 
.A(n_612),
.B(n_239),
.C(n_238),
.Y(n_680)
);

OAI22xp33_ASAP7_75t_L g681 ( 
.A1(n_574),
.A2(n_420),
.B1(n_413),
.B2(n_273),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_562),
.B(n_480),
.Y(n_682)
);

NAND2xp33_ASAP7_75t_L g683 ( 
.A(n_623),
.B(n_448),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_526),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_533),
.B(n_198),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_566),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_640),
.B(n_480),
.Y(n_687)
);

O2A1O1Ixp33_ASAP7_75t_L g688 ( 
.A1(n_531),
.A2(n_574),
.B(n_662),
.C(n_650),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_640),
.B(n_480),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_582),
.B(n_495),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_596),
.B(n_535),
.Y(n_691)
);

AND2x6_ASAP7_75t_L g692 ( 
.A(n_665),
.B(n_271),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_535),
.B(n_495),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_525),
.B(n_198),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_535),
.B(n_547),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_528),
.Y(n_696)
);

NOR2xp67_ASAP7_75t_L g697 ( 
.A(n_575),
.B(n_484),
.Y(n_697)
);

AND2x6_ASAP7_75t_L g698 ( 
.A(n_665),
.B(n_227),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_528),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_638),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_537),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_547),
.B(n_495),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_638),
.A2(n_448),
.B1(n_518),
.B2(n_509),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_547),
.B(n_495),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_SL g705 ( 
.A(n_541),
.B(n_304),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_537),
.Y(n_706)
);

NAND2xp33_ASAP7_75t_L g707 ( 
.A(n_625),
.B(n_448),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_654),
.Y(n_708)
);

OAI22xp5_ASAP7_75t_L g709 ( 
.A1(n_625),
.A2(n_232),
.B1(n_244),
.B2(n_246),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_543),
.B(n_201),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_594),
.Y(n_711)
);

AND2x6_ASAP7_75t_SL g712 ( 
.A(n_615),
.B(n_276),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_566),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_608),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_592),
.B(n_332),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_594),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_657),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_655),
.B(n_495),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_564),
.B(n_495),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_564),
.B(n_495),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_662),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_564),
.B(n_498),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_540),
.B(n_498),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_570),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_542),
.B(n_201),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_540),
.B(n_570),
.Y(n_726)
);

AND2x2_ASAP7_75t_SL g727 ( 
.A(n_666),
.B(n_250),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_655),
.B(n_602),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_540),
.B(n_498),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_658),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_608),
.B(n_498),
.Y(n_731)
);

A2O1A1Ixp33_ASAP7_75t_L g732 ( 
.A1(n_556),
.A2(n_338),
.B(n_522),
.C(n_268),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_639),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_639),
.B(n_498),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_552),
.B(n_498),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_592),
.B(n_332),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_569),
.B(n_498),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_602),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_573),
.B(n_507),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_655),
.B(n_507),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_576),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_572),
.B(n_208),
.Y(n_742)
);

INVxp67_ASAP7_75t_SL g743 ( 
.A(n_527),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_577),
.B(n_507),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_546),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_589),
.B(n_507),
.Y(n_746)
);

NAND2x1_ASAP7_75t_L g747 ( 
.A(n_557),
.B(n_499),
.Y(n_747)
);

INVxp67_ASAP7_75t_L g748 ( 
.A(n_546),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_661),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_593),
.B(n_507),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_576),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_666),
.B(n_583),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_583),
.B(n_507),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_611),
.B(n_507),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_620),
.B(n_494),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_627),
.B(n_494),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_629),
.B(n_634),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_561),
.B(n_208),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_631),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_529),
.B(n_332),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_606),
.A2(n_653),
.B1(n_548),
.B2(n_560),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_616),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_529),
.B(n_209),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_661),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_677),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_644),
.B(n_505),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_606),
.A2(n_345),
.B1(n_209),
.B2(n_216),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_677),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_555),
.A2(n_255),
.B1(n_256),
.B2(n_258),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_631),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_645),
.B(n_505),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_580),
.A2(n_356),
.B1(n_321),
.B2(n_324),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_617),
.A2(n_356),
.B1(n_321),
.B2(n_324),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_621),
.A2(n_264),
.B1(n_216),
.B2(n_325),
.Y(n_774)
);

INVxp67_ASAP7_75t_SL g775 ( 
.A(n_527),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_550),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_647),
.B(n_505),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_609),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_609),
.B(n_522),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_609),
.A2(n_448),
.B1(n_518),
.B2(n_509),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_649),
.B(n_518),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_652),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_536),
.B(n_264),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_553),
.B(n_353),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_584),
.B(n_586),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_651),
.B(n_509),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_664),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_557),
.B(n_600),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_667),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_557),
.B(n_449),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_534),
.A2(n_448),
.B1(n_262),
.B2(n_294),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_584),
.B(n_191),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_536),
.B(n_325),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_605),
.B(n_453),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_668),
.B(n_453),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_652),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_578),
.B(n_457),
.Y(n_797)
);

NAND2xp33_ASAP7_75t_L g798 ( 
.A(n_532),
.B(n_448),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_656),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_584),
.B(n_191),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_579),
.B(n_457),
.Y(n_801)
);

NOR3xp33_ASAP7_75t_L g802 ( 
.A(n_591),
.B(n_252),
.C(n_248),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_656),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_586),
.B(n_191),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_671),
.Y(n_805)
);

NAND2xp33_ASAP7_75t_L g806 ( 
.A(n_532),
.B(n_191),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_671),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_599),
.B(n_458),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_586),
.B(n_191),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_637),
.A2(n_331),
.B1(n_345),
.B2(n_328),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_619),
.B(n_328),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_656),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_553),
.B(n_614),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_614),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_656),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_633),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_636),
.Y(n_817)
);

OR2x6_ASAP7_75t_L g818 ( 
.A(n_633),
.B(n_300),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_646),
.B(n_191),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_646),
.B(n_191),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_646),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_558),
.B(n_309),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_637),
.B(n_331),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_599),
.B(n_624),
.Y(n_824)
);

NOR3xp33_ASAP7_75t_L g825 ( 
.A(n_554),
.B(n_241),
.C(n_257),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_636),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_642),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_642),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_643),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_553),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_553),
.B(n_341),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_633),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_624),
.B(n_459),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_527),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_672),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_558),
.B(n_310),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_643),
.Y(n_837)
);

OAI22xp5_ASAP7_75t_L g838 ( 
.A1(n_622),
.A2(n_330),
.B1(n_348),
.B2(n_355),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_648),
.Y(n_839)
);

AND2x4_ASAP7_75t_L g840 ( 
.A(n_633),
.B(n_437),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_558),
.B(n_341),
.Y(n_841)
);

INVxp67_ASAP7_75t_L g842 ( 
.A(n_534),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_648),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_530),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_565),
.B(n_342),
.Y(n_845)
);

BUFx8_ASAP7_75t_L g846 ( 
.A(n_550),
.Y(n_846)
);

O2A1O1Ixp5_ASAP7_75t_L g847 ( 
.A1(n_660),
.A2(n_468),
.B(n_488),
.C(n_478),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_L g848 ( 
.A1(n_691),
.A2(n_549),
.B1(n_618),
.B2(n_641),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_762),
.B(n_595),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_685),
.B(n_725),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_742),
.B(n_613),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_758),
.B(n_613),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_779),
.Y(n_853)
);

INVx1_ASAP7_75t_SL g854 ( 
.A(n_745),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_694),
.B(n_613),
.Y(n_855)
);

INVxp67_ASAP7_75t_L g856 ( 
.A(n_811),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_695),
.A2(n_549),
.B(n_610),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_710),
.B(n_613),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_788),
.A2(n_549),
.B(n_610),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_693),
.A2(n_549),
.B(n_610),
.Y(n_860)
);

NOR2x1_ASAP7_75t_L g861 ( 
.A(n_680),
.B(n_544),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_702),
.A2(n_670),
.B(n_587),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_721),
.B(n_565),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_716),
.B(n_558),
.Y(n_864)
);

NOR3xp33_ASAP7_75t_L g865 ( 
.A(n_681),
.B(n_601),
.C(n_581),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_704),
.A2(n_670),
.B(n_587),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_686),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_686),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_719),
.A2(n_670),
.B(n_587),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_779),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_716),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_720),
.A2(n_551),
.B(n_538),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_713),
.Y(n_873)
);

INVx4_ASAP7_75t_L g874 ( 
.A(n_716),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_721),
.B(n_565),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_722),
.A2(n_551),
.B(n_538),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_748),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_713),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_714),
.Y(n_879)
);

NAND2xp33_ASAP7_75t_L g880 ( 
.A(n_716),
.B(n_532),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_690),
.A2(n_551),
.B(n_538),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_683),
.A2(n_538),
.B(n_527),
.Y(n_882)
);

A2O1A1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_688),
.A2(n_676),
.B(n_663),
.C(n_675),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_714),
.Y(n_884)
);

A2O1A1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_732),
.A2(n_336),
.B(n_194),
.C(n_205),
.Y(n_885)
);

NOR2x1_ASAP7_75t_L g886 ( 
.A(n_752),
.B(n_565),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_733),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_760),
.B(n_626),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_701),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_733),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_683),
.A2(n_545),
.B(n_628),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_723),
.A2(n_729),
.B(n_790),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_682),
.A2(n_689),
.B(n_687),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_715),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_724),
.B(n_626),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_687),
.A2(n_545),
.B(n_628),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_724),
.B(n_626),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_727),
.A2(n_568),
.B1(n_626),
.B2(n_567),
.Y(n_898)
);

NAND2x1p5_ASAP7_75t_L g899 ( 
.A(n_821),
.B(n_558),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_749),
.B(n_669),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_749),
.B(n_672),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_727),
.A2(n_568),
.B1(n_567),
.B2(n_532),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_700),
.Y(n_903)
);

O2A1O1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_732),
.A2(n_659),
.B(n_590),
.C(n_607),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_761),
.B(n_632),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_764),
.B(n_673),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_689),
.A2(n_775),
.B(n_743),
.Y(n_907)
);

O2A1O1Ixp5_ASAP7_75t_L g908 ( 
.A1(n_682),
.A2(n_632),
.B(n_674),
.C(n_673),
.Y(n_908)
);

O2A1O1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_752),
.A2(n_659),
.B(n_590),
.C(n_607),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_701),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_718),
.A2(n_538),
.B(n_545),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_740),
.A2(n_545),
.B(n_527),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_740),
.A2(n_628),
.B(n_632),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_824),
.A2(n_628),
.B(n_630),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_814),
.B(n_571),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_708),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_701),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_706),
.B(n_711),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_726),
.A2(n_635),
.B(n_630),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_736),
.Y(n_920)
);

NAND2xp33_ASAP7_75t_L g921 ( 
.A(n_698),
.B(n_532),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_814),
.B(n_349),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_764),
.A2(n_568),
.B1(n_348),
.B2(n_342),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_717),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_678),
.B(n_588),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_728),
.A2(n_559),
.B(n_603),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_765),
.B(n_532),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_765),
.B(n_567),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_706),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_768),
.B(n_567),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_730),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_728),
.A2(n_539),
.B(n_603),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_785),
.A2(n_539),
.B(n_598),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_768),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_813),
.B(n_588),
.Y(n_935)
);

OAI21xp5_ASAP7_75t_L g936 ( 
.A1(n_753),
.A2(n_530),
.B(n_598),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_706),
.Y(n_937)
);

AO21x1_ASAP7_75t_L g938 ( 
.A1(n_819),
.A2(n_488),
.B(n_476),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_797),
.B(n_567),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_782),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_711),
.B(n_559),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_778),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_753),
.A2(n_567),
.B1(n_604),
.B2(n_568),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_842),
.B(n_265),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_782),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_783),
.B(n_353),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_L g947 ( 
.A1(n_711),
.A2(n_355),
.B1(n_597),
.B2(n_585),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_801),
.B(n_604),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_785),
.A2(n_597),
.B(n_585),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_793),
.B(n_679),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_796),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_794),
.B(n_604),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_707),
.A2(n_475),
.B(n_478),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_707),
.A2(n_475),
.B(n_476),
.Y(n_954)
);

AND3x4_ASAP7_75t_L g955 ( 
.A(n_802),
.B(n_353),
.C(n_350),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_763),
.B(n_604),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_792),
.A2(n_474),
.B(n_468),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_796),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_L g959 ( 
.A1(n_731),
.A2(n_604),
.B(n_499),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_684),
.B(n_437),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_738),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_792),
.A2(n_474),
.B(n_467),
.Y(n_962)
);

BUFx3_ASAP7_75t_L g963 ( 
.A(n_816),
.Y(n_963)
);

NAND2xp33_ASAP7_75t_L g964 ( 
.A(n_698),
.B(n_604),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_800),
.A2(n_467),
.B(n_499),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_696),
.B(n_699),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_821),
.B(n_467),
.Y(n_967)
);

OR2x6_ASAP7_75t_L g968 ( 
.A(n_832),
.B(n_467),
.Y(n_968)
);

INVx5_ASAP7_75t_L g969 ( 
.A(n_698),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_832),
.A2(n_301),
.B1(n_267),
.B2(n_272),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_821),
.B(n_274),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_834),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_741),
.A2(n_350),
.B(n_346),
.C(n_339),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_697),
.B(n_275),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_816),
.B(n_87),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_759),
.B(n_499),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_805),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_770),
.B(n_192),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_757),
.B(n_499),
.Y(n_979)
);

NOR3xp33_ASAP7_75t_L g980 ( 
.A(n_831),
.B(n_288),
.C(n_286),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_L g981 ( 
.A1(n_751),
.A2(n_194),
.B1(n_346),
.B2(n_339),
.Y(n_981)
);

O2A1O1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_769),
.A2(n_211),
.B(n_206),
.C(n_205),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_823),
.B(n_499),
.Y(n_983)
);

NAND2x1p5_ASAP7_75t_L g984 ( 
.A(n_747),
.B(n_91),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_800),
.A2(n_499),
.B(n_313),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_773),
.B(n_282),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_804),
.A2(n_809),
.B(n_819),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_787),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_709),
.A2(n_206),
.B(n_211),
.C(n_336),
.Y(n_989)
);

BUFx4f_ASAP7_75t_L g990 ( 
.A(n_818),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_774),
.B(n_285),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_789),
.B(n_499),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_804),
.A2(n_318),
.B(n_296),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_840),
.B(n_291),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_809),
.A2(n_297),
.B(n_302),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_820),
.A2(n_312),
.B(n_314),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_840),
.B(n_337),
.Y(n_997)
);

INVx4_ASAP7_75t_L g998 ( 
.A(n_834),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_805),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_840),
.B(n_337),
.Y(n_1000)
);

NOR2xp67_ASAP7_75t_SL g1001 ( 
.A(n_834),
.B(n_335),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_820),
.A2(n_335),
.B(n_329),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_735),
.A2(n_329),
.B(n_326),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_807),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_755),
.B(n_326),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_780),
.B(n_323),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_703),
.A2(n_323),
.B1(n_322),
.B2(n_169),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_807),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_799),
.B(n_157),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_835),
.Y(n_1010)
);

NOR3xp33_ASAP7_75t_L g1011 ( 
.A(n_825),
.B(n_322),
.C(n_13),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_835),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_756),
.B(n_6),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_766),
.B(n_13),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_737),
.A2(n_154),
.B(n_153),
.Y(n_1015)
);

INVx5_ASAP7_75t_L g1016 ( 
.A(n_698),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_739),
.A2(n_145),
.B(n_140),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_744),
.A2(n_132),
.B(n_130),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_771),
.B(n_15),
.Y(n_1019)
);

O2A1O1Ixp5_ASAP7_75t_L g1020 ( 
.A1(n_847),
.A2(n_128),
.B(n_124),
.C(n_121),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_844),
.Y(n_1021)
);

AOI221x1_ASAP7_75t_L g1022 ( 
.A1(n_734),
.A2(n_120),
.B1(n_110),
.B2(n_108),
.C(n_103),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_803),
.B(n_95),
.Y(n_1023)
);

INVxp67_ASAP7_75t_L g1024 ( 
.A(n_784),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_845),
.B(n_66),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_817),
.Y(n_1026)
);

O2A1O1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_838),
.A2(n_15),
.B(n_17),
.C(n_18),
.Y(n_1027)
);

OR2x6_ASAP7_75t_L g1028 ( 
.A(n_818),
.B(n_20),
.Y(n_1028)
);

NAND3xp33_ASAP7_75t_L g1029 ( 
.A(n_772),
.B(n_21),
.C(n_23),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_SL g1030 ( 
.A1(n_746),
.A2(n_66),
.B(n_27),
.C(n_28),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_750),
.A2(n_26),
.B(n_27),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_826),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_754),
.B(n_28),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_830),
.B(n_29),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_777),
.B(n_31),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_827),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_828),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_781),
.B(n_32),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_786),
.B(n_33),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_850),
.B(n_705),
.Y(n_1040)
);

AOI221xp5_ASAP7_75t_L g1041 ( 
.A1(n_981),
.A2(n_767),
.B1(n_810),
.B2(n_815),
.C(n_812),
.Y(n_1041)
);

HB1xp67_ASAP7_75t_L g1042 ( 
.A(n_854),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_892),
.A2(n_798),
.B(n_806),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_877),
.Y(n_1044)
);

O2A1O1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_856),
.A2(n_795),
.B(n_818),
.C(n_841),
.Y(n_1045)
);

NOR2x1_ASAP7_75t_L g1046 ( 
.A(n_874),
.B(n_818),
.Y(n_1046)
);

AOI22xp33_ASAP7_75t_L g1047 ( 
.A1(n_1011),
.A2(n_698),
.B1(n_806),
.B2(n_791),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_851),
.A2(n_808),
.B1(n_833),
.B2(n_839),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_859),
.A2(n_798),
.B(n_841),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_915),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_871),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_950),
.B(n_843),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_871),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_894),
.B(n_712),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_946),
.B(n_888),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_987),
.A2(n_836),
.B(n_822),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_881),
.A2(n_836),
.B(n_822),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_853),
.B(n_698),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_986),
.A2(n_837),
.B(n_829),
.C(n_39),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_871),
.Y(n_1060)
);

AOI21x1_ASAP7_75t_L g1061 ( 
.A1(n_905),
.A2(n_692),
.B(n_34),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_857),
.A2(n_692),
.B(n_776),
.Y(n_1062)
);

CKINVDCx20_ASAP7_75t_R g1063 ( 
.A(n_963),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_L g1064 ( 
.A1(n_872),
.A2(n_692),
.B(n_45),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_986),
.A2(n_33),
.B(n_46),
.C(n_47),
.Y(n_1065)
);

AOI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_980),
.A2(n_692),
.B1(n_776),
.B2(n_846),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_918),
.A2(n_692),
.B(n_48),
.Y(n_1067)
);

AOI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_980),
.A2(n_692),
.B1(n_846),
.B2(n_50),
.Y(n_1068)
);

BUFx10_ASAP7_75t_L g1069 ( 
.A(n_935),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_871),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_910),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_918),
.A2(n_46),
.B(n_49),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_920),
.B(n_846),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_991),
.A2(n_50),
.B(n_51),
.C(n_55),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_867),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_852),
.B(n_51),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_910),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_855),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_1078)
);

AOI21x1_ASAP7_75t_L g1079 ( 
.A1(n_905),
.A2(n_967),
.B(n_956),
.Y(n_1079)
);

NAND3xp33_ASAP7_75t_SL g1080 ( 
.A(n_1011),
.B(n_57),
.C(n_60),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_870),
.B(n_60),
.Y(n_1081)
);

OAI22x1_ASAP7_75t_L g1082 ( 
.A1(n_955),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_915),
.B(n_61),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_858),
.B(n_63),
.Y(n_1084)
);

AOI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_849),
.A2(n_65),
.B1(n_991),
.B2(n_865),
.Y(n_1085)
);

NOR2xp67_ASAP7_75t_SL g1086 ( 
.A(n_969),
.B(n_1016),
.Y(n_1086)
);

HB1xp67_ASAP7_75t_L g1087 ( 
.A(n_903),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_910),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_907),
.A2(n_860),
.B(n_882),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_867),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_903),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_849),
.B(n_922),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_893),
.A2(n_891),
.B(n_908),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_878),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_934),
.B(n_916),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_874),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_910),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_924),
.B(n_931),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_963),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_848),
.A2(n_876),
.B(n_866),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_922),
.B(n_944),
.Y(n_1101)
);

O2A1O1Ixp33_ASAP7_75t_SL g1102 ( 
.A1(n_883),
.A2(n_1038),
.B(n_1033),
.C(n_885),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_944),
.B(n_1024),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_889),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_966),
.B(n_1005),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_902),
.A2(n_898),
.B1(n_886),
.B2(n_937),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_942),
.B(n_988),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1025),
.B(n_884),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_975),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_884),
.Y(n_1110)
);

OR2x2_ASAP7_75t_L g1111 ( 
.A(n_997),
.B(n_1000),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_887),
.B(n_895),
.Y(n_1112)
);

O2A1O1Ixp5_ASAP7_75t_L g1113 ( 
.A1(n_938),
.A2(n_1033),
.B(n_1020),
.C(n_1038),
.Y(n_1113)
);

HB1xp67_ASAP7_75t_L g1114 ( 
.A(n_889),
.Y(n_1114)
);

AO32x1_ASAP7_75t_L g1115 ( 
.A1(n_923),
.A2(n_947),
.A3(n_873),
.B1(n_879),
.B2(n_890),
.Y(n_1115)
);

OAI22x1_ASAP7_75t_L g1116 ( 
.A1(n_955),
.A2(n_925),
.B1(n_1034),
.B2(n_935),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_1027),
.A2(n_885),
.B(n_973),
.C(n_982),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_862),
.A2(n_869),
.B(n_1016),
.Y(n_1118)
);

O2A1O1Ixp5_ASAP7_75t_L g1119 ( 
.A1(n_1001),
.A2(n_971),
.B(n_974),
.C(n_1039),
.Y(n_1119)
);

NOR3xp33_ASAP7_75t_SL g1120 ( 
.A(n_973),
.B(n_1029),
.C(n_989),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_897),
.A2(n_883),
.B(n_909),
.C(n_939),
.Y(n_1121)
);

HB1xp67_ASAP7_75t_L g1122 ( 
.A(n_917),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_969),
.A2(n_1016),
.B(n_964),
.Y(n_1123)
);

NOR2x1_ASAP7_75t_R g1124 ( 
.A(n_975),
.B(n_1009),
.Y(n_1124)
);

OAI21xp33_ASAP7_75t_SL g1125 ( 
.A1(n_902),
.A2(n_898),
.B(n_943),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_887),
.B(n_960),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_1009),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_961),
.B(n_868),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_969),
.A2(n_921),
.B(n_896),
.Y(n_1129)
);

AO22x1_ASAP7_75t_L g1130 ( 
.A1(n_865),
.A2(n_925),
.B1(n_1023),
.B2(n_861),
.Y(n_1130)
);

O2A1O1Ixp5_ASAP7_75t_L g1131 ( 
.A1(n_971),
.A2(n_974),
.B(n_1035),
.C(n_1019),
.Y(n_1131)
);

CKINVDCx16_ASAP7_75t_R g1132 ( 
.A(n_1028),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_880),
.A2(n_928),
.B(n_930),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_978),
.B(n_900),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_917),
.Y(n_1135)
);

O2A1O1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_1013),
.A2(n_1014),
.B(n_994),
.C(n_1030),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_929),
.B(n_937),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_863),
.B(n_875),
.Y(n_1138)
);

A2O1A1Ixp33_ASAP7_75t_SL g1139 ( 
.A1(n_983),
.A2(n_959),
.B(n_929),
.C(n_904),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_R g1140 ( 
.A(n_990),
.B(n_972),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_981),
.B(n_1023),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1021),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_927),
.A2(n_901),
.B(n_906),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1021),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_990),
.B(n_995),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1008),
.Y(n_1146)
);

NOR2x1p5_ASAP7_75t_SL g1147 ( 
.A(n_945),
.B(n_1004),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1008),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_1028),
.Y(n_1149)
);

BUFx8_ASAP7_75t_SL g1150 ( 
.A(n_1028),
.Y(n_1150)
);

AOI21x1_ASAP7_75t_L g1151 ( 
.A1(n_967),
.A2(n_933),
.B(n_949),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_972),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_970),
.B(n_1003),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_993),
.B(n_996),
.Y(n_1154)
);

OR2x6_ASAP7_75t_L g1155 ( 
.A(n_984),
.B(n_968),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_1032),
.B(n_1037),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_945),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1036),
.B(n_1026),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_958),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_958),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1026),
.B(n_1006),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1004),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_1030),
.A2(n_1007),
.B(n_1002),
.C(n_1006),
.Y(n_1163)
);

CKINVDCx11_ASAP7_75t_R g1164 ( 
.A(n_968),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_948),
.A2(n_941),
.B(n_952),
.Y(n_1165)
);

AND2x6_ASAP7_75t_SL g1166 ( 
.A(n_968),
.B(n_976),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_940),
.B(n_977),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_998),
.A2(n_1010),
.B1(n_1012),
.B2(n_899),
.Y(n_1168)
);

O2A1O1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1031),
.A2(n_979),
.B(n_941),
.C(n_951),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_999),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_998),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_864),
.B(n_992),
.Y(n_1172)
);

BUFx3_ASAP7_75t_L g1173 ( 
.A(n_984),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_919),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_864),
.B(n_954),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_953),
.A2(n_957),
.B(n_936),
.C(n_985),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_1015),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_899),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_1017),
.Y(n_1179)
);

INVx4_ASAP7_75t_L g1180 ( 
.A(n_913),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_911),
.B(n_912),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_926),
.B(n_932),
.Y(n_1182)
);

O2A1O1Ixp5_ASAP7_75t_L g1183 ( 
.A1(n_914),
.A2(n_962),
.B(n_1018),
.C(n_965),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1022),
.B(n_950),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_867),
.Y(n_1185)
);

AOI221xp5_ASAP7_75t_L g1186 ( 
.A1(n_981),
.A2(n_991),
.B1(n_986),
.B2(n_568),
.C(n_825),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_850),
.B(n_762),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_850),
.B(n_856),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_950),
.B(n_721),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_850),
.B(n_950),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_871),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_871),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_850),
.A2(n_691),
.B1(n_685),
.B2(n_851),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_892),
.A2(n_549),
.B(n_547),
.Y(n_1194)
);

OAI21xp33_ASAP7_75t_L g1195 ( 
.A1(n_850),
.A2(n_685),
.B(n_986),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_892),
.A2(n_549),
.B(n_547),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_850),
.A2(n_685),
.B1(n_742),
.B2(n_725),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_850),
.B(n_762),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_892),
.A2(n_549),
.B(n_547),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_963),
.B(n_853),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_SL g1201 ( 
.A1(n_1195),
.A2(n_1124),
.B(n_1121),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1092),
.B(n_1189),
.Y(n_1202)
);

OAI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1197),
.A2(n_1113),
.B(n_1165),
.Y(n_1203)
);

OAI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1113),
.A2(n_1175),
.B(n_1143),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1152),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1186),
.A2(n_1190),
.B1(n_1085),
.B2(n_1101),
.Y(n_1206)
);

CKINVDCx9p33_ASAP7_75t_R g1207 ( 
.A(n_1044),
.Y(n_1207)
);

AO31x2_ASAP7_75t_L g1208 ( 
.A1(n_1100),
.A2(n_1175),
.A3(n_1193),
.B(n_1089),
.Y(n_1208)
);

O2A1O1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1101),
.A2(n_1092),
.B(n_1198),
.C(n_1187),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1194),
.A2(n_1199),
.B(n_1196),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1129),
.A2(n_1118),
.B(n_1176),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1075),
.Y(n_1212)
);

AO31x2_ASAP7_75t_L g1213 ( 
.A1(n_1048),
.A2(n_1174),
.A3(n_1106),
.B(n_1180),
.Y(n_1213)
);

AOI31xp67_ASAP7_75t_L g1214 ( 
.A1(n_1181),
.A2(n_1154),
.A3(n_1182),
.B(n_1145),
.Y(n_1214)
);

AO31x2_ASAP7_75t_L g1215 ( 
.A1(n_1180),
.A2(n_1049),
.A3(n_1172),
.B(n_1168),
.Y(n_1215)
);

AO21x2_ASAP7_75t_L g1216 ( 
.A1(n_1093),
.A2(n_1184),
.B(n_1136),
.Y(n_1216)
);

OR2x2_ASAP7_75t_L g1217 ( 
.A(n_1105),
.B(n_1042),
.Y(n_1217)
);

O2A1O1Ixp5_ASAP7_75t_SL g1218 ( 
.A1(n_1078),
.A2(n_1076),
.B(n_1084),
.C(n_1040),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1090),
.Y(n_1219)
);

AOI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1187),
.A2(n_1198),
.B1(n_1083),
.B2(n_1103),
.Y(n_1220)
);

AO22x2_ASAP7_75t_L g1221 ( 
.A1(n_1080),
.A2(n_1141),
.B1(n_1072),
.B2(n_1149),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1134),
.B(n_1188),
.Y(n_1222)
);

AO32x2_ASAP7_75t_L g1223 ( 
.A1(n_1115),
.A2(n_1102),
.A3(n_1117),
.B1(n_1120),
.B2(n_1125),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1133),
.A2(n_1079),
.B(n_1183),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1183),
.A2(n_1123),
.B(n_1043),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1139),
.A2(n_1177),
.B(n_1056),
.Y(n_1226)
);

AO31x2_ASAP7_75t_L g1227 ( 
.A1(n_1172),
.A2(n_1057),
.A3(n_1161),
.B(n_1115),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1050),
.B(n_1103),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_SL g1229 ( 
.A1(n_1061),
.A2(n_1062),
.B(n_1163),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1131),
.A2(n_1179),
.B(n_1108),
.Y(n_1230)
);

AOI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1130),
.A2(n_1112),
.B(n_1153),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1131),
.A2(n_1169),
.B(n_1119),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1119),
.A2(n_1126),
.B(n_1045),
.Y(n_1233)
);

AOI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1058),
.A2(n_1064),
.B(n_1158),
.Y(n_1234)
);

NAND2xp33_ASAP7_75t_L g1235 ( 
.A(n_1109),
.B(n_1127),
.Y(n_1235)
);

NAND3x1_ASAP7_75t_L g1236 ( 
.A(n_1083),
.B(n_1054),
.C(n_1066),
.Y(n_1236)
);

A2O1A1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1120),
.A2(n_1059),
.B(n_1111),
.C(n_1138),
.Y(n_1237)
);

INVx5_ASAP7_75t_L g1238 ( 
.A(n_1051),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1138),
.A2(n_1055),
.B(n_1047),
.C(n_1065),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1110),
.Y(n_1240)
);

A2O1A1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1047),
.A2(n_1074),
.B(n_1156),
.C(n_1041),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1155),
.A2(n_1086),
.B(n_1137),
.Y(n_1242)
);

NAND3xp33_ASAP7_75t_L g1243 ( 
.A(n_1068),
.B(n_1054),
.C(n_1156),
.Y(n_1243)
);

NAND2x1p5_ASAP7_75t_L g1244 ( 
.A(n_1096),
.B(n_1099),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1087),
.B(n_1091),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1094),
.A2(n_1162),
.B(n_1160),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1095),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1098),
.B(n_1109),
.Y(n_1248)
);

HB1xp67_ASAP7_75t_L g1249 ( 
.A(n_1087),
.Y(n_1249)
);

A2O1A1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1081),
.A2(n_1173),
.B(n_1067),
.C(n_1147),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1091),
.B(n_1052),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1142),
.B(n_1144),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1200),
.B(n_1109),
.Y(n_1253)
);

AO31x2_ASAP7_75t_L g1254 ( 
.A1(n_1115),
.A2(n_1116),
.A3(n_1185),
.B(n_1157),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1155),
.A2(n_1128),
.B(n_1178),
.Y(n_1255)
);

A2O1A1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1127),
.A2(n_1109),
.B(n_1046),
.C(n_1080),
.Y(n_1256)
);

O2A1O1Ixp33_ASAP7_75t_SL g1257 ( 
.A1(n_1114),
.A2(n_1122),
.B(n_1170),
.C(n_1159),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1200),
.B(n_1127),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1167),
.A2(n_1122),
.B(n_1114),
.Y(n_1259)
);

O2A1O1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1073),
.A2(n_1155),
.B(n_1146),
.C(n_1148),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1127),
.B(n_1135),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1132),
.B(n_1063),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1171),
.A2(n_1135),
.B(n_1104),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1104),
.B(n_1140),
.Y(n_1264)
);

INVx2_ASAP7_75t_SL g1265 ( 
.A(n_1069),
.Y(n_1265)
);

AO31x2_ASAP7_75t_L g1266 ( 
.A1(n_1082),
.A2(n_1096),
.A3(n_1166),
.B(n_1152),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1088),
.A2(n_1097),
.B(n_1140),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1051),
.Y(n_1268)
);

AO31x2_ASAP7_75t_L g1269 ( 
.A1(n_1152),
.A2(n_1077),
.A3(n_1071),
.B(n_1088),
.Y(n_1269)
);

INVxp67_ASAP7_75t_L g1270 ( 
.A(n_1150),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1051),
.Y(n_1271)
);

O2A1O1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1097),
.A2(n_1069),
.B(n_1164),
.C(n_1152),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_SL g1273 ( 
.A1(n_1071),
.A2(n_1077),
.B(n_1053),
.Y(n_1273)
);

O2A1O1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_1071),
.A2(n_1077),
.B(n_1053),
.C(n_1060),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1071),
.B(n_1077),
.Y(n_1275)
);

NOR2xp67_ASAP7_75t_L g1276 ( 
.A(n_1053),
.B(n_1060),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1060),
.B(n_1070),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1070),
.A2(n_1191),
.B(n_1192),
.Y(n_1278)
);

OAI22x1_ASAP7_75t_L g1279 ( 
.A1(n_1070),
.A2(n_1191),
.B1(n_1192),
.B2(n_1085),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1191),
.B(n_1192),
.Y(n_1280)
);

INVx1_ASAP7_75t_SL g1281 ( 
.A(n_1191),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1194),
.A2(n_549),
.B(n_691),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1118),
.A2(n_1089),
.B(n_1151),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1118),
.A2(n_1089),
.B(n_1151),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1195),
.B(n_762),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1121),
.A2(n_1197),
.B(n_850),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1197),
.A2(n_850),
.B1(n_1195),
.B2(n_1186),
.Y(n_1287)
);

O2A1O1Ixp5_ASAP7_75t_SL g1288 ( 
.A1(n_1181),
.A2(n_1193),
.B(n_682),
.C(n_1078),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1194),
.A2(n_549),
.B(n_691),
.Y(n_1289)
);

NAND2x1p5_ASAP7_75t_L g1290 ( 
.A(n_1096),
.B(n_1086),
.Y(n_1290)
);

AOI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1195),
.A2(n_1092),
.B1(n_1101),
.B2(n_1186),
.Y(n_1291)
);

AO32x2_ASAP7_75t_L g1292 ( 
.A1(n_1078),
.A2(n_1193),
.A3(n_1106),
.B1(n_923),
.B2(n_769),
.Y(n_1292)
);

AOI31xp67_ASAP7_75t_L g1293 ( 
.A1(n_1181),
.A2(n_682),
.A3(n_905),
.B(n_1154),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1118),
.A2(n_1089),
.B(n_1151),
.Y(n_1294)
);

CKINVDCx11_ASAP7_75t_R g1295 ( 
.A(n_1063),
.Y(n_1295)
);

A2O1A1Ixp33_ASAP7_75t_L g1296 ( 
.A1(n_1195),
.A2(n_1197),
.B(n_1101),
.C(n_850),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1063),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1195),
.B(n_762),
.Y(n_1298)
);

A2O1A1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1195),
.A2(n_1197),
.B(n_1101),
.C(n_850),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1107),
.Y(n_1300)
);

AOI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1195),
.A2(n_1092),
.B1(n_1101),
.B2(n_1186),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_SL g1302 ( 
.A1(n_1101),
.A2(n_705),
.B1(n_541),
.B2(n_1092),
.Y(n_1302)
);

NOR2xp67_ASAP7_75t_L g1303 ( 
.A(n_1111),
.B(n_761),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1190),
.B(n_571),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1092),
.B(n_1189),
.Y(n_1305)
);

A2O1A1Ixp33_ASAP7_75t_L g1306 ( 
.A1(n_1195),
.A2(n_1197),
.B(n_1101),
.C(n_850),
.Y(n_1306)
);

AOI221x1_ASAP7_75t_L g1307 ( 
.A1(n_1195),
.A2(n_850),
.B1(n_1101),
.B2(n_1092),
.C(n_1193),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1075),
.Y(n_1308)
);

O2A1O1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1195),
.A2(n_1101),
.B(n_850),
.C(n_762),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1121),
.A2(n_1197),
.B(n_850),
.Y(n_1310)
);

O2A1O1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1195),
.A2(n_1101),
.B(n_850),
.C(n_762),
.Y(n_1311)
);

AOI31xp67_ASAP7_75t_L g1312 ( 
.A1(n_1181),
.A2(n_682),
.A3(n_905),
.B(n_1154),
.Y(n_1312)
);

AO31x2_ASAP7_75t_L g1313 ( 
.A1(n_1121),
.A2(n_1100),
.A3(n_1175),
.B(n_1193),
.Y(n_1313)
);

BUFx6f_ASAP7_75t_L g1314 ( 
.A(n_1051),
.Y(n_1314)
);

O2A1O1Ixp5_ASAP7_75t_L g1315 ( 
.A1(n_1101),
.A2(n_850),
.B(n_685),
.C(n_742),
.Y(n_1315)
);

NAND2x1p5_ASAP7_75t_L g1316 ( 
.A(n_1096),
.B(n_1086),
.Y(n_1316)
);

AO21x2_ASAP7_75t_L g1317 ( 
.A1(n_1100),
.A2(n_1089),
.B(n_1093),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1063),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1075),
.Y(n_1319)
);

BUFx2_ASAP7_75t_L g1320 ( 
.A(n_1044),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1118),
.A2(n_1089),
.B(n_1151),
.Y(n_1321)
);

NOR2xp67_ASAP7_75t_L g1322 ( 
.A(n_1111),
.B(n_761),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1107),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1118),
.A2(n_1089),
.B(n_1151),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1190),
.B(n_1198),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1118),
.A2(n_1089),
.B(n_1151),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1194),
.A2(n_549),
.B(n_691),
.Y(n_1327)
);

AO22x2_ASAP7_75t_L g1328 ( 
.A1(n_1080),
.A2(n_955),
.B1(n_1184),
.B2(n_1078),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1194),
.A2(n_549),
.B(n_691),
.Y(n_1329)
);

INVx5_ASAP7_75t_L g1330 ( 
.A(n_1051),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1107),
.Y(n_1331)
);

AO31x2_ASAP7_75t_L g1332 ( 
.A1(n_1121),
.A2(n_1100),
.A3(n_1175),
.B(n_1193),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1121),
.A2(n_1197),
.B(n_850),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1195),
.A2(n_1186),
.B1(n_1101),
.B2(n_1092),
.Y(n_1334)
);

OAI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1121),
.A2(n_1197),
.B(n_850),
.Y(n_1335)
);

INVx3_ASAP7_75t_L g1336 ( 
.A(n_1152),
.Y(n_1336)
);

INVxp67_ASAP7_75t_L g1337 ( 
.A(n_1042),
.Y(n_1337)
);

INVx3_ASAP7_75t_L g1338 ( 
.A(n_1152),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_L g1339 ( 
.A(n_1051),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1194),
.A2(n_549),
.B(n_691),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1092),
.B(n_1189),
.Y(n_1341)
);

AO31x2_ASAP7_75t_L g1342 ( 
.A1(n_1121),
.A2(n_1100),
.A3(n_1175),
.B(n_1193),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1107),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_1195),
.B(n_1050),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1118),
.A2(n_1089),
.B(n_1151),
.Y(n_1345)
);

AND2x6_ASAP7_75t_L g1346 ( 
.A(n_1109),
.B(n_1127),
.Y(n_1346)
);

AO31x2_ASAP7_75t_L g1347 ( 
.A1(n_1121),
.A2(n_1100),
.A3(n_1175),
.B(n_1193),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1107),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1118),
.A2(n_1089),
.B(n_1151),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1190),
.B(n_1198),
.Y(n_1350)
);

O2A1O1Ixp33_ASAP7_75t_SL g1351 ( 
.A1(n_1197),
.A2(n_850),
.B(n_1195),
.C(n_1186),
.Y(n_1351)
);

AOI221x1_ASAP7_75t_L g1352 ( 
.A1(n_1195),
.A2(n_850),
.B1(n_1101),
.B2(n_1092),
.C(n_1193),
.Y(n_1352)
);

AO21x2_ASAP7_75t_L g1353 ( 
.A1(n_1100),
.A2(n_1089),
.B(n_1093),
.Y(n_1353)
);

NAND3xp33_ASAP7_75t_L g1354 ( 
.A(n_1197),
.B(n_850),
.C(n_1195),
.Y(n_1354)
);

OR2x6_ASAP7_75t_L g1355 ( 
.A(n_1109),
.B(n_1127),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1118),
.A2(n_1089),
.B(n_1151),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1118),
.A2(n_1089),
.B(n_1151),
.Y(n_1357)
);

OR2x6_ASAP7_75t_L g1358 ( 
.A(n_1109),
.B(n_1127),
.Y(n_1358)
);

BUFx12f_ASAP7_75t_L g1359 ( 
.A(n_1295),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1212),
.Y(n_1360)
);

INVx6_ASAP7_75t_L g1361 ( 
.A(n_1238),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1219),
.Y(n_1362)
);

BUFx12f_ASAP7_75t_L g1363 ( 
.A(n_1320),
.Y(n_1363)
);

INVx4_ASAP7_75t_L g1364 ( 
.A(n_1238),
.Y(n_1364)
);

CKINVDCx6p67_ASAP7_75t_R g1365 ( 
.A(n_1207),
.Y(n_1365)
);

INVx4_ASAP7_75t_L g1366 ( 
.A(n_1238),
.Y(n_1366)
);

OAI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1220),
.A2(n_1301),
.B1(n_1291),
.B2(n_1287),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1259),
.Y(n_1368)
);

INVx4_ASAP7_75t_L g1369 ( 
.A(n_1330),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1206),
.A2(n_1334),
.B1(n_1287),
.B2(n_1301),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1325),
.B(n_1350),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1240),
.Y(n_1372)
);

CKINVDCx20_ASAP7_75t_R g1373 ( 
.A(n_1297),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_SL g1374 ( 
.A1(n_1206),
.A2(n_1243),
.B1(n_1285),
.B2(n_1298),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1308),
.Y(n_1375)
);

CKINVDCx11_ASAP7_75t_R g1376 ( 
.A(n_1318),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1291),
.A2(n_1354),
.B1(n_1335),
.B2(n_1333),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1265),
.Y(n_1378)
);

OAI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1354),
.A2(n_1243),
.B1(n_1307),
.B2(n_1352),
.Y(n_1379)
);

CKINVDCx20_ASAP7_75t_R g1380 ( 
.A(n_1262),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1319),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1246),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1286),
.A2(n_1335),
.B1(n_1310),
.B2(n_1333),
.Y(n_1383)
);

BUFx12f_ASAP7_75t_L g1384 ( 
.A(n_1217),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1302),
.A2(n_1296),
.B1(n_1299),
.B2(n_1306),
.Y(n_1385)
);

INVx4_ASAP7_75t_L g1386 ( 
.A(n_1330),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1209),
.A2(n_1241),
.B1(n_1228),
.B2(n_1310),
.Y(n_1387)
);

CKINVDCx11_ASAP7_75t_R g1388 ( 
.A(n_1355),
.Y(n_1388)
);

INVx5_ASAP7_75t_L g1389 ( 
.A(n_1346),
.Y(n_1389)
);

INVx1_ASAP7_75t_SL g1390 ( 
.A(n_1304),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1286),
.A2(n_1328),
.B1(n_1202),
.B2(n_1341),
.Y(n_1391)
);

BUFx5_ASAP7_75t_L g1392 ( 
.A(n_1346),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1305),
.B(n_1245),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1252),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1252),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1236),
.A2(n_1237),
.B1(n_1344),
.B2(n_1323),
.Y(n_1396)
);

BUFx12f_ASAP7_75t_L g1397 ( 
.A(n_1244),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1328),
.A2(n_1303),
.B1(n_1322),
.B2(n_1222),
.Y(n_1398)
);

CKINVDCx6p67_ASAP7_75t_R g1399 ( 
.A(n_1330),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1303),
.A2(n_1322),
.B1(n_1221),
.B2(n_1203),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1253),
.Y(n_1401)
);

AOI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1351),
.A2(n_1221),
.B1(n_1239),
.B2(n_1251),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1214),
.Y(n_1403)
);

OAI21xp33_ASAP7_75t_L g1404 ( 
.A1(n_1309),
.A2(n_1311),
.B(n_1201),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1293),
.Y(n_1405)
);

NAND2x1p5_ASAP7_75t_L g1406 ( 
.A(n_1267),
.B(n_1205),
.Y(n_1406)
);

CKINVDCx14_ASAP7_75t_R g1407 ( 
.A(n_1258),
.Y(n_1407)
);

BUFx4f_ASAP7_75t_L g1408 ( 
.A(n_1346),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1259),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1315),
.A2(n_1218),
.B(n_1233),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1312),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1203),
.A2(n_1279),
.B1(n_1348),
.B2(n_1300),
.Y(n_1412)
);

INVx11_ASAP7_75t_L g1413 ( 
.A(n_1346),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1331),
.Y(n_1414)
);

BUFx2_ASAP7_75t_SL g1415 ( 
.A(n_1276),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1270),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_SL g1417 ( 
.A1(n_1343),
.A2(n_1247),
.B1(n_1204),
.B2(n_1216),
.Y(n_1417)
);

BUFx8_ASAP7_75t_L g1418 ( 
.A(n_1314),
.Y(n_1418)
);

AOI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1264),
.A2(n_1248),
.B1(n_1337),
.B2(n_1256),
.Y(n_1419)
);

INVx6_ASAP7_75t_L g1420 ( 
.A(n_1355),
.Y(n_1420)
);

INVx8_ASAP7_75t_L g1421 ( 
.A(n_1355),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1204),
.A2(n_1216),
.B1(n_1226),
.B2(n_1249),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1257),
.Y(n_1423)
);

CKINVDCx11_ASAP7_75t_R g1424 ( 
.A(n_1358),
.Y(n_1424)
);

BUFx12f_ASAP7_75t_L g1425 ( 
.A(n_1314),
.Y(n_1425)
);

AOI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1235),
.A2(n_1255),
.B1(n_1358),
.B2(n_1261),
.Y(n_1426)
);

BUFx12f_ASAP7_75t_L g1427 ( 
.A(n_1314),
.Y(n_1427)
);

INVxp67_ASAP7_75t_SL g1428 ( 
.A(n_1274),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_SL g1429 ( 
.A1(n_1229),
.A2(n_1232),
.B1(n_1292),
.B2(n_1317),
.Y(n_1429)
);

OAI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1358),
.A2(n_1231),
.B1(n_1230),
.B2(n_1242),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_SL g1431 ( 
.A1(n_1292),
.A2(n_1317),
.B1(n_1353),
.B2(n_1290),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_SL g1432 ( 
.A1(n_1292),
.A2(n_1353),
.B1(n_1316),
.B2(n_1211),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1210),
.A2(n_1329),
.B(n_1289),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1313),
.B(n_1347),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1205),
.A2(n_1336),
.B1(n_1338),
.B2(n_1268),
.Y(n_1435)
);

OAI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1336),
.A2(n_1338),
.B1(n_1223),
.B2(n_1263),
.Y(n_1436)
);

BUFx4f_ASAP7_75t_SL g1437 ( 
.A(n_1339),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1271),
.A2(n_1223),
.B1(n_1224),
.B2(n_1339),
.Y(n_1438)
);

BUFx12f_ASAP7_75t_L g1439 ( 
.A(n_1339),
.Y(n_1439)
);

BUFx12f_ASAP7_75t_L g1440 ( 
.A(n_1272),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1275),
.Y(n_1441)
);

BUFx3_ASAP7_75t_L g1442 ( 
.A(n_1273),
.Y(n_1442)
);

BUFx10_ASAP7_75t_L g1443 ( 
.A(n_1260),
.Y(n_1443)
);

BUFx4_ASAP7_75t_R g1444 ( 
.A(n_1266),
.Y(n_1444)
);

OAI21xp5_ASAP7_75t_SL g1445 ( 
.A1(n_1250),
.A2(n_1234),
.B(n_1223),
.Y(n_1445)
);

BUFx12f_ASAP7_75t_L g1446 ( 
.A(n_1281),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1281),
.A2(n_1225),
.B1(n_1280),
.B2(n_1288),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1277),
.A2(n_1347),
.B1(n_1342),
.B2(n_1332),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1254),
.Y(n_1449)
);

BUFx2_ASAP7_75t_L g1450 ( 
.A(n_1269),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_SL g1451 ( 
.A1(n_1266),
.A2(n_1347),
.B1(n_1342),
.B2(n_1332),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1332),
.A2(n_1342),
.B1(n_1357),
.B2(n_1294),
.Y(n_1452)
);

INVxp67_ASAP7_75t_SL g1453 ( 
.A(n_1278),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1283),
.A2(n_1284),
.B1(n_1349),
.B2(n_1345),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_SL g1455 ( 
.A1(n_1266),
.A2(n_1321),
.B1(n_1326),
.B2(n_1324),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_SL g1456 ( 
.A1(n_1356),
.A2(n_1282),
.B1(n_1327),
.B2(n_1340),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1213),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1213),
.A2(n_1208),
.B1(n_1227),
.B2(n_1215),
.Y(n_1458)
);

BUFx12f_ASAP7_75t_L g1459 ( 
.A(n_1215),
.Y(n_1459)
);

BUFx2_ASAP7_75t_L g1460 ( 
.A(n_1215),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_1227),
.Y(n_1461)
);

INVx1_ASAP7_75t_SL g1462 ( 
.A(n_1320),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1246),
.Y(n_1463)
);

AOI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1302),
.A2(n_1195),
.B1(n_1101),
.B2(n_1092),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1325),
.B(n_1350),
.Y(n_1465)
);

BUFx2_ASAP7_75t_L g1466 ( 
.A(n_1320),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1320),
.Y(n_1467)
);

OAI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1220),
.A2(n_1197),
.B1(n_850),
.B2(n_1291),
.Y(n_1468)
);

OAI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1220),
.A2(n_1301),
.B1(n_1291),
.B2(n_1085),
.Y(n_1469)
);

CKINVDCx11_ASAP7_75t_R g1470 ( 
.A(n_1295),
.Y(n_1470)
);

NAND2x1p5_ASAP7_75t_L g1471 ( 
.A(n_1238),
.B(n_1330),
.Y(n_1471)
);

INVx5_ASAP7_75t_L g1472 ( 
.A(n_1346),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1212),
.Y(n_1473)
);

INVx6_ASAP7_75t_L g1474 ( 
.A(n_1238),
.Y(n_1474)
);

OAI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1220),
.A2(n_1301),
.B1(n_1291),
.B2(n_1085),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1212),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1220),
.A2(n_1197),
.B1(n_850),
.B2(n_1291),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1212),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1220),
.A2(n_1197),
.B1(n_850),
.B2(n_1291),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1325),
.B(n_1350),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1220),
.A2(n_1197),
.B1(n_850),
.B2(n_1291),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1212),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1212),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1246),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1206),
.A2(n_1195),
.B1(n_1334),
.B2(n_1287),
.Y(n_1485)
);

AOI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1211),
.A2(n_850),
.B(n_1204),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1220),
.A2(n_1197),
.B1(n_850),
.B2(n_1291),
.Y(n_1487)
);

OAI21xp33_ASAP7_75t_SL g1488 ( 
.A1(n_1291),
.A2(n_1301),
.B(n_1197),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1212),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1212),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1212),
.Y(n_1491)
);

INVx4_ASAP7_75t_SL g1492 ( 
.A(n_1346),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1374),
.A2(n_1469),
.B1(n_1475),
.B2(n_1479),
.Y(n_1493)
);

AO21x2_ASAP7_75t_L g1494 ( 
.A1(n_1410),
.A2(n_1433),
.B(n_1379),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1449),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1391),
.B(n_1393),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1370),
.A2(n_1485),
.B1(n_1383),
.B2(n_1464),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1434),
.B(n_1368),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1370),
.A2(n_1485),
.B1(n_1383),
.B2(n_1481),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1469),
.A2(n_1475),
.B1(n_1468),
.B2(n_1487),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1457),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_SL g1502 ( 
.A1(n_1477),
.A2(n_1385),
.B1(n_1387),
.B2(n_1488),
.Y(n_1502)
);

AO21x1_ASAP7_75t_SL g1503 ( 
.A1(n_1377),
.A2(n_1404),
.B(n_1402),
.Y(n_1503)
);

BUFx2_ASAP7_75t_L g1504 ( 
.A(n_1450),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1367),
.A2(n_1396),
.B1(n_1377),
.B2(n_1384),
.Y(n_1505)
);

OR2x6_ASAP7_75t_L g1506 ( 
.A(n_1486),
.B(n_1459),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1368),
.B(n_1409),
.Y(n_1507)
);

O2A1O1Ixp33_ASAP7_75t_SL g1508 ( 
.A1(n_1367),
.A2(n_1465),
.B(n_1371),
.C(n_1480),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1382),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1454),
.A2(n_1452),
.B(n_1484),
.Y(n_1510)
);

INVx2_ASAP7_75t_SL g1511 ( 
.A(n_1361),
.Y(n_1511)
);

OAI21x1_ASAP7_75t_L g1512 ( 
.A1(n_1454),
.A2(n_1452),
.B(n_1463),
.Y(n_1512)
);

AND2x4_ASAP7_75t_SL g1513 ( 
.A(n_1443),
.B(n_1426),
.Y(n_1513)
);

AOI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1423),
.A2(n_1403),
.B(n_1405),
.Y(n_1514)
);

INVx1_ASAP7_75t_SL g1515 ( 
.A(n_1441),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1451),
.B(n_1398),
.Y(n_1516)
);

AO21x2_ASAP7_75t_L g1517 ( 
.A1(n_1379),
.A2(n_1430),
.B(n_1445),
.Y(n_1517)
);

OAI21x1_ASAP7_75t_L g1518 ( 
.A1(n_1403),
.A2(n_1411),
.B(n_1447),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_1470),
.Y(n_1519)
);

OA21x2_ASAP7_75t_L g1520 ( 
.A1(n_1458),
.A2(n_1411),
.B(n_1400),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1408),
.A2(n_1414),
.B1(n_1390),
.B2(n_1412),
.Y(n_1521)
);

AO21x1_ASAP7_75t_L g1522 ( 
.A1(n_1428),
.A2(n_1430),
.B(n_1436),
.Y(n_1522)
);

OR2x6_ASAP7_75t_L g1523 ( 
.A(n_1460),
.B(n_1421),
.Y(n_1523)
);

INVx3_ASAP7_75t_L g1524 ( 
.A(n_1406),
.Y(n_1524)
);

A2O1A1Ixp33_ASAP7_75t_L g1525 ( 
.A1(n_1400),
.A2(n_1408),
.B(n_1419),
.C(n_1412),
.Y(n_1525)
);

OA21x2_ASAP7_75t_L g1526 ( 
.A1(n_1458),
.A2(n_1422),
.B(n_1447),
.Y(n_1526)
);

AO21x1_ASAP7_75t_SL g1527 ( 
.A1(n_1422),
.A2(n_1438),
.B(n_1448),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1440),
.A2(n_1443),
.B1(n_1401),
.B2(n_1466),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1461),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1395),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1453),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1359),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1394),
.B(n_1417),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1448),
.Y(n_1534)
);

INVx2_ASAP7_75t_SL g1535 ( 
.A(n_1361),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1429),
.B(n_1431),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1432),
.B(n_1438),
.Y(n_1537)
);

INVx2_ASAP7_75t_SL g1538 ( 
.A(n_1361),
.Y(n_1538)
);

OR2x6_ASAP7_75t_L g1539 ( 
.A(n_1421),
.B(n_1420),
.Y(n_1539)
);

BUFx3_ASAP7_75t_L g1540 ( 
.A(n_1420),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1436),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1360),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1362),
.Y(n_1543)
);

OAI21x1_ASAP7_75t_L g1544 ( 
.A1(n_1435),
.A2(n_1471),
.B(n_1491),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1444),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1372),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1462),
.B(n_1478),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1444),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1375),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1381),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1473),
.Y(n_1551)
);

NOR2x1p5_ASAP7_75t_L g1552 ( 
.A(n_1365),
.B(n_1359),
.Y(n_1552)
);

INVxp33_ASAP7_75t_L g1553 ( 
.A(n_1467),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1476),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1482),
.Y(n_1555)
);

BUFx6f_ASAP7_75t_L g1556 ( 
.A(n_1389),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1483),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1489),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1490),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1392),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1407),
.B(n_1380),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1392),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1455),
.Y(n_1563)
);

AO21x2_ASAP7_75t_L g1564 ( 
.A1(n_1456),
.A2(n_1392),
.B(n_1435),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1407),
.B(n_1373),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1442),
.Y(n_1566)
);

OAI21xp33_ASAP7_75t_SL g1567 ( 
.A1(n_1413),
.A2(n_1364),
.B(n_1366),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1389),
.Y(n_1568)
);

OAI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1471),
.A2(n_1472),
.B(n_1389),
.Y(n_1569)
);

INVx4_ASAP7_75t_L g1570 ( 
.A(n_1389),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1472),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1472),
.Y(n_1572)
);

NAND2x1p5_ASAP7_75t_L g1573 ( 
.A(n_1472),
.B(n_1364),
.Y(n_1573)
);

INVxp33_ASAP7_75t_L g1574 ( 
.A(n_1376),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1492),
.Y(n_1575)
);

INVxp67_ASAP7_75t_L g1576 ( 
.A(n_1378),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1446),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1492),
.Y(n_1578)
);

OAI21xp5_ASAP7_75t_L g1579 ( 
.A1(n_1502),
.A2(n_1366),
.B(n_1369),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1515),
.B(n_1421),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1496),
.B(n_1424),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1493),
.A2(n_1363),
.B1(n_1397),
.B2(n_1399),
.Y(n_1582)
);

AOI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1499),
.A2(n_1497),
.B1(n_1500),
.B2(n_1505),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1508),
.B(n_1388),
.Y(n_1584)
);

AOI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1499),
.A2(n_1386),
.B(n_1415),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1507),
.B(n_1416),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1515),
.B(n_1397),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1509),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1495),
.Y(n_1589)
);

A2O1A1Ixp33_ASAP7_75t_L g1590 ( 
.A1(n_1525),
.A2(n_1474),
.B(n_1418),
.C(n_1437),
.Y(n_1590)
);

A2O1A1Ixp33_ASAP7_75t_L g1591 ( 
.A1(n_1497),
.A2(n_1474),
.B(n_1418),
.C(n_1437),
.Y(n_1591)
);

OAI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1521),
.A2(n_1474),
.B(n_1427),
.Y(n_1592)
);

A2O1A1Ixp33_ASAP7_75t_L g1593 ( 
.A1(n_1521),
.A2(n_1425),
.B(n_1439),
.C(n_1516),
.Y(n_1593)
);

OAI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1528),
.A2(n_1544),
.B(n_1567),
.Y(n_1594)
);

INVx2_ASAP7_75t_SL g1595 ( 
.A(n_1566),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1513),
.B(n_1533),
.Y(n_1596)
);

AOI21xp33_ASAP7_75t_L g1597 ( 
.A1(n_1494),
.A2(n_1517),
.B(n_1533),
.Y(n_1597)
);

INVx3_ASAP7_75t_L g1598 ( 
.A(n_1524),
.Y(n_1598)
);

OR2x6_ASAP7_75t_L g1599 ( 
.A(n_1506),
.B(n_1522),
.Y(n_1599)
);

AO21x2_ASAP7_75t_L g1600 ( 
.A1(n_1514),
.A2(n_1494),
.B(n_1522),
.Y(n_1600)
);

OA21x2_ASAP7_75t_L g1601 ( 
.A1(n_1510),
.A2(n_1512),
.B(n_1518),
.Y(n_1601)
);

AO21x2_ASAP7_75t_L g1602 ( 
.A1(n_1514),
.A2(n_1494),
.B(n_1512),
.Y(n_1602)
);

CKINVDCx20_ASAP7_75t_R g1603 ( 
.A(n_1519),
.Y(n_1603)
);

A2O1A1Ixp33_ASAP7_75t_L g1604 ( 
.A1(n_1516),
.A2(n_1536),
.B(n_1513),
.C(n_1541),
.Y(n_1604)
);

AND2x4_ASAP7_75t_L g1605 ( 
.A(n_1560),
.B(n_1562),
.Y(n_1605)
);

AOI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1506),
.A2(n_1494),
.B(n_1564),
.Y(n_1606)
);

AOI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1506),
.A2(n_1552),
.B1(n_1576),
.B2(n_1517),
.Y(n_1607)
);

AOI21xp33_ASAP7_75t_L g1608 ( 
.A1(n_1517),
.A2(n_1563),
.B(n_1507),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_L g1609 ( 
.A(n_1553),
.B(n_1498),
.Y(n_1609)
);

A2O1A1Ixp33_ASAP7_75t_L g1610 ( 
.A1(n_1536),
.A2(n_1541),
.B(n_1537),
.C(n_1503),
.Y(n_1610)
);

OAI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1577),
.A2(n_1561),
.B1(n_1548),
.B2(n_1545),
.Y(n_1611)
);

AOI211xp5_ASAP7_75t_SL g1612 ( 
.A1(n_1563),
.A2(n_1534),
.B(n_1537),
.C(n_1571),
.Y(n_1612)
);

INVxp33_ASAP7_75t_L g1613 ( 
.A(n_1547),
.Y(n_1613)
);

OAI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1506),
.A2(n_1569),
.B(n_1571),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_1532),
.Y(n_1615)
);

INVxp67_ASAP7_75t_L g1616 ( 
.A(n_1565),
.Y(n_1616)
);

CKINVDCx6p67_ASAP7_75t_R g1617 ( 
.A(n_1577),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1504),
.B(n_1542),
.Y(n_1618)
);

A2O1A1Ixp33_ASAP7_75t_L g1619 ( 
.A1(n_1503),
.A2(n_1569),
.B(n_1556),
.C(n_1540),
.Y(n_1619)
);

O2A1O1Ixp33_ASAP7_75t_L g1620 ( 
.A1(n_1517),
.A2(n_1566),
.B(n_1572),
.C(n_1568),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1504),
.B(n_1543),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1546),
.B(n_1551),
.Y(n_1622)
);

OA21x2_ASAP7_75t_L g1623 ( 
.A1(n_1510),
.A2(n_1518),
.B(n_1501),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1551),
.B(n_1555),
.Y(n_1624)
);

AO32x2_ASAP7_75t_L g1625 ( 
.A1(n_1511),
.A2(n_1535),
.A3(n_1538),
.B1(n_1570),
.B2(n_1527),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1555),
.B(n_1557),
.Y(n_1626)
);

AO21x2_ASAP7_75t_L g1627 ( 
.A1(n_1501),
.A2(n_1531),
.B(n_1564),
.Y(n_1627)
);

NOR2x1_ASAP7_75t_SL g1628 ( 
.A(n_1539),
.B(n_1523),
.Y(n_1628)
);

AOI221xp5_ASAP7_75t_L g1629 ( 
.A1(n_1549),
.A2(n_1554),
.B1(n_1550),
.B2(n_1558),
.C(n_1531),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1549),
.B(n_1550),
.Y(n_1630)
);

NOR2x1_ASAP7_75t_SL g1631 ( 
.A(n_1539),
.B(n_1523),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1527),
.B(n_1520),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1588),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1583),
.A2(n_1539),
.B1(n_1526),
.B2(n_1556),
.Y(n_1634)
);

NAND2x1_ASAP7_75t_L g1635 ( 
.A(n_1599),
.B(n_1570),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1632),
.B(n_1623),
.Y(n_1636)
);

INVx2_ASAP7_75t_R g1637 ( 
.A(n_1589),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1613),
.B(n_1554),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1592),
.B(n_1556),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1605),
.B(n_1628),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1627),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1623),
.B(n_1529),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1605),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1618),
.B(n_1621),
.Y(n_1644)
);

HB1xp67_ASAP7_75t_L g1645 ( 
.A(n_1627),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1609),
.Y(n_1646)
);

BUFx6f_ASAP7_75t_L g1647 ( 
.A(n_1601),
.Y(n_1647)
);

AOI222xp33_ASAP7_75t_L g1648 ( 
.A1(n_1584),
.A2(n_1552),
.B1(n_1574),
.B2(n_1558),
.C1(n_1530),
.C2(n_1559),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1622),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1624),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1602),
.B(n_1520),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_1595),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1625),
.B(n_1600),
.Y(n_1653)
);

BUFx2_ASAP7_75t_L g1654 ( 
.A(n_1625),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1631),
.B(n_1562),
.Y(n_1655)
);

HB1xp67_ASAP7_75t_L g1656 ( 
.A(n_1595),
.Y(n_1656)
);

BUFx8_ASAP7_75t_SL g1657 ( 
.A(n_1603),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1625),
.B(n_1520),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1584),
.A2(n_1526),
.B1(n_1564),
.B2(n_1520),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1626),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1630),
.Y(n_1661)
);

BUFx3_ASAP7_75t_L g1662 ( 
.A(n_1635),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1636),
.B(n_1625),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1661),
.B(n_1609),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1636),
.B(n_1600),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1642),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1661),
.B(n_1630),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1655),
.B(n_1598),
.Y(n_1668)
);

NOR2x1_ASAP7_75t_L g1669 ( 
.A(n_1654),
.B(n_1599),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1636),
.B(n_1606),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1658),
.B(n_1599),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1658),
.B(n_1599),
.Y(n_1672)
);

INVx1_ASAP7_75t_SL g1673 ( 
.A(n_1652),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1652),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1658),
.B(n_1597),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1633),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1653),
.B(n_1608),
.Y(n_1677)
);

INVx2_ASAP7_75t_SL g1678 ( 
.A(n_1640),
.Y(n_1678)
);

OAI21xp33_ASAP7_75t_L g1679 ( 
.A1(n_1659),
.A2(n_1610),
.B(n_1604),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1643),
.B(n_1620),
.Y(n_1680)
);

OAI21xp33_ASAP7_75t_SL g1681 ( 
.A1(n_1653),
.A2(n_1607),
.B(n_1596),
.Y(n_1681)
);

BUFx3_ASAP7_75t_L g1682 ( 
.A(n_1635),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1656),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1633),
.Y(n_1684)
);

INVx3_ASAP7_75t_L g1685 ( 
.A(n_1647),
.Y(n_1685)
);

OAI21xp33_ASAP7_75t_SL g1686 ( 
.A1(n_1653),
.A2(n_1596),
.B(n_1629),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1644),
.B(n_1637),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1637),
.B(n_1614),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1660),
.B(n_1613),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1637),
.B(n_1526),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1644),
.B(n_1526),
.Y(n_1691)
);

INVxp67_ASAP7_75t_L g1692 ( 
.A(n_1656),
.Y(n_1692)
);

OAI221xp5_ASAP7_75t_L g1693 ( 
.A1(n_1659),
.A2(n_1610),
.B1(n_1593),
.B2(n_1590),
.C(n_1604),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1666),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1675),
.B(n_1641),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1674),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1663),
.B(n_1670),
.Y(n_1697)
);

OAI31xp33_ASAP7_75t_L g1698 ( 
.A1(n_1679),
.A2(n_1693),
.A3(n_1612),
.B(n_1634),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1675),
.B(n_1641),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1674),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1678),
.B(n_1640),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1663),
.B(n_1651),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1667),
.B(n_1646),
.Y(n_1703)
);

AND2x4_ASAP7_75t_L g1704 ( 
.A(n_1678),
.B(n_1640),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1676),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1683),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1676),
.Y(n_1707)
);

HB1xp67_ASAP7_75t_L g1708 ( 
.A(n_1683),
.Y(n_1708)
);

HB1xp67_ASAP7_75t_L g1709 ( 
.A(n_1692),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1663),
.B(n_1651),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1676),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1678),
.B(n_1640),
.Y(n_1712)
);

INVxp67_ASAP7_75t_SL g1713 ( 
.A(n_1692),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1670),
.B(n_1651),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1670),
.B(n_1649),
.Y(n_1715)
);

BUFx2_ASAP7_75t_L g1716 ( 
.A(n_1669),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1673),
.Y(n_1717)
);

NAND2x1p5_ASAP7_75t_L g1718 ( 
.A(n_1669),
.B(n_1635),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_L g1719 ( 
.A(n_1664),
.B(n_1646),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1666),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1671),
.B(n_1650),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1684),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_1664),
.Y(n_1723)
);

BUFx2_ASAP7_75t_L g1724 ( 
.A(n_1716),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1701),
.B(n_1662),
.Y(n_1725)
);

INVx1_ASAP7_75t_SL g1726 ( 
.A(n_1723),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1709),
.Y(n_1727)
);

AND2x4_ASAP7_75t_L g1728 ( 
.A(n_1701),
.B(n_1662),
.Y(n_1728)
);

NAND2x1p5_ASAP7_75t_L g1729 ( 
.A(n_1716),
.B(n_1669),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1719),
.B(n_1689),
.Y(n_1730)
);

BUFx2_ASAP7_75t_L g1731 ( 
.A(n_1716),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1703),
.B(n_1675),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1701),
.B(n_1662),
.Y(n_1733)
);

INVxp67_ASAP7_75t_L g1734 ( 
.A(n_1719),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1697),
.B(n_1671),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1709),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1708),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1697),
.B(n_1672),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1723),
.B(n_1689),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1703),
.B(n_1677),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1697),
.B(n_1672),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1717),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1705),
.Y(n_1743)
);

NAND4xp75_ASAP7_75t_L g1744 ( 
.A(n_1698),
.B(n_1686),
.C(n_1681),
.D(n_1639),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1708),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1698),
.B(n_1667),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1717),
.B(n_1680),
.Y(n_1747)
);

INVx2_ASAP7_75t_SL g1748 ( 
.A(n_1701),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1714),
.B(n_1672),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1714),
.B(n_1680),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1714),
.B(n_1701),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1701),
.B(n_1668),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1715),
.B(n_1680),
.Y(n_1753)
);

NAND2x1_ASAP7_75t_L g1754 ( 
.A(n_1704),
.B(n_1712),
.Y(n_1754)
);

AND2x4_ASAP7_75t_SL g1755 ( 
.A(n_1704),
.B(n_1617),
.Y(n_1755)
);

NOR2x1p5_ASAP7_75t_L g1756 ( 
.A(n_1713),
.B(n_1617),
.Y(n_1756)
);

INVx2_ASAP7_75t_SL g1757 ( 
.A(n_1704),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1695),
.B(n_1677),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1704),
.B(n_1668),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1713),
.B(n_1657),
.Y(n_1760)
);

NAND4xp25_ASAP7_75t_SL g1761 ( 
.A(n_1702),
.B(n_1686),
.C(n_1681),
.D(n_1693),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1695),
.B(n_1677),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1704),
.B(n_1668),
.Y(n_1763)
);

INVx1_ASAP7_75t_SL g1764 ( 
.A(n_1696),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_L g1765 ( 
.A(n_1715),
.B(n_1657),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1704),
.B(n_1668),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1734),
.B(n_1691),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_SL g1768 ( 
.A(n_1744),
.B(n_1679),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1735),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1746),
.B(n_1696),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1727),
.B(n_1700),
.Y(n_1771)
);

NAND2x1_ASAP7_75t_L g1772 ( 
.A(n_1724),
.B(n_1712),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1765),
.B(n_1721),
.Y(n_1773)
);

AOI22xp33_ASAP7_75t_L g1774 ( 
.A1(n_1761),
.A2(n_1679),
.B1(n_1634),
.B2(n_1686),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1727),
.B(n_1736),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1742),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1736),
.B(n_1700),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1730),
.B(n_1732),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1732),
.B(n_1740),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1740),
.B(n_1691),
.Y(n_1780)
);

OR2x2_ASAP7_75t_L g1781 ( 
.A(n_1747),
.B(n_1691),
.Y(n_1781)
);

AND2x4_ASAP7_75t_L g1782 ( 
.A(n_1756),
.B(n_1712),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1737),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1737),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1750),
.B(n_1706),
.Y(n_1785)
);

NAND2x1_ASAP7_75t_L g1786 ( 
.A(n_1724),
.B(n_1712),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1753),
.B(n_1706),
.Y(n_1787)
);

OR2x2_ASAP7_75t_L g1788 ( 
.A(n_1739),
.B(n_1695),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1764),
.B(n_1702),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1758),
.B(n_1699),
.Y(n_1790)
);

AOI211xp5_ASAP7_75t_L g1791 ( 
.A1(n_1760),
.A2(n_1681),
.B(n_1590),
.C(n_1639),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1745),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1745),
.B(n_1702),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1726),
.B(n_1721),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1756),
.B(n_1721),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1735),
.Y(n_1796)
);

OAI21xp5_ASAP7_75t_SL g1797 ( 
.A1(n_1729),
.A2(n_1648),
.B(n_1718),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1743),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1758),
.B(n_1699),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1762),
.B(n_1699),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1731),
.B(n_1710),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1755),
.B(n_1712),
.Y(n_1802)
);

NOR4xp25_ASAP7_75t_SL g1803 ( 
.A(n_1797),
.B(n_1731),
.C(n_1744),
.D(n_1729),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1768),
.A2(n_1729),
.B(n_1603),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1779),
.B(n_1770),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1783),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1794),
.B(n_1738),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1784),
.Y(n_1808)
);

OAI21xp5_ASAP7_75t_L g1809 ( 
.A1(n_1768),
.A2(n_1688),
.B(n_1718),
.Y(n_1809)
);

AOI21xp33_ASAP7_75t_L g1810 ( 
.A1(n_1770),
.A2(n_1762),
.B(n_1648),
.Y(n_1810)
);

OAI32xp33_ASAP7_75t_L g1811 ( 
.A1(n_1774),
.A2(n_1718),
.A3(n_1685),
.B1(n_1688),
.B2(n_1757),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1792),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1775),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1772),
.Y(n_1814)
);

AOI32xp33_ASAP7_75t_L g1815 ( 
.A1(n_1774),
.A2(n_1688),
.A3(n_1738),
.B1(n_1741),
.B2(n_1755),
.Y(n_1815)
);

NAND2x1p5_ASAP7_75t_L g1816 ( 
.A(n_1786),
.B(n_1754),
.Y(n_1816)
);

AOI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1782),
.A2(n_1755),
.B1(n_1725),
.B2(n_1728),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1775),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1776),
.B(n_1741),
.Y(n_1819)
);

NAND3xp33_ASAP7_75t_L g1820 ( 
.A(n_1791),
.B(n_1593),
.C(n_1645),
.Y(n_1820)
);

NOR2xp33_ASAP7_75t_L g1821 ( 
.A(n_1778),
.B(n_1615),
.Y(n_1821)
);

A2O1A1Ixp33_ASAP7_75t_L g1822 ( 
.A1(n_1788),
.A2(n_1594),
.B(n_1591),
.C(n_1581),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1773),
.B(n_1749),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1795),
.B(n_1782),
.Y(n_1824)
);

AOI31xp33_ASAP7_75t_L g1825 ( 
.A1(n_1790),
.A2(n_1615),
.A3(n_1582),
.B(n_1718),
.Y(n_1825)
);

INVxp67_ASAP7_75t_SL g1826 ( 
.A(n_1801),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_L g1827 ( 
.A(n_1769),
.B(n_1616),
.Y(n_1827)
);

OA21x2_ASAP7_75t_L g1828 ( 
.A1(n_1771),
.A2(n_1743),
.B(n_1707),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1826),
.B(n_1796),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1826),
.B(n_1789),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1805),
.B(n_1785),
.Y(n_1831)
);

OAI22xp5_ASAP7_75t_L g1832 ( 
.A1(n_1803),
.A2(n_1820),
.B1(n_1822),
.B2(n_1825),
.Y(n_1832)
);

AOI21xp5_ASAP7_75t_L g1833 ( 
.A1(n_1804),
.A2(n_1777),
.B(n_1771),
.Y(n_1833)
);

NAND2x1p5_ASAP7_75t_L g1834 ( 
.A(n_1821),
.B(n_1802),
.Y(n_1834)
);

OAI21xp5_ASAP7_75t_L g1835 ( 
.A1(n_1822),
.A2(n_1777),
.B(n_1801),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1806),
.Y(n_1836)
);

AOI21xp33_ASAP7_75t_SL g1837 ( 
.A1(n_1821),
.A2(n_1800),
.B(n_1799),
.Y(n_1837)
);

AOI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1810),
.A2(n_1789),
.B(n_1793),
.Y(n_1838)
);

O2A1O1Ixp33_ASAP7_75t_L g1839 ( 
.A1(n_1811),
.A2(n_1813),
.B(n_1818),
.C(n_1809),
.Y(n_1839)
);

AOI221xp5_ASAP7_75t_L g1840 ( 
.A1(n_1815),
.A2(n_1808),
.B1(n_1812),
.B2(n_1819),
.C(n_1823),
.Y(n_1840)
);

AOI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1814),
.A2(n_1793),
.B(n_1767),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1828),
.Y(n_1842)
);

NOR2xp33_ASAP7_75t_L g1843 ( 
.A(n_1824),
.B(n_1827),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1828),
.Y(n_1844)
);

O2A1O1Ixp33_ASAP7_75t_L g1845 ( 
.A1(n_1827),
.A2(n_1787),
.B(n_1798),
.C(n_1781),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1828),
.Y(n_1846)
);

INVxp67_ASAP7_75t_L g1847 ( 
.A(n_1807),
.Y(n_1847)
);

INVx1_ASAP7_75t_SL g1848 ( 
.A(n_1817),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1829),
.Y(n_1849)
);

OAI22xp33_ASAP7_75t_L g1850 ( 
.A1(n_1832),
.A2(n_1816),
.B1(n_1718),
.B2(n_1754),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1842),
.Y(n_1851)
);

XNOR2x1_ASAP7_75t_L g1852 ( 
.A(n_1848),
.B(n_1586),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1847),
.B(n_1749),
.Y(n_1853)
);

OAI21xp5_ASAP7_75t_SL g1854 ( 
.A1(n_1834),
.A2(n_1816),
.B(n_1802),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1844),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1846),
.Y(n_1856)
);

NAND3xp33_ASAP7_75t_L g1857 ( 
.A(n_1833),
.B(n_1780),
.C(n_1645),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1836),
.Y(n_1858)
);

NAND2x1_ASAP7_75t_L g1859 ( 
.A(n_1843),
.B(n_1725),
.Y(n_1859)
);

OAI221xp5_ASAP7_75t_L g1860 ( 
.A1(n_1835),
.A2(n_1757),
.B1(n_1748),
.B2(n_1662),
.C(n_1682),
.Y(n_1860)
);

AOI322xp5_ASAP7_75t_L g1861 ( 
.A1(n_1840),
.A2(n_1710),
.A3(n_1665),
.B1(n_1751),
.B2(n_1748),
.C1(n_1690),
.C2(n_1733),
.Y(n_1861)
);

AOI211xp5_ASAP7_75t_L g1862 ( 
.A1(n_1854),
.A2(n_1839),
.B(n_1837),
.C(n_1838),
.Y(n_1862)
);

INVxp67_ASAP7_75t_L g1863 ( 
.A(n_1852),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1853),
.B(n_1831),
.Y(n_1864)
);

AOI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1850),
.A2(n_1834),
.B1(n_1830),
.B2(n_1841),
.Y(n_1865)
);

INVx2_ASAP7_75t_SL g1866 ( 
.A(n_1859),
.Y(n_1866)
);

AND4x1_ASAP7_75t_SL g1867 ( 
.A(n_1861),
.B(n_1845),
.C(n_1587),
.D(n_1580),
.Y(n_1867)
);

NOR3x1_ASAP7_75t_L g1868 ( 
.A(n_1849),
.B(n_1579),
.C(n_1611),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1858),
.B(n_1751),
.Y(n_1869)
);

NOR2xp33_ASAP7_75t_SL g1870 ( 
.A(n_1860),
.B(n_1725),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1851),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1855),
.B(n_1710),
.Y(n_1872)
);

BUFx2_ASAP7_75t_L g1873 ( 
.A(n_1866),
.Y(n_1873)
);

AOI21xp33_ASAP7_75t_SL g1874 ( 
.A1(n_1863),
.A2(n_1857),
.B(n_1856),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1864),
.Y(n_1875)
);

AOI211x1_ASAP7_75t_SL g1876 ( 
.A1(n_1872),
.A2(n_1857),
.B(n_1720),
.C(n_1694),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1862),
.B(n_1665),
.Y(n_1877)
);

AOI221xp5_ASAP7_75t_L g1878 ( 
.A1(n_1874),
.A2(n_1871),
.B1(n_1865),
.B2(n_1869),
.C(n_1870),
.Y(n_1878)
);

AOI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1875),
.A2(n_1725),
.B1(n_1728),
.B2(n_1733),
.Y(n_1879)
);

OA211x2_ASAP7_75t_L g1880 ( 
.A1(n_1877),
.A2(n_1867),
.B(n_1868),
.C(n_1638),
.Y(n_1880)
);

AOI211xp5_ASAP7_75t_L g1881 ( 
.A1(n_1873),
.A2(n_1728),
.B(n_1733),
.C(n_1591),
.Y(n_1881)
);

AOI211xp5_ASAP7_75t_L g1882 ( 
.A1(n_1873),
.A2(n_1728),
.B(n_1733),
.C(n_1682),
.Y(n_1882)
);

HB1xp67_ASAP7_75t_L g1883 ( 
.A(n_1876),
.Y(n_1883)
);

INVx2_ASAP7_75t_SL g1884 ( 
.A(n_1879),
.Y(n_1884)
);

INVxp67_ASAP7_75t_L g1885 ( 
.A(n_1883),
.Y(n_1885)
);

AOI22xp33_ASAP7_75t_L g1886 ( 
.A1(n_1880),
.A2(n_1682),
.B1(n_1685),
.B2(n_1759),
.Y(n_1886)
);

NOR3xp33_ASAP7_75t_L g1887 ( 
.A(n_1878),
.B(n_1685),
.C(n_1585),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1881),
.B(n_1665),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1888),
.Y(n_1889)
);

OAI21xp5_ASAP7_75t_SL g1890 ( 
.A1(n_1885),
.A2(n_1882),
.B(n_1759),
.Y(n_1890)
);

OAI221xp5_ASAP7_75t_L g1891 ( 
.A1(n_1884),
.A2(n_1682),
.B1(n_1685),
.B2(n_1619),
.C(n_1687),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1889),
.Y(n_1892)
);

OAI22xp5_ASAP7_75t_L g1893 ( 
.A1(n_1892),
.A2(n_1891),
.B1(n_1886),
.B2(n_1890),
.Y(n_1893)
);

OAI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1893),
.A2(n_1887),
.B1(n_1694),
.B2(n_1720),
.Y(n_1894)
);

XNOR2x1_ASAP7_75t_L g1895 ( 
.A(n_1893),
.B(n_1573),
.Y(n_1895)
);

XNOR2xp5_ASAP7_75t_L g1896 ( 
.A(n_1895),
.B(n_1573),
.Y(n_1896)
);

OAI22xp5_ASAP7_75t_SL g1897 ( 
.A1(n_1894),
.A2(n_1573),
.B1(n_1538),
.B2(n_1535),
.Y(n_1897)
);

OAI22xp33_ASAP7_75t_L g1898 ( 
.A1(n_1896),
.A2(n_1720),
.B1(n_1694),
.B2(n_1685),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_SL g1899 ( 
.A(n_1897),
.B(n_1766),
.Y(n_1899)
);

AOI21xp5_ASAP7_75t_L g1900 ( 
.A1(n_1899),
.A2(n_1763),
.B(n_1752),
.Y(n_1900)
);

AO21x2_ASAP7_75t_L g1901 ( 
.A1(n_1900),
.A2(n_1898),
.B(n_1763),
.Y(n_1901)
);

AOI22x1_ASAP7_75t_L g1902 ( 
.A1(n_1901),
.A2(n_1511),
.B1(n_1570),
.B2(n_1556),
.Y(n_1902)
);

AOI221xp5_ASAP7_75t_L g1903 ( 
.A1(n_1902),
.A2(n_1711),
.B1(n_1707),
.B2(n_1722),
.C(n_1705),
.Y(n_1903)
);

AOI211xp5_ASAP7_75t_L g1904 ( 
.A1(n_1903),
.A2(n_1578),
.B(n_1575),
.C(n_1556),
.Y(n_1904)
);


endmodule