module real_jpeg_4941_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_525;
wire n_78;
wire n_288;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_324;
wire n_86;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_0),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_52)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_0),
.A2(n_56),
.B1(n_307),
.B2(n_309),
.Y(n_306)
);

OAI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_0),
.A2(n_56),
.B1(n_203),
.B2(n_393),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_SL g407 ( 
.A1(n_0),
.A2(n_56),
.B1(n_360),
.B2(n_406),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_1),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_1),
.Y(n_195)
);

INVx8_ASAP7_75t_L g214 ( 
.A(n_1),
.Y(n_214)
);

BUFx5_ASAP7_75t_L g273 ( 
.A(n_1),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_1),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_2),
.A2(n_169),
.B1(n_202),
.B2(n_204),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_2),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_2),
.A2(n_204),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_2),
.A2(n_204),
.B1(n_296),
.B2(n_298),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_2),
.A2(n_204),
.B1(n_433),
.B2(n_435),
.Y(n_432)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_3),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_3),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_3),
.Y(n_324)
);

BUFx5_ASAP7_75t_L g434 ( 
.A(n_3),
.Y(n_434)
);

INVx6_ASAP7_75t_L g436 ( 
.A(n_3),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_4),
.A2(n_60),
.B1(n_62),
.B2(n_64),
.Y(n_59)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g341 ( 
.A1(n_4),
.A2(n_64),
.B1(n_342),
.B2(n_345),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_4),
.A2(n_64),
.B1(n_164),
.B2(n_397),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_4),
.A2(n_64),
.B1(n_448),
.B2(n_449),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_5),
.A2(n_119),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_5),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_5),
.A2(n_171),
.B1(n_190),
.B2(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_5),
.A2(n_171),
.B1(n_259),
.B2(n_261),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_5),
.A2(n_53),
.B1(n_171),
.B2(n_356),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_6),
.A2(n_93),
.B1(n_95),
.B2(n_96),
.Y(n_92)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_6),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_6),
.A2(n_96),
.B1(n_139),
.B2(n_144),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_6),
.A2(n_96),
.B1(n_378),
.B2(n_380),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_6),
.A2(n_96),
.B1(n_118),
.B2(n_416),
.Y(n_415)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_9),
.Y(n_113)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_9),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_9),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_10),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_19)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_11),
.Y(n_87)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_12),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_12),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_12),
.Y(n_177)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_14),
.A2(n_162),
.B1(n_164),
.B2(n_166),
.Y(n_161)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_14),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_14),
.B(n_121),
.C(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_14),
.B(n_83),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_14),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_14),
.B(n_132),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_14),
.B(n_93),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_15),
.A2(n_181),
.B1(n_182),
.B2(n_186),
.Y(n_180)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_15),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_15),
.A2(n_118),
.B1(n_186),
.B2(n_248),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g359 ( 
.A1(n_15),
.A2(n_186),
.B1(n_360),
.B2(n_362),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_15),
.A2(n_186),
.B1(n_410),
.B2(n_411),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_16),
.A2(n_47),
.B1(n_99),
.B2(n_102),
.Y(n_98)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_16),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_16),
.A2(n_102),
.B1(n_134),
.B2(n_136),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_16),
.A2(n_62),
.B1(n_102),
.B2(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_16),
.A2(n_102),
.B1(n_219),
.B2(n_386),
.Y(n_385)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_18),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_18),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_18),
.A2(n_203),
.B1(n_269),
.B2(n_368),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_18),
.A2(n_269),
.B1(n_402),
.B2(n_404),
.Y(n_401)
);

OAI22xp33_ASAP7_75t_L g462 ( 
.A1(n_18),
.A2(n_269),
.B1(n_324),
.B2(n_433),
.Y(n_462)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_537),
.B(n_540),
.Y(n_24)
);

AO21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_151),
.B(n_536),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_148),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_27),
.B(n_148),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_137),
.C(n_145),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_28),
.A2(n_29),
.B1(n_532),
.B2(n_533),
.Y(n_531)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_65),
.C(n_103),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g523 ( 
.A(n_30),
.B(n_524),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_52),
.B1(n_57),
.B2(n_59),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_31),
.A2(n_57),
.B1(n_59),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_31),
.A2(n_57),
.B1(n_138),
.B2(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_31),
.A2(n_354),
.B(n_409),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_31),
.A2(n_42),
.B1(n_409),
.B2(n_432),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_31),
.A2(n_52),
.B1(n_57),
.B2(n_509),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_32),
.A2(n_352),
.B(n_353),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_32),
.B(n_355),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_32),
.A2(n_58),
.B(n_539),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_42),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_42),
.B(n_166),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_47),
.B2(n_50),
.Y(n_42)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_43),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_45),
.Y(n_260)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_45),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_46),
.Y(n_332)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_46),
.Y(n_403)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_46),
.Y(n_406)
);

OAI32xp33_ASAP7_75t_L g320 ( 
.A1(n_47),
.A2(n_321),
.A3(n_325),
.B1(n_327),
.B2(n_333),
.Y(n_320)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx5_ASAP7_75t_L g329 ( 
.A(n_51),
.Y(n_329)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp33_ASAP7_75t_SL g352 ( 
.A1(n_54),
.A2(n_166),
.B(n_333),
.Y(n_352)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_55),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_57),
.A2(n_432),
.B(n_463),
.Y(n_473)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_58),
.B(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_58),
.B(n_462),
.Y(n_461)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_61),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_61),
.Y(n_356)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_65),
.A2(n_103),
.B1(n_104),
.B2(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_65),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_92),
.B1(n_97),
.B2(n_98),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_66),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_66),
.A2(n_97),
.B1(n_295),
.B2(n_359),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_66),
.A2(n_97),
.B1(n_401),
.B2(n_407),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_66),
.A2(n_92),
.B1(n_97),
.B2(n_513),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_83),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_73),
.B1(n_76),
.B2(n_78),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx8_ASAP7_75t_L g278 ( 
.A(n_70),
.Y(n_278)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_72),
.Y(n_284)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

INVx6_ASAP7_75t_L g365 ( 
.A(n_75),
.Y(n_365)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_81),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g254 ( 
.A(n_82),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_82),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_82),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_82),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_83),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_83),
.A2(n_146),
.B(n_147),
.Y(n_145)
);

AOI22x1_ASAP7_75t_L g437 ( 
.A1(n_83),
.A2(n_146),
.B1(n_302),
.B2(n_438),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_83),
.A2(n_146),
.B1(n_446),
.B2(n_447),
.Y(n_445)
);

AO22x2_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_88),
.B2(n_90),
.Y(n_83)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_86),
.Y(n_203)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_87),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g281 ( 
.A(n_87),
.Y(n_281)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_87),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_89),
.Y(n_163)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_89),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_89),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_89),
.Y(n_398)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_97),
.B(n_258),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_97),
.A2(n_295),
.B(n_301),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_103),
.A2(n_104),
.B1(n_511),
.B2(n_512),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_103),
.B(n_508),
.C(n_511),
.Y(n_519)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_131),
.B(n_133),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_105),
.A2(n_161),
.B(n_167),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_105),
.A2(n_131),
.B1(n_201),
.B2(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_105),
.A2(n_167),
.B(n_247),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_105),
.A2(n_131),
.B1(n_367),
.B2(n_427),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_106),
.B(n_168),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_106),
.A2(n_132),
.B1(n_392),
.B2(n_396),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_106),
.A2(n_132),
.B1(n_396),
.B2(n_415),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_106),
.A2(n_132),
.B1(n_415),
.B2(n_453),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_120),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_111),
.B1(n_114),
.B2(n_118),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_110),
.Y(n_250)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_120),
.A2(n_201),
.B(n_205),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_123),
.B1(n_127),
.B2(n_129),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_125),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_126),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_126),
.Y(n_192)
);

INVx8_ASAP7_75t_L g310 ( 
.A(n_127),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_127),
.Y(n_345)
);

BUFx8_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_128),
.Y(n_390)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_131),
.A2(n_205),
.B(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_132),
.B(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_133),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_136),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_137),
.B(n_145),
.Y(n_533)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_144),
.B(n_166),
.Y(n_333)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_144),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_146),
.A2(n_253),
.B(n_257),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_146),
.B(n_302),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_146),
.A2(n_257),
.B(n_476),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_148),
.B(n_538),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_148),
.B(n_538),
.Y(n_541)
);

CKINVDCx16_ASAP7_75t_R g539 ( 
.A(n_149),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_530),
.B(n_535),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_502),
.B(n_527),
.Y(n_152)
);

OAI311xp33_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_371),
.A3(n_478),
.B1(n_496),
.C1(n_497),
.Y(n_153)
);

AOI21x1_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_314),
.B(n_370),
.Y(n_154)
);

AO21x1_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_286),
.B(n_313),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_241),
.B(n_285),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_208),
.B(n_240),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_178),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_159),
.B(n_178),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_172),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_160),
.A2(n_172),
.B1(n_173),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_160),
.Y(n_238)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_163),
.Y(n_165)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_166),
.A2(n_187),
.B(n_193),
.Y(n_215)
);

OAI21xp33_ASAP7_75t_SL g253 ( 
.A1(n_166),
.A2(n_254),
.B(n_255),
.Y(n_253)
);

INVx3_ASAP7_75t_SL g276 ( 
.A(n_169),
.Y(n_276)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_177),
.Y(n_223)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_177),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_177),
.Y(n_308)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_177),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_198),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_179),
.B(n_199),
.C(n_207),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_187),
.B(n_193),
.Y(n_179)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_180),
.Y(n_233)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_185),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_187),
.A2(n_336),
.B1(n_337),
.B2(n_340),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_187),
.A2(n_377),
.B1(n_382),
.B2(n_385),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_187),
.A2(n_385),
.B(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_188),
.B(n_196),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_188),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_188),
.A2(n_267),
.B1(n_306),
.B2(n_311),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_188),
.A2(n_341),
.B1(n_421),
.B2(n_429),
.Y(n_428)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_189),
.Y(n_236)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx8_ASAP7_75t_L g381 ( 
.A(n_192),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_195),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_212),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_206),
.B2(n_207),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_230),
.B(n_239),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_216),
.B(n_229),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_215),
.Y(n_210)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_214),
.Y(n_339)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_214),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_228),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_228),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_224),
.B(n_227),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_227),
.A2(n_266),
.B(n_273),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_237),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_237),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_235),
.Y(n_234)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_242),
.B(n_243),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_264),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_251),
.B2(n_252),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_246),
.B(n_251),
.C(n_264),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_250),
.Y(n_418)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVxp33_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

AOI32xp33_ASAP7_75t_L g274 ( 
.A1(n_256),
.A2(n_275),
.A3(n_276),
.B1(n_277),
.B2(n_279),
.Y(n_274)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_258),
.Y(n_302)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_274),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_274),
.Y(n_292)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp33_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_282),
.Y(n_279)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_287),
.B(n_288),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_293),
.B2(n_312),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_292),
.C(n_312),
.Y(n_315)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_293),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_303),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_294),
.B(n_304),
.C(n_305),
.Y(n_346)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

BUFx12f_ASAP7_75t_L g361 ( 
.A(n_297),
.Y(n_361)
);

INVx4_ASAP7_75t_SL g298 ( 
.A(n_299),
.Y(n_298)
);

INVx5_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_306),
.Y(n_336)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_315),
.B(n_316),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_349),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_346),
.B1(n_347),
.B2(n_348),
.Y(n_317)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_318),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_320),
.B1(n_334),
.B2(n_335),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_320),
.B(n_334),
.Y(n_474)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx8_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_330),
.Y(n_327)
);

INVx6_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_331),
.Y(n_330)
);

INVx6_ASAP7_75t_SL g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx6_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_346),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_346),
.B(n_347),
.C(n_349),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_350),
.A2(n_351),
.B1(n_357),
.B2(n_369),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_350),
.B(n_358),
.C(n_366),
.Y(n_487)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_357),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_358),
.B(n_366),
.Y(n_357)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_359),
.Y(n_476)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

NAND2xp33_ASAP7_75t_SL g371 ( 
.A(n_372),
.B(n_464),
.Y(n_371)
);

A2O1A1Ixp33_ASAP7_75t_SL g497 ( 
.A1(n_372),
.A2(n_464),
.B(n_498),
.C(n_501),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_439),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g496 ( 
.A(n_373),
.B(n_439),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_412),
.C(n_424),
.Y(n_373)
);

FAx1_ASAP7_75t_SL g477 ( 
.A(n_374),
.B(n_412),
.CI(n_424),
.CON(n_477),
.SN(n_477)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_399),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_375),
.B(n_400),
.C(n_408),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_391),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_376),
.B(n_391),
.Y(n_470)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_377),
.Y(n_429)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx4_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_387),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_392),
.Y(n_427)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_408),
.Y(n_399)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_401),
.Y(n_438)
);

INVx4_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_403),
.Y(n_450)
);

INVx4_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_407),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_413),
.A2(n_414),
.B1(n_419),
.B2(n_423),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_414),
.B(n_419),
.Y(n_457)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_419),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_419),
.A2(n_423),
.B1(n_459),
.B2(n_460),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_419),
.A2(n_457),
.B(n_460),
.Y(n_505)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_430),
.C(n_437),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_425),
.B(n_468),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_426),
.B(n_428),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_426),
.B(n_428),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_430),
.A2(n_431),
.B1(n_437),
.B2(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx8_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_437),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_441),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_440),
.B(n_443),
.C(n_455),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_442),
.A2(n_443),
.B1(n_455),
.B2(n_456),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_444),
.A2(n_451),
.B(n_454),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_445),
.B(n_452),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_447),
.Y(n_513)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

FAx1_ASAP7_75t_SL g504 ( 
.A(n_454),
.B(n_505),
.CI(n_506),
.CON(n_504),
.SN(n_504)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_454),
.B(n_505),
.C(n_506),
.Y(n_526)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_458),
.Y(n_456)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_463),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_462),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_477),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_465),
.B(n_477),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_470),
.C(n_471),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_466),
.A2(n_467),
.B1(n_470),
.B2(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_470),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_471),
.B(n_489),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_474),
.C(n_475),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_472),
.A2(n_473),
.B1(n_475),
.B2(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_474),
.B(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_475),
.Y(n_484)
);

BUFx24_ASAP7_75t_SL g542 ( 
.A(n_477),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_479),
.B(n_491),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_480),
.A2(n_499),
.B(n_500),
.Y(n_498)
);

NOR2x1_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_488),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_481),
.B(n_488),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_485),
.C(n_487),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_482),
.B(n_494),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_485),
.A2(n_486),
.B1(n_487),
.B2(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_487),
.Y(n_495)
);

OR2x2_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_493),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_492),
.B(n_493),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_516),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_504),
.B(n_515),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_504),
.B(n_515),
.Y(n_528)
);

BUFx24_ASAP7_75t_SL g543 ( 
.A(n_504),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_507),
.A2(n_508),
.B1(n_510),
.B2(n_514),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_507),
.A2(n_508),
.B1(n_522),
.B2(n_523),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_507),
.B(n_518),
.C(n_522),
.Y(n_534)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_510),
.Y(n_514)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_516),
.A2(n_528),
.B(n_529),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_517),
.B(n_526),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_517),
.B(n_526),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_518),
.A2(n_519),
.B1(n_520),
.B2(n_521),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_534),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_531),
.B(n_534),
.Y(n_535)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_541),
.Y(n_540)
);


endmodule