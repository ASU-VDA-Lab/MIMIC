module fake_jpeg_1188_n_142 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_142);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_25),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_53),
.Y(n_62)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_45),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_1),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_1),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NAND3xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_43),
.C(n_47),
.Y(n_77)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_66),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_51),
.A2(n_36),
.B1(n_47),
.B2(n_43),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_62),
.B(n_48),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_68),
.B(n_80),
.Y(n_93)
);

AO22x1_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_60),
.B1(n_67),
.B2(n_66),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_3),
.Y(n_87)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_58),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_72),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_48),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_40),
.B1(n_35),
.B2(n_41),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_41),
.B1(n_38),
.B2(n_42),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_42),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_74),
.B(n_6),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_2),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_49),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_82),
.B1(n_84),
.B2(n_87),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_76),
.A2(n_38),
.B1(n_44),
.B2(n_37),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_90),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_76),
.A2(n_37),
.B1(n_4),
.B2(n_5),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_37),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_85),
.B(n_91),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_89),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_3),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_4),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_94),
.B(n_95),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_70),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_102),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_69),
.B(n_79),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_108),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_87),
.A2(n_69),
.B1(n_7),
.B2(n_8),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_107),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_93),
.B(n_85),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_110),
.Y(n_122)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_6),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_111),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_21),
.C(n_32),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_114),
.Y(n_128)
);

AOI322xp5_ASAP7_75t_L g114 ( 
.A1(n_105),
.A2(n_19),
.A3(n_31),
.B1(n_30),
.B2(n_29),
.C1(n_26),
.C2(n_12),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_119),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_99),
.C(n_101),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_103),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_123)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_104),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_124),
.Y(n_126)
);

NOR2x1_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_103),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_125),
.A2(n_122),
.B(n_112),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_120),
.Y(n_130)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_132),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_119),
.C(n_129),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_127),
.A2(n_117),
.B1(n_107),
.B2(n_116),
.Y(n_133)
);

AOI322xp5_ASAP7_75t_L g136 ( 
.A1(n_133),
.A2(n_126),
.A3(n_129),
.B1(n_118),
.B2(n_112),
.C1(n_127),
.C2(n_128),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_132),
.B1(n_135),
.B2(n_134),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_137),
.A2(n_113),
.B(n_115),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_14),
.C(n_16),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_22),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_23),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_24),
.Y(n_142)
);


endmodule