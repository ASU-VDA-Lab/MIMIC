module fake_jpeg_5557_n_307 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_307);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_307;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_42),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_16),
.Y(n_53)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx2_ASAP7_75t_SL g73 ( 
.A(n_45),
.Y(n_73)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_46),
.B(n_61),
.Y(n_75)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_52),
.Y(n_71)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_33),
.B1(n_30),
.B2(n_26),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_64),
.B1(n_65),
.B2(n_69),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_31),
.B1(n_33),
.B2(n_17),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

NAND2xp33_ASAP7_75t_SL g55 ( 
.A(n_40),
.B(n_29),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_55),
.A2(n_26),
.B(n_29),
.C(n_25),
.Y(n_90)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_63),
.Y(n_82)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_43),
.A2(n_17),
.B1(n_19),
.B2(n_27),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_17),
.B1(n_19),
.B2(n_27),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_19),
.Y(n_66)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_37),
.A2(n_31),
.B1(n_33),
.B2(n_27),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_50),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_76),
.B(n_77),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_46),
.B(n_28),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_81),
.Y(n_98)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_44),
.B(n_28),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_85),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_86),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_31),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_67),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_87),
.A2(n_62),
.B1(n_57),
.B2(n_18),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_32),
.Y(n_89)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_92),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_45),
.B(n_68),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_95),
.B(n_96),
.Y(n_139)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_100),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_72),
.Y(n_99)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_55),
.B1(n_54),
.B2(n_48),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_101),
.A2(n_108),
.B1(n_89),
.B2(n_74),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_82),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_105),
.Y(n_129)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_44),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_107),
.A2(n_80),
.B(n_20),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_54),
.B1(n_58),
.B2(n_59),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_113),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_70),
.A2(n_29),
.B1(n_63),
.B2(n_52),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_73),
.Y(n_116)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_70),
.A2(n_49),
.B1(n_24),
.B2(n_20),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_118),
.A2(n_86),
.B1(n_81),
.B2(n_82),
.Y(n_134)
);

OR2x2_ASAP7_75t_SL g119 ( 
.A(n_103),
.B(n_76),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_SL g156 ( 
.A1(n_119),
.A2(n_114),
.B(n_77),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_90),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_140),
.C(n_141),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_104),
.A2(n_79),
.B1(n_74),
.B2(n_83),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_126),
.Y(n_163)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_127),
.B(n_133),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_131),
.A2(n_93),
.B1(n_109),
.B2(n_32),
.Y(n_166)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_134),
.A2(n_110),
.B1(n_113),
.B2(n_116),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_135),
.A2(n_137),
.B(n_18),
.Y(n_158)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_136),
.B(n_144),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_104),
.A2(n_96),
.B(n_95),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_138),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_79),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_87),
.C(n_84),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_103),
.A2(n_97),
.B(n_100),
.Y(n_143)
);

AO21x1_ASAP7_75t_L g162 ( 
.A1(n_143),
.A2(n_18),
.B(n_21),
.Y(n_162)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_94),
.Y(n_146)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_125),
.A2(n_112),
.B1(n_107),
.B2(n_94),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_147),
.A2(n_162),
.B(n_130),
.Y(n_176)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_148),
.B(n_149),
.Y(n_192)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_151),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_118),
.C(n_114),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_161),
.C(n_126),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_119),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_154),
.A2(n_158),
.B(n_159),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_156),
.A2(n_163),
.B1(n_167),
.B2(n_149),
.Y(n_185)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_157),
.A2(n_164),
.B1(n_165),
.B2(n_169),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_24),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_122),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_160),
.B(n_168),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_80),
.C(n_115),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_166),
.A2(n_128),
.B1(n_99),
.B2(n_130),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_135),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_167),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_134),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_125),
.A2(n_99),
.B1(n_93),
.B2(n_106),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_170),
.A2(n_121),
.B1(n_93),
.B2(n_122),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_171),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_178),
.C(n_180),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_169),
.A2(n_128),
.B(n_129),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_173),
.A2(n_175),
.B1(n_191),
.B2(n_157),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_162),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_124),
.C(n_121),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_170),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_186),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_154),
.B(n_24),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_181),
.A2(n_189),
.B1(n_196),
.B2(n_166),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_123),
.C(n_138),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_193),
.C(n_195),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_171),
.A2(n_123),
.B1(n_88),
.B2(n_78),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_184),
.A2(n_145),
.B1(n_102),
.B2(n_23),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_185),
.B(n_23),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_155),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_146),
.B(n_24),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_158),
.A2(n_16),
.B(n_20),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_152),
.C(n_153),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_60),
.C(n_88),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_163),
.A2(n_78),
.B1(n_28),
.B2(n_32),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_159),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_213),
.C(n_217),
.Y(n_230)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_192),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_202),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_159),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_205),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_181),
.Y(n_202)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_204),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_151),
.Y(n_205)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_206),
.Y(n_224)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_184),
.Y(n_207)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_207),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_148),
.Y(n_208)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_208),
.Y(n_229)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_165),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_211),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_193),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_219),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_164),
.C(n_147),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_214),
.A2(n_216),
.B1(n_196),
.B2(n_187),
.Y(n_228)
);

INVxp67_ASAP7_75t_SL g215 ( 
.A(n_189),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_215),
.A2(n_218),
.B1(n_21),
.B2(n_22),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_172),
.B(n_60),
.C(n_102),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_174),
.B(n_23),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_22),
.C(n_21),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_176),
.C(n_182),
.Y(n_231)
);

AND2x2_ASAP7_75t_SL g225 ( 
.A(n_205),
.B(n_189),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_SL g255 ( 
.A1(n_225),
.A2(n_234),
.B(n_0),
.C(n_2),
.Y(n_255)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_22),
.C(n_1),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_201),
.A2(n_177),
.B1(n_179),
.B2(n_185),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_232),
.A2(n_220),
.B1(n_209),
.B2(n_199),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_210),
.A2(n_177),
.B1(n_173),
.B2(n_191),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_233),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_213),
.A2(n_22),
.B1(n_16),
.B2(n_2),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_235),
.A2(n_214),
.B1(n_217),
.B2(n_209),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_200),
.B(n_22),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_199),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_22),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_0),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_241),
.A2(n_252),
.B1(n_233),
.B2(n_222),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_229),
.B(n_197),
.Y(n_243)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_244),
.A2(n_246),
.B(n_247),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_16),
.Y(n_245)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_22),
.C(n_1),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_7),
.Y(n_249)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

FAx1_ASAP7_75t_SL g261 ( 
.A(n_250),
.B(n_236),
.CI(n_231),
.CON(n_261),
.SN(n_261)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_238),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_251),
.A2(n_254),
.B(n_239),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_237),
.A2(n_15),
.B1(n_7),
.B2(n_8),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_224),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_253),
.A2(n_256),
.B1(n_255),
.B2(n_225),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_6),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_255),
.A2(n_226),
.B(n_223),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_255),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_248),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_266),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_263),
.C(n_260),
.Y(n_272)
);

MAJx2_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_221),
.C(n_244),
.Y(n_276)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_262),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_255),
.A2(n_225),
.B(n_230),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_3),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_256),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_4),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_5),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_264),
.A2(n_246),
.B1(n_247),
.B2(n_221),
.Y(n_271)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_279),
.C(n_274),
.Y(n_282)
);

NOR2x1_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_239),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_273),
.A2(n_275),
.B(n_276),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_268),
.B(n_250),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_240),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_278),
.A2(n_280),
.B(n_261),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_265),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_288),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_282),
.A2(n_287),
.B(n_276),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_269),
.Y(n_283)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_283),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_286),
.B(n_9),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_278),
.A2(n_261),
.B(n_6),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_9),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_5),
.Y(n_290)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_290),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_292),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_270),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_295),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_9),
.Y(n_295)
);

NAND4xp25_ASAP7_75t_SL g299 ( 
.A(n_296),
.B(n_10),
.C(n_12),
.D(n_13),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_299),
.B(n_296),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_301),
.B(n_302),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_300),
.A2(n_284),
.B(n_293),
.Y(n_302)
);

OAI321xp33_ASAP7_75t_L g304 ( 
.A1(n_303),
.A2(n_298),
.A3(n_291),
.B1(n_297),
.B2(n_15),
.C(n_10),
.Y(n_304)
);

NOR3xp33_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_10),
.C(n_12),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_12),
.C(n_15),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_306),
.Y(n_307)
);


endmodule