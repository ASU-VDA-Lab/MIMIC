module fake_jpeg_26964_n_168 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_168);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_33),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_11),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_32),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_4),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_48),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_4),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

BUFx8_ASAP7_75t_L g70 ( 
.A(n_0),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_0),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx6_ASAP7_75t_SL g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_78),
.Y(n_90)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_1),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_55),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_82),
.A2(n_65),
.B1(n_63),
.B2(n_72),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_69),
.B1(n_71),
.B2(n_68),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_89),
.B1(n_92),
.B2(n_66),
.Y(n_98)
);

BUFx10_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_82),
.A2(n_50),
.B1(n_74),
.B2(n_67),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_81),
.A2(n_79),
.B1(n_78),
.B2(n_55),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_58),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_96),
.B(n_99),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_83),
.A2(n_58),
.B1(n_61),
.B2(n_66),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_103),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_98),
.A2(n_104),
.B(n_59),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_90),
.B(n_61),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_90),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_100),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_88),
.B(n_64),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_102),
.Y(n_109)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_64),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_86),
.A2(n_59),
.B1(n_73),
.B2(n_60),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_1),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_2),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_112),
.Y(n_128)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_108),
.Y(n_111)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_2),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_113),
.A2(n_95),
.B1(n_87),
.B2(n_6),
.Y(n_126)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_118),
.Y(n_130)
);

INVx3_ASAP7_75t_SL g119 ( 
.A(n_106),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_122),
.Y(n_133)
);

AND2x6_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_36),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_23),
.Y(n_134)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_117),
.A2(n_95),
.B1(n_57),
.B2(n_75),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_124),
.A2(n_131),
.B1(n_3),
.B2(n_5),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_126),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_62),
.C(n_56),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_132),
.C(n_3),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_52),
.B1(n_51),
.B2(n_28),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_25),
.C(n_47),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_17),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_133),
.A2(n_109),
.B1(n_110),
.B2(n_7),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_138),
.Y(n_154)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_136),
.B(n_139),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_124),
.A2(n_115),
.B1(n_5),
.B2(n_7),
.Y(n_137)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_137),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_128),
.A2(n_26),
.B(n_45),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_131),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_123),
.Y(n_140)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_125),
.A2(n_21),
.B(n_44),
.Y(n_141)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_142),
.B(n_144),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_146),
.C(n_147),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_127),
.A2(n_39),
.B(n_49),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_145),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_129),
.Y(n_147)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_154),
.B(n_135),
.C(n_146),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_157),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_132),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_150),
.A2(n_140),
.B1(n_143),
.B2(n_13),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_155),
.C(n_148),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_160),
.B(n_158),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_149),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_152),
.C(n_154),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_163),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_151),
.C(n_34),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_42),
.C(n_15),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_41),
.B(n_30),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_40),
.Y(n_168)
);


endmodule