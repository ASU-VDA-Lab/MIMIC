module fake_jpeg_2629_n_694 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_694);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_694;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_514;
wire n_651;
wire n_242;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx11_ASAP7_75t_SL g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_58),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_59),
.Y(n_138)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_60),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_61),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_62),
.Y(n_191)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_63),
.Y(n_147)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx5_ASAP7_75t_SL g160 ( 
.A(n_64),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_52),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_65),
.B(n_69),
.Y(n_139)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_66),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_25),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_67),
.B(n_71),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_68),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_57),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_70),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_25),
.B(n_36),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_72),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_57),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_73),
.B(n_90),
.Y(n_174)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_75),
.Y(n_165)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_76),
.Y(n_171)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_77),
.Y(n_144)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_78),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_79),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_0),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_80),
.B(n_3),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_81),
.Y(n_224)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_82),
.Y(n_172)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_83),
.Y(n_164)
);

BUFx12_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_84),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_85),
.Y(n_168)
);

BUFx12_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g201 ( 
.A(n_86),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

BUFx12_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx6_ASAP7_75t_SL g219 ( 
.A(n_88),
.Y(n_219)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_89),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_26),
.B(n_2),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_91),
.Y(n_175)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_92),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_57),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_93),
.B(n_96),
.Y(n_180)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_22),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_31),
.B(n_2),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_97),
.B(n_100),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_29),
.Y(n_98)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_98),
.Y(n_149)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_28),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_99),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_22),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_35),
.Y(n_101)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_103),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_32),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_104),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_46),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_105),
.B(n_116),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_32),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_106),
.Y(n_195)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_38),
.Y(n_107)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_107),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_41),
.Y(n_108)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_108),
.Y(n_177)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_38),
.Y(n_109)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_109),
.Y(n_229)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_38),
.Y(n_110)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_110),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_32),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_111),
.Y(n_231)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_35),
.Y(n_112)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_113),
.Y(n_179)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_36),
.Y(n_114)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_114),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_37),
.Y(n_115)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_39),
.B(n_2),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_46),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_117),
.B(n_120),
.Y(n_193)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_39),
.Y(n_118)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_118),
.Y(n_205)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_37),
.Y(n_119)
);

INVx3_ASAP7_75t_SL g141 ( 
.A(n_119),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_23),
.B(n_3),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_121),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_23),
.B(n_3),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_122),
.B(n_124),
.Y(n_197)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_40),
.Y(n_123)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_123),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_37),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_125),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_42),
.Y(n_126)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_42),
.Y(n_127)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_127),
.Y(n_199)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_40),
.Y(n_128)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_128),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_42),
.Y(n_129)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_129),
.Y(n_202)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_40),
.Y(n_130)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_130),
.Y(n_212)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_47),
.Y(n_131)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_131),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_47),
.Y(n_132)
);

INVx8_ASAP7_75t_L g233 ( 
.A(n_132),
.Y(n_233)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_134),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_66),
.B(n_60),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_137),
.B(n_158),
.Y(n_305)
);

BUFx8_ASAP7_75t_L g145 ( 
.A(n_64),
.Y(n_145)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_145),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_64),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_155),
.B(n_206),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_63),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_157),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_79),
.A2(n_85),
.B1(n_91),
.B2(n_104),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_161),
.A2(n_232),
.B1(n_137),
.B2(n_141),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_125),
.B(n_49),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_173),
.B(n_178),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_77),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_72),
.B(n_49),
.C(n_53),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_183),
.B(n_226),
.C(n_88),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_61),
.Y(n_185)
);

INVx4_ASAP7_75t_SL g323 ( 
.A(n_185),
.Y(n_323)
);

INVx11_ASAP7_75t_SL g186 ( 
.A(n_58),
.Y(n_186)
);

INVx6_ASAP7_75t_SL g306 ( 
.A(n_186),
.Y(n_306)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_58),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_188),
.Y(n_240)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_62),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_189),
.Y(n_272)
);

INVx11_ASAP7_75t_L g192 ( 
.A(n_68),
.Y(n_192)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_192),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_62),
.B(n_34),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_198),
.B(n_200),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_89),
.B(n_53),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_78),
.B(n_51),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_203),
.B(n_211),
.Y(n_311)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_113),
.Y(n_204)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_204),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_83),
.Y(n_206)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_121),
.Y(n_207)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_207),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_103),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_208),
.B(n_214),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_102),
.B(n_51),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_103),
.B(n_33),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_213),
.B(n_216),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_81),
.B(n_50),
.Y(n_214)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_87),
.Y(n_215)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_215),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_131),
.B(n_50),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_95),
.B(n_34),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_218),
.B(n_221),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_108),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_220),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_129),
.B(n_33),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_99),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_232),
.Y(n_255)
);

BUFx12_ASAP7_75t_L g225 ( 
.A(n_84),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_84),
.B(n_54),
.C(n_48),
.Y(n_226)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_106),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_228),
.Y(n_241)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_119),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_230),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_111),
.B(n_3),
.Y(n_232)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_145),
.Y(n_235)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_235),
.Y(n_332)
);

OA22x2_ASAP7_75t_L g236 ( 
.A1(n_161),
.A2(n_132),
.B1(n_127),
.B2(n_126),
.Y(n_236)
);

OA22x2_ASAP7_75t_L g345 ( 
.A1(n_236),
.A2(n_295),
.B1(n_195),
.B2(n_231),
.Y(n_345)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_156),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_237),
.Y(n_351)
);

OAI22xp33_ASAP7_75t_L g243 ( 
.A1(n_140),
.A2(n_115),
.B1(n_54),
.B2(n_48),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_243),
.A2(n_259),
.B1(n_279),
.B2(n_288),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_139),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_245),
.B(n_246),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_180),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_180),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_247),
.B(n_264),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_156),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_248),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_214),
.A2(n_54),
.B1(n_48),
.B2(n_47),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_251),
.Y(n_355)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_168),
.Y(n_252)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_252),
.Y(n_325)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_172),
.Y(n_253)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_253),
.Y(n_357)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_187),
.Y(n_254)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_254),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_143),
.B(n_4),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_256),
.B(n_265),
.Y(n_339)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_222),
.Y(n_257)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_257),
.Y(n_342)
);

INVx11_ASAP7_75t_L g258 ( 
.A(n_186),
.Y(n_258)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_258),
.Y(n_378)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_260),
.Y(n_347)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_163),
.Y(n_261)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_261),
.Y(n_341)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_209),
.Y(n_263)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_263),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_219),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_143),
.B(n_4),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_266),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_173),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_267),
.Y(n_366)
);

INVx8_ASAP7_75t_L g268 ( 
.A(n_168),
.Y(n_268)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_268),
.Y(n_344)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_141),
.Y(n_269)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_269),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_182),
.B(n_5),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_270),
.B(n_277),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_271),
.B(n_298),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_133),
.B(n_88),
.C(n_86),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_274),
.B(n_176),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_175),
.Y(n_275)
);

INVx8_ASAP7_75t_L g333 ( 
.A(n_275),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_182),
.B(n_6),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_227),
.Y(n_278)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_278),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_190),
.A2(n_86),
.B1(n_9),
.B2(n_10),
.Y(n_279)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_191),
.Y(n_280)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_280),
.Y(n_370)
);

OAI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_193),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_281),
.A2(n_304),
.B1(n_170),
.B2(n_195),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_200),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_282),
.B(n_284),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_157),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_193),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_285),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_218),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_286),
.A2(n_291),
.B1(n_293),
.B2(n_297),
.Y(n_327)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_169),
.Y(n_287)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_287),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_190),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_146),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_289),
.Y(n_336)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_152),
.Y(n_290)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_290),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_197),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_221),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_197),
.A2(n_16),
.B(n_17),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_294),
.A2(n_295),
.B(n_274),
.Y(n_372)
);

OA22x2_ASAP7_75t_L g295 ( 
.A1(n_202),
.A2(n_16),
.B1(n_18),
.B2(n_171),
.Y(n_295)
);

INVx11_ASAP7_75t_L g296 ( 
.A(n_160),
.Y(n_296)
);

BUFx8_ASAP7_75t_L g385 ( 
.A(n_296),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_203),
.A2(n_18),
.B1(n_211),
.B2(n_166),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_144),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_166),
.B(n_147),
.Y(n_299)
);

NAND2xp33_ASAP7_75t_SL g381 ( 
.A(n_299),
.B(n_300),
.Y(n_381)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_177),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_210),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_301),
.B(n_312),
.Y(n_361)
);

BUFx12f_ASAP7_75t_L g302 ( 
.A(n_160),
.Y(n_302)
);

INVx8_ASAP7_75t_L g387 ( 
.A(n_302),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_198),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_303),
.B(n_309),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_174),
.A2(n_213),
.B1(n_135),
.B2(n_205),
.Y(n_304)
);

INVx6_ASAP7_75t_L g307 ( 
.A(n_175),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_307),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_174),
.B(n_154),
.Y(n_309)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_148),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_159),
.A2(n_165),
.B1(n_164),
.B2(n_144),
.Y(n_313)
);

AO22x1_ASAP7_75t_L g388 ( 
.A1(n_313),
.A2(n_296),
.B1(n_236),
.B2(n_299),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_185),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_314),
.B(n_316),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_220),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_164),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_317),
.B(n_319),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_162),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_151),
.B(n_153),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_320),
.B(n_322),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_167),
.B(n_212),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_162),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_324),
.B(n_194),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_249),
.A2(n_181),
.B1(n_179),
.B2(n_149),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_328),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_255),
.B(n_196),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_330),
.B(n_346),
.Y(n_396)
);

OAI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_250),
.A2(n_292),
.B1(n_311),
.B2(n_294),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_338),
.A2(n_367),
.B1(n_313),
.B2(n_278),
.Y(n_424)
);

FAx1_ASAP7_75t_SL g343 ( 
.A(n_271),
.B(n_217),
.CI(n_184),
.CON(n_343),
.SN(n_343)
);

AOI32xp33_ASAP7_75t_L g435 ( 
.A1(n_343),
.A2(n_321),
.A3(n_310),
.B1(n_262),
.B2(n_276),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_345),
.B(n_388),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_311),
.B(n_176),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_349),
.B(n_369),
.C(n_323),
.Y(n_403)
);

O2A1O1Ixp33_ASAP7_75t_SL g350 ( 
.A1(n_295),
.A2(n_142),
.B(n_201),
.C(n_233),
.Y(n_350)
);

AO22x1_ASAP7_75t_L g412 ( 
.A1(n_350),
.A2(n_365),
.B1(n_386),
.B2(n_302),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_299),
.A2(n_138),
.B1(n_224),
.B2(n_136),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_356),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_292),
.B(n_231),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_362),
.B(n_275),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_364),
.B(n_375),
.Y(n_399)
);

O2A1O1Ixp33_ASAP7_75t_L g365 ( 
.A1(n_273),
.A2(n_142),
.B(n_201),
.C(n_225),
.Y(n_365)
);

OAI22xp33_ASAP7_75t_L g367 ( 
.A1(n_236),
.A2(n_194),
.B1(n_150),
.B2(n_199),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_318),
.A2(n_150),
.B(n_199),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_368),
.A2(n_372),
.B(n_379),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_305),
.B(n_233),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_306),
.Y(n_375)
);

INVxp33_ASAP7_75t_L g437 ( 
.A(n_376),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_238),
.A2(n_263),
.B(n_301),
.Y(n_379)
);

BUFx24_ASAP7_75t_SL g380 ( 
.A(n_302),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_380),
.B(n_382),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_240),
.B(n_272),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_312),
.B(n_316),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_384),
.B(n_323),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_236),
.A2(n_295),
.B1(n_243),
.B2(n_298),
.Y(n_386)
);

NAND3xp33_ASAP7_75t_L g389 ( 
.A(n_335),
.B(n_235),
.C(n_308),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_389),
.B(n_416),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_371),
.A2(n_317),
.B1(n_283),
.B2(n_307),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_390),
.A2(n_394),
.B1(n_407),
.B2(n_388),
.Y(n_447)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_385),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_392),
.B(n_409),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_371),
.A2(n_372),
.B1(n_358),
.B2(n_346),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_354),
.Y(n_395)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_395),
.Y(n_445)
);

INVx11_ASAP7_75t_L g397 ( 
.A(n_385),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_SL g441 ( 
.A1(n_397),
.A2(n_258),
.B1(n_387),
.B2(n_332),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_387),
.Y(n_398)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_398),
.Y(n_450)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_354),
.Y(n_401)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_401),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_403),
.B(n_347),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_379),
.B(n_266),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_404),
.B(n_411),
.Y(n_446)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_361),
.Y(n_405)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_405),
.Y(n_449)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_361),
.Y(n_406)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_406),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_358),
.A2(n_283),
.B1(n_237),
.B2(n_252),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_361),
.Y(n_408)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_408),
.Y(n_457)
);

INVx6_ASAP7_75t_L g410 ( 
.A(n_351),
.Y(n_410)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_410),
.Y(n_442)
);

CKINVDCx12_ASAP7_75t_R g411 ( 
.A(n_385),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_412),
.B(n_434),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_340),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_413),
.B(n_422),
.Y(n_460)
);

INVx6_ASAP7_75t_L g414 ( 
.A(n_351),
.Y(n_414)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_414),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_415),
.B(n_421),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_348),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_358),
.B(n_257),
.C(n_260),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_417),
.B(n_429),
.C(n_374),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_381),
.B(n_283),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_418),
.B(n_435),
.Y(n_439)
);

AND2x6_ASAP7_75t_L g419 ( 
.A(n_343),
.B(n_306),
.Y(n_419)
);

AND2x6_ASAP7_75t_L g443 ( 
.A(n_419),
.B(n_428),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_352),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_420),
.B(n_359),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_362),
.B(n_254),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_326),
.B(n_334),
.Y(n_422)
);

BUFx5_ASAP7_75t_L g423 ( 
.A(n_365),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_423),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_424),
.A2(n_355),
.B1(n_345),
.B2(n_366),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_331),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_425),
.B(n_426),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_330),
.B(n_253),
.Y(n_426)
);

AND2x6_ASAP7_75t_L g428 ( 
.A(n_343),
.B(n_244),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_349),
.B(n_276),
.C(n_315),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_369),
.B(n_287),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_430),
.B(n_345),
.Y(n_469)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_360),
.Y(n_431)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_431),
.Y(n_470)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_377),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_432),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_374),
.Y(n_433)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_433),
.Y(n_478)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_360),
.Y(n_434)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_337),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_436),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_SL g438 ( 
.A1(n_355),
.A2(n_290),
.B1(n_289),
.B2(n_300),
.Y(n_438)
);

OAI21xp33_ASAP7_75t_SL g481 ( 
.A1(n_438),
.A2(n_315),
.B(n_341),
.Y(n_481)
);

AOI22xp33_ASAP7_75t_L g440 ( 
.A1(n_399),
.A2(n_345),
.B1(n_367),
.B2(n_350),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_440),
.A2(n_370),
.B1(n_341),
.B2(n_377),
.Y(n_523)
);

OAI21xp33_ASAP7_75t_SL g483 ( 
.A1(n_441),
.A2(n_469),
.B(n_471),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_444),
.B(n_458),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_447),
.B(n_461),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_391),
.A2(n_386),
.B1(n_388),
.B2(n_368),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_453),
.A2(n_465),
.B1(n_434),
.B2(n_431),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_454),
.A2(n_464),
.B1(n_475),
.B2(n_412),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_427),
.A2(n_383),
.B(n_327),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_455),
.A2(n_476),
.B(n_427),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_403),
.B(n_339),
.Y(n_458)
);

OAI32xp33_ASAP7_75t_L g459 ( 
.A1(n_396),
.A2(n_383),
.A3(n_366),
.B1(n_339),
.B2(n_329),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_459),
.B(n_480),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_391),
.A2(n_424),
.B1(n_396),
.B2(n_430),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_391),
.A2(n_394),
.B1(n_390),
.B2(n_412),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_425),
.A2(n_350),
.B1(n_363),
.B2(n_344),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_472),
.B(n_477),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g474 ( 
.A(n_435),
.B(n_337),
.Y(n_474)
);

NAND3xp33_ASAP7_75t_L g501 ( 
.A(n_474),
.B(n_417),
.C(n_418),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_416),
.A2(n_363),
.B1(n_344),
.B2(n_325),
.Y(n_475)
);

AOI22x1_ASAP7_75t_SL g476 ( 
.A1(n_419),
.A2(n_321),
.B1(n_310),
.B2(n_262),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_420),
.B(n_336),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_421),
.B(n_342),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_481),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_429),
.B(n_342),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_482),
.B(n_359),
.Y(n_519)
);

OAI22xp33_ASAP7_75t_SL g542 ( 
.A1(n_484),
.A2(n_450),
.B1(n_446),
.B2(n_462),
.Y(n_542)
);

INVx13_ASAP7_75t_L g486 ( 
.A(n_466),
.Y(n_486)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_486),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_487),
.A2(n_489),
.B(n_490),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_474),
.A2(n_428),
.B(n_400),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_468),
.A2(n_402),
.B(n_437),
.Y(n_490)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_445),
.Y(n_492)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_492),
.Y(n_527)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_445),
.Y(n_493)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_493),
.Y(n_531)
);

AND2x2_ASAP7_75t_SL g494 ( 
.A(n_464),
.B(n_418),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_494),
.Y(n_562)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_448),
.Y(n_495)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_495),
.Y(n_536)
);

CKINVDCx12_ASAP7_75t_R g496 ( 
.A(n_456),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_496),
.Y(n_528)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_448),
.Y(n_497)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_497),
.Y(n_546)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_470),
.Y(n_498)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_498),
.Y(n_550)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_470),
.Y(n_499)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_499),
.Y(n_552)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_480),
.Y(n_500)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_500),
.Y(n_553)
);

NAND3xp33_ASAP7_75t_L g537 ( 
.A(n_501),
.B(n_467),
.C(n_473),
.Y(n_537)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_479),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_502),
.B(n_503),
.Y(n_547)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_479),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_442),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_504),
.B(n_510),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_463),
.A2(n_402),
.B(n_423),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_505),
.A2(n_506),
.B(n_509),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_468),
.A2(n_405),
.B(n_406),
.Y(n_506)
);

AOI32xp33_ASAP7_75t_L g508 ( 
.A1(n_439),
.A2(n_415),
.A3(n_408),
.B1(n_407),
.B2(n_401),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_508),
.B(n_515),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_455),
.A2(n_395),
.B(n_432),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_466),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_451),
.B(n_436),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_511),
.Y(n_534)
);

INVx13_ASAP7_75t_L g512 ( 
.A(n_450),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_512),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_514),
.A2(n_523),
.B1(n_447),
.B2(n_452),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_451),
.B(n_398),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_449),
.B(n_414),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_516),
.B(n_517),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_449),
.B(n_457),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_478),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_518),
.B(n_520),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_519),
.B(n_347),
.Y(n_554)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_478),
.Y(n_520)
);

AND2x6_ASAP7_75t_L g521 ( 
.A(n_443),
.B(n_393),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_521),
.B(n_460),
.Y(n_543)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_452),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_SL g525 ( 
.A1(n_522),
.A2(n_469),
.B1(n_397),
.B2(n_463),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_484),
.A2(n_465),
.B1(n_453),
.B2(n_468),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_524),
.A2(n_525),
.B1(n_529),
.B2(n_533),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_507),
.B(n_461),
.C(n_444),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_532),
.B(n_535),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_500),
.A2(n_476),
.B1(n_457),
.B2(n_443),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_485),
.B(n_482),
.C(n_458),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_537),
.B(n_554),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_514),
.A2(n_439),
.B1(n_459),
.B2(n_462),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_539),
.A2(n_555),
.B1(n_494),
.B2(n_505),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_542),
.A2(n_513),
.B1(n_510),
.B2(n_502),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_543),
.B(n_548),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_491),
.B(n_336),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_491),
.B(n_373),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_549),
.B(n_558),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_509),
.A2(n_370),
.B(n_442),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_551),
.A2(n_489),
.B(n_517),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_483),
.A2(n_353),
.B1(n_325),
.B2(n_333),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_487),
.A2(n_373),
.B(n_378),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g584 ( 
.A(n_556),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_485),
.B(n_357),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_557),
.B(n_561),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_488),
.B(n_357),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_488),
.B(n_410),
.Y(n_560)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_560),
.Y(n_564)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_485),
.B(n_241),
.Y(n_561)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_547),
.Y(n_565)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_565),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_530),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_566),
.B(n_576),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_532),
.B(n_506),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g606 ( 
.A(n_569),
.B(n_589),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_570),
.A2(n_580),
.B1(n_591),
.B2(n_593),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_524),
.A2(n_523),
.B1(n_511),
.B2(n_515),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g599 ( 
.A1(n_571),
.A2(n_581),
.B1(n_582),
.B2(n_529),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_535),
.B(n_494),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g601 ( 
.A(n_572),
.B(n_577),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_SL g596 ( 
.A1(n_573),
.A2(n_551),
.B1(n_555),
.B2(n_556),
.Y(n_596)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_547),
.Y(n_574)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_574),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_530),
.Y(n_576)
);

XOR2xp5_ASAP7_75t_L g577 ( 
.A(n_557),
.B(n_508),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_530),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_578),
.B(n_585),
.Y(n_612)
);

XNOR2x1_ASAP7_75t_SL g579 ( 
.A(n_538),
.B(n_490),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_579),
.B(n_583),
.Y(n_602)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_541),
.Y(n_580)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_553),
.B(n_503),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_SL g583 ( 
.A(n_539),
.B(n_521),
.Y(n_583)
);

AOI21xp5_ASAP7_75t_L g585 ( 
.A1(n_544),
.A2(n_522),
.B(n_520),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_SL g587 ( 
.A(n_554),
.B(n_516),
.Y(n_587)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_587),
.B(n_492),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_534),
.B(n_518),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_559),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_SL g617 ( 
.A(n_590),
.B(n_495),
.Y(n_617)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_559),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_561),
.B(n_497),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g610 ( 
.A(n_592),
.B(n_594),
.Y(n_610)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_527),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_534),
.B(n_553),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_567),
.B(n_562),
.C(n_526),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_595),
.B(n_600),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_SL g627 ( 
.A1(n_596),
.A2(n_584),
.B1(n_589),
.B2(n_594),
.Y(n_627)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_599),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_567),
.B(n_562),
.C(n_526),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_569),
.B(n_533),
.C(n_544),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g637 ( 
.A(n_603),
.B(n_604),
.C(n_607),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_572),
.B(n_528),
.C(n_550),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_L g605 ( 
.A1(n_580),
.A2(n_528),
.B1(n_550),
.B2(n_546),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g635 ( 
.A1(n_605),
.A2(n_613),
.B1(n_615),
.B2(n_582),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_563),
.B(n_552),
.C(n_546),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_563),
.B(n_552),
.C(n_536),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_608),
.B(n_587),
.C(n_593),
.Y(n_642)
);

XOR2xp5_ASAP7_75t_L g631 ( 
.A(n_609),
.B(n_611),
.Y(n_631)
);

XOR2xp5_ASAP7_75t_L g611 ( 
.A(n_577),
.B(n_527),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_575),
.A2(n_531),
.B1(n_536),
.B2(n_545),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g614 ( 
.A(n_579),
.B(n_531),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_614),
.B(n_620),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_564),
.A2(n_540),
.B1(n_499),
.B2(n_493),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_617),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_SL g619 ( 
.A1(n_571),
.A2(n_498),
.B1(n_540),
.B2(n_545),
.Y(n_619)
);

INVxp67_ASAP7_75t_L g623 ( 
.A(n_619),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g620 ( 
.A(n_573),
.B(n_504),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_SL g621 ( 
.A(n_603),
.B(n_595),
.C(n_600),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g648 ( 
.A(n_621),
.B(n_636),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_618),
.A2(n_568),
.B1(n_570),
.B2(n_591),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_624),
.A2(n_635),
.B1(n_620),
.B2(n_610),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_SL g626 ( 
.A(n_614),
.B(n_588),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_626),
.B(n_628),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_627),
.B(n_610),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_SL g628 ( 
.A(n_604),
.B(n_586),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_597),
.Y(n_629)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_629),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_SL g632 ( 
.A(n_606),
.B(n_583),
.C(n_592),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_632),
.B(n_634),
.Y(n_647)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_598),
.Y(n_633)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_633),
.Y(n_657)
);

CKINVDCx16_ASAP7_75t_R g634 ( 
.A(n_612),
.Y(n_634)
);

XNOR2xp5_ASAP7_75t_L g636 ( 
.A(n_611),
.B(n_606),
.Y(n_636)
);

XNOR2x1_ASAP7_75t_SL g638 ( 
.A(n_602),
.B(n_578),
.Y(n_638)
);

XNOR2xp5_ASAP7_75t_L g650 ( 
.A(n_638),
.B(n_639),
.Y(n_650)
);

XNOR2xp5_ASAP7_75t_L g639 ( 
.A(n_607),
.B(n_581),
.Y(n_639)
);

OAI21xp5_ASAP7_75t_SL g640 ( 
.A1(n_616),
.A2(n_585),
.B(n_584),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_640),
.A2(n_601),
.B(n_486),
.Y(n_652)
);

XNOR2xp5_ASAP7_75t_L g651 ( 
.A(n_642),
.B(n_609),
.Y(n_651)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_644),
.Y(n_663)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_637),
.B(n_608),
.C(n_601),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_645),
.B(n_649),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_SL g664 ( 
.A1(n_646),
.A2(n_630),
.B1(n_638),
.B2(n_625),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_641),
.B(n_602),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_651),
.B(n_654),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_652),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_642),
.B(n_333),
.Y(n_653)
);

NOR2xp67_ASAP7_75t_L g666 ( 
.A(n_653),
.B(n_625),
.Y(n_666)
);

CKINVDCx16_ASAP7_75t_R g654 ( 
.A(n_627),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_637),
.B(n_512),
.C(n_353),
.Y(n_655)
);

MAJIxp5_ASAP7_75t_L g671 ( 
.A(n_655),
.B(n_658),
.C(n_631),
.Y(n_671)
);

MAJIxp5_ASAP7_75t_L g658 ( 
.A(n_621),
.B(n_378),
.C(n_248),
.Y(n_658)
);

CKINVDCx16_ASAP7_75t_R g659 ( 
.A(n_624),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_659),
.B(n_623),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g672 ( 
.A(n_661),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_643),
.A2(n_622),
.B1(n_623),
.B2(n_639),
.Y(n_662)
);

XOR2xp5_ASAP7_75t_L g675 ( 
.A(n_662),
.B(n_670),
.Y(n_675)
);

XNOR2xp5_ASAP7_75t_L g676 ( 
.A(n_664),
.B(n_666),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_648),
.B(n_640),
.Y(n_668)
);

NOR2xp67_ASAP7_75t_L g678 ( 
.A(n_668),
.B(n_669),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_656),
.B(n_636),
.Y(n_669)
);

XOR2xp5_ASAP7_75t_L g670 ( 
.A(n_650),
.B(n_631),
.Y(n_670)
);

XOR2xp5_ASAP7_75t_L g677 ( 
.A(n_671),
.B(n_658),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_SL g673 ( 
.A1(n_667),
.A2(n_647),
.B(n_646),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_673),
.B(n_674),
.Y(n_683)
);

MAJIxp5_ASAP7_75t_L g674 ( 
.A(n_663),
.B(n_645),
.C(n_648),
.Y(n_674)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_677),
.Y(n_681)
);

MAJIxp5_ASAP7_75t_L g679 ( 
.A(n_671),
.B(n_651),
.C(n_644),
.Y(n_679)
);

XNOR2xp5_ASAP7_75t_L g682 ( 
.A(n_679),
.B(n_664),
.Y(n_682)
);

XNOR2xp5_ASAP7_75t_L g680 ( 
.A(n_679),
.B(n_669),
.Y(n_680)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_680),
.A2(n_682),
.B(n_677),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_672),
.B(n_665),
.Y(n_684)
);

OAI21x1_ASAP7_75t_L g685 ( 
.A1(n_684),
.A2(n_678),
.B(n_657),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_685),
.A2(n_686),
.B(n_687),
.Y(n_688)
);

OAI21xp5_ASAP7_75t_L g687 ( 
.A1(n_683),
.A2(n_676),
.B(n_674),
.Y(n_687)
);

AOI322xp5_ASAP7_75t_L g689 ( 
.A1(n_687),
.A2(n_681),
.A3(n_660),
.B1(n_680),
.B2(n_662),
.C1(n_675),
.C2(n_650),
.Y(n_689)
);

OAI21x1_ASAP7_75t_L g690 ( 
.A1(n_689),
.A2(n_675),
.B(n_670),
.Y(n_690)
);

AOI322xp5_ASAP7_75t_L g691 ( 
.A1(n_690),
.A2(n_688),
.A3(n_655),
.B1(n_244),
.B2(n_280),
.C1(n_261),
.C2(n_268),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_691),
.A2(n_239),
.B1(n_242),
.B2(n_241),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_692),
.B(n_239),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g694 ( 
.A1(n_693),
.A2(n_242),
.B(n_269),
.Y(n_694)
);


endmodule