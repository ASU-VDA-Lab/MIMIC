module real_jpeg_2685_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx2_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_1),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_1),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_1),
.B(n_55),
.Y(n_65)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_1),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_1),
.B(n_44),
.Y(n_178)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_2),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_2),
.B(n_75),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_2),
.B(n_30),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_2),
.B(n_44),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_2),
.B(n_27),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_2),
.B(n_90),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_3),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_4),
.B(n_75),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_4),
.B(n_33),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_4),
.B(n_39),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_4),
.B(n_55),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_4),
.B(n_30),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_4),
.B(n_27),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_4),
.B(n_44),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_4),
.B(n_90),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_5),
.B(n_33),
.Y(n_161)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_5),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_5),
.B(n_39),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_5),
.B(n_55),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_5),
.B(n_30),
.Y(n_263)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_7),
.Y(n_76)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_10),
.B(n_30),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_10),
.B(n_27),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_10),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_10),
.B(n_55),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_10),
.B(n_39),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_10),
.B(n_44),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_10),
.B(n_90),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_11),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_11),
.B(n_30),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_11),
.B(n_39),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_11),
.B(n_44),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_11),
.B(n_27),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_11),
.B(n_90),
.Y(n_163)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_12),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_12),
.B(n_39),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_12),
.B(n_33),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_12),
.B(n_55),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_12),
.B(n_30),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_12),
.B(n_27),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_14),
.B(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_14),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_14),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_14),
.B(n_75),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_14),
.B(n_55),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_14),
.B(n_39),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_152),
.B1(n_347),
.B2(n_348),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g347 ( 
.A(n_18),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_151),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_123),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_21),
.B(n_123),
.Y(n_151)
);

BUFx24_ASAP7_75t_SL g354 ( 
.A(n_21),
.Y(n_354)
);

FAx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_58),
.CI(n_93),
.CON(n_21),
.SN(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_35),
.B1(n_56),
.B2(n_57),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_23),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_32),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_SL g36 ( 
.A(n_25),
.B(n_37),
.C(n_42),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_25),
.A2(n_26),
.B1(n_42),
.B2(n_43),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_25),
.A2(n_26),
.B1(n_187),
.B2(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_26),
.B(n_187),
.C(n_188),
.Y(n_186)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_27),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_28),
.A2(n_29),
.B1(n_66),
.B2(n_96),
.Y(n_169)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_29),
.B(n_66),
.C(n_167),
.Y(n_206)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_30),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_47),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_37),
.A2(n_38),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_39),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_42),
.A2(n_43),
.B1(n_89),
.B2(n_102),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_42),
.A2(n_43),
.B1(n_148),
.B2(n_227),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_43),
.B(n_87),
.C(n_89),
.Y(n_86)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_45),
.B(n_145),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.C(n_53),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_48),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_49),
.B(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_51),
.A2(n_52),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_52),
.B(n_134),
.C(n_135),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g174 ( 
.A(n_55),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_72),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_64),
.C(n_68),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_60),
.A2(n_61),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_64),
.B(n_68),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.C(n_67),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_65),
.B(n_67),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_84),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_77),
.B1(n_82),
.B2(n_83),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_74),
.Y(n_82)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_75),
.Y(n_146)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_78),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_79),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_79),
.B(n_116),
.C(n_118),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_79),
.A2(n_80),
.B1(n_116),
.B2(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_91),
.C(n_92),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_85),
.A2(n_86),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_101),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_89),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_89),
.A2(n_102),
.B1(n_244),
.B2(n_245),
.Y(n_257)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_90),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_91),
.A2(n_92),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_92),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_115),
.C(n_121),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_92),
.A2(n_112),
.B1(n_121),
.B2(n_122),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_109),
.C(n_114),
.Y(n_93)
);

FAx1_ASAP7_75t_SL g124 ( 
.A(n_94),
.B(n_109),
.CI(n_114),
.CON(n_124),
.SN(n_124)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.C(n_105),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_95),
.B(n_99),
.Y(n_333)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_102),
.B(n_103),
.C(n_104),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_100),
.B(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_100),
.A2(n_101),
.B1(n_183),
.B2(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_102),
.B(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_103),
.B(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_104),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_104),
.A2(n_159),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_105),
.B(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_140),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_117),
.B(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_117),
.B(n_209),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_120),
.B(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_120),
.B(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.C(n_128),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_124),
.B(n_125),
.Y(n_335)
);

BUFx24_ASAP7_75t_SL g353 ( 
.A(n_124),
.Y(n_353)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_126),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_128),
.B(n_335),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_139),
.C(n_141),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_129),
.A2(n_130),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.C(n_136),
.Y(n_130)
);

FAx1_ASAP7_75t_SL g309 ( 
.A(n_131),
.B(n_133),
.CI(n_136),
.CON(n_309),
.SN(n_309)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_134),
.A2(n_135),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_134),
.Y(n_217)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_135),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_139),
.B(n_141),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_149),
.C(n_150),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_142),
.A2(n_143),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.C(n_148),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_144),
.B(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_147),
.A2(n_148),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_147),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_148),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_149),
.A2(n_150),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_149),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_150),
.Y(n_321)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_152),
.Y(n_348)
);

OAI31xp33_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_323),
.A3(n_336),
.B(n_341),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_303),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_228),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_200),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_156),
.B(n_200),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_170),
.C(n_190),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_157),
.B(n_300),
.Y(n_299)
);

BUFx24_ASAP7_75t_SL g349 ( 
.A(n_157),
.Y(n_349)
);

FAx1_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_162),
.CI(n_166),
.CON(n_157),
.SN(n_157)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_158),
.B(n_162),
.C(n_166),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.C(n_161),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_160),
.B(n_161),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B(n_165),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_164),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_165),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_165),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_168),
.B(n_184),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_168),
.B(n_211),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_170),
.B(n_190),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_180),
.B2(n_189),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_181),
.C(n_186),
.Y(n_202)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_173),
.B(n_177),
.C(n_179),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_176),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_185),
.B2(n_186),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_183),
.Y(n_199)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_187),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_192),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.C(n_198),
.Y(n_190)
);

FAx1_ASAP7_75t_SL g290 ( 
.A(n_191),
.B(n_194),
.CI(n_198),
.CON(n_290),
.SN(n_290)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.C(n_197),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_195),
.B(n_197),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_196),
.B(n_239),
.Y(n_238)
);

BUFx24_ASAP7_75t_SL g352 ( 
.A(n_200),
.Y(n_352)
);

FAx1_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_218),
.CI(n_219),
.CON(n_200),
.SN(n_200)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_201),
.B(n_218),
.C(n_219),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_202),
.B(n_205),
.C(n_212),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_212),
.B2(n_213),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_206),
.B(n_208),
.C(n_210),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_224),
.Y(n_219)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_221),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_221),
.B(n_222),
.C(n_224),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_298),
.B(n_302),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_286),
.B(n_297),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_258),
.B(n_285),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_249),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_232),
.B(n_249),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_242),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_238),
.B1(n_240),
.B2(n_241),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_234),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.C(n_237),
.Y(n_234)
);

FAx1_ASAP7_75t_SL g250 ( 
.A(n_235),
.B(n_236),
.CI(n_237),
.CON(n_250),
.SN(n_250)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_238),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_238),
.B(n_240),
.C(n_242),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_243),
.B(n_247),
.C(n_248),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.C(n_257),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_250),
.B(n_282),
.Y(n_281)
);

BUFx24_ASAP7_75t_SL g355 ( 
.A(n_250),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_251),
.A2(n_252),
.B1(n_257),
.B2(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_253),
.A2(n_254),
.B1(n_255),
.B2(n_256),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_279),
.B(n_284),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_270),
.B(n_278),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_266),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_266),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_264),
.C(n_265),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_267),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_273),
.B(n_277),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_275),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_281),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_287),
.B(n_288),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_291),
.B2(n_292),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_293),
.C(n_294),
.Y(n_301)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

BUFx24_ASAP7_75t_SL g356 ( 
.A(n_290),
.Y(n_356)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_301),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_301),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_304),
.A2(n_343),
.B(n_344),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_322),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_305),
.B(n_322),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_306),
.B(n_308),
.C(n_311),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

BUFx24_ASAP7_75t_SL g351 ( 
.A(n_309),
.Y(n_351)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_312),
.B(n_316),
.C(n_317),
.Y(n_330)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVxp33_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g341 ( 
.A1(n_324),
.A2(n_337),
.B(n_342),
.C(n_345),
.D(n_346),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_334),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_325),
.B(n_334),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_330),
.C(n_331),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_326),
.A2(n_327),
.B1(n_331),
.B2(n_332),
.Y(n_339)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_330),
.B(n_339),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_338),
.B(n_340),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_338),
.B(n_340),
.Y(n_345)
);


endmodule