module fake_jpeg_4667_n_326 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_8),
.B(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_21),
.Y(n_42)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_46),
.B(n_47),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_56),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_29),
.B(n_0),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_52),
.B(n_59),
.Y(n_97)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_54),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_19),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_60),
.Y(n_76)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_64),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_2),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_22),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_61),
.B(n_62),
.Y(n_108)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_20),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_17),
.B(n_3),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_36),
.B1(n_40),
.B2(n_39),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_65),
.A2(n_70),
.B(n_78),
.Y(n_120)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_36),
.B1(n_40),
.B2(n_39),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_71),
.B(n_74),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_23),
.B1(n_33),
.B2(n_31),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_72),
.A2(n_85),
.B1(n_89),
.B2(n_99),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_73),
.B(n_86),
.Y(n_142)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_84),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_36),
.B1(n_41),
.B2(n_22),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_56),
.A2(n_23),
.B1(n_33),
.B2(n_31),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_83),
.A2(n_95),
.B1(n_102),
.B2(n_28),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_55),
.C(n_61),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_60),
.A2(n_25),
.B1(n_41),
.B2(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_25),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_58),
.A2(n_17),
.B1(n_34),
.B2(n_32),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_56),
.A2(n_34),
.B1(n_32),
.B2(n_24),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_92),
.A2(n_101),
.B1(n_30),
.B2(n_26),
.Y(n_117)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_94),
.Y(n_119)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_62),
.A2(n_27),
.B1(n_24),
.B2(n_35),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

NOR2x1_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_27),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_98),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_51),
.A2(n_30),
.B1(n_26),
.B2(n_35),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_51),
.A2(n_35),
.B1(n_30),
.B2(n_26),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_57),
.A2(n_35),
.B1(n_30),
.B2(n_26),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_106),
.Y(n_129)
);

CKINVDCx6p67_ASAP7_75t_R g104 ( 
.A(n_44),
.Y(n_104)
);

BUFx4f_ASAP7_75t_SL g139 ( 
.A(n_104),
.Y(n_139)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_4),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_45),
.B(n_28),
.Y(n_109)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_42),
.Y(n_110)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_110),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_111),
.A2(n_122),
.B1(n_91),
.B2(n_87),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_112),
.B(n_6),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_117),
.A2(n_145),
.B1(n_122),
.B2(n_146),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_67),
.B(n_76),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_118),
.A2(n_83),
.B(n_95),
.Y(n_158)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_123),
.Y(n_150)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_108),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_124),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_88),
.A2(n_93),
.B1(n_107),
.B2(n_100),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_125),
.Y(n_169)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_128),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_20),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_127),
.B(n_137),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_68),
.Y(n_128)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_138),
.Y(n_157)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

AND2x2_ASAP7_75t_SL g134 ( 
.A(n_69),
.B(n_20),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_143),
.Y(n_167)
);

OA22x2_ASAP7_75t_L g136 ( 
.A1(n_102),
.A2(n_70),
.B1(n_65),
.B2(n_78),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_136),
.A2(n_145),
.B1(n_6),
.B2(n_8),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_20),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_20),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_77),
.Y(n_171)
);

AND2x2_ASAP7_75t_SL g143 ( 
.A(n_79),
.B(n_4),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g145 ( 
.A1(n_90),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_87),
.Y(n_159)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_151),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_90),
.B1(n_84),
.B2(n_81),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_148),
.A2(n_113),
.B1(n_16),
.B2(n_15),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_153),
.B(n_155),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_141),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_119),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_156),
.B(n_160),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_158),
.A2(n_120),
.B(n_145),
.Y(n_188)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

AND2x6_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_127),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_161),
.B(n_175),
.C(n_177),
.Y(n_209)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_114),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_162),
.B(n_172),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_91),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_143),
.Y(n_184)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_120),
.A2(n_82),
.B(n_80),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_116),
.B(n_145),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_80),
.Y(n_168)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_170),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_174),
.Y(n_185)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

AND2x6_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_77),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_176),
.A2(n_180),
.B1(n_123),
.B2(n_130),
.Y(n_207)
);

AND2x6_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_82),
.Y(n_177)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_178),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_135),
.B(n_9),
.Y(n_179)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_124),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_142),
.B(n_10),
.Y(n_182)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_184),
.A2(n_195),
.B(n_196),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_188),
.A2(n_190),
.B(n_211),
.Y(n_221)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_189),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_144),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_193),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_132),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_161),
.A2(n_126),
.B(n_121),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_158),
.A2(n_138),
.B(n_112),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_166),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_197),
.B(n_199),
.Y(n_240)
);

NOR3xp33_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_133),
.C(n_12),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_157),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_203),
.Y(n_230)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_152),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_206),
.B(n_208),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_207),
.A2(n_169),
.B1(n_156),
.B2(n_163),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_117),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_166),
.B(n_115),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_210),
.B(n_213),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_165),
.A2(n_113),
.B(n_12),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_150),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_214),
.A2(n_176),
.B1(n_167),
.B2(n_169),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_151),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_172),
.C(n_174),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_220),
.C(n_190),
.Y(n_242)
);

MAJx2_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_185),
.C(n_210),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_217),
.B(n_240),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_175),
.C(n_148),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_222),
.A2(n_231),
.B1(n_232),
.B2(n_236),
.Y(n_249)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

INVx13_ASAP7_75t_L g252 ( 
.A(n_224),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_226),
.A2(n_184),
.B1(n_214),
.B2(n_201),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_189),
.B(n_167),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_231),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_194),
.Y(n_228)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_192),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_188),
.A2(n_167),
.B1(n_163),
.B2(n_162),
.Y(n_231)
);

A2O1A1Ixp33_ASAP7_75t_SL g232 ( 
.A1(n_211),
.A2(n_196),
.B(n_186),
.C(n_184),
.Y(n_232)
);

FAx1_ASAP7_75t_L g234 ( 
.A(n_195),
.B(n_153),
.CI(n_154),
.CON(n_234),
.SN(n_234)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_234),
.A2(n_221),
.B(n_240),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_212),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_235),
.B(n_238),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_208),
.A2(n_155),
.B1(n_160),
.B2(n_154),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_205),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_239),
.B(n_241),
.Y(n_258)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_205),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_246),
.C(n_251),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_260),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_191),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_246),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_250),
.A2(n_257),
.B1(n_262),
.B2(n_232),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_216),
.B(n_201),
.C(n_193),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_253),
.B(n_254),
.Y(n_264)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_207),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_256),
.C(n_261),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_192),
.C(n_213),
.Y(n_256)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_259),
.B(n_218),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_219),
.B(n_215),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_220),
.A2(n_183),
.B1(n_184),
.B2(n_199),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_276),
.Y(n_286)
);

AOI321xp33_ASAP7_75t_L g282 ( 
.A1(n_265),
.A2(n_258),
.A3(n_252),
.B1(n_248),
.B2(n_245),
.C(n_198),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_269),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_249),
.A2(n_233),
.B1(n_234),
.B2(n_217),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_268),
.A2(n_278),
.B1(n_279),
.B2(n_187),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_221),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_262),
.A2(n_232),
.B1(n_236),
.B2(n_222),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_271),
.A2(n_272),
.B1(n_248),
.B2(n_252),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_257),
.A2(n_232),
.B1(n_230),
.B2(n_234),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_244),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_277),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_250),
.B(n_233),
.Y(n_275)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_275),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_251),
.B(n_204),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_256),
.A2(n_206),
.B1(n_203),
.B2(n_229),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_255),
.A2(n_186),
.B(n_198),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_242),
.C(n_261),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_288),
.C(n_289),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_260),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_282),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_278),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_283),
.A2(n_279),
.B(n_275),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_284),
.A2(n_164),
.B1(n_170),
.B2(n_147),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_200),
.C(n_202),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_200),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_291),
.B(n_264),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_267),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_292),
.Y(n_296)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_293),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_283),
.A2(n_273),
.B(n_263),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_298),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_295),
.B(n_300),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_290),
.A2(n_268),
.B(n_269),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_187),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_299),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_286),
.B(n_204),
.Y(n_300)
);

AND2x2_ASAP7_75t_SL g302 ( 
.A(n_285),
.B(n_202),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_289),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_288),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_304),
.A2(n_302),
.B(n_301),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_178),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_311),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_285),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_281),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_312),
.B(n_314),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_317),
.Y(n_320)
);

MAJx2_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_280),
.C(n_297),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_301),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_316),
.A2(n_315),
.B1(n_307),
.B2(n_304),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_10),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_319),
.B(n_15),
.C(n_10),
.Y(n_322)
);

OAI21xp33_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_305),
.B(n_316),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_322),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_323),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_318),
.C(n_13),
.Y(n_325)
);

FAx1_ASAP7_75t_SL g326 ( 
.A(n_325),
.B(n_13),
.CI(n_15),
.CON(n_326),
.SN(n_326)
);


endmodule