module fake_netlist_6_5_n_1697 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1697);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1697;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_114),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_124),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_38),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_148),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_113),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_69),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_28),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_83),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_81),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_40),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_34),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_121),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_25),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_49),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_88),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_2),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_12),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_57),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_98),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_87),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_105),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_144),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_2),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_36),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_120),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_89),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_139),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_47),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_59),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_30),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_46),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_44),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_127),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_99),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_104),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_50),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_143),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_61),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_29),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_85),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_115),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_149),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_147),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_80),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_106),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_53),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_26),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_141),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_117),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_91),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_153),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_31),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_46),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_29),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_67),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_95),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_30),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_94),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_78),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_116),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_150),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_100),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_72),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_23),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_71),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_65),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_92),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_11),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_138),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_109),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_35),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_23),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_44),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_20),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_101),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_0),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_103),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_54),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_1),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_129),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_9),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_108),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_41),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_20),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_22),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_0),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_22),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_140),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_34),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_16),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_41),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_6),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_58),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_40),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_68),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_5),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_9),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_38),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_76),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_135),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_17),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_90),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_50),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_28),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_56),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_74),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_39),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_96),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_51),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_154),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_77),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_36),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_152),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_137),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_6),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_145),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_75),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_70),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_1),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_47),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_11),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_93),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_33),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_142),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_43),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_4),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_25),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_33),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_122),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_32),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_5),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_21),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_66),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_123),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_84),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_146),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_24),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_3),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_82),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_27),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_63),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_4),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_8),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_49),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_3),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_60),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_8),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_55),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_112),
.Y(n_307)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_195),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_155),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_222),
.Y(n_310)
);

INVxp33_ASAP7_75t_L g311 ( 
.A(n_284),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_158),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_222),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_226),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_226),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_222),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_222),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_222),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_230),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_230),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_187),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_161),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_247),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_195),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_247),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_232),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_232),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_157),
.B(n_7),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_262),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_262),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_177),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_278),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_162),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_169),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_190),
.B(n_173),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_278),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_289),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_220),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_172),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_289),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_176),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_210),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_210),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_215),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_215),
.Y(n_345)
);

INVxp33_ASAP7_75t_L g346 ( 
.A(n_229),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_229),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_179),
.Y(n_348)
);

INVxp33_ASAP7_75t_L g349 ( 
.A(n_231),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_183),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_185),
.Y(n_351)
);

BUFx6f_ASAP7_75t_SL g352 ( 
.A(n_177),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_231),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_157),
.B(n_7),
.Y(n_354)
);

INVxp33_ASAP7_75t_SL g355 ( 
.A(n_160),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_196),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_159),
.B(n_10),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_193),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_234),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_234),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_199),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_241),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_200),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_202),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_241),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_287),
.Y(n_366)
);

NOR2xp67_ASAP7_75t_L g367 ( 
.A(n_173),
.B(n_10),
.Y(n_367)
);

NOR2xp67_ASAP7_75t_L g368 ( 
.A(n_281),
.B(n_12),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_245),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_203),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_198),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_206),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_245),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_208),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_248),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_214),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_216),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_248),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_190),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_217),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_219),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_223),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_159),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_310),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_310),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_313),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_308),
.A2(n_243),
.B1(n_288),
.B2(n_239),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_324),
.B(n_201),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_321),
.B(n_167),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_335),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_335),
.B(n_379),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_313),
.Y(n_392)
);

OA21x2_ASAP7_75t_L g393 ( 
.A1(n_383),
.A2(n_165),
.B(n_163),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_383),
.Y(n_394)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_319),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_316),
.Y(n_396)
);

AND2x4_ASAP7_75t_L g397 ( 
.A(n_316),
.B(n_275),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_317),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_317),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_318),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_318),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_358),
.A2(n_249),
.B1(n_170),
.B2(n_164),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_319),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_355),
.B(n_314),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_342),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_320),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_342),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_343),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_320),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_331),
.B(n_163),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_328),
.B(n_307),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_343),
.B(n_275),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_344),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_323),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_323),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_325),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_325),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_329),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_329),
.B(n_165),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_354),
.B(n_227),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g421 ( 
.A(n_338),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_357),
.B(n_306),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_330),
.Y(n_423)
);

AND2x6_ASAP7_75t_L g424 ( 
.A(n_344),
.B(n_156),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_330),
.B(n_166),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_326),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_371),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_345),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_332),
.B(n_166),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_345),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_347),
.B(n_228),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_347),
.B(n_233),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_332),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_336),
.B(n_175),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_353),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_336),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_337),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_315),
.B(n_204),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_366),
.B(n_168),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_353),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_359),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_337),
.Y(n_442)
);

INVx6_ASAP7_75t_L g443 ( 
.A(n_371),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_367),
.B(n_232),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g445 ( 
.A(n_327),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_340),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_359),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_311),
.B(n_207),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_360),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_340),
.B(n_175),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_368),
.A2(n_305),
.B1(n_303),
.B2(n_302),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_346),
.A2(n_250),
.B1(n_252),
.B2(n_259),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_391),
.B(n_309),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_405),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_388),
.B(n_312),
.Y(n_455)
);

INVx2_ASAP7_75t_SL g456 ( 
.A(n_391),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_384),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_426),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_411),
.B(n_322),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g460 ( 
.A(n_390),
.B(n_333),
.Y(n_460)
);

AO22x2_ASAP7_75t_L g461 ( 
.A1(n_410),
.A2(n_281),
.B1(n_252),
.B2(n_259),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_391),
.B(n_360),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_388),
.B(n_334),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_384),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_405),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_384),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_390),
.B(n_411),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_407),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_410),
.B(n_362),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_420),
.B(n_339),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_394),
.Y(n_471)
);

OAI21xp33_ASAP7_75t_SL g472 ( 
.A1(n_410),
.A2(n_181),
.B(n_178),
.Y(n_472)
);

AND2x6_ASAP7_75t_L g473 ( 
.A(n_419),
.B(n_282),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_404),
.A2(n_382),
.B1(n_381),
.B2(n_372),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_389),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_407),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_426),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_408),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_408),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_386),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g481 ( 
.A(n_431),
.B(n_341),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_394),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_420),
.B(n_348),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_394),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_413),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_394),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_413),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_386),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_428),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_422),
.B(n_350),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_394),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_438),
.B(n_351),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_422),
.B(n_356),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_393),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_419),
.B(n_362),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_404),
.B(n_361),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_393),
.Y(n_497)
);

NAND2xp33_ASAP7_75t_L g498 ( 
.A(n_424),
.B(n_156),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_438),
.B(n_363),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_386),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_443),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_431),
.B(n_364),
.Y(n_502)
);

INVx5_ASAP7_75t_L g503 ( 
.A(n_424),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_394),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_393),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_393),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_396),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_432),
.B(n_370),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_448),
.B(n_374),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_448),
.B(n_376),
.Y(n_510)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_389),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_426),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_432),
.B(n_380),
.Y(n_513)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_445),
.B(n_349),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_451),
.B(n_377),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_394),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_395),
.B(n_299),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_428),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_394),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_395),
.B(n_238),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_419),
.B(n_365),
.Y(n_521)
);

BUFx4f_ASAP7_75t_L g522 ( 
.A(n_393),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_395),
.B(n_240),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_430),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_396),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_443),
.A2(n_352),
.B1(n_251),
.B2(n_304),
.Y(n_526)
);

BUFx10_ASAP7_75t_L g527 ( 
.A(n_443),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_430),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_435),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_403),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_395),
.B(n_246),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_435),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_403),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_396),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_403),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_425),
.B(n_365),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_385),
.Y(n_537)
);

AND3x1_ASAP7_75t_L g538 ( 
.A(n_387),
.B(n_286),
.C(n_250),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_425),
.B(n_178),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_403),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_451),
.B(n_257),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_399),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_403),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_440),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_395),
.B(n_263),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_440),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_403),
.Y(n_547)
);

OAI22xp33_ASAP7_75t_SL g548 ( 
.A1(n_444),
.A2(n_209),
.B1(n_235),
.B2(n_225),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_441),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g550 ( 
.A(n_445),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_425),
.B(n_181),
.Y(n_551)
);

INVx5_ASAP7_75t_L g552 ( 
.A(n_424),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_399),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_399),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_429),
.B(n_369),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_443),
.Y(n_556)
);

AND2x2_ASAP7_75t_SL g557 ( 
.A(n_427),
.B(n_282),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_385),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_403),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_401),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_397),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_392),
.B(n_264),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_392),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_SL g564 ( 
.A1(n_402),
.A2(n_352),
.B1(n_279),
.B2(n_265),
.Y(n_564)
);

INVx2_ASAP7_75t_SL g565 ( 
.A(n_443),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_397),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_397),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_443),
.A2(n_352),
.B1(n_276),
.B2(n_267),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_427),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_389),
.B(n_171),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_429),
.B(n_184),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_445),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_441),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_397),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_444),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_398),
.B(n_400),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_401),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_398),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_400),
.B(n_268),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_447),
.Y(n_580)
);

AND2x6_ASAP7_75t_L g581 ( 
.A(n_429),
.B(n_184),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_434),
.B(n_369),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_397),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_387),
.A2(n_197),
.B1(n_212),
.B2(n_211),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_401),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_447),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_406),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_434),
.B(n_373),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_452),
.A2(n_194),
.B1(n_301),
.B2(n_300),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_421),
.B(n_269),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_421),
.B(n_271),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_406),
.Y(n_592)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_439),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_406),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_406),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_449),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_SL g597 ( 
.A(n_421),
.B(n_272),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_449),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_439),
.Y(n_599)
);

INVx4_ASAP7_75t_L g600 ( 
.A(n_412),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_402),
.B(n_274),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_459),
.B(n_409),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_456),
.B(n_156),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_467),
.B(n_452),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_566),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_495),
.B(n_521),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_456),
.A2(n_277),
.B1(n_265),
.B2(n_270),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_470),
.B(n_493),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_566),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_583),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_513),
.B(n_483),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_583),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_490),
.B(n_409),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_502),
.B(n_409),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_561),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_453),
.A2(n_224),
.B1(n_191),
.B2(n_192),
.Y(n_616)
);

OAI22xp33_ASAP7_75t_L g617 ( 
.A1(n_575),
.A2(n_224),
.B1(n_236),
.B2(n_235),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_537),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_514),
.B(n_439),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_494),
.A2(n_279),
.B1(n_270),
.B2(n_273),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_508),
.B(n_409),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_598),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_598),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_458),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_454),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_L g626 ( 
.A1(n_575),
.A2(n_213),
.B1(n_191),
.B2(n_266),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_465),
.Y(n_627)
);

INVxp33_ASAP7_75t_L g628 ( 
.A(n_514),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_537),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_600),
.B(n_156),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_501),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_494),
.A2(n_286),
.B1(n_273),
.B2(n_277),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_561),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_468),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_458),
.B(n_434),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_476),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_460),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_478),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_481),
.A2(n_209),
.B1(n_192),
.B2(n_266),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_558),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_469),
.B(n_409),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_479),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_485),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_462),
.B(n_450),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_558),
.Y(n_645)
);

INVxp67_ASAP7_75t_L g646 ( 
.A(n_477),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_460),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_487),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_563),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_489),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_518),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_469),
.B(n_437),
.Y(n_652)
);

OAI22xp33_ASAP7_75t_L g653 ( 
.A1(n_481),
.A2(n_213),
.B1(n_218),
.B2(n_221),
.Y(n_653)
);

NOR3xp33_ASAP7_75t_L g654 ( 
.A(n_515),
.B(n_450),
.C(n_189),
.Y(n_654)
);

NAND2x1p5_ASAP7_75t_L g655 ( 
.A(n_501),
.B(n_218),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_524),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_528),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_462),
.B(n_437),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_529),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_563),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_495),
.B(n_437),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_521),
.B(n_437),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_578),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_557),
.B(n_280),
.Y(n_664)
);

NAND2xp33_ASAP7_75t_SL g665 ( 
.A(n_477),
.B(n_512),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_536),
.B(n_437),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_561),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_496),
.B(n_174),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_578),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_536),
.B(n_412),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_555),
.B(n_412),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_512),
.B(n_450),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_492),
.B(n_180),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_556),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_561),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_497),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_499),
.B(n_182),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_497),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_600),
.B(n_156),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_555),
.B(n_412),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_532),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_582),
.B(n_412),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_550),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_544),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_505),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_582),
.B(n_406),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_588),
.B(n_406),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_588),
.B(n_406),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_600),
.B(n_522),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_546),
.B(n_549),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_522),
.B(n_297),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_573),
.B(n_406),
.Y(n_692)
);

INVx4_ASAP7_75t_L g693 ( 
.A(n_561),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_505),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_567),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_506),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_567),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_522),
.B(n_297),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_567),
.B(n_297),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_580),
.B(n_436),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_506),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_556),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_455),
.B(n_186),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_463),
.B(n_188),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_586),
.B(n_436),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_509),
.B(n_510),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_596),
.B(n_436),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_557),
.A2(n_294),
.B1(n_293),
.B2(n_292),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_517),
.B(n_436),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_461),
.A2(n_298),
.B1(n_256),
.B2(n_254),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_576),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_541),
.B(n_205),
.Y(n_712)
);

NAND3xp33_ASAP7_75t_L g713 ( 
.A(n_472),
.B(n_295),
.C(n_237),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_539),
.B(n_436),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_539),
.B(n_551),
.Y(n_715)
);

OR2x2_ASAP7_75t_SL g716 ( 
.A(n_538),
.B(n_298),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_457),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_539),
.B(n_436),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_551),
.B(n_436),
.Y(n_719)
);

OAI22x1_ASAP7_75t_SL g720 ( 
.A1(n_599),
.A2(n_261),
.B1(n_255),
.B2(n_285),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_567),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_551),
.B(n_436),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_567),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_461),
.A2(n_221),
.B1(n_225),
.B2(n_236),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_571),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_571),
.B(n_446),
.Y(n_726)
);

INVxp33_ASAP7_75t_L g727 ( 
.A(n_570),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_601),
.B(n_242),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_571),
.B(n_373),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_562),
.B(n_579),
.Y(n_730)
);

NAND2xp33_ASAP7_75t_L g731 ( 
.A(n_473),
.B(n_291),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_461),
.A2(n_253),
.B1(n_260),
.B2(n_297),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_574),
.B(n_297),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_581),
.B(n_446),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_597),
.B(n_244),
.Y(n_735)
);

OR2x6_ASAP7_75t_L g736 ( 
.A(n_550),
.B(n_253),
.Y(n_736)
);

INVx6_ASAP7_75t_L g737 ( 
.A(n_527),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_581),
.B(n_446),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_464),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_464),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_574),
.B(n_258),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_574),
.B(n_446),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_466),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_572),
.B(n_584),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_581),
.B(n_520),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_572),
.B(n_375),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_466),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_474),
.B(n_375),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_480),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_527),
.B(n_565),
.Y(n_750)
);

NAND3xp33_ASAP7_75t_L g751 ( 
.A(n_564),
.B(n_283),
.C(n_290),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_565),
.Y(n_752)
);

OR2x2_ASAP7_75t_L g753 ( 
.A(n_475),
.B(n_378),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_590),
.B(n_591),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_581),
.B(n_446),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_461),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_581),
.B(n_446),
.Y(n_757)
);

AND2x6_ASAP7_75t_SL g758 ( 
.A(n_570),
.B(n_378),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_581),
.B(n_446),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_569),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_526),
.B(n_296),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_523),
.B(n_531),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_527),
.B(n_446),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_511),
.B(n_260),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_545),
.B(n_442),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_480),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_473),
.B(n_535),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_488),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_473),
.B(n_442),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_473),
.B(n_442),
.Y(n_770)
);

OR2x6_ASAP7_75t_SL g771 ( 
.A(n_569),
.B(n_433),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_473),
.B(n_433),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_488),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_691),
.A2(n_698),
.B(n_689),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_608),
.B(n_473),
.Y(n_775)
);

OAI21xp5_ASAP7_75t_L g776 ( 
.A1(n_691),
.A2(n_486),
.B(n_471),
.Y(n_776)
);

A2O1A1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_604),
.A2(n_568),
.B(n_595),
.C(n_594),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_698),
.A2(n_533),
.B(n_595),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_611),
.B(n_548),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_672),
.B(n_746),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_605),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_711),
.B(n_577),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_730),
.B(n_577),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_730),
.B(n_577),
.Y(n_784)
);

OAI21xp33_ASAP7_75t_L g785 ( 
.A1(n_604),
.A2(n_589),
.B(n_593),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_618),
.Y(n_786)
);

AO21x1_ASAP7_75t_L g787 ( 
.A1(n_668),
.A2(n_594),
.B(n_592),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_644),
.B(n_668),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_606),
.B(n_599),
.Y(n_789)
);

A2O1A1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_706),
.A2(n_592),
.B(n_516),
.C(n_471),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_689),
.A2(n_533),
.B(n_535),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_686),
.A2(n_688),
.B(n_687),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_606),
.B(n_414),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_605),
.Y(n_794)
);

A2O1A1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_706),
.A2(n_491),
.B(n_471),
.C(n_484),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_622),
.B(n_535),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_623),
.B(n_540),
.Y(n_797)
);

O2A1O1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_756),
.A2(n_498),
.B(n_585),
.C(n_560),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_676),
.B(n_540),
.Y(n_799)
);

NOR3xp33_ASAP7_75t_L g800 ( 
.A(n_735),
.B(n_498),
.C(n_415),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_676),
.B(n_540),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_715),
.A2(n_533),
.B(n_543),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_678),
.B(n_543),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_605),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_618),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_658),
.A2(n_559),
.B(n_543),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_629),
.Y(n_807)
);

AOI22x1_ASAP7_75t_SL g808 ( 
.A1(n_758),
.A2(n_414),
.B1(n_415),
.B2(n_416),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_637),
.B(n_647),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_629),
.Y(n_810)
);

NOR2xp67_ASAP7_75t_L g811 ( 
.A(n_760),
.B(n_559),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_748),
.B(n_414),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_678),
.B(n_559),
.Y(n_813)
);

OAI21xp5_ASAP7_75t_L g814 ( 
.A1(n_641),
.A2(n_491),
.B(n_516),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_614),
.A2(n_621),
.B(n_652),
.Y(n_815)
);

NOR2xp67_ASAP7_75t_L g816 ( 
.A(n_646),
.B(n_484),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_624),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_754),
.A2(n_516),
.B1(n_491),
.B2(n_486),
.Y(n_818)
);

NAND2x1p5_ASAP7_75t_L g819 ( 
.A(n_615),
.B(n_503),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_729),
.B(n_484),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_613),
.A2(n_486),
.B(n_587),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_685),
.B(n_587),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_635),
.B(n_415),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_605),
.B(n_503),
.Y(n_824)
);

HB1xp67_ASAP7_75t_L g825 ( 
.A(n_683),
.Y(n_825)
);

AOI21xp33_ASAP7_75t_L g826 ( 
.A1(n_728),
.A2(n_525),
.B(n_560),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_709),
.A2(n_587),
.B(n_585),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_640),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_612),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_640),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_628),
.B(n_416),
.Y(n_831)
);

OAI21x1_ASAP7_75t_L g832 ( 
.A1(n_767),
.A2(n_554),
.B(n_553),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_754),
.A2(n_554),
.B1(n_553),
.B2(n_500),
.Y(n_833)
);

OAI21xp5_ASAP7_75t_L g834 ( 
.A1(n_661),
.A2(n_500),
.B(n_542),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_685),
.B(n_507),
.Y(n_835)
);

O2A1O1Ixp5_ASAP7_75t_L g836 ( 
.A1(n_630),
.A2(n_507),
.B(n_525),
.C(n_542),
.Y(n_836)
);

AOI22x1_ASAP7_75t_L g837 ( 
.A1(n_694),
.A2(n_534),
.B1(n_482),
.B2(n_519),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_694),
.B(n_534),
.Y(n_838)
);

CKINVDCx20_ASAP7_75t_R g839 ( 
.A(n_665),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_696),
.B(n_482),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_670),
.A2(n_547),
.B(n_530),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_771),
.Y(n_842)
);

OAI21xp5_ASAP7_75t_L g843 ( 
.A1(n_662),
.A2(n_666),
.B(n_762),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_696),
.B(n_482),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_671),
.A2(n_547),
.B(n_530),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_735),
.B(n_530),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_701),
.B(n_482),
.Y(n_847)
);

BUFx4f_ASAP7_75t_L g848 ( 
.A(n_753),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_645),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_744),
.B(n_530),
.Y(n_850)
);

BUFx2_ASAP7_75t_L g851 ( 
.A(n_736),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_645),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_701),
.B(n_482),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_602),
.B(n_504),
.Y(n_854)
);

OR2x2_ASAP7_75t_L g855 ( 
.A(n_764),
.B(n_416),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_703),
.A2(n_504),
.B1(n_519),
.B2(n_530),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_725),
.B(n_504),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_680),
.A2(n_547),
.B(n_519),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_682),
.B(n_649),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_612),
.B(n_503),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_612),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_649),
.B(n_504),
.Y(n_862)
);

AO21x1_ASAP7_75t_L g863 ( 
.A1(n_728),
.A2(n_417),
.B(n_418),
.Y(n_863)
);

INVxp67_ASAP7_75t_L g864 ( 
.A(n_619),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_660),
.B(n_504),
.Y(n_865)
);

A2O1A1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_703),
.A2(n_433),
.B(n_418),
.C(n_423),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_765),
.A2(n_718),
.B(n_714),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_609),
.A2(n_519),
.B1(n_547),
.B2(n_552),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_719),
.A2(n_547),
.B(n_519),
.Y(n_869)
);

NOR2xp67_ASAP7_75t_L g870 ( 
.A(n_708),
.B(n_64),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_729),
.B(n_417),
.Y(n_871)
);

NOR2x1_ASAP7_75t_L g872 ( 
.A(n_751),
.B(n_423),
.Y(n_872)
);

INVx4_ASAP7_75t_L g873 ( 
.A(n_612),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_673),
.B(n_417),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_609),
.Y(n_875)
);

AND2x2_ASAP7_75t_SL g876 ( 
.A(n_761),
.B(n_418),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_631),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_744),
.B(n_13),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_660),
.B(n_423),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_736),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_722),
.A2(n_552),
.B(n_503),
.Y(n_881)
);

INVx4_ASAP7_75t_L g882 ( 
.A(n_737),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_663),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_625),
.B(n_52),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_663),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_726),
.A2(n_552),
.B(n_503),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_669),
.B(n_424),
.Y(n_887)
);

OAI21xp5_ASAP7_75t_L g888 ( 
.A1(n_745),
.A2(n_552),
.B(n_424),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_669),
.B(n_424),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_673),
.B(n_13),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_627),
.B(n_424),
.Y(n_891)
);

O2A1O1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_616),
.A2(n_424),
.B(n_15),
.C(n_16),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_634),
.B(n_424),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_636),
.B(n_424),
.Y(n_894)
);

INVx1_ASAP7_75t_SL g895 ( 
.A(n_736),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_769),
.A2(n_552),
.B(n_62),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_L g897 ( 
.A1(n_712),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_638),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_770),
.A2(n_73),
.B(n_134),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_SL g900 ( 
.A(n_704),
.B(n_151),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_642),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_643),
.B(n_14),
.Y(n_902)
);

A2O1A1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_704),
.A2(n_18),
.B(n_19),
.C(n_21),
.Y(n_903)
);

O2A1O1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_639),
.A2(n_18),
.B(n_19),
.C(n_24),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_648),
.B(n_26),
.Y(n_905)
);

NOR3xp33_ASAP7_75t_L g906 ( 
.A(n_761),
.B(n_27),
.C(n_31),
.Y(n_906)
);

AOI21xp33_ASAP7_75t_L g907 ( 
.A1(n_712),
.A2(n_32),
.B(n_35),
.Y(n_907)
);

AO22x1_ASAP7_75t_L g908 ( 
.A1(n_677),
.A2(n_37),
.B1(n_39),
.B2(n_42),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_677),
.B(n_37),
.Y(n_909)
);

BUFx8_ASAP7_75t_L g910 ( 
.A(n_650),
.Y(n_910)
);

AO21x2_ASAP7_75t_L g911 ( 
.A1(n_741),
.A2(n_733),
.B(n_630),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_651),
.Y(n_912)
);

A2O1A1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_656),
.A2(n_42),
.B(n_43),
.C(n_45),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_657),
.B(n_45),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_615),
.B(n_111),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_659),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_681),
.B(n_48),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_684),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_690),
.B(n_48),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_734),
.A2(n_79),
.B(n_86),
.Y(n_920)
);

INVxp67_ASAP7_75t_SL g921 ( 
.A(n_615),
.Y(n_921)
);

A2O1A1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_654),
.A2(n_97),
.B(n_102),
.C(n_107),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_664),
.B(n_110),
.Y(n_923)
);

AO21x1_ASAP7_75t_L g924 ( 
.A1(n_603),
.A2(n_741),
.B(n_733),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_615),
.B(n_633),
.Y(n_925)
);

AND2x2_ASAP7_75t_SL g926 ( 
.A(n_607),
.B(n_119),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_610),
.A2(n_126),
.B1(n_128),
.B2(n_130),
.Y(n_927)
);

AO21x1_ASAP7_75t_L g928 ( 
.A1(n_603),
.A2(n_132),
.B(n_133),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_631),
.B(n_752),
.Y(n_929)
);

OAI22xp5_ASAP7_75t_L g930 ( 
.A1(n_620),
.A2(n_632),
.B1(n_752),
.B2(n_674),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_717),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_772),
.A2(n_750),
.B(n_763),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_653),
.B(n_716),
.Y(n_933)
);

NOR2x1p5_ASAP7_75t_SL g934 ( 
.A(n_740),
.B(n_768),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_740),
.Y(n_935)
);

O2A1O1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_617),
.A2(n_626),
.B(n_710),
.C(n_620),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_674),
.B(n_702),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_632),
.A2(n_699),
.B(n_679),
.C(n_724),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_633),
.B(n_697),
.Y(n_939)
);

NOR3xp33_ASAP7_75t_L g940 ( 
.A(n_713),
.B(n_731),
.C(n_721),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_633),
.B(n_697),
.Y(n_941)
);

INVx1_ASAP7_75t_SL g942 ( 
.A(n_720),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_633),
.Y(n_943)
);

NAND2x1_ASAP7_75t_L g944 ( 
.A(n_737),
.B(n_697),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_750),
.A2(n_763),
.B(n_755),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_702),
.B(n_697),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_655),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_738),
.A2(n_759),
.B(n_757),
.Y(n_948)
);

OR2x2_ASAP7_75t_L g949 ( 
.A(n_727),
.B(n_607),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_747),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_742),
.A2(n_705),
.B(n_707),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_747),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_675),
.B(n_723),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_742),
.A2(n_700),
.B(n_692),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_667),
.B(n_675),
.Y(n_955)
);

AOI21xp33_ASAP7_75t_L g956 ( 
.A1(n_724),
.A2(n_710),
.B(n_732),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_768),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_679),
.A2(n_693),
.B(n_723),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_667),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_695),
.B(n_693),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_667),
.B(n_695),
.Y(n_961)
);

AND3x1_ASAP7_75t_SL g962 ( 
.A(n_898),
.B(n_739),
.C(n_766),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_774),
.A2(n_667),
.B(n_699),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_774),
.A2(n_655),
.B(n_743),
.Y(n_964)
);

AOI21x1_ASAP7_75t_L g965 ( 
.A1(n_932),
.A2(n_749),
.B(n_773),
.Y(n_965)
);

BUFx2_ASAP7_75t_L g966 ( 
.A(n_789),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_788),
.B(n_732),
.Y(n_967)
);

CKINVDCx20_ASAP7_75t_R g968 ( 
.A(n_839),
.Y(n_968)
);

O2A1O1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_878),
.A2(n_737),
.B(n_909),
.C(n_907),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_785),
.B(n_864),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_876),
.A2(n_850),
.B1(n_926),
.B2(n_779),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_843),
.A2(n_775),
.B(n_859),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_930),
.A2(n_784),
.B1(n_783),
.B2(n_846),
.Y(n_973)
);

AOI22xp33_ASAP7_75t_L g974 ( 
.A1(n_890),
.A2(n_933),
.B1(n_956),
.B2(n_923),
.Y(n_974)
);

OA21x2_ASAP7_75t_L g975 ( 
.A1(n_863),
.A2(n_787),
.B(n_814),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_L g976 ( 
.A1(n_780),
.A2(n_900),
.B1(n_812),
.B2(n_820),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_L g977 ( 
.A1(n_929),
.A2(n_937),
.B1(n_875),
.B2(n_946),
.Y(n_977)
);

BUFx2_ASAP7_75t_L g978 ( 
.A(n_817),
.Y(n_978)
);

O2A1O1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_903),
.A2(n_906),
.B(n_904),
.C(n_919),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_949),
.B(n_855),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_848),
.B(n_877),
.Y(n_981)
);

NAND3xp33_ASAP7_75t_SL g982 ( 
.A(n_897),
.B(n_904),
.C(n_895),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_815),
.A2(n_792),
.B(n_867),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_815),
.A2(n_792),
.B(n_867),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_808),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_854),
.A2(n_948),
.B(n_932),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_848),
.B(n_877),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_877),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_825),
.B(n_809),
.Y(n_989)
);

O2A1O1Ixp5_ASAP7_75t_SL g990 ( 
.A1(n_826),
.A2(n_920),
.B(n_915),
.C(n_885),
.Y(n_990)
);

AOI22x1_ASAP7_75t_L g991 ( 
.A1(n_874),
.A2(n_945),
.B1(n_958),
.B2(n_951),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_948),
.A2(n_858),
.B(n_845),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_820),
.B(n_884),
.Y(n_993)
);

NAND2xp33_ASAP7_75t_L g994 ( 
.A(n_781),
.B(n_794),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_823),
.B(n_793),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_781),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_880),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_858),
.A2(n_845),
.B(n_841),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_842),
.Y(n_999)
);

O2A1O1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_777),
.A2(n_902),
.B(n_917),
.C(n_914),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_905),
.A2(n_913),
.B(n_936),
.C(n_918),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_831),
.B(n_871),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_851),
.B(n_901),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_786),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_938),
.A2(n_945),
.B(n_870),
.C(n_916),
.Y(n_1005)
);

OAI21xp33_ASAP7_75t_SL g1006 ( 
.A1(n_912),
.A2(n_782),
.B(n_810),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_875),
.A2(n_856),
.B1(n_818),
.B2(n_805),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_828),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_830),
.B(n_849),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_884),
.B(n_947),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_882),
.B(n_955),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_910),
.Y(n_1012)
);

INVxp67_ASAP7_75t_SL g1013 ( 
.A(n_781),
.Y(n_1013)
);

NOR2x1_ASAP7_75t_L g1014 ( 
.A(n_882),
.B(n_873),
.Y(n_1014)
);

AO32x1_ASAP7_75t_L g1015 ( 
.A1(n_852),
.A2(n_883),
.A3(n_935),
.B1(n_950),
.B2(n_952),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_816),
.B(n_960),
.Y(n_1016)
);

BUFx4f_ASAP7_75t_SL g1017 ( 
.A(n_942),
.Y(n_1017)
);

NAND2xp33_ASAP7_75t_L g1018 ( 
.A(n_794),
.B(n_804),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_841),
.A2(n_951),
.B(n_954),
.Y(n_1019)
);

BUFx4f_ASAP7_75t_SL g1020 ( 
.A(n_794),
.Y(n_1020)
);

INVx4_ASAP7_75t_L g1021 ( 
.A(n_804),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_921),
.A2(n_938),
.B1(n_961),
.B2(n_857),
.Y(n_1022)
);

AND2x2_ASAP7_75t_SL g1023 ( 
.A(n_873),
.B(n_804),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_931),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_960),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_958),
.A2(n_953),
.B1(n_829),
.B2(n_861),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_829),
.B(n_861),
.Y(n_1027)
);

O2A1O1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_892),
.A2(n_795),
.B(n_790),
.C(n_922),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_954),
.A2(n_776),
.B(n_869),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_829),
.A2(n_861),
.B1(n_943),
.B2(n_959),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_811),
.B(n_959),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_943),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_940),
.A2(n_800),
.B(n_798),
.C(n_872),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_957),
.B(n_835),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_925),
.B(n_939),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_869),
.A2(n_924),
.B(n_778),
.Y(n_1036)
);

AOI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_911),
.A2(n_941),
.B1(n_894),
.B2(n_891),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_R g1038 ( 
.A(n_893),
.B(n_796),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_797),
.B(n_847),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_892),
.A2(n_798),
.B(n_866),
.C(n_865),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_838),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_833),
.B(n_862),
.Y(n_1042)
);

OR2x2_ASAP7_75t_L g1043 ( 
.A(n_879),
.B(n_813),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_799),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_778),
.A2(n_802),
.B(n_844),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_840),
.A2(n_853),
.B1(n_944),
.B2(n_803),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_822),
.B(n_801),
.Y(n_1047)
);

INVx3_ASAP7_75t_L g1048 ( 
.A(n_819),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_908),
.Y(n_1049)
);

BUFx3_ASAP7_75t_L g1050 ( 
.A(n_928),
.Y(n_1050)
);

BUFx2_ASAP7_75t_L g1051 ( 
.A(n_927),
.Y(n_1051)
);

HB1xp67_ASAP7_75t_L g1052 ( 
.A(n_887),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_802),
.A2(n_821),
.B(n_834),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_911),
.B(n_806),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_821),
.A2(n_791),
.B(n_806),
.Y(n_1055)
);

INVx1_ASAP7_75t_SL g1056 ( 
.A(n_899),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_934),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_791),
.A2(n_827),
.B(n_888),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_819),
.Y(n_1059)
);

NOR2x1_ASAP7_75t_SL g1060 ( 
.A(n_868),
.B(n_824),
.Y(n_1060)
);

O2A1O1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_899),
.A2(n_889),
.B(n_896),
.C(n_836),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_827),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_832),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_860),
.B(n_896),
.Y(n_1064)
);

CKINVDCx6p67_ASAP7_75t_R g1065 ( 
.A(n_837),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_R g1066 ( 
.A(n_881),
.B(n_886),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_881),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_886),
.B(n_608),
.Y(n_1068)
);

BUFx8_ASAP7_75t_SL g1069 ( 
.A(n_839),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_788),
.B(n_608),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_909),
.A2(n_608),
.B(n_878),
.C(n_604),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_788),
.B(n_608),
.Y(n_1072)
);

NAND2x1p5_ASAP7_75t_L g1073 ( 
.A(n_882),
.B(n_873),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_780),
.B(n_672),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_788),
.B(n_608),
.Y(n_1075)
);

AND2x2_ASAP7_75t_SL g1076 ( 
.A(n_926),
.B(n_608),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_R g1077 ( 
.A(n_839),
.B(n_569),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_788),
.B(n_608),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_909),
.A2(n_608),
.B(n_788),
.C(n_878),
.Y(n_1079)
);

NAND2x1_ASAP7_75t_L g1080 ( 
.A(n_873),
.B(n_737),
.Y(n_1080)
);

AOI22xp33_ASAP7_75t_L g1081 ( 
.A1(n_926),
.A2(n_608),
.B1(n_909),
.B2(n_878),
.Y(n_1081)
);

O2A1O1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_878),
.A2(n_608),
.B(n_909),
.C(n_668),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_788),
.B(n_608),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_877),
.Y(n_1084)
);

AO32x1_ASAP7_75t_L g1085 ( 
.A1(n_890),
.A2(n_616),
.A3(n_626),
.B1(n_639),
.B2(n_756),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_774),
.A2(n_843),
.B(n_608),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_789),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_774),
.A2(n_843),
.B(n_608),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_788),
.B(n_608),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_807),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_877),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_877),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_774),
.A2(n_843),
.B(n_608),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_788),
.B(n_608),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_774),
.A2(n_843),
.B(n_608),
.Y(n_1095)
);

INVx1_ASAP7_75t_SL g1096 ( 
.A(n_817),
.Y(n_1096)
);

OAI22x1_ASAP7_75t_L g1097 ( 
.A1(n_878),
.A2(n_604),
.B1(n_933),
.B2(n_570),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_788),
.B(n_608),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_807),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_774),
.A2(n_843),
.B(n_608),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_788),
.B(n_608),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_780),
.B(n_672),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_807),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_1081),
.A2(n_1071),
.B1(n_1076),
.B2(n_974),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_1069),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_1072),
.A2(n_1078),
.B1(n_1089),
.B2(n_1101),
.Y(n_1106)
);

NAND2x1p5_ASAP7_75t_L g1107 ( 
.A(n_1023),
.B(n_1080),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1086),
.A2(n_1093),
.B(n_1088),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_1070),
.B(n_1094),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1086),
.A2(n_1093),
.B(n_1088),
.Y(n_1110)
);

AOI211x1_ASAP7_75t_L g1111 ( 
.A1(n_1098),
.A2(n_1075),
.B(n_1083),
.C(n_967),
.Y(n_1111)
);

INVx2_ASAP7_75t_SL g1112 ( 
.A(n_978),
.Y(n_1112)
);

AOI221x1_ASAP7_75t_L g1113 ( 
.A1(n_971),
.A2(n_1097),
.B1(n_983),
.B2(n_984),
.C(n_973),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_998),
.A2(n_965),
.B(n_963),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_1082),
.B(n_1074),
.Y(n_1115)
);

AO31x2_ASAP7_75t_L g1116 ( 
.A1(n_1019),
.A2(n_998),
.A3(n_1053),
.B(n_992),
.Y(n_1116)
);

OR2x6_ASAP7_75t_L g1117 ( 
.A(n_1010),
.B(n_981),
.Y(n_1117)
);

NOR2xp67_ASAP7_75t_L g1118 ( 
.A(n_1025),
.B(n_976),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_1079),
.A2(n_969),
.B(n_979),
.C(n_1001),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1004),
.Y(n_1120)
);

O2A1O1Ixp5_ASAP7_75t_SL g1121 ( 
.A1(n_1062),
.A2(n_1054),
.B(n_1057),
.C(n_1022),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1008),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_1079),
.A2(n_970),
.B(n_1049),
.C(n_982),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1102),
.B(n_1002),
.Y(n_1124)
);

OAI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1095),
.A2(n_1100),
.B(n_972),
.Y(n_1125)
);

NAND3xp33_ASAP7_75t_L g1126 ( 
.A(n_1005),
.B(n_1100),
.C(n_1095),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_1000),
.A2(n_1028),
.B(n_1051),
.C(n_1006),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_980),
.B(n_989),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_995),
.B(n_1041),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_963),
.A2(n_1045),
.B(n_1055),
.Y(n_1130)
);

OA21x2_ASAP7_75t_L g1131 ( 
.A1(n_1036),
.A2(n_992),
.B(n_1053),
.Y(n_1131)
);

O2A1O1Ixp5_ASAP7_75t_L g1132 ( 
.A1(n_983),
.A2(n_984),
.B(n_1055),
.C(n_1019),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_972),
.A2(n_1068),
.B(n_986),
.Y(n_1133)
);

BUFx4f_ASAP7_75t_SL g1134 ( 
.A(n_968),
.Y(n_1134)
);

AO31x2_ASAP7_75t_L g1135 ( 
.A1(n_1036),
.A2(n_1033),
.A3(n_986),
.B(n_1058),
.Y(n_1135)
);

BUFx4f_ASAP7_75t_SL g1136 ( 
.A(n_1096),
.Y(n_1136)
);

INVx2_ASAP7_75t_SL g1137 ( 
.A(n_997),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1029),
.A2(n_1058),
.B(n_1056),
.Y(n_1138)
);

AOI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_993),
.A2(n_1087),
.B1(n_966),
.B2(n_1003),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_1040),
.A2(n_1050),
.B(n_1039),
.C(n_1035),
.Y(n_1140)
);

NAND3xp33_ASAP7_75t_L g1141 ( 
.A(n_990),
.B(n_991),
.C(n_1029),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_1045),
.A2(n_964),
.B(n_1063),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_1025),
.Y(n_1143)
);

O2A1O1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_987),
.A2(n_1007),
.B(n_977),
.C(n_1042),
.Y(n_1144)
);

OAI21xp33_ASAP7_75t_SL g1145 ( 
.A1(n_1044),
.A2(n_1009),
.B(n_1034),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1024),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_964),
.A2(n_1061),
.B(n_1067),
.Y(n_1147)
);

NOR2x1_ASAP7_75t_SL g1148 ( 
.A(n_1030),
.B(n_1016),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1064),
.A2(n_1031),
.B(n_1052),
.C(n_1026),
.Y(n_1149)
);

AO21x2_ASAP7_75t_L g1150 ( 
.A1(n_1066),
.A2(n_1037),
.B(n_1060),
.Y(n_1150)
);

AO21x1_ASAP7_75t_L g1151 ( 
.A1(n_1046),
.A2(n_1047),
.B(n_1011),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_999),
.B(n_985),
.Y(n_1152)
);

OR2x2_ASAP7_75t_L g1153 ( 
.A(n_1103),
.B(n_1099),
.Y(n_1153)
);

O2A1O1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1090),
.A2(n_1043),
.B(n_994),
.C(n_1018),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_SL g1155 ( 
.A1(n_1027),
.A2(n_1013),
.B(n_1032),
.C(n_1048),
.Y(n_1155)
);

INVx3_ASAP7_75t_L g1156 ( 
.A(n_1048),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_996),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_SL g1158 ( 
.A1(n_1073),
.A2(n_996),
.B(n_975),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_1014),
.A2(n_962),
.B(n_1065),
.Y(n_1159)
);

AO32x2_ASAP7_75t_L g1160 ( 
.A1(n_1085),
.A2(n_1015),
.A3(n_1021),
.B1(n_1038),
.B2(n_1020),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_1059),
.Y(n_1161)
);

A2O1A1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_988),
.A2(n_1092),
.B(n_1091),
.C(n_1084),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1085),
.A2(n_1015),
.B(n_1021),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_996),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_988),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1084),
.A2(n_1091),
.B(n_1077),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_1017),
.A2(n_1071),
.B(n_608),
.C(n_1082),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1012),
.A2(n_608),
.B(n_1095),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_1071),
.B(n_848),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1004),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_978),
.Y(n_1171)
);

INVx1_ASAP7_75t_SL g1172 ( 
.A(n_1096),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_978),
.Y(n_1173)
);

NAND2x1p5_ASAP7_75t_L g1174 ( 
.A(n_1023),
.B(n_882),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1072),
.B(n_1078),
.Y(n_1175)
);

AOI21x1_ASAP7_75t_L g1176 ( 
.A1(n_963),
.A2(n_964),
.B(n_965),
.Y(n_1176)
);

OA21x2_ASAP7_75t_L g1177 ( 
.A1(n_1036),
.A2(n_992),
.B(n_998),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1086),
.A2(n_608),
.B(n_1095),
.Y(n_1178)
);

INVx3_ASAP7_75t_SL g1179 ( 
.A(n_999),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1086),
.A2(n_608),
.B(n_1095),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1086),
.A2(n_608),
.B(n_1095),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1086),
.A2(n_608),
.B(n_1095),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_978),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1004),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_998),
.A2(n_832),
.B(n_965),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_1071),
.B(n_848),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_998),
.A2(n_832),
.B(n_965),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1086),
.A2(n_608),
.B(n_1095),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_998),
.A2(n_832),
.B(n_965),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1082),
.A2(n_608),
.B(n_1071),
.C(n_1081),
.Y(n_1190)
);

AO31x2_ASAP7_75t_L g1191 ( 
.A1(n_1019),
.A2(n_787),
.A3(n_863),
.B(n_998),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_SL g1192 ( 
.A1(n_1005),
.A2(n_608),
.B(n_1082),
.Y(n_1192)
);

OR2x2_ASAP7_75t_L g1193 ( 
.A(n_980),
.B(n_949),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1074),
.B(n_1102),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_998),
.A2(n_832),
.B(n_965),
.Y(n_1195)
);

AO31x2_ASAP7_75t_L g1196 ( 
.A1(n_1019),
.A2(n_787),
.A3(n_863),
.B(n_998),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1074),
.B(n_1102),
.Y(n_1197)
);

AO32x2_ASAP7_75t_L g1198 ( 
.A1(n_971),
.A2(n_973),
.A3(n_1022),
.B1(n_1007),
.B2(n_756),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1071),
.B(n_608),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_SL g1200 ( 
.A(n_1076),
.B(n_926),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1086),
.A2(n_608),
.B(n_1095),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1086),
.A2(n_608),
.B(n_1095),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1086),
.A2(n_608),
.B(n_1095),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_978),
.Y(n_1204)
);

INVx4_ASAP7_75t_L g1205 ( 
.A(n_1020),
.Y(n_1205)
);

AOI21xp33_ASAP7_75t_L g1206 ( 
.A1(n_1082),
.A2(n_1079),
.B(n_1071),
.Y(n_1206)
);

OAI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1071),
.A2(n_1082),
.B(n_974),
.Y(n_1207)
);

HB1xp67_ASAP7_75t_L g1208 ( 
.A(n_978),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1071),
.B(n_608),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1086),
.A2(n_608),
.B(n_1095),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_1010),
.B(n_981),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1086),
.A2(n_608),
.B(n_1095),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1072),
.B(n_1078),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1072),
.B(n_1078),
.Y(n_1214)
);

NAND3xp33_ASAP7_75t_L g1215 ( 
.A(n_1082),
.B(n_608),
.C(n_1071),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1072),
.B(n_1078),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1004),
.Y(n_1217)
);

AO22x2_ASAP7_75t_L g1218 ( 
.A1(n_971),
.A2(n_982),
.B1(n_1049),
.B2(n_906),
.Y(n_1218)
);

O2A1O1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_1071),
.A2(n_608),
.B(n_1082),
.C(n_878),
.Y(n_1219)
);

AO32x2_ASAP7_75t_L g1220 ( 
.A1(n_971),
.A2(n_973),
.A3(n_1022),
.B1(n_1007),
.B2(n_756),
.Y(n_1220)
);

O2A1O1Ixp5_ASAP7_75t_L g1221 ( 
.A1(n_1071),
.A2(n_608),
.B(n_909),
.C(n_668),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1072),
.B(n_1078),
.Y(n_1222)
);

OAI22x1_ASAP7_75t_L g1223 ( 
.A1(n_1049),
.A2(n_878),
.B1(n_909),
.B2(n_604),
.Y(n_1223)
);

O2A1O1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1071),
.A2(n_608),
.B(n_1082),
.C(n_878),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1004),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_998),
.A2(n_832),
.B(n_965),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1086),
.A2(n_608),
.B(n_1095),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1072),
.B(n_1078),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1086),
.A2(n_608),
.B(n_1095),
.Y(n_1229)
);

O2A1O1Ixp33_ASAP7_75t_SL g1230 ( 
.A1(n_1071),
.A2(n_1082),
.B(n_608),
.C(n_956),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_998),
.A2(n_832),
.B(n_965),
.Y(n_1231)
);

OR2x2_ASAP7_75t_L g1232 ( 
.A(n_980),
.B(n_949),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1004),
.Y(n_1233)
);

AOI221xp5_ASAP7_75t_SL g1234 ( 
.A1(n_1071),
.A2(n_1082),
.B1(n_1081),
.B2(n_878),
.C(n_1079),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_R g1235 ( 
.A1(n_971),
.A2(n_639),
.B(n_584),
.Y(n_1235)
);

CKINVDCx8_ASAP7_75t_R g1236 ( 
.A(n_999),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1120),
.Y(n_1237)
);

BUFx5_ASAP7_75t_L g1238 ( 
.A(n_1122),
.Y(n_1238)
);

CKINVDCx6p67_ASAP7_75t_R g1239 ( 
.A(n_1179),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1199),
.A2(n_1209),
.B1(n_1104),
.B2(n_1207),
.Y(n_1240)
);

BUFx2_ASAP7_75t_L g1241 ( 
.A(n_1204),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1104),
.A2(n_1207),
.B1(n_1223),
.B2(n_1215),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1215),
.A2(n_1206),
.B1(n_1218),
.B2(n_1228),
.Y(n_1243)
);

AOI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1109),
.A2(n_1200),
.B1(n_1222),
.B2(n_1175),
.Y(n_1244)
);

OR2x2_ASAP7_75t_L g1245 ( 
.A(n_1193),
.B(n_1232),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1206),
.A2(n_1218),
.B1(n_1213),
.B2(n_1216),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1170),
.Y(n_1247)
);

BUFx10_ASAP7_75t_L g1248 ( 
.A(n_1152),
.Y(n_1248)
);

BUFx3_ASAP7_75t_L g1249 ( 
.A(n_1136),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1173),
.Y(n_1250)
);

CKINVDCx11_ASAP7_75t_R g1251 ( 
.A(n_1236),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1214),
.A2(n_1106),
.B1(n_1200),
.B2(n_1186),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1184),
.Y(n_1253)
);

CKINVDCx11_ASAP7_75t_R g1254 ( 
.A(n_1105),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_1134),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1153),
.Y(n_1256)
);

OR2x2_ASAP7_75t_L g1257 ( 
.A(n_1124),
.B(n_1128),
.Y(n_1257)
);

BUFx12f_ASAP7_75t_L g1258 ( 
.A(n_1183),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_SL g1259 ( 
.A1(n_1106),
.A2(n_1235),
.B1(n_1126),
.B2(n_1197),
.Y(n_1259)
);

CKINVDCx6p67_ASAP7_75t_R g1260 ( 
.A(n_1172),
.Y(n_1260)
);

CKINVDCx8_ASAP7_75t_R g1261 ( 
.A(n_1211),
.Y(n_1261)
);

OAI22x1_ASAP7_75t_L g1262 ( 
.A1(n_1139),
.A2(n_1169),
.B1(n_1115),
.B2(n_1211),
.Y(n_1262)
);

OAI21xp33_ASAP7_75t_L g1263 ( 
.A1(n_1190),
.A2(n_1119),
.B(n_1224),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1139),
.A2(n_1140),
.B1(n_1127),
.B2(n_1117),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1126),
.A2(n_1168),
.B1(n_1129),
.B2(n_1194),
.Y(n_1265)
);

BUFx3_ASAP7_75t_L g1266 ( 
.A(n_1112),
.Y(n_1266)
);

INVxp67_ASAP7_75t_SL g1267 ( 
.A(n_1144),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1118),
.A2(n_1188),
.B1(n_1178),
.B2(n_1180),
.Y(n_1268)
);

CKINVDCx20_ASAP7_75t_R g1269 ( 
.A(n_1171),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1118),
.A2(n_1212),
.B1(n_1181),
.B2(n_1182),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1201),
.A2(n_1202),
.B1(n_1210),
.B2(n_1203),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_SL g1272 ( 
.A1(n_1234),
.A2(n_1150),
.B1(n_1141),
.B2(n_1125),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_1208),
.Y(n_1273)
);

OAI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1113),
.A2(n_1233),
.B1(n_1225),
.B2(n_1217),
.Y(n_1274)
);

CKINVDCx6p67_ASAP7_75t_R g1275 ( 
.A(n_1157),
.Y(n_1275)
);

INVx1_ASAP7_75t_SL g1276 ( 
.A(n_1137),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1146),
.B(n_1123),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_SL g1278 ( 
.A1(n_1234),
.A2(n_1150),
.B1(n_1141),
.B2(n_1125),
.Y(n_1278)
);

OAI221xp5_ASAP7_75t_L g1279 ( 
.A1(n_1219),
.A2(n_1221),
.B1(n_1167),
.B2(n_1192),
.C(n_1230),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1174),
.A2(n_1111),
.B1(n_1107),
.B2(n_1161),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1165),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1164),
.Y(n_1282)
);

BUFx10_ASAP7_75t_L g1283 ( 
.A(n_1166),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1154),
.A2(n_1143),
.B1(n_1162),
.B2(n_1156),
.Y(n_1284)
);

INVx5_ASAP7_75t_L g1285 ( 
.A(n_1143),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1227),
.B(n_1229),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1159),
.Y(n_1287)
);

BUFx2_ASAP7_75t_SL g1288 ( 
.A(n_1151),
.Y(n_1288)
);

OAI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1108),
.A2(n_1110),
.B1(n_1138),
.B2(n_1131),
.Y(n_1289)
);

BUFx12f_ASAP7_75t_L g1290 ( 
.A(n_1148),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1145),
.A2(n_1131),
.B1(n_1177),
.B2(n_1133),
.Y(n_1291)
);

INVxp67_ASAP7_75t_L g1292 ( 
.A(n_1177),
.Y(n_1292)
);

OAI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1163),
.A2(n_1220),
.B1(n_1198),
.B2(n_1176),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_SL g1294 ( 
.A1(n_1145),
.A2(n_1163),
.B1(n_1220),
.B2(n_1198),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1130),
.A2(n_1147),
.B1(n_1114),
.B2(n_1142),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1198),
.A2(n_1220),
.B1(n_1231),
.B2(n_1187),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1185),
.A2(n_1226),
.B1(n_1195),
.B2(n_1189),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1135),
.A2(n_1149),
.B1(n_1121),
.B2(n_1132),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1160),
.A2(n_1116),
.B1(n_1191),
.B2(n_1196),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_1160),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1158),
.A2(n_1155),
.B1(n_1160),
.B2(n_1116),
.Y(n_1301)
);

CKINVDCx11_ASAP7_75t_R g1302 ( 
.A(n_1191),
.Y(n_1302)
);

INVx6_ASAP7_75t_L g1303 ( 
.A(n_1191),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1196),
.A2(n_1081),
.B1(n_608),
.B2(n_1175),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1153),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1199),
.A2(n_878),
.B1(n_1081),
.B2(n_1209),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1199),
.A2(n_878),
.B1(n_1081),
.B2(n_1209),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1175),
.A2(n_1081),
.B1(n_608),
.B2(n_1213),
.Y(n_1308)
);

BUFx3_ASAP7_75t_L g1309 ( 
.A(n_1136),
.Y(n_1309)
);

BUFx4f_ASAP7_75t_SL g1310 ( 
.A(n_1105),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1175),
.A2(n_1081),
.B1(n_608),
.B2(n_1213),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1175),
.B(n_1213),
.Y(n_1312)
);

INVx1_ASAP7_75t_SL g1313 ( 
.A(n_1136),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1153),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1175),
.A2(n_1081),
.B1(n_608),
.B2(n_1213),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1175),
.B(n_1213),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1211),
.B(n_1117),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_SL g1318 ( 
.A1(n_1200),
.A2(n_1076),
.B1(n_926),
.B2(n_878),
.Y(n_1318)
);

BUFx4_ASAP7_75t_R g1319 ( 
.A(n_1204),
.Y(n_1319)
);

CKINVDCx11_ASAP7_75t_R g1320 ( 
.A(n_1236),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1135),
.Y(n_1321)
);

BUFx2_ASAP7_75t_R g1322 ( 
.A(n_1236),
.Y(n_1322)
);

BUFx10_ASAP7_75t_L g1323 ( 
.A(n_1152),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1175),
.B(n_1213),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1153),
.Y(n_1325)
);

INVx4_ASAP7_75t_L g1326 ( 
.A(n_1136),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1199),
.A2(n_878),
.B1(n_1081),
.B2(n_1209),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1105),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1105),
.Y(n_1329)
);

CKINVDCx11_ASAP7_75t_R g1330 ( 
.A(n_1236),
.Y(n_1330)
);

INVx6_ASAP7_75t_L g1331 ( 
.A(n_1205),
.Y(n_1331)
);

INVx8_ASAP7_75t_L g1332 ( 
.A(n_1117),
.Y(n_1332)
);

CKINVDCx6p67_ASAP7_75t_R g1333 ( 
.A(n_1179),
.Y(n_1333)
);

CKINVDCx6p67_ASAP7_75t_R g1334 ( 
.A(n_1179),
.Y(n_1334)
);

AOI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1199),
.A2(n_608),
.B1(n_668),
.B2(n_1081),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1175),
.A2(n_1081),
.B1(n_608),
.B2(n_1213),
.Y(n_1336)
);

NAND2xp33_ASAP7_75t_SL g1337 ( 
.A(n_1175),
.B(n_608),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1199),
.A2(n_878),
.B1(n_1081),
.B2(n_1209),
.Y(n_1338)
);

CKINVDCx20_ASAP7_75t_R g1339 ( 
.A(n_1105),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1153),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1245),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1321),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1246),
.B(n_1267),
.Y(n_1343)
);

INVx4_ASAP7_75t_SL g1344 ( 
.A(n_1303),
.Y(n_1344)
);

BUFx12f_ASAP7_75t_L g1345 ( 
.A(n_1330),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1303),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1238),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1286),
.A2(n_1271),
.B(n_1297),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1306),
.A2(n_1327),
.B1(n_1338),
.B2(n_1307),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1290),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1242),
.B(n_1299),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1292),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1237),
.Y(n_1353)
);

INVx4_ASAP7_75t_L g1354 ( 
.A(n_1332),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1274),
.Y(n_1355)
);

OR2x6_ASAP7_75t_L g1356 ( 
.A(n_1288),
.B(n_1332),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1274),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1294),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1294),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1271),
.A2(n_1297),
.B(n_1295),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1256),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1312),
.B(n_1316),
.Y(n_1362)
);

OAI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1335),
.A2(n_1307),
.B(n_1338),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1247),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1253),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1246),
.B(n_1267),
.Y(n_1366)
);

BUFx3_ASAP7_75t_L g1367 ( 
.A(n_1317),
.Y(n_1367)
);

INVx2_ASAP7_75t_SL g1368 ( 
.A(n_1283),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1306),
.A2(n_1327),
.B1(n_1318),
.B2(n_1240),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1287),
.B(n_1285),
.Y(n_1370)
);

INVxp67_ASAP7_75t_L g1371 ( 
.A(n_1277),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1293),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1318),
.A2(n_1263),
.B1(n_1311),
.B2(n_1308),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1302),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1300),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1293),
.Y(n_1376)
);

INVxp67_ASAP7_75t_SL g1377 ( 
.A(n_1289),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1301),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1300),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1300),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1295),
.A2(n_1268),
.B(n_1270),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1305),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_1261),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1289),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1272),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1272),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1268),
.A2(n_1270),
.B(n_1291),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1291),
.A2(n_1298),
.B(n_1296),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1278),
.B(n_1243),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1278),
.Y(n_1390)
);

AO21x2_ASAP7_75t_L g1391 ( 
.A1(n_1279),
.A2(n_1304),
.B(n_1264),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1262),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1298),
.A2(n_1296),
.B(n_1299),
.Y(n_1393)
);

AO21x2_ASAP7_75t_L g1394 ( 
.A1(n_1284),
.A2(n_1336),
.B(n_1315),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1243),
.B(n_1257),
.Y(n_1395)
);

CKINVDCx20_ASAP7_75t_R g1396 ( 
.A(n_1254),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1265),
.A2(n_1280),
.B(n_1252),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1265),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1259),
.Y(n_1399)
);

AOI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1281),
.A2(n_1282),
.B(n_1314),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1259),
.B(n_1252),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1325),
.B(n_1340),
.Y(n_1402)
);

CKINVDCx6p67_ASAP7_75t_R g1403 ( 
.A(n_1251),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1244),
.B(n_1324),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1337),
.A2(n_1269),
.B1(n_1250),
.B2(n_1258),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_1275),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1273),
.B(n_1260),
.Y(n_1407)
);

CKINVDCx20_ASAP7_75t_R g1408 ( 
.A(n_1339),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1341),
.B(n_1241),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1363),
.A2(n_1276),
.B(n_1266),
.Y(n_1410)
);

AOI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1349),
.A2(n_1369),
.B1(n_1363),
.B2(n_1373),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1362),
.B(n_1255),
.Y(n_1412)
);

AOI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1400),
.A2(n_1319),
.B(n_1248),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1404),
.B(n_1319),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1375),
.B(n_1323),
.Y(n_1415)
);

AOI221xp5_ASAP7_75t_L g1416 ( 
.A1(n_1389),
.A2(n_1313),
.B1(n_1326),
.B2(n_1249),
.C(n_1309),
.Y(n_1416)
);

INVx2_ASAP7_75t_SL g1417 ( 
.A(n_1370),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1404),
.B(n_1323),
.Y(n_1418)
);

CKINVDCx6p67_ASAP7_75t_R g1419 ( 
.A(n_1345),
.Y(n_1419)
);

OR2x6_ASAP7_75t_L g1420 ( 
.A(n_1356),
.B(n_1331),
.Y(n_1420)
);

CKINVDCx20_ASAP7_75t_R g1421 ( 
.A(n_1396),
.Y(n_1421)
);

INVx4_ASAP7_75t_L g1422 ( 
.A(n_1406),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1353),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1372),
.B(n_1239),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1376),
.B(n_1334),
.Y(n_1425)
);

AND2x4_ASAP7_75t_SL g1426 ( 
.A(n_1406),
.B(n_1333),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1391),
.A2(n_1329),
.B(n_1328),
.Y(n_1427)
);

AND4x1_ASAP7_75t_L g1428 ( 
.A(n_1405),
.B(n_1322),
.C(n_1320),
.D(n_1251),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1379),
.B(n_1320),
.Y(n_1429)
);

OR2x2_ASAP7_75t_L g1430 ( 
.A(n_1371),
.B(n_1310),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1364),
.Y(n_1431)
);

AO32x1_ASAP7_75t_L g1432 ( 
.A1(n_1389),
.A2(n_1401),
.A3(n_1390),
.B1(n_1386),
.B2(n_1385),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1380),
.B(n_1358),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1361),
.B(n_1382),
.Y(n_1434)
);

CKINVDCx16_ASAP7_75t_R g1435 ( 
.A(n_1345),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1391),
.A2(n_1387),
.B(n_1377),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1401),
.A2(n_1399),
.B1(n_1394),
.B2(n_1391),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_SL g1438 ( 
.A1(n_1391),
.A2(n_1394),
.B1(n_1399),
.B2(n_1366),
.Y(n_1438)
);

AND3x1_ASAP7_75t_L g1439 ( 
.A(n_1374),
.B(n_1407),
.C(n_1402),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1358),
.B(n_1359),
.Y(n_1440)
);

INVx5_ASAP7_75t_SL g1441 ( 
.A(n_1403),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1359),
.B(n_1385),
.Y(n_1442)
);

OA21x2_ASAP7_75t_L g1443 ( 
.A1(n_1388),
.A2(n_1360),
.B(n_1381),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1374),
.B(n_1402),
.Y(n_1444)
);

O2A1O1Ixp33_ASAP7_75t_L g1445 ( 
.A1(n_1343),
.A2(n_1366),
.B(n_1394),
.C(n_1392),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1386),
.B(n_1390),
.Y(n_1446)
);

AO21x2_ASAP7_75t_L g1447 ( 
.A1(n_1360),
.A2(n_1348),
.B(n_1384),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1378),
.B(n_1353),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_SL g1449 ( 
.A1(n_1343),
.A2(n_1374),
.B(n_1354),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1378),
.B(n_1353),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1344),
.B(n_1368),
.Y(n_1451)
);

AND2x6_ASAP7_75t_L g1452 ( 
.A(n_1392),
.B(n_1346),
.Y(n_1452)
);

A2O1A1Ixp33_ASAP7_75t_L g1453 ( 
.A1(n_1387),
.A2(n_1397),
.B(n_1381),
.C(n_1398),
.Y(n_1453)
);

NOR2xp67_ASAP7_75t_L g1454 ( 
.A(n_1427),
.B(n_1423),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1446),
.B(n_1355),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1411),
.A2(n_1392),
.B1(n_1395),
.B2(n_1367),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1449),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1443),
.B(n_1384),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1437),
.A2(n_1351),
.B1(n_1355),
.B2(n_1357),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1423),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_SL g1461 ( 
.A1(n_1438),
.A2(n_1345),
.B1(n_1357),
.B2(n_1383),
.Y(n_1461)
);

BUFx2_ASAP7_75t_L g1462 ( 
.A(n_1452),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1453),
.B(n_1447),
.Y(n_1463)
);

NOR2x1_ASAP7_75t_SL g1464 ( 
.A(n_1420),
.B(n_1356),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1447),
.B(n_1393),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1445),
.B(n_1352),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1453),
.B(n_1393),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1448),
.B(n_1393),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1417),
.B(n_1347),
.Y(n_1469)
);

CKINVDCx20_ASAP7_75t_R g1470 ( 
.A(n_1421),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1450),
.B(n_1433),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1442),
.B(n_1365),
.Y(n_1472)
);

BUFx2_ASAP7_75t_L g1473 ( 
.A(n_1452),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1431),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1434),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1467),
.B(n_1436),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1466),
.B(n_1442),
.Y(n_1477)
);

AND2x2_ASAP7_75t_SL g1478 ( 
.A(n_1462),
.B(n_1439),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1466),
.B(n_1440),
.Y(n_1479)
);

AOI221xp5_ASAP7_75t_L g1480 ( 
.A1(n_1461),
.A2(n_1410),
.B1(n_1416),
.B2(n_1414),
.C(n_1440),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1458),
.Y(n_1481)
);

AND2x4_ASAP7_75t_L g1482 ( 
.A(n_1464),
.B(n_1451),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1458),
.B(n_1342),
.Y(n_1483)
);

OAI221xp5_ASAP7_75t_L g1484 ( 
.A1(n_1461),
.A2(n_1418),
.B1(n_1428),
.B2(n_1414),
.C(n_1412),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1454),
.B(n_1413),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1460),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1467),
.B(n_1444),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1458),
.Y(n_1488)
);

NOR2x1_ASAP7_75t_L g1489 ( 
.A(n_1454),
.B(n_1420),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1468),
.B(n_1415),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_L g1491 ( 
.A(n_1475),
.B(n_1430),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1456),
.A2(n_1425),
.B1(n_1424),
.B2(n_1383),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_L g1493 ( 
.A(n_1460),
.Y(n_1493)
);

NAND3xp33_ASAP7_75t_L g1494 ( 
.A(n_1463),
.B(n_1459),
.C(n_1465),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1468),
.B(n_1415),
.Y(n_1495)
);

INVx3_ASAP7_75t_L g1496 ( 
.A(n_1469),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1474),
.Y(n_1497)
);

NOR2x1_ASAP7_75t_L g1498 ( 
.A(n_1457),
.B(n_1420),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1477),
.B(n_1471),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1482),
.B(n_1473),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1497),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_SL g1502 ( 
.A(n_1478),
.B(n_1457),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1478),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1483),
.B(n_1463),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1486),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1477),
.B(n_1471),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1497),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1477),
.B(n_1471),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1497),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1481),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1479),
.B(n_1455),
.Y(n_1511)
);

BUFx2_ASAP7_75t_L g1512 ( 
.A(n_1489),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1486),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1484),
.B(n_1435),
.Y(n_1514)
);

AND2x4_ASAP7_75t_L g1515 ( 
.A(n_1482),
.B(n_1473),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1479),
.B(n_1455),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1481),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1496),
.B(n_1476),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1479),
.B(n_1472),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1481),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1481),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1488),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1488),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1493),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1511),
.B(n_1491),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1505),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1505),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1510),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1513),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1499),
.B(n_1494),
.Y(n_1530)
);

INVx1_ASAP7_75t_SL g1531 ( 
.A(n_1502),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1513),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1511),
.B(n_1491),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1524),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1524),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_SL g1536 ( 
.A(n_1502),
.B(n_1478),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1510),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1503),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1501),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1501),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1501),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1499),
.B(n_1506),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1506),
.B(n_1494),
.Y(n_1543)
);

INVx2_ASAP7_75t_SL g1544 ( 
.A(n_1503),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1507),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1508),
.B(n_1516),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1507),
.Y(n_1547)
);

NAND2x1p5_ASAP7_75t_L g1548 ( 
.A(n_1512),
.B(n_1489),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1516),
.B(n_1487),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1507),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1510),
.Y(n_1551)
);

INVxp67_ASAP7_75t_L g1552 ( 
.A(n_1514),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1509),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1503),
.B(n_1482),
.Y(n_1554)
);

NAND4xp25_ASAP7_75t_L g1555 ( 
.A(n_1503),
.B(n_1480),
.C(n_1492),
.D(n_1484),
.Y(n_1555)
);

AOI211xp5_ASAP7_75t_SL g1556 ( 
.A1(n_1514),
.A2(n_1480),
.B(n_1459),
.C(n_1476),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1519),
.B(n_1487),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1500),
.B(n_1482),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1510),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1509),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1508),
.B(n_1483),
.Y(n_1561)
);

INVx2_ASAP7_75t_SL g1562 ( 
.A(n_1500),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1519),
.B(n_1483),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1517),
.Y(n_1564)
);

INVxp67_ASAP7_75t_L g1565 ( 
.A(n_1512),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1504),
.B(n_1487),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1536),
.B(n_1500),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1556),
.B(n_1490),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1536),
.B(n_1500),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1554),
.B(n_1500),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1554),
.B(n_1500),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1538),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1539),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1531),
.B(n_1515),
.Y(n_1574)
);

AOI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1555),
.A2(n_1552),
.B(n_1544),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1525),
.B(n_1504),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1540),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1533),
.B(n_1504),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1541),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1530),
.B(n_1517),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1545),
.Y(n_1581)
);

NAND4xp25_ASAP7_75t_SL g1582 ( 
.A(n_1530),
.B(n_1476),
.C(n_1498),
.D(n_1492),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1544),
.B(n_1490),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1543),
.B(n_1490),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1562),
.B(n_1512),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1543),
.B(n_1495),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1547),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1562),
.B(n_1515),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_1526),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1550),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1528),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1546),
.B(n_1517),
.Y(n_1592)
);

AOI22x1_ASAP7_75t_L g1593 ( 
.A1(n_1548),
.A2(n_1350),
.B1(n_1406),
.B2(n_1403),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1558),
.B(n_1515),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1527),
.B(n_1488),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1546),
.B(n_1517),
.Y(n_1596)
);

INVxp67_ASAP7_75t_L g1597 ( 
.A(n_1529),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1528),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1532),
.B(n_1488),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1534),
.B(n_1509),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1558),
.B(n_1515),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1568),
.A2(n_1478),
.B1(n_1548),
.B2(n_1498),
.Y(n_1602)
);

AOI31xp33_ASAP7_75t_L g1603 ( 
.A1(n_1575),
.A2(n_1548),
.A3(n_1565),
.B(n_1498),
.Y(n_1603)
);

AOI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1582),
.A2(n_1485),
.B(n_1421),
.Y(n_1604)
);

O2A1O1Ixp33_ASAP7_75t_SL g1605 ( 
.A1(n_1572),
.A2(n_1597),
.B(n_1470),
.C(n_1485),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1573),
.Y(n_1606)
);

NOR3xp33_ASAP7_75t_L g1607 ( 
.A(n_1589),
.B(n_1535),
.C(n_1425),
.Y(n_1607)
);

AOI31xp33_ASAP7_75t_L g1608 ( 
.A1(n_1567),
.A2(n_1489),
.A3(n_1424),
.B(n_1403),
.Y(n_1608)
);

OAI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1593),
.A2(n_1542),
.B(n_1515),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1589),
.B(n_1549),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1573),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1589),
.B(n_1557),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1577),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1593),
.A2(n_1566),
.B(n_1432),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1585),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1585),
.Y(n_1616)
);

INVx2_ASAP7_75t_SL g1617 ( 
.A(n_1585),
.Y(n_1617)
);

AOI21xp33_ASAP7_75t_L g1618 ( 
.A1(n_1580),
.A2(n_1542),
.B(n_1457),
.Y(n_1618)
);

OAI21xp33_ASAP7_75t_L g1619 ( 
.A1(n_1567),
.A2(n_1561),
.B(n_1563),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1569),
.B(n_1515),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1569),
.B(n_1518),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1576),
.B(n_1563),
.Y(n_1622)
);

AOI221xp5_ASAP7_75t_L g1623 ( 
.A1(n_1576),
.A2(n_1553),
.B1(n_1560),
.B2(n_1564),
.C(n_1559),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1570),
.B(n_1518),
.Y(n_1624)
);

XOR2x2_ASAP7_75t_L g1625 ( 
.A(n_1584),
.B(n_1419),
.Y(n_1625)
);

O2A1O1Ixp33_ASAP7_75t_L g1626 ( 
.A1(n_1578),
.A2(n_1409),
.B(n_1561),
.C(n_1559),
.Y(n_1626)
);

OAI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1604),
.A2(n_1585),
.B(n_1578),
.Y(n_1627)
);

XOR2x2_ASAP7_75t_L g1628 ( 
.A(n_1625),
.B(n_1602),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1607),
.B(n_1574),
.Y(n_1629)
);

OAI21xp33_ASAP7_75t_SL g1630 ( 
.A1(n_1603),
.A2(n_1571),
.B(n_1570),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1606),
.Y(n_1631)
);

AOI221xp5_ASAP7_75t_L g1632 ( 
.A1(n_1605),
.A2(n_1586),
.B1(n_1574),
.B2(n_1579),
.C(n_1587),
.Y(n_1632)
);

AOI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1605),
.A2(n_1571),
.B1(n_1588),
.B2(n_1583),
.Y(n_1633)
);

AOI21xp33_ASAP7_75t_L g1634 ( 
.A1(n_1617),
.A2(n_1608),
.B(n_1615),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1620),
.B(n_1621),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1611),
.Y(n_1636)
);

OA21x2_ASAP7_75t_L g1637 ( 
.A1(n_1615),
.A2(n_1598),
.B(n_1591),
.Y(n_1637)
);

NOR2xp67_ASAP7_75t_L g1638 ( 
.A(n_1617),
.B(n_1580),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1613),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1619),
.B(n_1419),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1616),
.Y(n_1641)
);

OAI31xp33_ASAP7_75t_L g1642 ( 
.A1(n_1618),
.A2(n_1588),
.A3(n_1601),
.B(n_1594),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1620),
.B(n_1594),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1616),
.Y(n_1644)
);

INVxp67_ASAP7_75t_SL g1645 ( 
.A(n_1610),
.Y(n_1645)
);

NAND3xp33_ASAP7_75t_L g1646 ( 
.A(n_1623),
.B(n_1579),
.C(n_1577),
.Y(n_1646)
);

OAI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1645),
.A2(n_1625),
.B(n_1612),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1645),
.B(n_1621),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1641),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1635),
.B(n_1601),
.Y(n_1650)
);

XOR2x2_ASAP7_75t_L g1651 ( 
.A(n_1628),
.B(n_1609),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1640),
.B(n_1622),
.Y(n_1652)
);

AOI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1628),
.A2(n_1626),
.B(n_1614),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1641),
.Y(n_1654)
);

INVxp67_ASAP7_75t_L g1655 ( 
.A(n_1640),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1644),
.Y(n_1656)
);

OAI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1653),
.A2(n_1633),
.B1(n_1629),
.B2(n_1627),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1655),
.B(n_1634),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1648),
.Y(n_1659)
);

INVxp67_ASAP7_75t_L g1660 ( 
.A(n_1649),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_SL g1661 ( 
.A(n_1647),
.B(n_1638),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1652),
.B(n_1630),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1654),
.Y(n_1663)
);

NAND4xp75_ASAP7_75t_L g1664 ( 
.A(n_1647),
.B(n_1632),
.C(n_1642),
.D(n_1637),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1650),
.B(n_1643),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1657),
.A2(n_1651),
.B1(n_1646),
.B2(n_1656),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1665),
.B(n_1631),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1661),
.B(n_1636),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1663),
.Y(n_1669)
);

OAI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1664),
.A2(n_1639),
.B(n_1637),
.Y(n_1670)
);

CKINVDCx20_ASAP7_75t_R g1671 ( 
.A(n_1667),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1670),
.A2(n_1662),
.B(n_1658),
.Y(n_1672)
);

INVxp67_ASAP7_75t_SL g1673 ( 
.A(n_1668),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1666),
.A2(n_1659),
.B1(n_1660),
.B2(n_1624),
.Y(n_1674)
);

AOI31xp33_ASAP7_75t_L g1675 ( 
.A1(n_1669),
.A2(n_1660),
.A3(n_1407),
.B(n_1581),
.Y(n_1675)
);

O2A1O1Ixp33_ASAP7_75t_L g1676 ( 
.A1(n_1670),
.A2(n_1637),
.B(n_1581),
.C(n_1587),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1671),
.Y(n_1677)
);

OAI322xp33_ASAP7_75t_L g1678 ( 
.A1(n_1672),
.A2(n_1590),
.A3(n_1591),
.B1(n_1598),
.B2(n_1596),
.C1(n_1592),
.C2(n_1600),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1674),
.A2(n_1590),
.B1(n_1600),
.B2(n_1595),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_SL g1680 ( 
.A(n_1675),
.B(n_1591),
.Y(n_1680)
);

AND3x4_ASAP7_75t_L g1681 ( 
.A(n_1673),
.B(n_1598),
.C(n_1441),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1677),
.B(n_1624),
.Y(n_1682)
);

AND4x1_ASAP7_75t_L g1683 ( 
.A(n_1681),
.B(n_1676),
.C(n_1441),
.D(n_1595),
.Y(n_1683)
);

OAI222xp33_ASAP7_75t_L g1684 ( 
.A1(n_1679),
.A2(n_1596),
.B1(n_1592),
.B2(n_1599),
.C1(n_1537),
.C2(n_1564),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1682),
.Y(n_1685)
);

NAND4xp25_ASAP7_75t_L g1686 ( 
.A(n_1685),
.B(n_1680),
.C(n_1683),
.D(n_1678),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1686),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1686),
.B(n_1408),
.Y(n_1688)
);

AO22x2_ASAP7_75t_L g1689 ( 
.A1(n_1687),
.A2(n_1684),
.B1(n_1537),
.B2(n_1551),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1688),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1689),
.Y(n_1691)
);

AO21x2_ASAP7_75t_L g1692 ( 
.A1(n_1690),
.A2(n_1599),
.B(n_1551),
.Y(n_1692)
);

AOI221xp5_ASAP7_75t_L g1693 ( 
.A1(n_1691),
.A2(n_1523),
.B1(n_1522),
.B2(n_1520),
.C(n_1521),
.Y(n_1693)
);

AOI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1693),
.A2(n_1692),
.B(n_1426),
.Y(n_1694)
);

OAI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1694),
.A2(n_1692),
.B1(n_1523),
.B2(n_1522),
.Y(n_1695)
);

OAI221xp5_ASAP7_75t_L g1696 ( 
.A1(n_1695),
.A2(n_1350),
.B1(n_1406),
.B2(n_1441),
.C(n_1422),
.Y(n_1696)
);

AOI211xp5_ASAP7_75t_L g1697 ( 
.A1(n_1696),
.A2(n_1350),
.B(n_1406),
.C(n_1429),
.Y(n_1697)
);


endmodule