module fake_jpeg_2606_n_599 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_599);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_599;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_8),
.B(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_6),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_3),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_7),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_57),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_59),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_61),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_62),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_63),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_30),
.B(n_18),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_64),
.B(n_69),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_65),
.Y(n_202)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_68),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_30),
.B(n_18),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_71),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

BUFx4f_ASAP7_75t_SL g142 ( 
.A(n_72),
.Y(n_142)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_73),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_0),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_74),
.B(n_75),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_0),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_76),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_77),
.Y(n_178)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_79),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g164 ( 
.A(n_80),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_17),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_81),
.B(n_127),
.Y(n_143)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_82),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_31),
.B(n_1),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_83),
.B(n_86),
.Y(n_163)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_84),
.Y(n_149)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_85),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_20),
.B(n_1),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_33),
.B(n_1),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_87),
.B(n_88),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_31),
.B(n_29),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_91),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_31),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_92),
.A2(n_107),
.B1(n_83),
.B2(n_88),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_93),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_94),
.Y(n_172)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_35),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_95),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_96),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_20),
.B(n_2),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_97),
.B(n_98),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_23),
.B(n_2),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_99),
.Y(n_181)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_102),
.Y(n_212)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_103),
.Y(n_175)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_104),
.Y(n_193)
);

BUFx12_ASAP7_75t_L g105 ( 
.A(n_35),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g194 ( 
.A(n_105),
.Y(n_194)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_106),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_22),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_35),
.A2(n_5),
.B(n_6),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_108),
.B(n_109),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_23),
.B(n_6),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_35),
.Y(n_110)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_110),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_26),
.B(n_7),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_111),
.B(n_120),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_32),
.Y(n_112)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_112),
.Y(n_198)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_22),
.Y(n_113)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_113),
.Y(n_199)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_40),
.Y(n_114)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_114),
.Y(n_186)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_38),
.Y(n_115)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_115),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_32),
.Y(n_116)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_116),
.Y(n_200)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_40),
.Y(n_117)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_117),
.Y(n_195)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_38),
.Y(n_118)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_118),
.Y(n_203)
);

BUFx12f_ASAP7_75t_SL g119 ( 
.A(n_38),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_119),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_26),
.B(n_7),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_45),
.Y(n_121)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_121),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_32),
.Y(n_122)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_122),
.Y(n_201)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_25),
.Y(n_123)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_123),
.Y(n_205)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_45),
.Y(n_124)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_124),
.Y(n_196)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_25),
.Y(n_125)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_37),
.Y(n_126)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_126),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_27),
.B(n_56),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_69),
.B(n_64),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_129),
.B(n_169),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_58),
.A2(n_54),
.B1(n_53),
.B2(n_51),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_137),
.A2(n_165),
.B1(n_167),
.B2(n_208),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_138),
.A2(n_48),
.B1(n_14),
.B2(n_16),
.Y(n_252)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_146),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_SL g147 ( 
.A(n_105),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_147),
.Y(n_285)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_74),
.Y(n_151)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_151),
.Y(n_235)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_72),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_154),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_75),
.B(n_98),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_155),
.B(n_157),
.Y(n_283)
);

INVx5_ASAP7_75t_SL g156 ( 
.A(n_112),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g247 ( 
.A(n_156),
.B(n_206),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_109),
.B(n_54),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_111),
.B(n_37),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_160),
.B(n_185),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_120),
.A2(n_45),
.B1(n_22),
.B2(n_53),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_60),
.A2(n_46),
.B1(n_39),
.B2(n_55),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_116),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_87),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_177),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_122),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_184),
.B(n_176),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_61),
.B(n_51),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_62),
.Y(n_187)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_187),
.Y(n_251)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_63),
.Y(n_188)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_188),
.Y(n_263)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_65),
.Y(n_192)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_192),
.Y(n_266)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_67),
.Y(n_204)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_204),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_68),
.B(n_46),
.Y(n_206)
);

AND2x2_ASAP7_75t_SL g207 ( 
.A(n_76),
.B(n_28),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_207),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_77),
.A2(n_55),
.B1(n_44),
.B2(n_39),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_80),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_34),
.Y(n_222)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_91),
.Y(n_211)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_211),
.Y(n_224)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_102),
.Y(n_215)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_93),
.Y(n_216)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_94),
.Y(n_217)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_217),
.Y(n_243)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_96),
.Y(n_218)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_218),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_99),
.A2(n_46),
.B1(n_27),
.B2(n_44),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_219),
.A2(n_166),
.B1(n_139),
.B2(n_197),
.Y(n_299)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_123),
.Y(n_220)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_220),
.Y(n_257)
);

INVx5_ASAP7_75t_SL g221 ( 
.A(n_105),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_221),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_222),
.Y(n_307)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_147),
.Y(n_223)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_223),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_213),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_225),
.Y(n_338)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_144),
.Y(n_226)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_226),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_131),
.Y(n_227)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_227),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_170),
.B(n_28),
.C(n_34),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_228),
.B(n_301),
.C(n_270),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_213),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_229),
.B(n_238),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_159),
.B(n_29),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_230),
.B(n_231),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_133),
.B(n_11),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_145),
.Y(n_232)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_232),
.Y(n_318)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_189),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_236),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_152),
.B(n_12),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_237),
.B(n_245),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_153),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_182),
.B(n_13),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_239),
.B(n_269),
.Y(n_354)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_191),
.Y(n_240)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_240),
.Y(n_306)
);

OAI22xp33_ASAP7_75t_L g241 ( 
.A1(n_165),
.A2(n_28),
.B1(n_48),
.B2(n_15),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_241),
.A2(n_293),
.B1(n_299),
.B2(n_246),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_152),
.B(n_141),
.Y(n_245)
);

AND2x4_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_28),
.Y(n_246)
);

BUFx24_ASAP7_75t_L g355 ( 
.A(n_246),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_173),
.A2(n_28),
.B1(n_48),
.B2(n_16),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_248),
.A2(n_250),
.B1(n_285),
.B2(n_298),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_182),
.A2(n_48),
.B1(n_14),
.B2(n_16),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_249),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_252),
.A2(n_276),
.B1(n_277),
.B2(n_300),
.Y(n_336)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_131),
.Y(n_253)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_253),
.Y(n_309)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_210),
.Y(n_254)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_254),
.Y(n_323)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_175),
.Y(n_256)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_256),
.Y(n_326)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_193),
.Y(n_258)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_258),
.Y(n_327)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_203),
.Y(n_259)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_259),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_177),
.A2(n_13),
.B1(n_14),
.B2(n_17),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_260),
.B(n_262),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_132),
.Y(n_261)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_261),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_170),
.A2(n_13),
.B1(n_14),
.B2(n_17),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_163),
.A2(n_174),
.B1(n_141),
.B2(n_150),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_264),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_163),
.B(n_143),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_268),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_174),
.B(n_180),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_207),
.B(n_171),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_135),
.B(n_136),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_271),
.B(n_272),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_140),
.B(n_158),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_206),
.B(n_199),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_273),
.B(n_282),
.Y(n_330)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_198),
.Y(n_274)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_274),
.Y(n_345)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_200),
.Y(n_275)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_275),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_156),
.A2(n_201),
.B1(n_164),
.B2(n_202),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_164),
.A2(n_197),
.B1(n_202),
.B2(n_183),
.Y(n_277)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_279),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_161),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_280),
.Y(n_346)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_130),
.Y(n_281)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_281),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_172),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_168),
.A2(n_162),
.B1(n_214),
.B2(n_195),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_284),
.A2(n_297),
.B1(n_250),
.B2(n_285),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_221),
.B(n_186),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_287),
.B(n_290),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_137),
.B(n_208),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_288),
.B(n_289),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_130),
.B(n_178),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_181),
.Y(n_290)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_132),
.Y(n_291)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_291),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_149),
.A2(n_178),
.B1(n_166),
.B2(n_139),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_134),
.Y(n_295)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_295),
.Y(n_356)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_179),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_298),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_196),
.A2(n_212),
.B1(n_190),
.B2(n_128),
.Y(n_297)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_194),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_134),
.A2(n_148),
.B1(n_183),
.B2(n_142),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_148),
.B(n_142),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_154),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_302),
.B(n_294),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_310),
.B(n_311),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_255),
.A2(n_288),
.B1(n_239),
.B2(n_267),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_228),
.B(n_286),
.C(n_269),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_312),
.B(n_333),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_225),
.Y(n_313)
);

NAND3xp33_ASAP7_75t_L g400 ( 
.A(n_313),
.B(n_316),
.C(n_317),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_271),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_272),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_252),
.A2(n_247),
.B1(n_273),
.B2(n_289),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_321),
.A2(n_322),
.B1(n_348),
.B2(n_352),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_247),
.A2(n_235),
.B1(n_262),
.B2(n_283),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_328),
.A2(n_337),
.B1(n_242),
.B2(n_224),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_329),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_SL g333 ( 
.A(n_260),
.B(n_241),
.C(n_278),
.Y(n_333)
);

NOR2x1_ASAP7_75t_R g334 ( 
.A(n_246),
.B(n_254),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_334),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_246),
.A2(n_293),
.B1(n_301),
.B2(n_276),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_256),
.B(n_258),
.C(n_233),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_341),
.B(n_342),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_257),
.B(n_296),
.C(n_266),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_343),
.Y(n_396)
);

OAI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_277),
.A2(n_240),
.B1(n_259),
.B2(n_226),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_285),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_349),
.B(n_352),
.Y(n_394)
);

OAI22xp33_ASAP7_75t_L g352 ( 
.A1(n_253),
.A2(n_281),
.B1(n_263),
.B2(n_292),
.Y(n_352)
);

AO22x1_ASAP7_75t_SL g357 ( 
.A1(n_257),
.A2(n_275),
.B1(n_274),
.B2(n_243),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_357),
.B(n_295),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_359),
.A2(n_223),
.B1(n_261),
.B2(n_338),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_347),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_360),
.Y(n_416)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_331),
.Y(n_361)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_361),
.Y(n_429)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_339),
.Y(n_362)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_362),
.Y(n_419)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_331),
.Y(n_363)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_363),
.Y(n_431)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_323),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_365),
.Y(n_405)
);

INVx5_ASAP7_75t_L g366 ( 
.A(n_358),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_366),
.Y(n_436)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_323),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_367),
.B(n_371),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_347),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_368),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_369),
.A2(n_391),
.B1(n_395),
.B2(n_342),
.Y(n_408)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_309),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_370),
.B(n_373),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_319),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_357),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_321),
.A2(n_251),
.B1(n_224),
.B2(n_242),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_375),
.A2(n_380),
.B1(n_381),
.B2(n_390),
.Y(n_426)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_326),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_376),
.B(n_377),
.Y(n_418)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_326),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_335),
.A2(n_291),
.B(n_232),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_378),
.A2(n_355),
.B(n_324),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_307),
.B(n_236),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_379),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_314),
.A2(n_234),
.B1(n_243),
.B2(n_244),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_314),
.A2(n_234),
.B1(n_244),
.B2(n_227),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_382),
.B(n_383),
.Y(n_411)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_357),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g385 ( 
.A(n_356),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_385),
.B(n_386),
.Y(n_424)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_309),
.Y(n_386)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_327),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_388),
.B(n_397),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_305),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_389),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_336),
.A2(n_328),
.B1(n_337),
.B2(n_320),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_356),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_392),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_394),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_335),
.A2(n_322),
.B1(n_311),
.B2(n_330),
.Y(n_395)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_327),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_345),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_398),
.B(n_399),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_303),
.B(n_312),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_310),
.B(n_354),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_401),
.B(n_354),
.Y(n_407)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_345),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_402),
.Y(n_430)
);

OAI22xp33_ASAP7_75t_SL g403 ( 
.A1(n_340),
.A2(n_324),
.B1(n_315),
.B2(n_355),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_403),
.A2(n_338),
.B1(n_344),
.B2(n_358),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_406),
.A2(n_425),
.B(n_434),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_407),
.B(n_414),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_408),
.A2(n_393),
.B1(n_364),
.B2(n_381),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_391),
.A2(n_351),
.B1(n_355),
.B2(n_333),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_409),
.A2(n_415),
.B1(n_432),
.B2(n_433),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_401),
.B(n_341),
.C(n_334),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_412),
.B(n_413),
.C(n_420),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_384),
.B(n_307),
.C(n_350),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_SL g414 ( 
.A(n_384),
.B(n_351),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_373),
.A2(n_351),
.B1(n_332),
.B2(n_339),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_374),
.A2(n_350),
.B(n_344),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_417),
.A2(n_378),
.B(n_396),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_384),
.B(n_304),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_399),
.B(n_346),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_421),
.B(n_439),
.C(n_308),
.Y(n_470)
);

NAND2x1_ASAP7_75t_SL g425 ( 
.A(n_374),
.B(n_346),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_383),
.A2(n_306),
.B1(n_325),
.B2(n_318),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_395),
.A2(n_306),
.B1(n_325),
.B2(n_318),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_387),
.B(n_353),
.Y(n_439)
);

XNOR2x1_ASAP7_75t_L g440 ( 
.A(n_387),
.B(n_353),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_440),
.B(n_393),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_406),
.A2(n_425),
.B(n_417),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_441),
.A2(n_456),
.B(n_469),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_443),
.A2(n_448),
.B1(n_467),
.B2(n_432),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g494 ( 
.A(n_444),
.B(n_419),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_422),
.B(n_372),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_445),
.B(n_452),
.Y(n_490)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_418),
.Y(n_446)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_446),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_408),
.A2(n_364),
.B1(n_382),
.B2(n_400),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g449 ( 
.A(n_434),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_449),
.B(n_450),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_435),
.B(n_388),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_428),
.Y(n_451)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_451),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_422),
.B(n_372),
.Y(n_452)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_428),
.Y(n_454)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_454),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_411),
.A2(n_380),
.B1(n_375),
.B2(n_396),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_455),
.A2(n_457),
.B1(n_405),
.B2(n_419),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_411),
.A2(n_385),
.B1(n_392),
.B2(n_386),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_435),
.B(n_385),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_458),
.B(n_464),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_407),
.B(n_398),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_459),
.B(n_470),
.Y(n_475)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_429),
.Y(n_460)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_460),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_439),
.B(n_370),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_461),
.B(n_463),
.C(n_470),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_404),
.B(n_362),
.Y(n_462)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_462),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_424),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_410),
.Y(n_465)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_465),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_424),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_466),
.B(n_471),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_410),
.A2(n_360),
.B1(n_368),
.B2(n_366),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_429),
.Y(n_468)
);

INVxp33_ASAP7_75t_L g487 ( 
.A(n_468),
.Y(n_487)
);

A2O1A1O1Ixp25_ASAP7_75t_L g469 ( 
.A1(n_412),
.A2(n_438),
.B(n_409),
.C(n_414),
.D(n_413),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_437),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_404),
.B(n_308),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_472),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_438),
.B(n_421),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_473),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_425),
.A2(n_415),
.B(n_433),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_474),
.A2(n_453),
.B(n_455),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_444),
.B(n_440),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_477),
.B(n_481),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_479),
.B(n_489),
.Y(n_528)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_446),
.Y(n_480)
);

CKINVDCx14_ASAP7_75t_R g525 ( 
.A(n_480),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_447),
.B(n_420),
.C(n_431),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_483),
.B(n_463),
.C(n_459),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_441),
.A2(n_453),
.B(n_456),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_484),
.A2(n_491),
.B(n_504),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_443),
.A2(n_426),
.B1(n_405),
.B2(n_423),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_485),
.B(n_497),
.Y(n_508)
);

A2O1A1Ixp33_ASAP7_75t_SL g486 ( 
.A1(n_442),
.A2(n_431),
.B(n_423),
.C(n_430),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_486),
.A2(n_457),
.B(n_467),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_489),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_449),
.A2(n_427),
.B1(n_436),
.B2(n_416),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_442),
.A2(n_448),
.B1(n_465),
.B2(n_454),
.Y(n_492)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_492),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_494),
.B(n_492),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_474),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_451),
.A2(n_427),
.B1(n_436),
.B2(n_416),
.Y(n_498)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_498),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_464),
.A2(n_466),
.B1(n_458),
.B2(n_450),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_500),
.B(n_495),
.Y(n_522)
);

NAND3xp33_ASAP7_75t_L g506 ( 
.A(n_476),
.B(n_471),
.C(n_447),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_506),
.B(n_507),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_475),
.B(n_461),
.Y(n_507)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_509),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_511),
.B(n_516),
.C(n_520),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_484),
.A2(n_469),
.B(n_468),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_512),
.A2(n_479),
.B(n_502),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_480),
.B(n_460),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_513),
.Y(n_532)
);

XNOR2x1_ASAP7_75t_L g515 ( 
.A(n_494),
.B(n_499),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_SL g541 ( 
.A(n_515),
.B(n_521),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_475),
.B(n_483),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_481),
.B(n_477),
.C(n_499),
.Y(n_520)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_522),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_478),
.B(n_488),
.C(n_482),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_523),
.B(n_527),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_495),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_524),
.Y(n_548)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_496),
.Y(n_526)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_526),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_485),
.B(n_505),
.C(n_496),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_528),
.A2(n_497),
.B1(n_504),
.B2(n_493),
.Y(n_533)
);

CKINVDCx14_ASAP7_75t_R g529 ( 
.A(n_490),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_529),
.B(n_530),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_500),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_533),
.A2(n_543),
.B1(n_509),
.B2(n_510),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_525),
.B(n_487),
.Y(n_537)
);

OAI21xp33_ASAP7_75t_SL g561 ( 
.A1(n_537),
.A2(n_539),
.B(n_517),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_522),
.B(n_487),
.Y(n_539)
);

FAx1_ASAP7_75t_L g540 ( 
.A(n_514),
.B(n_486),
.CI(n_493),
.CON(n_540),
.SN(n_540)
);

OAI21xp5_ASAP7_75t_SL g551 ( 
.A1(n_540),
.A2(n_508),
.B(n_514),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_L g563 ( 
.A1(n_542),
.A2(n_503),
.B(n_520),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_527),
.A2(n_486),
.B1(n_491),
.B2(n_498),
.Y(n_543)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_523),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_526),
.Y(n_547)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_547),
.Y(n_559)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_519),
.Y(n_549)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_549),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_546),
.B(n_501),
.Y(n_550)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_550),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_551),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_542),
.A2(n_517),
.B1(n_510),
.B2(n_528),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_552),
.Y(n_568)
);

OAI21x1_ASAP7_75t_L g553 ( 
.A1(n_531),
.A2(n_512),
.B(n_521),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_553),
.B(n_558),
.C(n_560),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_537),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_554),
.B(n_557),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_555),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_545),
.B(n_516),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_545),
.B(n_507),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_SL g560 ( 
.A1(n_543),
.A2(n_528),
.B1(n_519),
.B2(n_508),
.Y(n_560)
);

AOI211xp5_ASAP7_75t_L g573 ( 
.A1(n_561),
.A2(n_562),
.B(n_540),
.C(n_533),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_548),
.A2(n_486),
.B1(n_515),
.B2(n_503),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_563),
.B(n_564),
.C(n_536),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_535),
.A2(n_511),
.B1(n_518),
.B2(n_548),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_557),
.B(n_531),
.C(n_518),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_566),
.B(n_573),
.Y(n_583)
);

OAI21xp5_ASAP7_75t_SL g569 ( 
.A1(n_564),
.A2(n_534),
.B(n_536),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_569),
.A2(n_551),
.B(n_540),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_574),
.B(n_535),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_558),
.B(n_532),
.C(n_549),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_575),
.B(n_563),
.Y(n_576)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_576),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_571),
.B(n_532),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_577),
.B(n_559),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_566),
.B(n_570),
.C(n_572),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_578),
.B(n_568),
.Y(n_589)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_565),
.B(n_555),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_579),
.B(n_580),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_580),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_L g584 ( 
.A1(n_581),
.A2(n_582),
.B(n_567),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_SL g582 ( 
.A1(n_567),
.A2(n_540),
.B(n_556),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_L g592 ( 
.A1(n_584),
.A2(n_583),
.B(n_586),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_585),
.B(n_587),
.Y(n_591)
);

CKINVDCx14_ASAP7_75t_R g590 ( 
.A(n_589),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_592),
.B(n_588),
.Y(n_593)
);

OAI21x1_ASAP7_75t_SL g595 ( 
.A1(n_593),
.A2(n_594),
.B(n_590),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_SL g594 ( 
.A1(n_591),
.A2(n_587),
.B(n_556),
.Y(n_594)
);

OAI321xp33_ASAP7_75t_L g596 ( 
.A1(n_595),
.A2(n_547),
.A3(n_544),
.B1(n_539),
.B2(n_538),
.C(n_579),
.Y(n_596)
);

OAI21xp5_ASAP7_75t_L g597 ( 
.A1(n_596),
.A2(n_544),
.B(n_538),
.Y(n_597)
);

XOR2xp5_ASAP7_75t_L g598 ( 
.A(n_597),
.B(n_562),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_598),
.A2(n_552),
.B(n_541),
.Y(n_599)
);


endmodule