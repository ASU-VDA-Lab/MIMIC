module fake_jpeg_8164_n_76 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_76);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_76;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_67;
wire n_75;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx11_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx5p33_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_11),
.B(n_1),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_27),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_18),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_24),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_21),
.B(n_26),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_29),
.B(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_25),
.A2(n_15),
.B(n_20),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_22),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_39),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_28),
.C(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_40),
.B(n_39),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_18),
.B1(n_20),
.B2(n_19),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_13),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_12),
.B1(n_19),
.B2(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_45),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_32),
.A2(n_12),
.B1(n_17),
.B2(n_14),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_14),
.Y(n_53)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_48),
.A2(n_46),
.B1(n_40),
.B2(n_37),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_SL g60 ( 
.A(n_49),
.B(n_8),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_51),
.A2(n_53),
.B1(n_2),
.B2(n_3),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_54),
.B(n_55),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_33),
.Y(n_55)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_61),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_48),
.A2(n_37),
.B1(n_22),
.B2(n_8),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_50),
.A2(n_6),
.B1(n_7),
.B2(n_52),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_49),
.B(n_57),
.Y(n_66)
);

NOR3xp33_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_62),
.C(n_6),
.Y(n_70)
);

BUFx24_ASAP7_75t_SL g67 ( 
.A(n_63),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_68),
.C(n_59),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_60),
.C(n_57),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_70),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_7),
.C(n_65),
.Y(n_71)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_72),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_74),
.B(n_72),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);


endmodule