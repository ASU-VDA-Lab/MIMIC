module fake_jpeg_30706_n_118 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_118);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_118;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_32),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_20),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_25),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_52),
.Y(n_57)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_42),
.B(n_0),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_63),
.Y(n_69)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_42),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_36),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_54),
.A2(n_41),
.B1(n_43),
.B2(n_46),
.Y(n_66)
);

OR2x6_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_1),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_57),
.B(n_65),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_67),
.B(n_5),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_45),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_72),
.C(n_3),
.Y(n_81)
);

MAJx2_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_40),
.C(n_36),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_55),
.B(n_39),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_75),
.Y(n_85)
);

NAND2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_40),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_74),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_33),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_78),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_56),
.B(n_35),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_1),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_80),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_2),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_90),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_4),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_84),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_16),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_6),
.C(n_7),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_74),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_71),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_87),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_5),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_73),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_95),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_67),
.B(n_6),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_93),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_100),
.B(n_85),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_97),
.C(n_105),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_92),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_103),
.A2(n_104),
.B(n_13),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_89),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_106),
.A2(n_109),
.B1(n_89),
.B2(n_88),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_108),
.A2(n_98),
.B1(n_94),
.B2(n_96),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_110),
.B(n_111),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_107),
.B(n_101),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_113),
.B(n_99),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_114),
.A2(n_102),
.B1(n_17),
.B2(n_18),
.Y(n_115)
);

NAND3xp33_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_15),
.C(n_21),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_22),
.B(n_23),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_27),
.Y(n_118)
);


endmodule