module real_aes_5738_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_971, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_969, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_973, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_972, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_970, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_971;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_969;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_973;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_972;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_970;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_919;
wire n_857;
wire n_461;
wire n_908;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_955;
wire n_889;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_961;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_281;
wire n_496;
wire n_962;
wire n_693;
wire n_468;
wire n_755;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_725;
wire n_504;
wire n_455;
wire n_960;
wire n_671;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_940;
wire n_770;
wire n_808;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_296;
wire n_702;
wire n_954;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_749;
wire n_358;
wire n_275;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_939;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_926;
wire n_922;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_959;
wire n_715;
wire n_946;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_967;
wire n_566;
wire n_719;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_259;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_0), .A2(n_446), .B(n_449), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_1), .A2(n_136), .B1(n_378), .B2(n_379), .Y(n_377) );
INVx1_ASAP7_75t_L g473 ( .A(n_2), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_3), .A2(n_51), .B1(n_732), .B2(n_735), .Y(n_740) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_4), .A2(n_7), .B1(n_398), .B2(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g513 ( .A(n_5), .Y(n_513) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_6), .Y(n_690) );
AND2x4_ASAP7_75t_L g705 ( .A(n_6), .B(n_706), .Y(n_705) );
AND2x4_ASAP7_75t_L g715 ( .A(n_6), .B(n_242), .Y(n_715) );
AOI221x1_ASAP7_75t_L g540 ( .A1(n_8), .A2(n_70), .B1(n_448), .B2(n_541), .C(n_542), .Y(n_540) );
INVx1_ASAP7_75t_L g638 ( .A(n_9), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_10), .A2(n_55), .B1(n_317), .B2(n_433), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_11), .A2(n_99), .B1(n_506), .B2(n_507), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_12), .A2(n_202), .B1(n_396), .B2(n_428), .Y(n_930) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_13), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_14), .A2(n_79), .B1(n_260), .B2(n_437), .Y(n_931) );
AOI22xp5_ASAP7_75t_L g738 ( .A1(n_15), .A2(n_77), .B1(n_725), .B2(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g330 ( .A(n_16), .Y(n_330) );
INVx1_ASAP7_75t_L g712 ( .A(n_17), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_18), .A2(n_80), .B1(n_371), .B2(n_374), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_19), .A2(n_237), .B1(n_452), .B2(n_587), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_20), .A2(n_82), .B1(n_430), .B2(n_491), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g302 ( .A1(n_21), .A2(n_87), .B1(n_303), .B2(n_310), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_22), .A2(n_147), .B1(n_454), .B2(n_456), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g558 ( .A(n_23), .Y(n_558) );
INVx1_ASAP7_75t_L g679 ( .A(n_24), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_25), .B(n_590), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_26), .A2(n_218), .B1(n_365), .B2(n_366), .Y(n_364) );
AOI22xp33_ASAP7_75t_SL g547 ( .A1(n_27), .A2(n_58), .B1(n_430), .B2(n_491), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_28), .A2(n_104), .B1(n_357), .B2(n_408), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_29), .A2(n_68), .B1(n_647), .B2(n_648), .Y(n_646) );
INVx1_ASAP7_75t_SL g781 ( .A(n_30), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_31), .A2(n_76), .B1(n_718), .B2(n_748), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_32), .A2(n_161), .B1(n_590), .B2(n_650), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_33), .A2(n_157), .B1(n_283), .B2(n_488), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_34), .A2(n_84), .B1(n_398), .B2(n_668), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_35), .A2(n_245), .B1(n_357), .B2(n_515), .Y(n_674) );
INVx1_ASAP7_75t_L g925 ( .A(n_36), .Y(n_925) );
INVx1_ASAP7_75t_L g280 ( .A(n_37), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_37), .B(n_186), .Y(n_337) );
INVxp67_ASAP7_75t_L g356 ( .A(n_37), .Y(n_356) );
AOI221xp5_ASAP7_75t_L g635 ( .A1(n_38), .A2(n_41), .B1(n_441), .B2(n_636), .C(n_637), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_39), .A2(n_206), .B1(n_593), .B2(n_594), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_40), .A2(n_85), .B1(n_702), .B2(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g476 ( .A(n_42), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_43), .A2(n_45), .B1(n_401), .B2(n_403), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g427 ( .A1(n_44), .A2(n_201), .B1(n_428), .B2(n_429), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_46), .B(n_454), .Y(n_611) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_47), .B(n_265), .Y(n_275) );
INVx1_ASAP7_75t_L g464 ( .A(n_48), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_49), .A2(n_162), .B1(n_466), .B2(n_583), .Y(n_582) );
AOI21xp33_ASAP7_75t_L g414 ( .A1(n_50), .A2(n_342), .B(n_415), .Y(n_414) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_52), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_53), .A2(n_248), .B1(n_714), .B2(n_749), .Y(n_769) );
INVxp67_ASAP7_75t_R g716 ( .A(n_54), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_56), .A2(n_244), .B1(n_283), .B2(n_438), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_57), .A2(n_148), .B1(n_310), .B2(n_428), .Y(n_651) );
INVx2_ASAP7_75t_L g688 ( .A(n_59), .Y(n_688) );
INVx1_ASAP7_75t_L g704 ( .A(n_60), .Y(n_704) );
AND2x4_ASAP7_75t_L g709 ( .A(n_60), .B(n_688), .Y(n_709) );
INVx1_ASAP7_75t_SL g726 ( .A(n_60), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_61), .A2(n_173), .B1(n_408), .B2(n_413), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_62), .A2(n_180), .B1(n_260), .B2(n_283), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_63), .A2(n_235), .B1(n_405), .B2(n_486), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_64), .A2(n_158), .B1(n_408), .B2(n_921), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_65), .A2(n_144), .B1(n_625), .B2(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g470 ( .A(n_66), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g314 ( .A1(n_67), .A2(n_214), .B1(n_315), .B2(n_317), .Y(n_314) );
INVx1_ASAP7_75t_L g613 ( .A(n_69), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_71), .A2(n_191), .B1(n_298), .B2(n_435), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_72), .A2(n_210), .B1(n_433), .B2(n_625), .Y(n_624) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_73), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_74), .A2(n_126), .B1(n_283), .B2(n_433), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_75), .A2(n_176), .B1(n_725), .B2(n_739), .Y(n_743) );
INVx1_ASAP7_75t_L g457 ( .A(n_77), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_78), .B(n_381), .Y(n_380) );
AOI21xp5_ASAP7_75t_L g922 ( .A1(n_81), .A2(n_923), .B(n_924), .Y(n_922) );
XOR2x2_ASAP7_75t_L g579 ( .A(n_83), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_SL g539 ( .A(n_85), .Y(n_539) );
NOR3xp33_ASAP7_75t_L g566 ( .A(n_85), .B(n_567), .C(n_568), .Y(n_566) );
OAI22xp5_ASAP7_75t_R g939 ( .A1(n_86), .A2(n_940), .B1(n_941), .B2(n_942), .Y(n_939) );
CKINVDCx5p33_ASAP7_75t_R g940 ( .A(n_86), .Y(n_940) );
CKINVDCx16_ASAP7_75t_R g710 ( .A(n_88), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_89), .A2(n_163), .B1(n_702), .B2(n_800), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_90), .A2(n_156), .B1(n_647), .B2(n_919), .Y(n_918) );
AOI22xp5_ASAP7_75t_L g341 ( .A1(n_91), .A2(n_170), .B1(n_342), .B2(n_344), .Y(n_341) );
INVx1_ASAP7_75t_L g266 ( .A(n_92), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_92), .B(n_184), .Y(n_353) );
AOI33xp33_ASAP7_75t_R g598 ( .A1(n_93), .A2(n_216), .A3(n_262), .B1(n_286), .B2(n_599), .B3(n_971), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_94), .A2(n_212), .B1(n_524), .B2(n_525), .Y(n_523) );
INVx1_ASAP7_75t_L g467 ( .A(n_95), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_96), .A2(n_229), .B1(n_961), .B2(n_962), .Y(n_960) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_97), .A2(n_174), .B1(n_303), .B2(n_396), .Y(n_671) );
AOI21xp5_ASAP7_75t_SL g324 ( .A1(n_98), .A2(n_325), .B(n_329), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_100), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_101), .A2(n_227), .B1(n_303), .B2(n_530), .Y(n_595) );
INVx1_ASAP7_75t_L g633 ( .A(n_102), .Y(n_633) );
OAI222xp33_ASAP7_75t_L g644 ( .A1(n_102), .A2(n_645), .B1(n_651), .B2(n_652), .C1(n_972), .C2(n_973), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_102), .B(n_652), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g359 ( .A(n_103), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_105), .A2(n_238), .B1(n_317), .B2(n_433), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_106), .A2(n_195), .B1(n_405), .B2(n_486), .Y(n_672) );
INVx1_ASAP7_75t_L g957 ( .A(n_107), .Y(n_957) );
INVx1_ASAP7_75t_L g392 ( .A(n_108), .Y(n_392) );
INVx1_ASAP7_75t_L g727 ( .A(n_109), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_110), .A2(n_164), .B1(n_748), .B2(n_749), .Y(n_747) );
INVx1_ASAP7_75t_L g955 ( .A(n_111), .Y(n_955) );
AOI21xp33_ASAP7_75t_L g677 ( .A1(n_112), .A2(n_383), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g388 ( .A(n_113), .Y(n_388) );
INVx1_ASAP7_75t_L g618 ( .A(n_114), .Y(n_618) );
AOI21xp33_ASAP7_75t_L g385 ( .A1(n_115), .A2(n_386), .B(n_387), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_116), .A2(n_138), .B1(n_372), .B2(n_375), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_117), .A2(n_239), .B1(n_371), .B2(n_372), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_118), .A2(n_199), .B1(n_396), .B2(n_428), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_119), .A2(n_142), .B1(n_298), .B2(n_398), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_120), .A2(n_137), .B1(n_403), .B2(n_438), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_121), .A2(n_226), .B1(n_260), .B2(n_283), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_122), .A2(n_197), .B1(n_298), .B2(n_524), .Y(n_928) );
AOI22x1_ASAP7_75t_L g602 ( .A1(n_123), .A2(n_603), .B1(n_604), .B2(n_627), .Y(n_602) );
INVx1_ASAP7_75t_L g627 ( .A(n_123), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_124), .A2(n_219), .B1(n_298), .B2(n_435), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_125), .A2(n_188), .B1(n_348), .B2(n_413), .Y(n_412) );
AO22x1_ASAP7_75t_L g643 ( .A1(n_127), .A2(n_129), .B1(n_435), .B2(n_438), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_128), .A2(n_172), .B1(n_374), .B2(n_375), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_130), .A2(n_135), .B1(n_310), .B2(n_428), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_131), .A2(n_146), .B1(n_368), .B2(n_369), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_132), .A2(n_139), .B1(n_528), .B2(n_529), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_133), .B(n_590), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_134), .A2(n_166), .B1(n_714), .B2(n_718), .Y(n_783) );
INVx1_ASAP7_75t_L g450 ( .A(n_140), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_141), .A2(n_321), .B(n_608), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_143), .A2(n_160), .B1(n_488), .B2(n_670), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_145), .A2(n_217), .B1(n_520), .B2(n_522), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_149), .A2(n_243), .B1(n_294), .B2(n_298), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_150), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g730 ( .A(n_151), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_152), .A2(n_179), .B1(n_315), .B2(n_405), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_153), .A2(n_224), .B1(n_732), .B2(n_735), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_154), .B(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g728 ( .A(n_155), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_159), .A2(n_200), .B1(n_480), .B2(n_481), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_165), .A2(n_187), .B1(n_357), .B2(n_585), .Y(n_584) );
XOR2xp5_ASAP7_75t_L g915 ( .A(n_166), .B(n_916), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_166), .A2(n_937), .B1(n_939), .B2(n_963), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_167), .B(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_168), .B(n_452), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_169), .A2(n_247), .B1(n_437), .B2(n_438), .Y(n_436) );
OA22x2_ASAP7_75t_L g270 ( .A1(n_171), .A2(n_186), .B1(n_265), .B2(n_269), .Y(n_270) );
INVx1_ASAP7_75t_L g290 ( .A(n_171), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g553 ( .A(n_175), .Y(n_553) );
AO22x2_ASAP7_75t_L g458 ( .A1(n_176), .A2(n_459), .B1(n_460), .B2(n_461), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_176), .Y(n_459) );
AND2x2_ASAP7_75t_L g542 ( .A(n_177), .B(n_543), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_178), .A2(n_198), .B1(n_433), .B2(n_625), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_181), .A2(n_228), .B1(n_344), .B2(n_504), .Y(n_503) );
CKINVDCx6p67_ASAP7_75t_R g707 ( .A(n_182), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_183), .B(n_481), .Y(n_926) );
INVx1_ASAP7_75t_L g282 ( .A(n_184), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_184), .B(n_288), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_185), .A2(n_209), .B1(n_383), .B2(n_384), .Y(n_382) );
OAI21xp33_ASAP7_75t_L g291 ( .A1(n_186), .A2(n_205), .B(n_292), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_189), .A2(n_204), .B1(n_298), .B2(n_398), .Y(n_622) );
XNOR2x1_ASAP7_75t_L g361 ( .A(n_190), .B(n_362), .Y(n_361) );
XNOR2x2_ASAP7_75t_SL g389 ( .A(n_190), .B(n_362), .Y(n_389) );
INVx1_ASAP7_75t_L g500 ( .A(n_192), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_193), .A2(n_222), .B1(n_365), .B2(n_398), .Y(n_538) );
INVx1_ASAP7_75t_L g664 ( .A(n_194), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_196), .A2(n_246), .B1(n_702), .B2(n_751), .Y(n_770) );
INVx1_ASAP7_75t_L g950 ( .A(n_203), .Y(n_950) );
INVx1_ASAP7_75t_L g268 ( .A(n_205), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_205), .B(n_236), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_207), .A2(n_232), .B1(n_486), .B2(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g951 ( .A(n_208), .Y(n_951) );
INVx1_ASAP7_75t_L g782 ( .A(n_211), .Y(n_782) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_213), .A2(n_509), .B(n_512), .Y(n_508) );
INVx1_ASAP7_75t_L g959 ( .A(n_215), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_220), .A2(n_233), .B1(n_303), .B2(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_221), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g615 ( .A(n_223), .Y(n_615) );
INVx1_ASAP7_75t_L g609 ( .A(n_225), .Y(n_609) );
INVx1_ASAP7_75t_L g416 ( .A(n_230), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_231), .A2(n_240), .B1(n_441), .B2(n_442), .Y(n_440) );
AOI22x1_ASAP7_75t_L g347 ( .A1(n_234), .A2(n_241), .B1(n_348), .B2(n_357), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_236), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g706 ( .A(n_242), .Y(n_706) );
HB1xp67_ASAP7_75t_L g966 ( .A(n_242), .Y(n_966) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_683), .B(n_691), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_419), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AOI21xp33_ASAP7_75t_L g683 ( .A1(n_252), .A2(n_420), .B(n_684), .Y(n_683) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
XOR2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_390), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_256), .B1(n_360), .B2(n_389), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
XNOR2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_359), .Y(n_256) );
NOR3xp33_ASAP7_75t_SL g257 ( .A(n_258), .B(n_301), .C(n_319), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_293), .Y(n_258) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
BUFx8_ASAP7_75t_L g438 ( .A(n_261), .Y(n_438) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_271), .Y(n_261) );
AND2x4_ASAP7_75t_L g295 ( .A(n_262), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g323 ( .A(n_262), .B(n_312), .Y(n_323) );
AND2x2_ASAP7_75t_L g358 ( .A(n_262), .B(n_308), .Y(n_358) );
AND2x4_ASAP7_75t_L g365 ( .A(n_262), .B(n_271), .Y(n_365) );
AND2x4_ASAP7_75t_L g366 ( .A(n_262), .B(n_300), .Y(n_366) );
AND2x4_ASAP7_75t_L g378 ( .A(n_262), .B(n_308), .Y(n_378) );
AND2x2_ASAP7_75t_L g383 ( .A(n_262), .B(n_312), .Y(n_383) );
AND2x2_ASAP7_75t_L g402 ( .A(n_262), .B(n_271), .Y(n_402) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_270), .Y(n_262) );
INVx1_ASAP7_75t_L g306 ( .A(n_263), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_267), .Y(n_263) );
NAND2xp33_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g269 ( .A(n_265), .Y(n_269) );
INVx3_ASAP7_75t_L g274 ( .A(n_265), .Y(n_274) );
NAND2xp33_ASAP7_75t_L g281 ( .A(n_265), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g292 ( .A(n_265), .Y(n_292) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_265), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_266), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
OAI21xp5_ASAP7_75t_L g355 ( .A1(n_268), .A2(n_292), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g307 ( .A(n_270), .Y(n_307) );
AND2x2_ASAP7_75t_L g328 ( .A(n_270), .B(n_306), .Y(n_328) );
AND2x2_ASAP7_75t_L g354 ( .A(n_270), .B(n_355), .Y(n_354) );
AND2x4_ASAP7_75t_L g285 ( .A(n_271), .B(n_286), .Y(n_285) );
AND2x4_ASAP7_75t_L g316 ( .A(n_271), .B(n_305), .Y(n_316) );
AND2x4_ASAP7_75t_L g371 ( .A(n_271), .B(n_305), .Y(n_371) );
AND2x4_ASAP7_75t_L g374 ( .A(n_271), .B(n_286), .Y(n_374) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_271), .Y(n_599) );
AND2x4_ASAP7_75t_L g271 ( .A(n_272), .B(n_276), .Y(n_271) );
OR2x2_ASAP7_75t_L g297 ( .A(n_272), .B(n_277), .Y(n_297) );
AND2x4_ASAP7_75t_L g308 ( .A(n_272), .B(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g313 ( .A(n_272), .Y(n_313) );
AND2x2_ASAP7_75t_L g351 ( .A(n_272), .B(n_352), .Y(n_351) );
AND2x4_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_274), .B(n_280), .Y(n_279) );
INVxp67_ASAP7_75t_L g288 ( .A(n_274), .Y(n_288) );
NAND3xp33_ASAP7_75t_L g339 ( .A(n_275), .B(n_287), .C(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g309 ( .A(n_278), .Y(n_309) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
INVx4_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx4_ASAP7_75t_L g403 ( .A(n_284), .Y(n_403) );
INVx4_ASAP7_75t_L g437 ( .A(n_284), .Y(n_437) );
INVx2_ASAP7_75t_SL g670 ( .A(n_284), .Y(n_670) );
INVx8_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x4_ASAP7_75t_L g299 ( .A(n_286), .B(n_300), .Y(n_299) );
AND2x4_ASAP7_75t_L g346 ( .A(n_286), .B(n_312), .Y(n_346) );
AND2x4_ASAP7_75t_L g375 ( .A(n_286), .B(n_300), .Y(n_375) );
AND2x4_ASAP7_75t_L g384 ( .A(n_286), .B(n_312), .Y(n_384) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_291), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
BUFx12f_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_295), .Y(n_398) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_295), .Y(n_435) );
BUFx3_ASAP7_75t_L g524 ( .A(n_295), .Y(n_524) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_295), .Y(n_594) );
AND2x4_ASAP7_75t_L g372 ( .A(n_296), .B(n_305), .Y(n_372) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g300 ( .A(n_297), .Y(n_300) );
BUFx12f_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx6_ASAP7_75t_L g495 ( .A(n_299), .Y(n_495) );
AND2x4_ASAP7_75t_L g318 ( .A(n_300), .B(n_305), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_314), .Y(n_301) );
BUFx12f_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_304), .Y(n_428) );
INVx3_ASAP7_75t_L g492 ( .A(n_304), .Y(n_492) );
AND2x4_ASAP7_75t_L g304 ( .A(n_305), .B(n_308), .Y(n_304) );
AND2x2_ASAP7_75t_L g311 ( .A(n_305), .B(n_312), .Y(n_311) );
AND2x4_ASAP7_75t_L g368 ( .A(n_305), .B(n_308), .Y(n_368) );
AND2x4_ASAP7_75t_L g369 ( .A(n_305), .B(n_312), .Y(n_369) );
AND2x4_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
AND2x4_ASAP7_75t_L g327 ( .A(n_308), .B(n_328), .Y(n_327) );
AND2x4_ASAP7_75t_L g386 ( .A(n_308), .B(n_328), .Y(n_386) );
AND2x4_ASAP7_75t_L g312 ( .A(n_309), .B(n_313), .Y(n_312) );
BUFx5_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_311), .Y(n_396) );
INVx1_ASAP7_75t_L g431 ( .A(n_311), .Y(n_431) );
BUFx3_ASAP7_75t_L g530 ( .A(n_311), .Y(n_530) );
AND2x4_ASAP7_75t_L g343 ( .A(n_312), .B(n_328), .Y(n_343) );
AND2x2_ASAP7_75t_L g381 ( .A(n_312), .B(n_328), .Y(n_381) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_316), .Y(n_433) );
BUFx12f_ASAP7_75t_L g486 ( .A(n_316), .Y(n_486) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_318), .Y(n_405) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_318), .Y(n_597) );
BUFx6f_ASAP7_75t_L g625 ( .A(n_318), .Y(n_625) );
NAND4xp25_ASAP7_75t_L g319 ( .A(n_320), .B(n_324), .C(n_341), .D(n_347), .Y(n_319) );
INVx3_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g410 ( .A(n_322), .Y(n_410) );
INVx2_ASAP7_75t_L g448 ( .A(n_322), .Y(n_448) );
INVx2_ASAP7_75t_L g511 ( .A(n_322), .Y(n_511) );
INVx3_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
BUFx3_ASAP7_75t_L g478 ( .A(n_323), .Y(n_478) );
INVx2_ASAP7_75t_L g588 ( .A(n_323), .Y(n_588) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g919 ( .A(n_326), .Y(n_919) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx3_ASAP7_75t_L g413 ( .A(n_327), .Y(n_413) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_327), .Y(n_441) );
BUFx3_ASAP7_75t_L g466 ( .A(n_327), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_331), .B(n_679), .Y(n_678) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_332), .B(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g452 ( .A(n_332), .Y(n_452) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_332), .Y(n_482) );
INVx2_ASAP7_75t_SL g962 ( .A(n_332), .Y(n_962) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx3_ASAP7_75t_L g418 ( .A(n_333), .Y(n_418) );
AO21x2_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_336), .B(n_339), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_335), .B(n_353), .Y(n_352) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_336), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g455 ( .A(n_343), .Y(n_455) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_343), .Y(n_472) );
BUFx8_ASAP7_75t_SL g541 ( .A(n_343), .Y(n_541) );
BUFx3_ASAP7_75t_L g590 ( .A(n_343), .Y(n_590) );
INVx2_ASAP7_75t_L g956 ( .A(n_343), .Y(n_956) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx3_ASAP7_75t_L g456 ( .A(n_345), .Y(n_456) );
INVx2_ASAP7_75t_L g583 ( .A(n_345), .Y(n_583) );
INVx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_346), .Y(n_408) );
BUFx6f_ASAP7_75t_L g650 ( .A(n_346), .Y(n_650) );
INVx4_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OAI21xp5_ASAP7_75t_L g449 ( .A1(n_349), .A2(n_450), .B(n_451), .Y(n_449) );
INVx3_ASAP7_75t_L g620 ( .A(n_349), .Y(n_620) );
INVx2_ASAP7_75t_L g648 ( .A(n_349), .Y(n_648) );
INVx2_ASAP7_75t_L g961 ( .A(n_349), .Y(n_961) );
INVx5_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx4f_ASAP7_75t_L g515 ( .A(n_350), .Y(n_515) );
BUFx2_ASAP7_75t_L g585 ( .A(n_350), .Y(n_585) );
AND2x4_ASAP7_75t_L g350 ( .A(n_351), .B(n_354), .Y(n_350) );
AND2x4_ASAP7_75t_L g379 ( .A(n_351), .B(n_354), .Y(n_379) );
AND2x2_ASAP7_75t_L g480 ( .A(n_351), .B(n_354), .Y(n_480) );
INVx3_ASAP7_75t_L g468 ( .A(n_357), .Y(n_468) );
BUFx3_ASAP7_75t_L g507 ( .A(n_357), .Y(n_507) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g444 ( .A(n_358), .Y(n_444) );
BUFx3_ASAP7_75t_L g647 ( .A(n_358), .Y(n_647) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_376), .Y(n_362) );
NAND4xp25_ASAP7_75t_L g363 ( .A(n_364), .B(n_367), .C(n_370), .D(n_373), .Y(n_363) );
NAND4xp25_ASAP7_75t_L g376 ( .A(n_377), .B(n_380), .C(n_382), .D(n_385), .Y(n_376) );
INVx2_ASAP7_75t_L g561 ( .A(n_378), .Y(n_561) );
INVx4_ASAP7_75t_L g554 ( .A(n_379), .Y(n_554) );
INVx2_ASAP7_75t_L g556 ( .A(n_384), .Y(n_556) );
INVx2_ASAP7_75t_L g559 ( .A(n_386), .Y(n_559) );
BUFx3_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
XNOR2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
NOR4xp75_ASAP7_75t_L g393 ( .A(n_394), .B(n_399), .C(n_406), .D(n_411), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_397), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_404), .Y(n_399) );
BUFx6f_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx4f_ASAP7_75t_L g488 ( .A(n_402), .Y(n_488) );
BUFx3_ASAP7_75t_L g522 ( .A(n_405), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_407), .B(n_409), .Y(n_406) );
INVx3_ASAP7_75t_L g474 ( .A(n_408), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_412), .B(n_414), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
INVx1_ASAP7_75t_L g517 ( .A(n_417), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_417), .B(n_638), .Y(n_637) );
INVx4_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx3_ASAP7_75t_L g544 ( .A(n_418), .Y(n_544) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
XNOR2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_573), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_498), .B1(n_571), .B2(n_572), .Y(n_421) );
BUFx2_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
INVxp67_ASAP7_75t_L g572 ( .A(n_423), .Y(n_572) );
AO22x2_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_458), .B1(n_496), .B2(n_497), .Y(n_423) );
INVx1_ASAP7_75t_L g496 ( .A(n_424), .Y(n_496) );
XOR2x2_ASAP7_75t_L g424 ( .A(n_425), .B(n_457), .Y(n_424) );
NOR2x1_ASAP7_75t_L g425 ( .A(n_426), .B(n_439), .Y(n_425) );
NAND4xp25_ASAP7_75t_L g426 ( .A(n_427), .B(n_432), .C(n_434), .D(n_436), .Y(n_426) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NAND3xp33_ASAP7_75t_L g439 ( .A(n_440), .B(n_445), .C(n_453), .Y(n_439) );
INVx4_ASAP7_75t_L g614 ( .A(n_441), .Y(n_614) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OAI21xp33_ASAP7_75t_L g617 ( .A1(n_443), .A2(n_618), .B(n_619), .Y(n_617) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g953 ( .A(n_444), .Y(n_953) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx3_ASAP7_75t_L g610 ( .A(n_452), .Y(n_610) );
INVx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g921 ( .A(n_455), .Y(n_921) );
INVx1_ASAP7_75t_L g616 ( .A(n_456), .Y(n_616) );
INVx2_ASAP7_75t_L g497 ( .A(n_458), .Y(n_497) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_483), .Y(n_461) );
NOR3xp33_ASAP7_75t_SL g462 ( .A(n_463), .B(n_469), .C(n_475), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B1(n_467), .B2(n_468), .Y(n_463) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
BUFx2_ASAP7_75t_L g506 ( .A(n_466), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_471), .B1(n_473), .B2(n_474), .Y(n_469) );
INVx1_ASAP7_75t_L g504 ( .A(n_471), .Y(n_504) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
OAI21xp33_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_477), .B(n_479), .Y(n_475) );
INVx2_ASAP7_75t_L g636 ( .A(n_477), .Y(n_636) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_484), .B(n_489), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_487), .Y(n_484) );
INVx1_ASAP7_75t_L g521 ( .A(n_486), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_493), .Y(n_489) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g528 ( .A(n_492), .Y(n_528) );
INVx3_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g526 ( .A(n_495), .Y(n_526) );
INVx5_ASAP7_75t_L g593 ( .A(n_495), .Y(n_593) );
INVx1_ASAP7_75t_L g642 ( .A(n_495), .Y(n_642) );
INVx2_ASAP7_75t_L g668 ( .A(n_495), .Y(n_668) );
INVx1_ASAP7_75t_L g571 ( .A(n_498), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_532), .B1(n_569), .B2(n_570), .Y(n_498) );
INVx2_ASAP7_75t_SL g569 ( .A(n_499), .Y(n_569) );
XNOR2x1_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
OR2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_518), .Y(n_501) );
NAND3xp33_ASAP7_75t_SL g502 ( .A(n_503), .B(n_505), .C(n_508), .Y(n_502) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OAI21xp33_ASAP7_75t_L g958 ( .A1(n_510), .A2(n_959), .B(n_960), .Y(n_958) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
OAI21xp33_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B(n_516), .Y(n_512) );
INVx2_ASAP7_75t_SL g514 ( .A(n_515), .Y(n_514) );
NAND4xp25_ASAP7_75t_L g518 ( .A(n_519), .B(n_523), .C(n_527), .D(n_531), .Y(n_518) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
BUFx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g570 ( .A(n_532), .Y(n_570) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
BUFx3_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
NAND2x1_ASAP7_75t_L g535 ( .A(n_536), .B(n_562), .Y(n_535) );
NOR3xp33_ASAP7_75t_L g536 ( .A(n_537), .B(n_545), .C(n_549), .Y(n_536) );
OAI22xp33_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_539), .B1(n_540), .B2(n_969), .Y(n_537) );
INVx1_ASAP7_75t_L g567 ( .A(n_538), .Y(n_567) );
NOR2xp67_ASAP7_75t_L g545 ( .A(n_539), .B(n_546), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_539), .A2(n_550), .B1(n_551), .B2(n_970), .Y(n_549) );
INVx1_ASAP7_75t_L g564 ( .A(n_540), .Y(n_564) );
INVx4_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NAND3xp33_ASAP7_75t_L g562 ( .A(n_546), .B(n_563), .C(n_566), .Y(n_562) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
INVx1_ASAP7_75t_L g568 ( .A(n_550), .Y(n_568) );
INVx1_ASAP7_75t_L g565 ( .A(n_551), .Y(n_565) );
NOR2x1_ASAP7_75t_L g551 ( .A(n_552), .B(n_557), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_554), .B1(n_555), .B2(n_556), .Y(n_552) );
OAI21xp5_ASAP7_75t_L g924 ( .A1(n_554), .A2(n_925), .B(n_926), .Y(n_924) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_559), .B1(n_560), .B2(n_561), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_629), .B1(n_681), .B2(n_682), .Y(n_573) );
INVx1_ASAP7_75t_L g682 ( .A(n_574), .Y(n_682) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OAI21x1_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_600), .B(n_628), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_579), .B(n_602), .Y(n_628) );
NOR2x1_ASAP7_75t_L g580 ( .A(n_581), .B(n_591), .Y(n_580) );
NAND4xp25_ASAP7_75t_L g581 ( .A(n_582), .B(n_584), .C(n_586), .D(n_589), .Y(n_581) );
BUFx3_ASAP7_75t_L g923 ( .A(n_587), .Y(n_923) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NAND4xp25_ASAP7_75t_L g591 ( .A(n_592), .B(n_595), .C(n_596), .D(n_598), .Y(n_591) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_621), .Y(n_604) );
NOR3xp33_ASAP7_75t_L g605 ( .A(n_606), .B(n_612), .C(n_617), .Y(n_605) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_607), .B(n_611), .Y(n_606) );
NOR2xp33_ASAP7_75t_SL g608 ( .A(n_609), .B(n_610), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_614), .B1(n_615), .B2(n_616), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g949 ( .A1(n_614), .A2(n_950), .B1(n_951), .B2(n_952), .Y(n_949) );
OAI22xp5_ASAP7_75t_L g954 ( .A1(n_616), .A2(n_955), .B1(n_956), .B2(n_957), .Y(n_954) );
AND4x1_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .C(n_624), .D(n_626), .Y(n_621) );
INVx2_ASAP7_75t_SL g681 ( .A(n_629), .Y(n_681) );
OA22x2_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_631), .B1(n_660), .B2(n_680), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x4_ASAP7_75t_L g631 ( .A(n_632), .B(n_653), .Y(n_631) );
AOI21x1_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B(n_644), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_639), .Y(n_634) );
BUFx2_ASAP7_75t_L g654 ( .A(n_635), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_640), .B(n_643), .Y(n_639) );
INVxp67_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g658 ( .A(n_641), .B(n_651), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_643), .Y(n_659) );
INVx1_ASAP7_75t_L g657 ( .A(n_645), .Y(n_657) );
AND2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_649), .Y(n_645) );
NAND4xp75_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .C(n_658), .D(n_659), .Y(n_653) );
NOR2x1_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
INVx1_ASAP7_75t_L g680 ( .A(n_660), .Y(n_680) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
BUFx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
XNOR2x1_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .Y(n_662) );
CKINVDCx5p33_ASAP7_75t_R g663 ( .A(n_664), .Y(n_663) );
NOR2x1_ASAP7_75t_L g665 ( .A(n_666), .B(n_673), .Y(n_665) );
NAND4xp25_ASAP7_75t_L g666 ( .A(n_667), .B(n_669), .C(n_671), .D(n_672), .Y(n_666) );
NAND4xp25_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .C(n_676), .D(n_677), .Y(n_673) );
BUFx4_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
NAND3xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_689), .C(n_690), .Y(n_685) );
AND2x2_ASAP7_75t_L g933 ( .A(n_686), .B(n_934), .Y(n_933) );
AND2x2_ASAP7_75t_L g938 ( .A(n_686), .B(n_935), .Y(n_938) );
AOI21xp5_ASAP7_75t_L g967 ( .A1(n_686), .A2(n_690), .B(n_726), .Y(n_967) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AO21x1_ASAP7_75t_L g964 ( .A1(n_687), .A2(n_965), .B(n_967), .Y(n_964) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g703 ( .A(n_688), .B(n_704), .Y(n_703) );
AND3x4_ASAP7_75t_L g725 ( .A(n_688), .B(n_705), .C(n_726), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g934 ( .A(n_689), .B(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g935 ( .A(n_690), .Y(n_935) );
OAI221xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_912), .B1(n_914), .B2(n_932), .C(n_936), .Y(n_691) );
AND5x1_ASAP7_75t_L g692 ( .A(n_693), .B(n_856), .C(n_873), .D(n_882), .E(n_902), .Y(n_692) );
AOI222xp33_ASAP7_75t_SL g693 ( .A1(n_694), .A2(n_779), .B1(n_793), .B2(n_802), .C1(n_835), .C2(n_855), .Y(n_693) );
OAI221xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_773), .B1(n_779), .B2(n_784), .C(n_789), .Y(n_694) );
NOR3xp33_ASAP7_75t_L g695 ( .A(n_696), .B(n_752), .C(n_765), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_697), .B(n_719), .Y(n_696) );
AND2x2_ASAP7_75t_L g907 ( .A(n_697), .B(n_908), .Y(n_907) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
OAI221xp5_ASAP7_75t_L g752 ( .A1(n_698), .A2(n_753), .B1(n_758), .B2(n_762), .C(n_764), .Y(n_752) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_698), .B(n_830), .Y(n_829) );
BUFx2_ASAP7_75t_L g852 ( .A(n_698), .Y(n_852) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx3_ASAP7_75t_L g760 ( .A(n_699), .Y(n_760) );
AND2x2_ASAP7_75t_L g776 ( .A(n_699), .B(n_774), .Y(n_776) );
OR2x2_ASAP7_75t_L g810 ( .A(n_699), .B(n_768), .Y(n_810) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_699), .B(n_722), .Y(n_812) );
AND2x2_ASAP7_75t_L g824 ( .A(n_699), .B(n_768), .Y(n_824) );
OR2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_711), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_707), .B1(n_708), .B2(n_710), .Y(n_700) );
OAI221xp5_ASAP7_75t_L g780 ( .A1(n_701), .A2(n_708), .B1(n_781), .B2(n_782), .C(n_783), .Y(n_780) );
INVx3_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AND2x4_ASAP7_75t_L g702 ( .A(n_703), .B(n_705), .Y(n_702) );
AND2x4_ASAP7_75t_L g714 ( .A(n_703), .B(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g735 ( .A(n_703), .B(n_715), .Y(n_735) );
AND2x2_ASAP7_75t_L g748 ( .A(n_703), .B(n_715), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_705), .B(n_709), .Y(n_708) );
AND2x4_ASAP7_75t_L g739 ( .A(n_705), .B(n_709), .Y(n_739) );
AND2x4_ASAP7_75t_L g751 ( .A(n_705), .B(n_709), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_708), .A2(n_724), .B1(n_727), .B2(n_728), .Y(n_723) );
AND2x4_ASAP7_75t_L g718 ( .A(n_709), .B(n_715), .Y(n_718) );
AND2x2_ASAP7_75t_L g732 ( .A(n_709), .B(n_715), .Y(n_732) );
AND2x2_ASAP7_75t_L g749 ( .A(n_709), .B(n_715), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_713), .B1(n_716), .B2(n_717), .Y(n_711) );
INVx3_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
BUFx2_ASAP7_75t_L g913 ( .A(n_714), .Y(n_913) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NOR2xp33_ASAP7_75t_L g878 ( .A(n_719), .B(n_818), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_720), .B(n_736), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_720), .B(n_755), .Y(n_764) );
NOR2xp33_ASAP7_75t_L g831 ( .A(n_720), .B(n_818), .Y(n_831) );
NOR2xp33_ASAP7_75t_L g894 ( .A(n_720), .B(n_797), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_720), .B(n_754), .Y(n_911) );
INVx3_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
CKINVDCx6p67_ASAP7_75t_R g761 ( .A(n_722), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_722), .B(n_772), .Y(n_771) );
AND2x2_ASAP7_75t_L g805 ( .A(n_722), .B(n_778), .Y(n_805) );
AND2x2_ASAP7_75t_L g815 ( .A(n_722), .B(n_760), .Y(n_815) );
NOR2xp33_ASAP7_75t_L g843 ( .A(n_722), .B(n_760), .Y(n_843) );
AND2x2_ASAP7_75t_L g862 ( .A(n_722), .B(n_828), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_722), .B(n_757), .Y(n_898) );
OR2x6_ASAP7_75t_SL g722 ( .A(n_723), .B(n_729), .Y(n_722) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_731), .B1(n_733), .B2(n_734), .Y(n_729) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g817 ( .A(n_736), .Y(n_817) );
NOR2xp33_ASAP7_75t_L g877 ( .A(n_736), .B(n_754), .Y(n_877) );
AND2x2_ASAP7_75t_L g736 ( .A(n_737), .B(n_741), .Y(n_736) );
CKINVDCx6p67_ASAP7_75t_R g757 ( .A(n_737), .Y(n_757) );
INVx1_ASAP7_75t_L g788 ( .A(n_737), .Y(n_788) );
OR2x2_ASAP7_75t_L g792 ( .A(n_737), .B(n_742), .Y(n_792) );
OAI32xp33_ASAP7_75t_L g808 ( .A1(n_737), .A2(n_792), .A3(n_809), .B1(n_810), .B2(n_811), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_737), .B(n_742), .Y(n_826) );
AND2x2_ASAP7_75t_L g828 ( .A(n_737), .B(n_755), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g892 ( .A(n_737), .B(n_756), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_737), .B(n_778), .Y(n_906) );
AND2x2_ASAP7_75t_L g737 ( .A(n_738), .B(n_740), .Y(n_737) );
INVx2_ASAP7_75t_SL g801 ( .A(n_739), .Y(n_801) );
OR2x2_ASAP7_75t_L g809 ( .A(n_741), .B(n_755), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_741), .B(n_815), .Y(n_814) );
AND2x2_ASAP7_75t_L g859 ( .A(n_741), .B(n_757), .Y(n_859) );
INVx1_ASAP7_75t_L g897 ( .A(n_741), .Y(n_897) );
AND2x2_ASAP7_75t_L g741 ( .A(n_742), .B(n_745), .Y(n_741) );
CKINVDCx5p33_ASAP7_75t_R g756 ( .A(n_742), .Y(n_756) );
AND2x2_ASAP7_75t_L g848 ( .A(n_742), .B(n_746), .Y(n_848) );
AND2x4_ASAP7_75t_SL g742 ( .A(n_743), .B(n_744), .Y(n_742) );
INVx1_ASAP7_75t_L g763 ( .A(n_745), .Y(n_763) );
AND2x2_ASAP7_75t_L g772 ( .A(n_745), .B(n_757), .Y(n_772) );
AND2x2_ASAP7_75t_L g778 ( .A(n_745), .B(n_756), .Y(n_778) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
AND2x2_ASAP7_75t_L g755 ( .A(n_746), .B(n_756), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_750), .Y(n_746) );
OAI211xp5_ASAP7_75t_SL g860 ( .A1(n_753), .A2(n_811), .B(n_861), .C(n_863), .Y(n_860) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_SL g754 ( .A(n_755), .B(n_757), .Y(n_754) );
AND2x2_ASAP7_75t_L g820 ( .A(n_755), .B(n_821), .Y(n_820) );
OAI21xp33_ASAP7_75t_L g850 ( .A1(n_755), .A2(n_759), .B(n_772), .Y(n_850) );
AND2x2_ASAP7_75t_L g889 ( .A(n_755), .B(n_865), .Y(n_889) );
OAI222xp33_ASAP7_75t_L g765 ( .A1(n_756), .A2(n_766), .B1(n_771), .B2(n_773), .C1(n_775), .C2(n_777), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_756), .B(n_787), .Y(n_786) );
AOI22xp33_ASAP7_75t_SL g836 ( .A1(n_756), .A2(n_824), .B1(n_837), .B2(n_838), .Y(n_836) );
AND2x2_ASAP7_75t_L g821 ( .A(n_757), .B(n_761), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_757), .B(n_778), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_757), .B(n_848), .Y(n_847) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_757), .B(n_869), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_757), .B(n_805), .Y(n_884) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_759), .B(n_794), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
AND2x2_ASAP7_75t_L g767 ( .A(n_760), .B(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g790 ( .A(n_760), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g845 ( .A(n_760), .B(n_816), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_760), .B(n_864), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_760), .B(n_889), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_761), .B(n_767), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g785 ( .A(n_761), .B(n_786), .Y(n_785) );
NOR2x1p5_ASAP7_75t_L g791 ( .A(n_761), .B(n_792), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_761), .B(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g840 ( .A(n_761), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_761), .B(n_859), .Y(n_858) );
AND2x2_ASAP7_75t_L g865 ( .A(n_761), .B(n_787), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_761), .B(n_776), .Y(n_875) );
NOR2xp33_ASAP7_75t_L g881 ( .A(n_761), .B(n_810), .Y(n_881) );
INVx1_ASAP7_75t_L g842 ( .A(n_762), .Y(n_842) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVxp67_ASAP7_75t_L g903 ( .A(n_766), .Y(n_903) );
INVx1_ASAP7_75t_L g849 ( .A(n_767), .Y(n_849) );
INVx2_ASAP7_75t_L g774 ( .A(n_768), .Y(n_774) );
AND2x2_ASAP7_75t_L g887 ( .A(n_768), .B(n_797), .Y(n_887) );
AND2x2_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
AOI221xp5_ASAP7_75t_L g827 ( .A1(n_772), .A2(n_828), .B1(n_829), .B2(n_831), .C(n_832), .Y(n_827) );
AOI211xp5_ASAP7_75t_L g844 ( .A1(n_772), .A2(n_845), .B(n_846), .C(n_853), .Y(n_844) );
OAI211xp5_ASAP7_75t_SL g802 ( .A1(n_773), .A2(n_803), .B(n_806), .C(n_827), .Y(n_802) );
INVx3_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
OR2x2_ASAP7_75t_L g816 ( .A(n_774), .B(n_797), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_774), .B(n_796), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_774), .B(n_797), .Y(n_909) );
OAI221xp5_ASAP7_75t_L g890 ( .A1(n_775), .A2(n_891), .B1(n_893), .B2(n_895), .C(n_899), .Y(n_890) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
BUFx3_ASAP7_75t_L g855 ( .A(n_780), .Y(n_855) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
AND2x2_ASAP7_75t_L g804 ( .A(n_787), .B(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
INVx3_ASAP7_75t_L g807 ( .A(n_793), .Y(n_807) );
OAI311xp33_ASAP7_75t_L g846 ( .A1(n_793), .A2(n_847), .A3(n_849), .B1(n_850), .C1(n_851), .Y(n_846) );
INVx3_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx3_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_795), .B(n_854), .Y(n_853) );
INVx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_796), .B(n_820), .Y(n_819) );
INVx3_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g830 ( .A(n_797), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_797), .B(n_824), .Y(n_834) );
AND2x2_ASAP7_75t_L g871 ( .A(n_797), .B(n_872), .Y(n_871) );
AND2x4_ASAP7_75t_L g797 ( .A(n_798), .B(n_799), .Y(n_797) );
INVx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
AOI211xp5_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_808), .B(n_813), .C(n_822), .Y(n_806) );
INVx1_ASAP7_75t_L g872 ( .A(n_810), .Y(n_872) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
OAI221xp5_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_816), .B1(n_817), .B2(n_818), .C(n_819), .Y(n_813) );
INVx1_ASAP7_75t_L g838 ( .A(n_816), .Y(n_838) );
OAI221xp5_ASAP7_75t_SL g835 ( .A1(n_818), .A2(n_836), .B1(n_839), .B2(n_841), .C(n_844), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_821), .B(n_848), .Y(n_901) );
AOI21xp33_ASAP7_75t_SL g822 ( .A1(n_823), .A2(n_825), .B(n_826), .Y(n_822) );
AOI211xp5_ASAP7_75t_SL g882 ( .A1(n_824), .A2(n_883), .B(n_885), .C(n_890), .Y(n_882) );
NOR2xp33_ASAP7_75t_L g879 ( .A(n_826), .B(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g904 ( .A(n_826), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_828), .B(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g854 ( .A(n_828), .Y(n_854) );
NOR2xp33_ASAP7_75t_L g891 ( .A(n_828), .B(n_892), .Y(n_891) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_833), .B(n_834), .Y(n_832) );
INVx1_ASAP7_75t_L g837 ( .A(n_833), .Y(n_837) );
AOI221xp5_ASAP7_75t_L g856 ( .A1(n_838), .A2(n_845), .B1(n_857), .B2(n_860), .C(n_866), .Y(n_856) );
CKINVDCx14_ASAP7_75t_R g839 ( .A(n_840), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_842), .B(n_843), .Y(n_841) );
AND2x2_ASAP7_75t_L g864 ( .A(n_848), .B(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g869 ( .A(n_848), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_852), .B(n_862), .Y(n_861) );
AOI322xp5_ASAP7_75t_L g902 ( .A1(n_855), .A2(n_887), .A3(n_903), .B1(n_904), .B2(n_905), .C1(n_907), .C2(n_910), .Y(n_902) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
NOR2xp33_ASAP7_75t_L g866 ( .A(n_867), .B(n_870), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_872), .B(n_894), .Y(n_893) );
OAI21xp33_ASAP7_75t_L g899 ( .A1(n_872), .A2(n_887), .B(n_900), .Y(n_899) );
AOI211xp5_ASAP7_75t_L g873 ( .A1(n_874), .A2(n_876), .B(n_878), .C(n_879), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
INVxp67_ASAP7_75t_SL g876 ( .A(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
NOR2xp33_ASAP7_75t_L g885 ( .A(n_886), .B(n_888), .Y(n_885) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVx1_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
NOR2xp33_ASAP7_75t_L g896 ( .A(n_897), .B(n_898), .Y(n_896) );
INVx1_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
INVx1_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
CKINVDCx5p33_ASAP7_75t_R g912 ( .A(n_913), .Y(n_912) );
HB1xp67_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
NOR2x1_ASAP7_75t_SL g916 ( .A(n_917), .B(n_927), .Y(n_916) );
NAND3xp33_ASAP7_75t_L g917 ( .A(n_918), .B(n_920), .C(n_922), .Y(n_917) );
NAND4xp25_ASAP7_75t_SL g927 ( .A(n_928), .B(n_929), .C(n_930), .D(n_931), .Y(n_927) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
BUFx2_ASAP7_75t_SL g937 ( .A(n_938), .Y(n_937) );
INVxp67_ASAP7_75t_SL g941 ( .A(n_942), .Y(n_941) );
AND2x2_ASAP7_75t_L g942 ( .A(n_943), .B(n_948), .Y(n_942) );
AND4x1_ASAP7_75t_L g943 ( .A(n_944), .B(n_945), .C(n_946), .D(n_947), .Y(n_943) );
NOR3xp33_ASAP7_75t_L g948 ( .A(n_949), .B(n_954), .C(n_958), .Y(n_948) );
INVx2_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
BUFx3_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
CKINVDCx5p33_ASAP7_75t_R g965 ( .A(n_966), .Y(n_965) );
endmodule