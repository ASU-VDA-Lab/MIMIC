module fake_jpeg_29888_n_230 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_230);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_22),
.B(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_12),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_22),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_30),
.Y(n_61)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_20),
.B1(n_16),
.B2(n_29),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_47),
.A2(n_49),
.B1(n_16),
.B2(n_21),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_31),
.B1(n_29),
.B2(n_20),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_50),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_23),
.B(n_25),
.C(n_34),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_25),
.B(n_23),
.C(n_32),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_24),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_60),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_57),
.B(n_14),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_61),
.B(n_30),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_68),
.Y(n_91)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_21),
.B1(n_44),
.B2(n_39),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_72),
.A2(n_75),
.B1(n_77),
.B2(n_98),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_35),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_31),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_21),
.B1(n_29),
.B2(n_20),
.Y(n_75)
);

NAND2x1_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_45),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_21),
.B1(n_16),
.B2(n_27),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_86),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_79),
.B(n_85),
.Y(n_124)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_52),
.B(n_26),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_88),
.B(n_100),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_89),
.A2(n_64),
.B1(n_54),
.B2(n_31),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_32),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_69),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_R g93 ( 
.A(n_64),
.B(n_24),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_33),
.B(n_2),
.C(n_3),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_26),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_47),
.B(n_43),
.C(n_27),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_28),
.Y(n_118)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_62),
.A2(n_45),
.B(n_24),
.C(n_18),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_97),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_58),
.A2(n_27),
.B1(n_28),
.B2(n_45),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_58),
.A2(n_28),
.B1(n_45),
.B2(n_31),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_99),
.A2(n_59),
.B1(n_54),
.B2(n_67),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_62),
.B(n_24),
.Y(n_100)
);

OA21x2_ASAP7_75t_L g101 ( 
.A1(n_59),
.A2(n_24),
.B(n_28),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_101),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_103),
.B(n_108),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_104),
.A2(n_107),
.B1(n_112),
.B2(n_84),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_66),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_66),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_109),
.B(n_123),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_89),
.A2(n_28),
.B1(n_33),
.B2(n_3),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_114),
.Y(n_136)
);

BUFx4f_ASAP7_75t_SL g115 ( 
.A(n_70),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_73),
.Y(n_149)
);

AOI32xp33_ASAP7_75t_L g119 ( 
.A1(n_93),
.A2(n_71),
.A3(n_79),
.B1(n_95),
.B2(n_76),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_SL g153 ( 
.A(n_119),
.B(n_120),
.C(n_115),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_33),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_100),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_129),
.Y(n_143)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_128),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_80),
.B(n_33),
.Y(n_129)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_82),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_80),
.C(n_81),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_131),
.B(n_132),
.C(n_148),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_81),
.C(n_76),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_109),
.B(n_101),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_149),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_113),
.B(n_124),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_135),
.A2(n_105),
.B(n_128),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_125),
.A2(n_122),
.B1(n_119),
.B2(n_103),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_101),
.B1(n_91),
.B2(n_97),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_126),
.A2(n_91),
.B1(n_96),
.B2(n_83),
.Y(n_140)
);

AND2x6_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_70),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_146),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_112),
.A2(n_86),
.B1(n_78),
.B2(n_84),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_130),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_33),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_73),
.C(n_13),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_120),
.B(n_1),
.Y(n_152)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_153),
.B(n_138),
.Y(n_158)
);

A2O1A1Ixp33_ASAP7_75t_SL g155 ( 
.A1(n_153),
.A2(n_104),
.B(n_107),
.C(n_105),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_155),
.A2(n_134),
.B(n_147),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_110),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_156),
.B(n_157),
.Y(n_177)
);

NAND3xp33_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_165),
.C(n_167),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_115),
.Y(n_159)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_160),
.Y(n_185)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_161),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_162),
.A2(n_171),
.B1(n_147),
.B2(n_4),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_114),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_166),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_127),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_136),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_116),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_169),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_116),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_106),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_149),
.C(n_132),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_173),
.B(n_176),
.Y(n_191)
);

AO32x1_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_142),
.A3(n_131),
.B1(n_150),
.B2(n_141),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_178),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_179),
.A2(n_160),
.B(n_170),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_106),
.C(n_147),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_180),
.B(n_181),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_147),
.C(n_4),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_187),
.Y(n_196)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_168),
.A2(n_2),
.B(n_5),
.C(n_6),
.Y(n_187)
);

NOR3xp33_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_2),
.C(n_5),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_188),
.B(n_6),
.Y(n_190)
);

BUFx12_ASAP7_75t_L g189 ( 
.A(n_176),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_189),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_190),
.B(n_6),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_193),
.A2(n_195),
.B1(n_174),
.B2(n_186),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_172),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_175),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_184),
.A2(n_170),
.B1(n_155),
.B2(n_157),
.Y(n_195)
);

AO221x1_ASAP7_75t_L g197 ( 
.A1(n_183),
.A2(n_166),
.B1(n_155),
.B2(n_9),
.C(n_10),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_197),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_162),
.Y(n_198)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_198),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_185),
.A2(n_155),
.B1(n_172),
.B2(n_9),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_179),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_180),
.C(n_177),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_201),
.B(n_202),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_199),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_181),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_206),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_174),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_205),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_210),
.B(n_191),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_212),
.Y(n_219)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_213),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_192),
.C(n_189),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_216),
.A2(n_217),
.B(n_214),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_204),
.A2(n_202),
.B(n_210),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_220),
.B(n_221),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_215),
.A2(n_193),
.B(n_196),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_211),
.C(n_203),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_224),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_200),
.Y(n_224)
);

AO21x1_ASAP7_75t_L g226 ( 
.A1(n_222),
.A2(n_208),
.B(n_196),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_195),
.B(n_207),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_228),
.Y(n_229)
);

AOI322xp5_ASAP7_75t_L g228 ( 
.A1(n_225),
.A2(n_7),
.A3(n_9),
.B1(n_187),
.B2(n_200),
.C1(n_209),
.C2(n_222),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_7),
.Y(n_230)
);


endmodule