module real_jpeg_5650_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_2),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_2),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_2),
.B(n_80),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_3),
.B(n_102),
.Y(n_101)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_4),
.Y(n_77)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_5),
.Y(n_105)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_6),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_7),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_7),
.B(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_8),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_8),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_8),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_8),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_18),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_9),
.B(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_9),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_9),
.B(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_10),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_21),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_11),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_11),
.B(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_11),
.B(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_85),
.Y(n_12)
);

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_56),
.B(n_84),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_43),
.B(n_55),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_23),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_16),
.B(n_23),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_20),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_17),
.B(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_19),
.Y(n_99)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_36),
.B2(n_37),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_26),
.B(n_30),
.C(n_36),
.Y(n_83)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_34),
.Y(n_117)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_41),
.Y(n_66)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_50),
.B(n_54),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_46),
.Y(n_54)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_83),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_83),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_67),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_66),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_66),
.C(n_89),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_60),
.B(n_63),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_72),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_68),
.B(n_78),
.C(n_82),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_78),
.B1(n_79),
.B2(n_82),
.Y(n_72)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_129),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_90),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_90),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_107),
.B2(n_108),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_100),
.B1(n_101),
.B2(n_106),
.Y(n_96)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_118),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_124),
.B2(n_128),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_124),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);


endmodule