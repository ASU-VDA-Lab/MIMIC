module fake_netlist_1_12596_n_651 (n_117, n_44, n_133, n_149, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_125, n_9, n_161, n_10, n_130, n_103, n_19, n_87, n_137, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_165, n_146, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_169, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_46, n_31, n_58, n_122, n_138, n_126, n_118, n_32, n_0, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_166, n_162, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_68, n_144, n_27, n_53, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_15, n_173, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_651);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_125;
input n_9;
input n_161;
input n_10;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_165;
input n_146;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_169;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_46;
input n_31;
input n_58;
input n_122;
input n_138;
input n_126;
input n_118;
input n_32;
input n_0;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_166;
input n_162;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_68;
input n_144;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_15;
input n_173;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_651;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_431;
wire n_484;
wire n_496;
wire n_177;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_612;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_202;
wire n_386;
wire n_432;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_205;
wire n_330;
wire n_587;
wire n_387;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_178;
wire n_616;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_295;
wire n_263;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_553;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_524;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_602;
wire n_198;
wire n_424;
wire n_629;
wire n_569;
wire n_297;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_187;
wire n_375;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_421;
wire n_175;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g175 ( .A(n_120), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_154), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_63), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_107), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_147), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_8), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_128), .Y(n_181) );
CKINVDCx5p33_ASAP7_75t_R g182 ( .A(n_43), .Y(n_182) );
INVxp67_ASAP7_75t_L g183 ( .A(n_161), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_40), .Y(n_184) );
INVx1_ASAP7_75t_SL g185 ( .A(n_56), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_72), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_36), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_38), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_114), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_167), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_9), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_135), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_143), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_39), .Y(n_194) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_30), .Y(n_195) );
INVx1_ASAP7_75t_SL g196 ( .A(n_78), .Y(n_196) );
INVx1_ASAP7_75t_SL g197 ( .A(n_47), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_41), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_125), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_156), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_174), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_109), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_20), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_4), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_69), .Y(n_205) );
CKINVDCx16_ASAP7_75t_R g206 ( .A(n_15), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_53), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_145), .Y(n_208) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_16), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_158), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_87), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_49), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_130), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_51), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_116), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_144), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_115), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_122), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_94), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_160), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_166), .Y(n_221) );
BUFx10_ASAP7_75t_L g222 ( .A(n_165), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_173), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_55), .Y(n_224) );
NOR2xp67_ASAP7_75t_L g225 ( .A(n_97), .B(n_3), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_113), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_28), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_71), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_151), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_1), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_17), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_164), .Y(n_232) );
INVx1_ASAP7_75t_SL g233 ( .A(n_0), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_91), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_33), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_44), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_162), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_60), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_11), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_153), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_24), .Y(n_241) );
CKINVDCx16_ASAP7_75t_R g242 ( .A(n_155), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_34), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_46), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_21), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_48), .Y(n_246) );
INVxp67_ASAP7_75t_SL g247 ( .A(n_64), .Y(n_247) );
INVxp67_ASAP7_75t_L g248 ( .A(n_75), .Y(n_248) );
BUFx3_ASAP7_75t_L g249 ( .A(n_157), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_170), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g251 ( .A(n_68), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g252 ( .A(n_22), .Y(n_252) );
INVxp67_ASAP7_75t_SL g253 ( .A(n_98), .Y(n_253) );
BUFx10_ASAP7_75t_L g254 ( .A(n_18), .Y(n_254) );
CKINVDCx20_ASAP7_75t_R g255 ( .A(n_142), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_52), .Y(n_256) );
BUFx10_ASAP7_75t_L g257 ( .A(n_50), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_138), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_106), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_77), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_104), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_159), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_150), .Y(n_263) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_4), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_152), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_54), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_148), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_85), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_149), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_126), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_171), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_58), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_139), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_141), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_163), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_168), .Y(n_276) );
CKINVDCx20_ASAP7_75t_R g277 ( .A(n_70), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_209), .B(n_0), .Y(n_278) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_204), .Y(n_279) );
OAI22x1_ASAP7_75t_L g280 ( .A1(n_230), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_280) );
AND2x4_ASAP7_75t_L g281 ( .A(n_214), .B(n_2), .Y(n_281) );
OA21x2_ASAP7_75t_L g282 ( .A1(n_175), .A2(n_101), .B(n_169), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_206), .B(n_5), .Y(n_283) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_242), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_284) );
BUFx12f_ASAP7_75t_L g285 ( .A(n_222), .Y(n_285) );
BUFx3_ASAP7_75t_L g286 ( .A(n_249), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_222), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_234), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_254), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_220), .Y(n_290) );
BUFx8_ASAP7_75t_SL g291 ( .A(n_235), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_223), .Y(n_292) );
BUFx3_ASAP7_75t_L g293 ( .A(n_273), .Y(n_293) );
AND2x4_ASAP7_75t_L g294 ( .A(n_238), .B(n_6), .Y(n_294) );
AOI22x1_ASAP7_75t_SL g295 ( .A1(n_251), .A2(n_7), .B1(n_10), .B2(n_12), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_245), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_254), .Y(n_297) );
AND2x4_ASAP7_75t_L g298 ( .A(n_176), .B(n_13), .Y(n_298) );
BUFx2_ASAP7_75t_L g299 ( .A(n_264), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_177), .B(n_14), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_264), .Y(n_301) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_287), .B(n_257), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_281), .Y(n_303) );
NAND2xp33_ASAP7_75t_R g304 ( .A(n_288), .B(n_178), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_286), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_281), .Y(n_306) );
AO21x2_ASAP7_75t_L g307 ( .A1(n_300), .A2(n_181), .B(n_179), .Y(n_307) );
OR2x6_ASAP7_75t_L g308 ( .A(n_285), .B(n_225), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_286), .Y(n_309) );
INVx3_ASAP7_75t_L g310 ( .A(n_294), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_293), .B(n_186), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_294), .Y(n_312) );
INVx3_ASAP7_75t_L g313 ( .A(n_298), .Y(n_313) );
OAI22xp33_ASAP7_75t_L g314 ( .A1(n_284), .A2(n_233), .B1(n_277), .B2(n_252), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_293), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_290), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_289), .B(n_183), .Y(n_317) );
NAND2xp5_ASAP7_75t_SL g318 ( .A(n_297), .B(n_257), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g319 ( .A(n_313), .B(n_298), .Y(n_319) );
INVx8_ASAP7_75t_L g320 ( .A(n_308), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_305), .Y(n_321) );
OR2x6_ASAP7_75t_L g322 ( .A(n_308), .B(n_280), .Y(n_322) );
NAND2xp33_ASAP7_75t_L g323 ( .A(n_313), .B(n_300), .Y(n_323) );
NAND2xp5_ASAP7_75t_SL g324 ( .A(n_303), .B(n_278), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_310), .B(n_279), .Y(n_325) );
BUFx3_ASAP7_75t_L g326 ( .A(n_309), .Y(n_326) );
NAND2xp33_ASAP7_75t_L g327 ( .A(n_306), .B(n_279), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_310), .B(n_283), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_315), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_316), .Y(n_330) );
NOR2xp67_ASAP7_75t_L g331 ( .A(n_317), .B(n_283), .Y(n_331) );
A2O1A1Ixp33_ASAP7_75t_L g332 ( .A1(n_312), .A2(n_292), .B(n_296), .C(n_262), .Y(n_332) );
NAND2xp5_ASAP7_75t_SL g333 ( .A(n_302), .B(n_180), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_328), .A2(n_288), .B1(n_255), .B2(n_311), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_326), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_331), .B(n_307), .Y(n_336) );
OA22x2_ASAP7_75t_L g337 ( .A1(n_322), .A2(n_291), .B1(n_308), .B2(n_314), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_325), .B(n_311), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_324), .B(n_307), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_327), .B(n_318), .Y(n_340) );
AOI22xp5_ASAP7_75t_L g341 ( .A1(n_323), .A2(n_304), .B1(n_319), .B2(n_322), .Y(n_341) );
NAND2x1p5_ASAP7_75t_L g342 ( .A(n_330), .B(n_299), .Y(n_342) );
AOI21xp5_ASAP7_75t_L g343 ( .A1(n_321), .A2(n_282), .B(n_253), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_332), .B(n_248), .Y(n_344) );
A2O1A1Ixp33_ASAP7_75t_L g345 ( .A1(n_329), .A2(n_256), .B(n_226), .C(n_187), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_333), .A2(n_282), .B(n_247), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_320), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_320), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_338), .B(n_295), .Y(n_349) );
O2A1O1Ixp5_ASAP7_75t_L g350 ( .A1(n_346), .A2(n_227), .B(n_190), .C(n_191), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_334), .B(n_291), .Y(n_351) );
AO31x2_ASAP7_75t_L g352 ( .A1(n_343), .A2(n_219), .A3(n_271), .B(n_268), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_341), .B(n_264), .Y(n_353) );
O2A1O1Ixp33_ASAP7_75t_L g354 ( .A1(n_345), .A2(n_208), .B(n_231), .C(n_192), .Y(n_354) );
NOR2x1_ASAP7_75t_L g355 ( .A(n_336), .B(n_193), .Y(n_355) );
A2O1A1Ixp33_ASAP7_75t_L g356 ( .A1(n_339), .A2(n_211), .B(n_232), .C(n_194), .Y(n_356) );
O2A1O1Ixp5_ASAP7_75t_L g357 ( .A1(n_344), .A2(n_229), .B(n_199), .C(n_200), .Y(n_357) );
OAI21x1_ASAP7_75t_SL g358 ( .A1(n_340), .A2(n_205), .B(n_202), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_342), .B(n_185), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_335), .Y(n_360) );
OAI22xp5_ASAP7_75t_L g361 ( .A1(n_335), .A2(n_196), .B1(n_197), .B2(n_275), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_347), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_348), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_337), .B(n_301), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g365 ( .A1(n_334), .A2(n_207), .B1(n_210), .B2(n_213), .Y(n_365) );
AND2x4_ASAP7_75t_SL g366 ( .A(n_347), .B(n_216), .Y(n_366) );
AOI21xp5_ASAP7_75t_L g367 ( .A1(n_336), .A2(n_217), .B(n_215), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_339), .Y(n_368) );
NAND2xp5_ASAP7_75t_SL g369 ( .A(n_338), .B(n_276), .Y(n_369) );
AOI21xp33_ASAP7_75t_L g370 ( .A1(n_334), .A2(n_184), .B(n_182), .Y(n_370) );
OAI21x1_ASAP7_75t_L g371 ( .A1(n_350), .A2(n_236), .B(n_221), .Y(n_371) );
OAI21x1_ASAP7_75t_L g372 ( .A1(n_358), .A2(n_244), .B(n_243), .Y(n_372) );
NAND2xp5_ASAP7_75t_SL g373 ( .A(n_359), .B(n_188), .Y(n_373) );
OR2x6_ASAP7_75t_L g374 ( .A(n_349), .B(n_246), .Y(n_374) );
BUFx2_ASAP7_75t_L g375 ( .A(n_355), .Y(n_375) );
OR2x6_ASAP7_75t_L g376 ( .A(n_351), .B(n_250), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_365), .B(n_266), .Y(n_377) );
INVx4_ASAP7_75t_L g378 ( .A(n_366), .Y(n_378) );
OR2x6_ASAP7_75t_L g379 ( .A(n_362), .B(n_363), .Y(n_379) );
OAI21x1_ASAP7_75t_L g380 ( .A1(n_368), .A2(n_267), .B(n_216), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_356), .B(n_274), .Y(n_381) );
OAI21x1_ASAP7_75t_L g382 ( .A1(n_355), .A2(n_216), .B(n_23), .Y(n_382) );
OAI21x1_ASAP7_75t_L g383 ( .A1(n_353), .A2(n_19), .B(n_25), .Y(n_383) );
AOI21x1_ASAP7_75t_L g384 ( .A1(n_367), .A2(n_272), .B(n_270), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_352), .Y(n_385) );
OAI21x1_ASAP7_75t_L g386 ( .A1(n_357), .A2(n_26), .B(n_27), .Y(n_386) );
AO31x2_ASAP7_75t_L g387 ( .A1(n_352), .A2(n_29), .A3(n_31), .B(n_32), .Y(n_387) );
AO21x2_ASAP7_75t_L g388 ( .A1(n_354), .A2(n_35), .B(n_37), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_370), .B(n_269), .Y(n_389) );
BUFx12f_ASAP7_75t_L g390 ( .A(n_364), .Y(n_390) );
AOI21xp5_ASAP7_75t_L g391 ( .A1(n_369), .A2(n_265), .B(n_263), .Y(n_391) );
NOR2xp67_ASAP7_75t_L g392 ( .A(n_361), .B(n_42), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_352), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_360), .Y(n_394) );
BUFx12f_ASAP7_75t_L g395 ( .A(n_364), .Y(n_395) );
OA21x2_ASAP7_75t_L g396 ( .A1(n_350), .A2(n_261), .B(n_260), .Y(n_396) );
NAND2x1p5_ASAP7_75t_L g397 ( .A(n_362), .B(n_45), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_362), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g399 ( .A1(n_350), .A2(n_259), .B(n_258), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_349), .B(n_189), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_362), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_368), .Y(n_402) );
OAI21x1_ASAP7_75t_L g403 ( .A1(n_350), .A2(n_57), .B(n_59), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_349), .B(n_241), .Y(n_404) );
OAI21x1_ASAP7_75t_L g405 ( .A1(n_350), .A2(n_61), .B(n_62), .Y(n_405) );
OR2x6_ASAP7_75t_L g406 ( .A(n_349), .B(n_65), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_349), .B(n_240), .Y(n_407) );
BUFx2_ASAP7_75t_L g408 ( .A(n_355), .Y(n_408) );
NAND3xp33_ASAP7_75t_L g409 ( .A(n_357), .B(n_239), .C(n_237), .Y(n_409) );
INVx3_ASAP7_75t_L g410 ( .A(n_366), .Y(n_410) );
BUFx2_ASAP7_75t_L g411 ( .A(n_378), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_385), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_398), .Y(n_413) );
AND2x4_ASAP7_75t_L g414 ( .A(n_402), .B(n_66), .Y(n_414) );
INVx3_ASAP7_75t_L g415 ( .A(n_379), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_379), .B(n_228), .Y(n_416) );
CKINVDCx11_ASAP7_75t_R g417 ( .A(n_390), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_401), .Y(n_418) );
INVx2_ASAP7_75t_SL g419 ( .A(n_410), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_374), .B(n_195), .Y(n_420) );
INVx3_ASAP7_75t_L g421 ( .A(n_406), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_394), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_406), .Y(n_423) );
AOI21xp33_ASAP7_75t_L g424 ( .A1(n_375), .A2(n_218), .B(n_212), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_393), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_397), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_374), .B(n_198), .Y(n_427) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_372), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_387), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_387), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_376), .B(n_201), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_376), .B(n_203), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_380), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_375), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_408), .Y(n_435) );
INVx3_ASAP7_75t_L g436 ( .A(n_408), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_373), .B(n_224), .Y(n_437) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_392), .Y(n_438) );
BUFx3_ASAP7_75t_L g439 ( .A(n_395), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_377), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_382), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_371), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_400), .B(n_67), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_384), .Y(n_444) );
AO21x2_ASAP7_75t_L g445 ( .A1(n_403), .A2(n_73), .B(n_74), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_386), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_409), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_389), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_381), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_404), .Y(n_450) );
INVx3_ASAP7_75t_L g451 ( .A(n_388), .Y(n_451) );
NAND2x1p5_ASAP7_75t_L g452 ( .A(n_396), .B(n_76), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_396), .B(n_79), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_407), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_391), .B(n_80), .Y(n_455) );
OAI21x1_ASAP7_75t_L g456 ( .A1(n_405), .A2(n_81), .B(n_82), .Y(n_456) );
NAND2x1_ASAP7_75t_L g457 ( .A(n_399), .B(n_83), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_383), .B(n_84), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_379), .B(n_86), .Y(n_459) );
BUFx3_ASAP7_75t_L g460 ( .A(n_410), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_402), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_402), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_398), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_374), .B(n_88), .Y(n_464) );
CKINVDCx5p33_ASAP7_75t_R g465 ( .A(n_390), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_398), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_398), .Y(n_467) );
INVx4_ASAP7_75t_L g468 ( .A(n_378), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_402), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_379), .B(n_89), .Y(n_470) );
BUFx3_ASAP7_75t_L g471 ( .A(n_411), .Y(n_471) );
AND2x4_ASAP7_75t_SL g472 ( .A(n_468), .B(n_90), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_440), .B(n_92), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_413), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_461), .B(n_93), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_462), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_418), .B(n_95), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_469), .B(n_96), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_448), .B(n_99), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_422), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_463), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_466), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_467), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_412), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_450), .B(n_100), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_412), .Y(n_486) );
INVxp67_ASAP7_75t_L g487 ( .A(n_438), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_454), .B(n_102), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_434), .B(n_103), .Y(n_489) );
BUFx3_ASAP7_75t_L g490 ( .A(n_468), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_435), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_415), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_421), .B(n_172), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_415), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_425), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_425), .Y(n_496) );
BUFx3_ASAP7_75t_L g497 ( .A(n_460), .Y(n_497) );
AO21x2_ASAP7_75t_L g498 ( .A1(n_446), .A2(n_105), .B(n_108), .Y(n_498) );
BUFx6f_ASAP7_75t_L g499 ( .A(n_460), .Y(n_499) );
AND2x4_ASAP7_75t_L g500 ( .A(n_436), .B(n_110), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_423), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_436), .B(n_111), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_421), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_459), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_438), .B(n_112), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_416), .B(n_117), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_470), .B(n_118), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_426), .Y(n_508) );
NOR2x1p5_ASAP7_75t_L g509 ( .A(n_439), .B(n_119), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_414), .Y(n_510) );
INVx1_ASAP7_75t_SL g511 ( .A(n_428), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_464), .B(n_121), .Y(n_512) );
AND2x4_ASAP7_75t_L g513 ( .A(n_428), .B(n_123), .Y(n_513) );
INVxp67_ASAP7_75t_SL g514 ( .A(n_428), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_464), .B(n_124), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_444), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_417), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_449), .B(n_127), .Y(n_518) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_447), .A2(n_129), .B(n_131), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_431), .B(n_132), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_420), .B(n_133), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_432), .B(n_134), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_419), .B(n_136), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_427), .B(n_137), .Y(n_524) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_442), .Y(n_525) );
INVxp67_ASAP7_75t_L g526 ( .A(n_441), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_452), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_490), .B(n_439), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_480), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_501), .B(n_429), .Y(n_530) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_486), .Y(n_531) );
INVxp67_ASAP7_75t_L g532 ( .A(n_471), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_476), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_481), .B(n_430), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_474), .Y(n_535) );
BUFx2_ASAP7_75t_L g536 ( .A(n_490), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_486), .B(n_451), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_504), .B(n_508), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_484), .B(n_465), .Y(n_539) );
NOR2x1_ASAP7_75t_L g540 ( .A(n_509), .B(n_453), .Y(n_540) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_495), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_482), .B(n_443), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_483), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_517), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_503), .B(n_451), .Y(n_545) );
NOR2xp33_ASAP7_75t_SL g546 ( .A(n_500), .B(n_452), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_491), .B(n_458), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_516), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_492), .B(n_455), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_496), .B(n_433), .Y(n_550) );
AND2x4_ASAP7_75t_SL g551 ( .A(n_499), .B(n_417), .Y(n_551) );
INVx1_ASAP7_75t_SL g552 ( .A(n_497), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_487), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_494), .B(n_465), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_497), .B(n_424), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_487), .B(n_424), .Y(n_556) );
AND2x4_ASAP7_75t_L g557 ( .A(n_510), .B(n_445), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_525), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_525), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_499), .B(n_437), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_493), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_506), .B(n_456), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_526), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_526), .B(n_457), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_477), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_505), .B(n_140), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_505), .B(n_146), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_541), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_548), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_536), .B(n_511), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_529), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_552), .B(n_511), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_552), .B(n_514), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_533), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_531), .B(n_514), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_538), .B(n_527), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_535), .B(n_500), .Y(n_577) );
NOR2x1_ASAP7_75t_L g578 ( .A(n_528), .B(n_502), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_543), .B(n_524), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_553), .B(n_522), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_547), .B(n_521), .Y(n_581) );
INVx3_ASAP7_75t_L g582 ( .A(n_563), .Y(n_582) );
AND2x4_ASAP7_75t_L g583 ( .A(n_558), .B(n_472), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_559), .Y(n_584) );
AND2x4_ASAP7_75t_L g585 ( .A(n_545), .B(n_513), .Y(n_585) );
AND2x4_ASAP7_75t_SL g586 ( .A(n_544), .B(n_520), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_532), .B(n_507), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_555), .B(n_479), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_550), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_556), .B(n_489), .Y(n_590) );
NAND2x1_ASAP7_75t_L g591 ( .A(n_540), .B(n_513), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_565), .B(n_489), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_539), .B(n_485), .Y(n_593) );
AND2x4_ASAP7_75t_L g594 ( .A(n_530), .B(n_498), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_568), .B(n_561), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_589), .B(n_537), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_590), .B(n_542), .Y(n_597) );
OR2x6_ASAP7_75t_L g598 ( .A(n_583), .B(n_560), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_576), .B(n_554), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_569), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_570), .B(n_534), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_569), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_588), .B(n_557), .Y(n_603) );
INVx1_ASAP7_75t_SL g604 ( .A(n_586), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_584), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_571), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_583), .B(n_551), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_571), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_572), .B(n_557), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_589), .B(n_549), .Y(n_610) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_582), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_611), .Y(n_612) );
AOI21xp5_ASAP7_75t_L g613 ( .A1(n_604), .A2(n_578), .B(n_591), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_600), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_601), .B(n_573), .Y(n_615) );
NAND3xp33_ASAP7_75t_SL g616 ( .A(n_607), .B(n_546), .C(n_517), .Y(n_616) );
INVx1_ASAP7_75t_SL g617 ( .A(n_598), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_598), .A2(n_580), .B1(n_577), .B2(n_579), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_600), .Y(n_619) );
INVx2_ASAP7_75t_SL g620 ( .A(n_599), .Y(n_620) );
AOI21xp33_ASAP7_75t_L g621 ( .A1(n_595), .A2(n_592), .B(n_575), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_596), .B(n_582), .Y(n_622) );
AOI221x1_ASAP7_75t_SL g623 ( .A1(n_621), .A2(n_597), .B1(n_610), .B2(n_605), .C(n_602), .Y(n_623) );
NAND3xp33_ASAP7_75t_SL g624 ( .A(n_613), .B(n_546), .C(n_587), .Y(n_624) );
AOI211xp5_ASAP7_75t_L g625 ( .A1(n_616), .A2(n_617), .B(n_618), .C(n_612), .Y(n_625) );
AND2x4_ASAP7_75t_L g626 ( .A(n_620), .B(n_603), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_614), .Y(n_627) );
NOR2xp67_ASAP7_75t_L g628 ( .A(n_618), .B(n_609), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_619), .Y(n_629) );
NAND3xp33_ASAP7_75t_L g630 ( .A(n_625), .B(n_608), .C(n_606), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_627), .Y(n_631) );
OAI211xp5_ASAP7_75t_L g632 ( .A1(n_624), .A2(n_628), .B(n_623), .C(n_622), .Y(n_632) );
INVx2_ASAP7_75t_SL g633 ( .A(n_626), .Y(n_633) );
NOR3xp33_ASAP7_75t_L g634 ( .A(n_632), .B(n_567), .C(n_566), .Y(n_634) );
NAND3xp33_ASAP7_75t_L g635 ( .A(n_630), .B(n_629), .C(n_519), .Y(n_635) );
NAND4xp25_ASAP7_75t_L g636 ( .A(n_631), .B(n_515), .C(n_512), .D(n_523), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_635), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_634), .B(n_633), .Y(n_638) );
NOR3xp33_ASAP7_75t_L g639 ( .A(n_637), .B(n_636), .C(n_519), .Y(n_639) );
NAND3xp33_ASAP7_75t_SL g640 ( .A(n_638), .B(n_566), .C(n_567), .Y(n_640) );
XNOR2x1_ASAP7_75t_L g641 ( .A(n_640), .B(n_488), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_639), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_642), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_641), .A2(n_615), .B1(n_581), .B2(n_593), .Y(n_644) );
AOI21xp33_ASAP7_75t_L g645 ( .A1(n_643), .A2(n_473), .B(n_477), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_644), .A2(n_518), .B1(n_562), .B2(n_594), .Y(n_646) );
AOI22x1_ASAP7_75t_L g647 ( .A1(n_645), .A2(n_478), .B1(n_475), .B2(n_594), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_647), .A2(n_646), .B(n_473), .Y(n_648) );
OAI21x1_ASAP7_75t_L g649 ( .A1(n_648), .A2(n_564), .B(n_537), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_649), .B(n_498), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_650), .A2(n_585), .B1(n_574), .B2(n_564), .Y(n_651) );
endmodule