module fake_jpeg_6846_n_258 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_258);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_258;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_5),
.B(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_37),
.Y(n_44)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_17),
.B1(n_18),
.B2(n_22),
.Y(n_52)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_39),
.B(n_20),
.Y(n_51)
);

CKINVDCx6p67_ASAP7_75t_R g40 ( 
.A(n_26),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_24),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_27),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_52),
.Y(n_64)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_53),
.Y(n_66)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_55),
.Y(n_67)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_56),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_78)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_36),
.A2(n_22),
.B1(n_17),
.B2(n_31),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_31),
.B1(n_22),
.B2(n_24),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_65),
.A2(n_83),
.B1(n_19),
.B2(n_26),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_25),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_72),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_27),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_79),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_25),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_42),
.B(n_20),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_73),
.B(n_75),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_25),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_81),
.Y(n_105)
);

OR2x2_ASAP7_75t_SL g76 ( 
.A(n_63),
.B(n_14),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_76),
.A2(n_77),
.B(n_26),
.C(n_21),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_18),
.B1(n_23),
.B2(n_15),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_27),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_43),
.B(n_25),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_54),
.A2(n_23),
.B1(n_28),
.B2(n_30),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_25),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_85),
.B(n_45),
.Y(n_108)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_89),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_63),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_72),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_94),
.Y(n_125)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_93),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_67),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_64),
.A2(n_56),
.B1(n_53),
.B2(n_62),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_95),
.A2(n_99),
.B1(n_103),
.B2(n_65),
.Y(n_126)
);

AOI21xp33_ASAP7_75t_L g97 ( 
.A1(n_75),
.A2(n_19),
.B(n_45),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_97),
.A2(n_73),
.B(n_79),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_75),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_100),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_64),
.A2(n_58),
.B1(n_57),
.B2(n_18),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_101),
.B(n_102),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_57),
.B1(n_15),
.B2(n_30),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_84),
.A2(n_50),
.B1(n_16),
.B2(n_21),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_79),
.Y(n_131)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_74),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_114),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_94),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_113),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_81),
.C(n_67),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_93),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_126),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_100),
.A2(n_78),
.B1(n_77),
.B2(n_80),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_127),
.A2(n_134),
.B1(n_95),
.B2(n_99),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_128),
.B(n_88),
.Y(n_140)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_133),
.Y(n_148)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_92),
.B(n_90),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_88),
.Y(n_146)
);

OA21x2_ASAP7_75t_L g133 ( 
.A1(n_89),
.A2(n_49),
.B(n_80),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_107),
.A2(n_86),
.B1(n_70),
.B2(n_49),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_139),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_117),
.A2(n_88),
.B1(n_87),
.B2(n_101),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_137),
.A2(n_149),
.B1(n_119),
.B2(n_131),
.Y(n_158)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_141),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_116),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_146),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_123),
.A2(n_111),
.B(n_96),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_128),
.Y(n_159)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_106),
.B1(n_98),
.B2(n_109),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_93),
.Y(n_150)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

INVxp33_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_129),
.A2(n_86),
.B1(n_104),
.B2(n_91),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_152),
.A2(n_153),
.B1(n_122),
.B2(n_118),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_70),
.B1(n_66),
.B2(n_33),
.Y(n_153)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_154),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_114),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g163 ( 
.A1(n_155),
.A2(n_146),
.B(n_137),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_110),
.Y(n_156)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_159),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_133),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_160),
.A2(n_143),
.B(n_133),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_154),
.Y(n_162)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_169),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_145),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_168),
.B(n_173),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_112),
.Y(n_169)
);

OAI22x1_ASAP7_75t_L g170 ( 
.A1(n_135),
.A2(n_133),
.B1(n_127),
.B2(n_134),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_170),
.A2(n_175),
.B1(n_176),
.B2(n_149),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_144),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_172),
.B(n_174),
.Y(n_179)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_152),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_153),
.A2(n_155),
.B1(n_136),
.B2(n_140),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_130),
.Y(n_178)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_164),
.A2(n_142),
.B(n_147),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_181),
.A2(n_187),
.B(n_188),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_160),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_SL g196 ( 
.A(n_182),
.B(n_189),
.C(n_177),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_183),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_170),
.B1(n_175),
.B2(n_176),
.Y(n_186)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_166),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_158),
.A2(n_155),
.B1(n_136),
.B2(n_118),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_190),
.A2(n_194),
.B1(n_195),
.B2(n_115),
.Y(n_205)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_167),
.Y(n_192)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_192),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_161),
.B(n_122),
.Y(n_193)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_177),
.A2(n_115),
.B1(n_139),
.B2(n_141),
.Y(n_194)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_169),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_203),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_202),
.A2(n_208),
.B(n_210),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_138),
.Y(n_203)
);

FAx1_ASAP7_75t_SL g213 ( 
.A(n_205),
.B(n_206),
.CI(n_187),
.CON(n_213),
.SN(n_213)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_190),
.A2(n_163),
.B1(n_159),
.B2(n_171),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_120),
.C(n_33),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_178),
.B(n_76),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_209),
.B(n_26),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_195),
.B(n_181),
.C(n_194),
.Y(n_212)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_219),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_201),
.A2(n_198),
.B1(n_202),
.B2(n_197),
.Y(n_215)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_192),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_217),
.C(n_220),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_188),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_207),
.B(n_180),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_218),
.B(n_0),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_209),
.A2(n_180),
.B1(n_110),
.B2(n_16),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_34),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_214),
.C(n_211),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_204),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_223),
.A2(n_225),
.B(n_227),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_1),
.Y(n_240)
);

AOI221xp5_ASAP7_75t_L g225 ( 
.A1(n_212),
.A2(n_66),
.B1(n_1),
.B2(n_2),
.C(n_3),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_222),
.B(n_0),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_228),
.A2(n_231),
.B(n_211),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_216),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_238),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_229),
.Y(n_234)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_234),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_232),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_236),
.B(n_240),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_239),
.C(n_2),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_220),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_230),
.B(n_231),
.Y(n_239)
);

AOI322xp5_ASAP7_75t_L g242 ( 
.A1(n_236),
.A2(n_213),
.A3(n_66),
.B1(n_16),
.B2(n_21),
.C1(n_32),
.C2(n_34),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_243),
.C(n_245),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_2),
.C(n_3),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_26),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_247),
.A2(n_248),
.B(n_249),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_244),
.A2(n_21),
.B(n_4),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_241),
.A2(n_3),
.B(n_6),
.Y(n_249)
);

OAI321xp33_ASAP7_75t_L g251 ( 
.A1(n_250),
.A2(n_242),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C(n_6),
.Y(n_251)
);

OAI21xp33_ASAP7_75t_L g255 ( 
.A1(n_251),
.A2(n_253),
.B(n_13),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_13),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_252),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_254),
.B(n_255),
.Y(n_256)
);

AOI321xp33_ASAP7_75t_L g257 ( 
.A1(n_256),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C(n_237),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_11),
.Y(n_258)
);


endmodule