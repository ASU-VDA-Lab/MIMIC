module real_jpeg_23051_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_1),
.A2(n_38),
.B1(n_56),
.B2(n_58),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_1),
.A2(n_25),
.B1(n_30),
.B2(n_38),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_3),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_3),
.B(n_55),
.Y(n_190)
);

O2A1O1Ixp33_ASAP7_75t_L g231 ( 
.A1(n_3),
.A2(n_58),
.B(n_69),
.C(n_232),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_3),
.A2(n_56),
.B1(n_58),
.B2(n_172),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_3),
.B(n_25),
.C(n_28),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_172),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_3),
.A2(n_102),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_3),
.B(n_72),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_5),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_5),
.A2(n_45),
.B1(n_56),
.B2(n_58),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_45),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_5),
.A2(n_25),
.B1(n_30),
.B2(n_45),
.Y(n_192)
);

INVx8_ASAP7_75t_SL g52 ( 
.A(n_6),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_7),
.A2(n_44),
.B1(n_49),
.B2(n_145),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_7),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_7),
.A2(n_56),
.B1(n_58),
.B2(n_145),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_145),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_7),
.A2(n_25),
.B1(n_30),
.B2(n_145),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_10),
.A2(n_44),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_10),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_10),
.A2(n_56),
.B1(n_58),
.B2(n_61),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_61),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_10),
.A2(n_25),
.B1(n_30),
.B2(n_61),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_11),
.A2(n_56),
.B1(n_58),
.B2(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_75),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_11),
.A2(n_25),
.B1(n_30),
.B2(n_75),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_12),
.A2(n_49),
.B1(n_53),
.B2(n_118),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_12),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_118),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_12),
.A2(n_56),
.B1(n_58),
.B2(n_118),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_12),
.A2(n_25),
.B1(n_30),
.B2(n_118),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_13),
.A2(n_56),
.B1(n_58),
.B2(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_13),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_13),
.A2(n_43),
.B1(n_44),
.B2(n_162),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_13),
.A2(n_33),
.B1(n_34),
.B2(n_162),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_13),
.A2(n_25),
.B1(n_30),
.B2(n_162),
.Y(n_259)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_15),
.A2(n_56),
.B1(n_58),
.B2(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_15),
.A2(n_49),
.B1(n_50),
.B2(n_65),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_15),
.A2(n_33),
.B1(n_34),
.B2(n_65),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_15),
.A2(n_25),
.B1(n_30),
.B2(n_65),
.Y(n_180)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_16),
.Y(n_105)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_16),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_16),
.A2(n_103),
.B1(n_178),
.B2(n_180),
.Y(n_177)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_16),
.Y(n_195)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_16),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_16),
.A2(n_103),
.B1(n_258),
.B2(n_260),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_121),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_119),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_87),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_20),
.B(n_87),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_76),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_39),
.C(n_62),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_22),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_22),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_22),
.A2(n_62),
.B1(n_85),
.B2(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_31),
.B(n_36),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_23),
.A2(n_31),
.B1(n_99),
.B2(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_23),
.A2(n_31),
.B1(n_112),
.B2(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_23),
.B(n_168),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_23),
.A2(n_31),
.B1(n_227),
.B2(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_24),
.A2(n_37),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_24),
.A2(n_166),
.B(n_167),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_24),
.A2(n_97),
.B1(n_139),
.B2(n_166),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_24),
.B(n_172),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_24),
.A2(n_167),
.B(n_242),
.Y(n_280)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_25),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp33_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_30),
.B(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_30),
.B(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_31),
.B(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_33),
.A2(n_34),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

OAI21xp33_ASAP7_75t_L g232 ( 
.A1(n_33),
.A2(n_70),
.B(n_172),
.Y(n_232)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_34),
.B(n_253),
.Y(n_252)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_39),
.A2(n_77),
.B1(n_78),
.B2(n_86),
.Y(n_76)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_39),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_46),
.B1(n_54),
.B2(n_59),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_40),
.A2(n_54),
.B(n_115),
.Y(n_114)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_41),
.Y(n_171)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND3xp33_ASAP7_75t_SL g183 ( 
.A(n_42),
.B(n_52),
.C(n_58),
.Y(n_183)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_46),
.A2(n_54),
.B1(n_59),
.B2(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_46),
.A2(n_143),
.B(n_146),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_47),
.B(n_116),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_47),
.A2(n_147),
.B(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_47),
.A2(n_55),
.B1(n_144),
.B2(n_204),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_54),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_50),
.B(n_172),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_51),
.A2(n_52),
.B1(n_56),
.B2(n_58),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_51),
.A2(n_56),
.B(n_173),
.C(n_183),
.Y(n_182)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_54),
.B(n_117),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_54),
.A2(n_115),
.B(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_56),
.A2(n_58),
.B1(n_69),
.B2(n_70),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_62),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_66),
.B1(n_72),
.B2(n_73),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_64),
.A2(n_67),
.B1(n_68),
.B2(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_66),
.A2(n_72),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_66),
.B(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_68),
.B1(n_74),
.B2(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_67),
.A2(n_68),
.B1(n_95),
.B2(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_67),
.A2(n_200),
.B(n_201),
.Y(n_199)
);

OAI21xp33_ASAP7_75t_L g244 ( 
.A1(n_67),
.A2(n_201),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_68),
.A2(n_186),
.B(n_187),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_68),
.A2(n_141),
.B(n_187),
.Y(n_311)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_72),
.B(n_188),
.Y(n_201)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_92),
.C(n_100),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_88),
.A2(n_92),
.B1(n_93),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_88),
.Y(n_150)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_93),
.A2(n_94),
.B(n_96),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_97),
.A2(n_226),
.B(n_228),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_97),
.A2(n_228),
.B(n_256),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_100),
.B(n_149),
.Y(n_148)
);

AOI21xp33_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_109),
.B(n_113),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_101),
.A2(n_113),
.B1(n_114),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_101),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_101),
.A2(n_110),
.B1(n_111),
.B2(n_126),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_106),
.B(n_108),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_102),
.A2(n_108),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_102),
.A2(n_179),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_102),
.A2(n_105),
.B1(n_134),
.B2(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_102),
.A2(n_261),
.B(n_267),
.Y(n_281)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_103),
.B(n_236),
.Y(n_235)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_106),
.B(n_172),
.Y(n_265)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_151),
.B(n_332),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_148),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_123),
.B(n_148),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.C(n_129),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_124),
.A2(n_127),
.B1(n_128),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_124),
.Y(n_328)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_129),
.A2(n_130),
.B1(n_327),
.B2(n_329),
.Y(n_326)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_140),
.C(n_142),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_131),
.A2(n_132),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_133),
.A2(n_136),
.B1(n_137),
.B2(n_304),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_133),
.Y(n_304)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_135),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_135),
.A2(n_235),
.B(n_259),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_140),
.B(n_142),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_325),
.B(n_331),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_315),
.B(n_324),
.Y(n_152)
);

O2A1O1Ixp33_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_213),
.B(n_298),
.C(n_314),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_196),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_155),
.B(n_196),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_174),
.C(n_184),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_156),
.A2(n_157),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_169),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_164),
.B2(n_165),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_160),
.B(n_164),
.C(n_169),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_161),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_163),
.Y(n_200)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B(n_173),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_174),
.A2(n_175),
.B1(n_184),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_181),
.B2(n_182),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_181),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_180),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_184),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_189),
.C(n_191),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_221),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_222),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_191),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_192),
.A2(n_234),
.B(n_235),
.Y(n_233)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_205),
.B1(n_206),
.B2(n_212),
.Y(n_196)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

BUFx24_ASAP7_75t_SL g334 ( 
.A(n_197),
.Y(n_334)
);

FAx1_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_199),
.CI(n_202),
.CON(n_197),
.SN(n_197)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_198),
.B(n_199),
.C(n_202),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_211),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_207),
.B(n_211),
.C(n_212),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_208),
.B(n_210),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_291),
.B(n_297),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_246),
.B(n_290),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_238),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_218),
.B(n_238),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_223),
.B2(n_237),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_219),
.B(n_225),
.C(n_229),
.Y(n_296)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_223),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_229),
.B2(n_230),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_231),
.B(n_233),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_268),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.C(n_243),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_239),
.B(n_286),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_240),
.A2(n_243),
.B1(n_244),
.B2(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_240),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_284),
.B(n_289),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_274),
.B(n_283),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_262),
.B(n_273),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_257),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_257),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_254),
.Y(n_282)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_269),
.B(n_272),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_270),
.B(n_271),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_282),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_282),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_281),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_280),
.C(n_281),
.Y(n_288)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_288),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_288),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_296),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_296),
.Y(n_297)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_313),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_313),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_303),
.C(n_305),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_305),
.B2(n_306),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_312),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_310),
.C(n_312),
.Y(n_323)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_317),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_323),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_319),
.B(n_320),
.C(n_323),
.Y(n_330)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_330),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_330),
.Y(n_331)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_327),
.Y(n_329)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);


endmodule