module fake_jpeg_10464_n_248 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_248);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_248;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_21),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_23),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_20),
.B1(n_32),
.B2(n_27),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_44),
.A2(n_45),
.B1(n_51),
.B2(n_57),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_20),
.B1(n_32),
.B2(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_50),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_33),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_59),
.Y(n_69)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_33),
.B1(n_29),
.B2(n_27),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_55),
.B(n_24),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_30),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_20),
.B1(n_29),
.B2(n_32),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_23),
.B1(n_16),
.B2(n_26),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_58),
.A2(n_60),
.B1(n_22),
.B2(n_17),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_24),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_23),
.B1(n_26),
.B2(n_28),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_24),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_43),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_50),
.A2(n_30),
.B1(n_28),
.B2(n_22),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_64),
.A2(n_66),
.B1(n_44),
.B2(n_58),
.Y(n_98)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_68),
.Y(n_92)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_70),
.Y(n_107)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_72),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_49),
.B(n_56),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_74),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_18),
.Y(n_75)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_77),
.Y(n_102)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_18),
.Y(n_78)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_45),
.A2(n_43),
.B(n_40),
.C(n_16),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_54),
.B1(n_48),
.B2(n_46),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_17),
.Y(n_81)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_1),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_83),
.C(n_86),
.Y(n_109)
);

AOI21xp33_ASAP7_75t_L g83 ( 
.A1(n_62),
.A2(n_24),
.B(n_15),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_61),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_1),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_15),
.Y(n_85)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_46),
.B(n_40),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_55),
.B(n_16),
.Y(n_87)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_65),
.B(n_60),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_90),
.B(n_98),
.Y(n_123)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_96),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_95),
.A2(n_99),
.B1(n_103),
.B2(n_110),
.Y(n_124)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_77),
.A2(n_57),
.B1(n_48),
.B2(n_54),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_68),
.A2(n_48),
.B1(n_52),
.B2(n_24),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_105),
.B(n_111),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_85),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_67),
.B1(n_75),
.B2(n_81),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_80),
.A2(n_52),
.B1(n_3),
.B2(n_5),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_86),
.Y(n_125)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_113),
.B(n_116),
.Y(n_162)
);

AND2x4_ASAP7_75t_SL g114 ( 
.A(n_112),
.B(n_73),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_114),
.A2(n_119),
.B(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_118),
.Y(n_150)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_76),
.C(n_84),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_137),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_69),
.Y(n_121)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

OAI21xp33_ASAP7_75t_SL g140 ( 
.A1(n_122),
.A2(n_125),
.B(n_132),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_93),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_133),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_69),
.Y(n_127)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_129),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_74),
.Y(n_130)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_100),
.A2(n_79),
.B1(n_66),
.B2(n_80),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_110),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_82),
.Y(n_134)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_111),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_135),
.A2(n_114),
.B1(n_113),
.B2(n_116),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_101),
.Y(n_136)
);

NOR3xp33_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_78),
.C(n_86),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_65),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_133),
.A2(n_100),
.B1(n_79),
.B2(n_109),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_138),
.A2(n_145),
.B1(n_148),
.B2(n_152),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_141),
.A2(n_7),
.B(n_10),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_107),
.B1(n_70),
.B2(n_71),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_115),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_146),
.B(n_149),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_117),
.A2(n_94),
.B1(n_91),
.B2(n_89),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_131),
.Y(n_149)
);

AOI221xp5_ASAP7_75t_L g179 ( 
.A1(n_151),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.C(n_9),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_119),
.A2(n_118),
.B1(n_123),
.B2(n_130),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_122),
.B(n_91),
.Y(n_153)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

AO22x1_ASAP7_75t_SL g154 ( 
.A1(n_114),
.A2(n_82),
.B1(n_63),
.B2(n_89),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_154),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_126),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_157),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_135),
.Y(n_158)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_144),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_137),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_165),
.C(n_166),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_120),
.C(n_121),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_114),
.C(n_134),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_135),
.C(n_124),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_170),
.C(n_172),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_94),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_147),
.C(n_161),
.Y(n_172)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_173),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_136),
.C(n_128),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_175),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_150),
.A2(n_63),
.B(n_97),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_147),
.A2(n_97),
.B(n_3),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_176),
.A2(n_181),
.B1(n_154),
.B2(n_156),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_162),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_177),
.B(n_180),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_178),
.A2(n_148),
.B1(n_138),
.B2(n_154),
.Y(n_191)
);

AOI322xp5_ASAP7_75t_L g194 ( 
.A1(n_179),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_14),
.C2(n_139),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_159),
.B(n_156),
.Y(n_181)
);

INVxp33_ASAP7_75t_L g184 ( 
.A(n_182),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_186),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_183),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_144),
.Y(n_188)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_181),
.Y(n_189)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_197),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_176),
.A2(n_145),
.B1(n_140),
.B2(n_159),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_178),
.Y(n_201)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_174),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_152),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_199),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_183),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_200),
.A2(n_186),
.B1(n_193),
.B2(n_187),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_164),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_163),
.C(n_165),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_204),
.C(n_205),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_167),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_172),
.C(n_166),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_170),
.C(n_169),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_209),
.C(n_185),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_164),
.Y(n_209)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_210),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_213),
.A2(n_189),
.B1(n_187),
.B2(n_191),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_221),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_203),
.C(n_215),
.Y(n_225)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_211),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_200),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_223),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_212),
.A2(n_195),
.B(n_168),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_220),
.A2(n_202),
.B(n_188),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_206),
.A2(n_190),
.B(n_169),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_207),
.A2(n_180),
.B(n_192),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_185),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_212),
.B(n_199),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_227),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_209),
.C(n_205),
.Y(n_227)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_228),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_230),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_216),
.B(n_208),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_231),
.A2(n_221),
.B1(n_223),
.B2(n_214),
.Y(n_233)
);

INVxp67_ASAP7_75t_SL g232 ( 
.A(n_226),
.Y(n_232)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_232),
.Y(n_238)
);

AOI21x1_ASAP7_75t_SL g239 ( 
.A1(n_233),
.A2(n_217),
.B(n_227),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_224),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_236),
.B(n_143),
.Y(n_241)
);

OAI21xp33_ASAP7_75t_L g242 ( 
.A1(n_239),
.A2(n_241),
.B(n_232),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_225),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_234),
.Y(n_243)
);

AO21x1_ASAP7_75t_L g245 ( 
.A1(n_242),
.A2(n_244),
.B(n_238),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_237),
.C(n_12),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_239),
.Y(n_244)
);

AO21x1_ASAP7_75t_L g247 ( 
.A1(n_245),
.A2(n_246),
.B(n_11),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_14),
.Y(n_248)
);


endmodule