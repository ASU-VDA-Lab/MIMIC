module fake_netlist_6_163_n_1818 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1818);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1818;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g166 ( 
.A(n_44),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_102),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_47),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_16),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_63),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_58),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_110),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_42),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_96),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_16),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_141),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_118),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_104),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_138),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_127),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_142),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_139),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_89),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_76),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_6),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_54),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_98),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_87),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_91),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_103),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_79),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_28),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_144),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_117),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_68),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_35),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_93),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_38),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_109),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_13),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_69),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_97),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_72),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_159),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_15),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_121),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_44),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_75),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_35),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_40),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_24),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_0),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_84),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_135),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_24),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_13),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_136),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_17),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_29),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_53),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_43),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_60),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_55),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_130),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_83),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_0),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_9),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_164),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_143),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_149),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_132),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_150),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_61),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_48),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_125),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_41),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_29),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_28),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_131),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_86),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_9),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_106),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_108),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_21),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_26),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_47),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_30),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_115),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_77),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_82),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_95),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_23),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_100),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_3),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_88),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_30),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_4),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_128),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_19),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_52),
.Y(n_264)
);

BUFx2_ASAP7_75t_SL g265 ( 
.A(n_152),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_25),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_52),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_40),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_15),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_6),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_113),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_105),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_154),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_71),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_81),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_101),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_14),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_120),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_46),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_59),
.Y(n_280)
);

CKINVDCx12_ASAP7_75t_R g281 ( 
.A(n_85),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_54),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_156),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_80),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_1),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_37),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_160),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_27),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_163),
.Y(n_289)
);

BUFx10_ASAP7_75t_L g290 ( 
.A(n_17),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_65),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_70),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_27),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_64),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g295 ( 
.A(n_119),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_92),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_73),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_158),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_94),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_99),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_21),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_3),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_90),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_162),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_41),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_123),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_157),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_161),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_49),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_20),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_112),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_165),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_38),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_4),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_129),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_55),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_14),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_74),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_7),
.Y(n_319)
);

BUFx10_ASAP7_75t_L g320 ( 
.A(n_137),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_46),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_153),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_2),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_18),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_33),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_22),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_33),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_8),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_39),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_25),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_111),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_140),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_78),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_66),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_7),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_5),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_205),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_175),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_167),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_196),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_193),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_181),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_192),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_196),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_196),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_205),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_178),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_196),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_211),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_169),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_196),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_205),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_195),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_197),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_222),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_222),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_199),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_178),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_222),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_222),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_228),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_205),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_222),
.Y(n_363)
);

BUFx6f_ASAP7_75t_SL g364 ( 
.A(n_207),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_238),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_238),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_229),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_238),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_238),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_206),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_201),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_238),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_233),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_279),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_290),
.Y(n_375)
);

CKINVDCx14_ASAP7_75t_R g376 ( 
.A(n_290),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_200),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_205),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_232),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_203),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_212),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_252),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_206),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_286),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_278),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_256),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_169),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_304),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_286),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_286),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_308),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_218),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_286),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_286),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_172),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_226),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_313),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_313),
.Y(n_398)
);

CKINVDCx14_ASAP7_75t_R g399 ( 
.A(n_290),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_313),
.Y(n_400)
);

INVxp33_ASAP7_75t_SL g401 ( 
.A(n_189),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_210),
.Y(n_402)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_279),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_189),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_313),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_168),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_190),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_313),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_317),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_234),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_317),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_317),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_237),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_317),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_190),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_317),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_166),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_235),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_242),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_173),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_254),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_235),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_244),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_340),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_340),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_344),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_344),
.Y(n_427)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_346),
.Y(n_428)
);

AND3x2_ASAP7_75t_L g429 ( 
.A(n_375),
.B(n_267),
.C(n_241),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_346),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_346),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_395),
.A2(n_216),
.B1(n_258),
.B2(n_215),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_358),
.B(n_276),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_345),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_343),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_353),
.Y(n_436)
);

NOR2x1_ASAP7_75t_L g437 ( 
.A(n_358),
.B(n_273),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_354),
.B(n_176),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_349),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_346),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_360),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_345),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_348),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_360),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_357),
.B(n_176),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_339),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_349),
.A2(n_288),
.B1(n_324),
.B2(n_242),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_346),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_348),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_421),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_408),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_371),
.Y(n_452)
);

BUFx8_ASAP7_75t_L g453 ( 
.A(n_364),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_351),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_355),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_341),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_346),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_338),
.A2(n_293),
.B1(n_335),
.B2(n_377),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_352),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_358),
.B(n_276),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_370),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_380),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_395),
.B(n_402),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_381),
.B(n_177),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_392),
.B(n_396),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_376),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_355),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g468 ( 
.A(n_370),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_356),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_408),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_356),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_359),
.Y(n_472)
);

AND2x6_ASAP7_75t_L g473 ( 
.A(n_352),
.B(n_273),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_352),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_359),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_347),
.B(n_285),
.Y(n_476)
);

BUFx8_ASAP7_75t_L g477 ( 
.A(n_364),
.Y(n_477)
);

NAND2xp33_ASAP7_75t_L g478 ( 
.A(n_352),
.B(n_285),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_410),
.B(n_413),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_361),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_363),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_386),
.A2(n_293),
.B1(n_335),
.B2(n_314),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_418),
.B(n_166),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_352),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_423),
.B(n_191),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_367),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_342),
.A2(n_269),
.B1(n_266),
.B2(n_264),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_370),
.B(n_209),
.Y(n_488)
);

NAND2xp33_ASAP7_75t_L g489 ( 
.A(n_352),
.B(n_209),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_363),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_373),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_365),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_362),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_365),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_402),
.B(n_207),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_383),
.B(n_191),
.Y(n_496)
);

INVx4_ASAP7_75t_L g497 ( 
.A(n_362),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_382),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_366),
.Y(n_499)
);

INVx4_ASAP7_75t_L g500 ( 
.A(n_473),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_434),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_441),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_441),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_468),
.B(n_366),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_468),
.B(n_368),
.Y(n_505)
);

BUFx8_ASAP7_75t_SL g506 ( 
.A(n_446),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_466),
.B(n_401),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_444),
.Y(n_508)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_488),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_444),
.Y(n_510)
);

BUFx10_ASAP7_75t_L g511 ( 
.A(n_435),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_456),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_451),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_464),
.B(n_399),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_449),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_451),
.Y(n_516)
);

NAND3xp33_ASAP7_75t_L g517 ( 
.A(n_483),
.B(n_369),
.C(n_368),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_470),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_438),
.B(n_207),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_470),
.Y(n_520)
);

INVx2_ASAP7_75t_SL g521 ( 
.A(n_461),
.Y(n_521)
);

INVx5_ASAP7_75t_L g522 ( 
.A(n_473),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_445),
.B(n_320),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_483),
.B(n_422),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_476),
.A2(n_273),
.B1(n_316),
.B2(n_319),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_454),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_435),
.B(n_436),
.Y(n_527)
);

AO22x2_ASAP7_75t_L g528 ( 
.A1(n_495),
.A2(n_221),
.B1(n_194),
.B2(n_295),
.Y(n_528)
);

INVx4_ASAP7_75t_L g529 ( 
.A(n_473),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_461),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_486),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_485),
.B(n_364),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_476),
.A2(n_460),
.B1(n_433),
.B2(n_488),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_436),
.B(n_320),
.Y(n_534)
);

NOR3xp33_ASAP7_75t_L g535 ( 
.A(n_458),
.B(n_387),
.C(n_350),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_433),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_430),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_471),
.Y(n_538)
);

BUFx10_ASAP7_75t_L g539 ( 
.A(n_452),
.Y(n_539)
);

OA22x2_ASAP7_75t_L g540 ( 
.A1(n_432),
.A2(n_374),
.B1(n_403),
.B2(n_316),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_433),
.B(n_460),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_460),
.A2(n_261),
.B1(n_225),
.B2(n_319),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_430),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g544 ( 
.A(n_437),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_471),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_486),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_455),
.Y(n_547)
);

AND2x6_ASAP7_75t_L g548 ( 
.A(n_465),
.B(n_182),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_490),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_490),
.Y(n_550)
);

XNOR2x2_ASAP7_75t_R g551 ( 
.A(n_447),
.B(n_385),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_475),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_494),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_492),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_494),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_424),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_479),
.B(n_404),
.Y(n_557)
);

NOR2x1p5_ASAP7_75t_L g558 ( 
.A(n_452),
.B(n_225),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_424),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_425),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_425),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_426),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_496),
.B(n_383),
.Y(n_563)
);

OAI22xp33_ASAP7_75t_L g564 ( 
.A1(n_463),
.A2(n_227),
.B1(n_220),
.B2(n_323),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_439),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_426),
.Y(n_566)
);

INVx1_ASAP7_75t_SL g567 ( 
.A(n_491),
.Y(n_567)
);

NAND2xp33_ASAP7_75t_L g568 ( 
.A(n_473),
.B(n_232),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_427),
.B(n_369),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_427),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_442),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_442),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_491),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_443),
.Y(n_574)
);

NAND2xp33_ASAP7_75t_L g575 ( 
.A(n_473),
.B(n_232),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_443),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_467),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_467),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_462),
.B(n_453),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_430),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_469),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_462),
.B(n_320),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_469),
.Y(n_583)
);

INVx5_ASAP7_75t_L g584 ( 
.A(n_473),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g585 ( 
.A1(n_487),
.A2(n_224),
.B1(n_310),
.B2(n_309),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_472),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_472),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_482),
.A2(n_261),
.B1(n_248),
.B2(n_305),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_481),
.Y(n_589)
);

AOI21x1_ASAP7_75t_L g590 ( 
.A1(n_481),
.A2(n_378),
.B(n_337),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_430),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_499),
.A2(n_214),
.B1(n_245),
.B2(n_325),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_499),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_489),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_428),
.B(n_407),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_428),
.B(n_415),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_430),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_431),
.Y(n_598)
);

OR2x6_ASAP7_75t_L g599 ( 
.A(n_450),
.B(n_265),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_489),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_448),
.B(n_372),
.Y(n_601)
);

NAND3xp33_ASAP7_75t_L g602 ( 
.A(n_478),
.B(n_384),
.C(n_372),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_450),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_431),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_448),
.B(n_384),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_431),
.Y(n_606)
);

INVx1_ASAP7_75t_SL g607 ( 
.A(n_480),
.Y(n_607)
);

OAI22xp33_ASAP7_75t_L g608 ( 
.A1(n_453),
.A2(n_329),
.B1(n_213),
.B2(n_302),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_448),
.B(n_383),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_453),
.B(n_170),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_477),
.B(n_170),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_431),
.Y(n_612)
);

OR2x6_ASAP7_75t_L g613 ( 
.A(n_477),
.B(n_194),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_484),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_431),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_440),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_477),
.B(n_171),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_484),
.B(n_389),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_484),
.B(n_389),
.Y(n_619)
);

BUFx8_ASAP7_75t_SL g620 ( 
.A(n_498),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_429),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_428),
.B(n_390),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_440),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_497),
.B(n_390),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_497),
.B(n_171),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_440),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_440),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_440),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_457),
.Y(n_629)
);

INVxp67_ASAP7_75t_L g630 ( 
.A(n_478),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_473),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_497),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_457),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_457),
.Y(n_634)
);

AND2x2_ASAP7_75t_SL g635 ( 
.A(n_457),
.B(n_182),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_493),
.B(n_180),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_493),
.B(n_180),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_459),
.Y(n_638)
);

NAND2xp33_ASAP7_75t_SL g639 ( 
.A(n_459),
.B(n_419),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_459),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_459),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_459),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_474),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_474),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_474),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_474),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_474),
.Y(n_647)
);

AND3x2_ASAP7_75t_L g648 ( 
.A(n_493),
.B(n_217),
.C(n_236),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_493),
.A2(n_305),
.B1(n_248),
.B2(n_221),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_541),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_509),
.B(n_295),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_509),
.B(n_374),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_635),
.B(n_232),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_530),
.Y(n_654)
);

BUFx6f_ASAP7_75t_SL g655 ( 
.A(n_511),
.Y(n_655)
);

O2A1O1Ixp33_ASAP7_75t_L g656 ( 
.A1(n_630),
.A2(n_406),
.B(n_420),
.C(n_394),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_632),
.A2(n_493),
.B(n_362),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_635),
.B(n_232),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_541),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_635),
.B(n_259),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_524),
.B(n_403),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_558),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_548),
.A2(n_250),
.B1(n_202),
.B2(n_336),
.Y(n_663)
);

NAND3xp33_ASAP7_75t_L g664 ( 
.A(n_533),
.B(n_422),
.C(n_249),
.Y(n_664)
);

AND2x2_ASAP7_75t_SL g665 ( 
.A(n_588),
.B(n_236),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_567),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_609),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_558),
.Y(n_668)
);

NAND2xp33_ASAP7_75t_SL g669 ( 
.A(n_534),
.B(n_388),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_502),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_557),
.B(n_198),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_563),
.B(n_306),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_536),
.A2(n_391),
.B1(n_257),
.B2(n_262),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_561),
.Y(n_674)
);

OR2x6_ASAP7_75t_L g675 ( 
.A(n_565),
.B(n_422),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_563),
.B(n_174),
.Y(n_676)
);

NOR3xp33_ASAP7_75t_L g677 ( 
.A(n_603),
.B(n_270),
.C(n_204),
.Y(n_677)
);

NAND3xp33_ASAP7_75t_L g678 ( 
.A(n_595),
.B(n_321),
.C(n_326),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_502),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_536),
.B(n_179),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_524),
.B(n_183),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_501),
.B(n_186),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_503),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_503),
.Y(n_684)
);

XOR2x2_ASAP7_75t_L g685 ( 
.A(n_582),
.B(n_1),
.Y(n_685)
);

BUFx2_ASAP7_75t_L g686 ( 
.A(n_512),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_530),
.B(n_417),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_599),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_508),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_501),
.B(n_187),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_548),
.A2(n_251),
.B1(n_219),
.B2(n_223),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_508),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_506),
.Y(n_693)
);

OAI22xp33_ASAP7_75t_L g694 ( 
.A1(n_540),
.A2(n_255),
.B1(n_334),
.B2(n_333),
.Y(n_694)
);

O2A1O1Ixp5_ASAP7_75t_L g695 ( 
.A1(n_594),
.A2(n_337),
.B(n_378),
.C(n_379),
.Y(n_695)
);

AO221x1_ASAP7_75t_L g696 ( 
.A1(n_528),
.A2(n_312),
.B1(n_259),
.B2(n_231),
.C(n_240),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_596),
.A2(n_298),
.B1(n_247),
.B2(n_300),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_521),
.B(n_519),
.Y(n_698)
);

INVx4_ASAP7_75t_L g699 ( 
.A(n_530),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_521),
.B(n_184),
.Y(n_700)
);

NAND2x1p5_ASAP7_75t_L g701 ( 
.A(n_500),
.B(n_208),
.Y(n_701)
);

O2A1O1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_594),
.A2(n_600),
.B(n_570),
.C(n_574),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_510),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_510),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_548),
.A2(n_230),
.B1(n_330),
.B2(n_328),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_515),
.B(n_239),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_500),
.B(n_259),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_500),
.B(n_259),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_500),
.B(n_259),
.Y(n_709)
);

INVx4_ASAP7_75t_L g710 ( 
.A(n_522),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_566),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_523),
.B(n_184),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_540),
.A2(n_303),
.B1(n_307),
.B2(n_311),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_580),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_567),
.B(n_260),
.Y(n_715)
);

OR2x6_ASAP7_75t_L g716 ( 
.A(n_599),
.B(n_263),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_515),
.B(n_246),
.Y(n_717)
);

NOR2x1p5_ASAP7_75t_L g718 ( 
.A(n_531),
.B(n_546),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_570),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_514),
.B(n_185),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_576),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_620),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_564),
.B(n_185),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_540),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_513),
.Y(n_725)
);

A2O1A1Ixp33_ASAP7_75t_L g726 ( 
.A1(n_517),
.A2(n_253),
.B(n_284),
.C(n_275),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_544),
.B(n_188),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_513),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_576),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_526),
.B(n_299),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_548),
.A2(n_301),
.B1(n_327),
.B2(n_282),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_528),
.Y(n_732)
);

NAND3xp33_ASAP7_75t_L g733 ( 
.A(n_535),
.B(n_585),
.C(n_542),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_607),
.B(n_268),
.Y(n_734)
);

NAND3x1_ASAP7_75t_L g735 ( 
.A(n_551),
.B(n_277),
.C(n_414),
.Y(n_735)
);

NAND2xp33_ASAP7_75t_L g736 ( 
.A(n_548),
.B(n_271),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_544),
.B(n_188),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_511),
.B(n_243),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_529),
.B(n_312),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_526),
.B(n_243),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_529),
.B(n_312),
.Y(n_741)
);

CKINVDCx20_ASAP7_75t_R g742 ( 
.A(n_531),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_528),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_577),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_547),
.B(n_272),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_547),
.B(n_272),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_552),
.B(n_274),
.Y(n_747)
);

BUFx3_ASAP7_75t_L g748 ( 
.A(n_552),
.Y(n_748)
);

NOR2xp67_ASAP7_75t_SL g749 ( 
.A(n_522),
.B(n_362),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_632),
.A2(n_362),
.B(n_337),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_554),
.B(n_315),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_516),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_554),
.B(n_577),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_589),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_518),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_631),
.B(n_318),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_589),
.B(n_322),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_532),
.B(n_280),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_556),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_511),
.B(n_280),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_504),
.B(n_505),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_556),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_608),
.B(n_283),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_625),
.B(n_283),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_631),
.B(n_287),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_517),
.B(n_610),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_539),
.B(n_287),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_520),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_SL g769 ( 
.A1(n_607),
.A2(n_281),
.B1(n_289),
.B2(n_291),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_559),
.B(n_393),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_560),
.B(n_562),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_560),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_562),
.B(n_571),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_631),
.B(n_289),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_599),
.B(n_393),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_520),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_571),
.B(n_394),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_572),
.B(n_397),
.Y(n_778)
);

AND2x6_ASAP7_75t_SL g779 ( 
.A(n_599),
.B(n_397),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_631),
.B(n_291),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_611),
.B(n_292),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_572),
.B(n_416),
.Y(n_782)
);

HB1xp67_ASAP7_75t_L g783 ( 
.A(n_621),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_617),
.B(n_292),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_538),
.Y(n_785)
);

AND2x4_ASAP7_75t_L g786 ( 
.A(n_578),
.B(n_412),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_522),
.B(n_294),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_592),
.B(n_294),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_578),
.B(n_411),
.Y(n_789)
);

NOR2x1p5_ASAP7_75t_L g790 ( 
.A(n_546),
.B(n_296),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_621),
.B(n_296),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_581),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_581),
.B(n_411),
.Y(n_793)
);

OAI22xp5_ASAP7_75t_L g794 ( 
.A1(n_528),
.A2(n_297),
.B1(n_331),
.B2(n_332),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_636),
.B(n_332),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_538),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_637),
.B(n_331),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_522),
.B(n_297),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_583),
.B(n_2),
.Y(n_799)
);

NAND2xp33_ASAP7_75t_SL g800 ( 
.A(n_579),
.B(n_409),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_583),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_586),
.B(n_409),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_586),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_587),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_671),
.B(n_672),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_667),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_SL g807 ( 
.A(n_666),
.B(n_573),
.Y(n_807)
);

BUFx2_ASAP7_75t_L g808 ( 
.A(n_675),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_714),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_652),
.B(n_527),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_766),
.B(n_573),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_650),
.Y(n_812)
);

NAND3xp33_ASAP7_75t_SL g813 ( 
.A(n_720),
.B(n_525),
.C(n_639),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_659),
.B(n_613),
.Y(n_814)
);

OR2x2_ASAP7_75t_L g815 ( 
.A(n_734),
.B(n_507),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_672),
.B(n_593),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_766),
.B(n_522),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_761),
.B(n_548),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_661),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_738),
.B(n_760),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_674),
.B(n_548),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_693),
.Y(n_822)
);

AND2x6_ASAP7_75t_SL g823 ( 
.A(n_763),
.B(n_613),
.Y(n_823)
);

BUFx3_ASAP7_75t_L g824 ( 
.A(n_686),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_670),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_675),
.Y(n_826)
);

OR2x6_ASAP7_75t_SL g827 ( 
.A(n_722),
.B(n_551),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_748),
.B(n_613),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_L g829 ( 
.A1(n_651),
.A2(n_649),
.B1(n_613),
.B2(n_614),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_723),
.B(n_613),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_748),
.Y(n_831)
);

INVx5_ASAP7_75t_L g832 ( 
.A(n_714),
.Y(n_832)
);

HB1xp67_ASAP7_75t_L g833 ( 
.A(n_675),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_742),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_723),
.B(n_614),
.Y(n_835)
);

BUFx12f_ASAP7_75t_L g836 ( 
.A(n_718),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_715),
.B(n_569),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_759),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_733),
.B(n_522),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_714),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_679),
.Y(n_841)
);

BUFx8_ASAP7_75t_L g842 ( 
.A(n_655),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_711),
.B(n_622),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_707),
.A2(n_709),
.B(n_708),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_698),
.B(n_584),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_698),
.B(n_584),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_719),
.B(n_624),
.Y(n_847)
);

BUFx8_ASAP7_75t_SL g848 ( 
.A(n_655),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_654),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_683),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_684),
.Y(n_851)
);

BUFx2_ASAP7_75t_L g852 ( 
.A(n_783),
.Y(n_852)
);

NOR3xp33_ASAP7_75t_SL g853 ( 
.A(n_694),
.B(n_602),
.C(n_400),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_732),
.B(n_623),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_762),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_724),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_743),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_721),
.B(n_615),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_729),
.B(n_615),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_689),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_692),
.Y(n_861)
);

OR2x6_ASAP7_75t_L g862 ( 
.A(n_716),
.B(n_688),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_665),
.A2(n_696),
.B1(n_691),
.B2(n_663),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_687),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_720),
.A2(n_764),
.B1(n_758),
.B2(n_795),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_R g866 ( 
.A(n_669),
.B(n_568),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_744),
.B(n_615),
.Y(n_867)
);

NAND2x1p5_ASAP7_75t_L g868 ( 
.A(n_699),
.B(n_584),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_687),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_754),
.B(n_615),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_753),
.B(n_623),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_758),
.B(n_626),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_772),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_662),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_703),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_699),
.Y(n_876)
);

INVx5_ASAP7_75t_L g877 ( 
.A(n_710),
.Y(n_877)
);

OR2x6_ASAP7_75t_L g878 ( 
.A(n_716),
.B(n_602),
.Y(n_878)
);

NAND2x1p5_ASAP7_75t_L g879 ( 
.A(n_710),
.B(n_584),
.Y(n_879)
);

OAI221xp5_ASAP7_75t_L g880 ( 
.A1(n_788),
.A2(n_605),
.B1(n_618),
.B2(n_619),
.C(n_601),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_792),
.Y(n_881)
);

OAI21xp5_ASAP7_75t_L g882 ( 
.A1(n_702),
.A2(n_708),
.B(n_707),
.Y(n_882)
);

INVx4_ASAP7_75t_L g883 ( 
.A(n_786),
.Y(n_883)
);

INVx5_ASAP7_75t_L g884 ( 
.A(n_775),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_668),
.Y(n_885)
);

BUFx2_ASAP7_75t_L g886 ( 
.A(n_716),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_775),
.Y(n_887)
);

INVx1_ASAP7_75t_SL g888 ( 
.A(n_685),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_SL g889 ( 
.A(n_781),
.B(n_648),
.Y(n_889)
);

OAI22xp33_ASAP7_75t_L g890 ( 
.A1(n_713),
.A2(n_545),
.B1(n_549),
.B2(n_555),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_700),
.B(n_647),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_801),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_779),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_788),
.B(n_626),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_700),
.B(n_676),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_727),
.B(n_628),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_665),
.B(n_646),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_664),
.B(n_597),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_727),
.B(n_549),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_737),
.B(n_740),
.Y(n_900)
);

AND3x2_ASAP7_75t_SL g901 ( 
.A(n_763),
.B(n_8),
.C(n_10),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_704),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_786),
.Y(n_903)
);

OR2x6_ASAP7_75t_L g904 ( 
.A(n_735),
.B(n_550),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_803),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_725),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_804),
.Y(n_907)
);

NOR3xp33_ASAP7_75t_L g908 ( 
.A(n_769),
.B(n_575),
.C(n_550),
.Y(n_908)
);

NOR3xp33_ASAP7_75t_L g909 ( 
.A(n_781),
.B(n_555),
.C(n_553),
.Y(n_909)
);

OAI22xp33_ASAP7_75t_L g910 ( 
.A1(n_681),
.A2(n_553),
.B1(n_400),
.B2(n_405),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_790),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_728),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_673),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_677),
.B(n_597),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_737),
.B(n_580),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_740),
.B(n_628),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_745),
.B(n_646),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_771),
.B(n_598),
.Y(n_918)
);

AND2x6_ASAP7_75t_SL g919 ( 
.A(n_784),
.B(n_398),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_678),
.B(n_598),
.Y(n_920)
);

AOI22xp33_ASAP7_75t_SL g921 ( 
.A1(n_784),
.A2(n_362),
.B1(n_11),
.B2(n_12),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_767),
.B(n_604),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_773),
.Y(n_923)
);

INVx5_ASAP7_75t_L g924 ( 
.A(n_785),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_701),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_796),
.Y(n_926)
);

OR2x6_ASAP7_75t_L g927 ( 
.A(n_656),
.B(n_680),
.Y(n_927)
);

BUFx12f_ASAP7_75t_SL g928 ( 
.A(n_800),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_791),
.B(n_629),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_752),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_682),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_701),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_764),
.B(n_580),
.Y(n_933)
);

NAND2x1p5_ASAP7_75t_L g934 ( 
.A(n_749),
.B(n_537),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_SL g935 ( 
.A(n_712),
.B(n_645),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_690),
.B(n_604),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_755),
.Y(n_937)
);

BUFx3_ASAP7_75t_L g938 ( 
.A(n_706),
.Y(n_938)
);

BUFx4f_ASAP7_75t_L g939 ( 
.A(n_768),
.Y(n_939)
);

NOR2x1_ASAP7_75t_L g940 ( 
.A(n_751),
.B(n_634),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_745),
.B(n_634),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_799),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_776),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_770),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_746),
.B(n_633),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_797),
.A2(n_633),
.B(n_640),
.C(n_641),
.Y(n_946)
);

BUFx8_ASAP7_75t_L g947 ( 
.A(n_791),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_697),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_777),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_778),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_717),
.Y(n_951)
);

AOI22xp33_ASAP7_75t_L g952 ( 
.A1(n_663),
.A2(n_398),
.B1(n_643),
.B2(n_642),
.Y(n_952)
);

AOI22xp33_ASAP7_75t_L g953 ( 
.A1(n_691),
.A2(n_612),
.B1(n_643),
.B2(n_642),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_746),
.B(n_640),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_747),
.B(n_641),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_757),
.B(n_537),
.Y(n_956)
);

XOR2x2_ASAP7_75t_L g957 ( 
.A(n_794),
.B(n_10),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_797),
.A2(n_644),
.B1(n_543),
.B2(n_537),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_782),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_789),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_793),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_747),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_765),
.A2(n_644),
.B1(n_543),
.B2(n_627),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_802),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_765),
.A2(n_543),
.B1(n_627),
.B2(n_616),
.Y(n_965)
);

NAND3xp33_ASAP7_75t_SL g966 ( 
.A(n_705),
.B(n_638),
.C(n_616),
.Y(n_966)
);

NOR2x1p5_ASAP7_75t_L g967 ( 
.A(n_730),
.B(n_638),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_799),
.B(n_612),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_695),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_774),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_653),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_774),
.A2(n_606),
.B1(n_591),
.B2(n_580),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_726),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_653),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_780),
.A2(n_606),
.B1(n_591),
.B2(n_379),
.Y(n_975)
);

INVx1_ASAP7_75t_SL g976 ( 
.A(n_658),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_856),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_877),
.A2(n_756),
.B(n_780),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_876),
.Y(n_979)
);

INVx2_ASAP7_75t_SL g980 ( 
.A(n_852),
.Y(n_980)
);

BUFx4f_ASAP7_75t_SL g981 ( 
.A(n_836),
.Y(n_981)
);

BUFx2_ASAP7_75t_L g982 ( 
.A(n_824),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_865),
.A2(n_756),
.B1(n_736),
.B2(n_787),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_805),
.B(n_660),
.Y(n_984)
);

NOR3xp33_ASAP7_75t_L g985 ( 
.A(n_811),
.B(n_798),
.C(n_787),
.Y(n_985)
);

O2A1O1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_900),
.A2(n_942),
.B(n_895),
.C(n_830),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_962),
.B(n_705),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_863),
.A2(n_731),
.B1(n_741),
.B2(n_739),
.Y(n_988)
);

NOR2xp67_ASAP7_75t_L g989 ( 
.A(n_822),
.B(n_798),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_885),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_820),
.B(n_731),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_830),
.A2(n_739),
.B(n_750),
.C(n_657),
.Y(n_992)
);

NAND3xp33_ASAP7_75t_L g993 ( 
.A(n_894),
.B(n_379),
.C(n_378),
.Y(n_993)
);

INVx4_ASAP7_75t_L g994 ( 
.A(n_884),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_R g995 ( 
.A(n_911),
.B(n_122),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_810),
.B(n_11),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_894),
.A2(n_12),
.B(n_18),
.C(n_19),
.Y(n_997)
);

CKINVDCx20_ASAP7_75t_R g998 ( 
.A(n_834),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_856),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_819),
.B(n_20),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_819),
.B(n_837),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_863),
.A2(n_590),
.B1(n_23),
.B2(n_26),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_815),
.B(n_22),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_835),
.A2(n_31),
.B(n_32),
.C(n_34),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_831),
.B(n_148),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_857),
.Y(n_1006)
);

OAI21xp33_ASAP7_75t_L g1007 ( 
.A1(n_807),
.A2(n_31),
.B(n_32),
.Y(n_1007)
);

AOI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_948),
.A2(n_62),
.B1(n_146),
.B2(n_145),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_825),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_857),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_923),
.B(n_147),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_809),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_905),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_931),
.B(n_34),
.Y(n_1014)
);

NAND2xp33_ASAP7_75t_SL g1015 ( 
.A(n_866),
.B(n_36),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_832),
.A2(n_134),
.B(n_126),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_R g1017 ( 
.A(n_913),
.B(n_116),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_SL g1018 ( 
.A(n_884),
.B(n_114),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_816),
.B(n_107),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_905),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_835),
.A2(n_36),
.B(n_37),
.C(n_39),
.Y(n_1021)
);

INVx4_ASAP7_75t_L g1022 ( 
.A(n_884),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_812),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_R g1024 ( 
.A(n_928),
.B(n_67),
.Y(n_1024)
);

INVx3_ASAP7_75t_SL g1025 ( 
.A(n_893),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_938),
.B(n_951),
.Y(n_1026)
);

INVx6_ASAP7_75t_L g1027 ( 
.A(n_842),
.Y(n_1027)
);

O2A1O1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_813),
.A2(n_43),
.B(n_45),
.C(n_48),
.Y(n_1028)
);

AO32x2_ASAP7_75t_L g1029 ( 
.A1(n_829),
.A2(n_45),
.A3(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_806),
.Y(n_1030)
);

NAND3xp33_ASAP7_75t_L g1031 ( 
.A(n_921),
.B(n_50),
.C(n_51),
.Y(n_1031)
);

OAI22x1_ASAP7_75t_L g1032 ( 
.A1(n_888),
.A2(n_53),
.B1(n_56),
.B2(n_57),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_L g1033 ( 
.A1(n_813),
.A2(n_56),
.B1(n_57),
.B2(n_973),
.Y(n_1033)
);

AND2x2_ASAP7_75t_SL g1034 ( 
.A(n_889),
.B(n_828),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_899),
.B(n_944),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_929),
.A2(n_896),
.B(n_882),
.C(n_818),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_838),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_959),
.B(n_961),
.Y(n_1038)
);

INVx4_ASAP7_75t_L g1039 ( 
.A(n_876),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_841),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_855),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_828),
.B(n_887),
.Y(n_1042)
);

NOR3xp33_ASAP7_75t_SL g1043 ( 
.A(n_901),
.B(n_957),
.C(n_890),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_826),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_896),
.B(n_950),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_869),
.B(n_887),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_832),
.A2(n_844),
.B(n_817),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_844),
.A2(n_817),
.B(n_933),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_850),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_809),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_848),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_826),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_851),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_964),
.B(n_843),
.Y(n_1054)
);

BUFx8_ASAP7_75t_L g1055 ( 
.A(n_808),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_847),
.B(n_974),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_809),
.Y(n_1057)
);

INVxp67_ASAP7_75t_SL g1058 ( 
.A(n_876),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_974),
.B(n_872),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_860),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_919),
.B(n_869),
.Y(n_1061)
);

INVxp67_ASAP7_75t_L g1062 ( 
.A(n_833),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_876),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_864),
.B(n_833),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_SL g1065 ( 
.A(n_862),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_921),
.A2(n_976),
.B1(n_853),
.B2(n_897),
.Y(n_1066)
);

INVxp33_ASAP7_75t_SL g1067 ( 
.A(n_866),
.Y(n_1067)
);

NOR3xp33_ASAP7_75t_SL g1068 ( 
.A(n_901),
.B(n_890),
.C(n_854),
.Y(n_1068)
);

AND2x4_ASAP7_75t_L g1069 ( 
.A(n_814),
.B(n_874),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_916),
.B(n_917),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_941),
.B(n_945),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_809),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_861),
.Y(n_1073)
);

AOI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_927),
.A2(n_914),
.B1(n_967),
.B2(n_920),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_954),
.B(n_955),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_871),
.B(n_891),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_918),
.A2(n_969),
.B(n_972),
.Y(n_1077)
);

O2A1O1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_946),
.A2(n_908),
.B(n_927),
.C(n_839),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_873),
.Y(n_1079)
);

AOI21x1_ASAP7_75t_L g1080 ( 
.A1(n_915),
.A2(n_846),
.B(n_845),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_862),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_849),
.A2(n_879),
.B(n_956),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_875),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_881),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_902),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_853),
.A2(n_971),
.B(n_956),
.C(n_898),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_854),
.B(n_949),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_879),
.A2(n_839),
.B(n_868),
.Y(n_1088)
);

O2A1O1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_908),
.A2(n_927),
.B(n_907),
.C(n_892),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_926),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_898),
.A2(n_821),
.B(n_914),
.C(n_922),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_922),
.A2(n_909),
.B(n_920),
.C(n_940),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_949),
.B(n_960),
.Y(n_1093)
);

AO32x1_ASAP7_75t_L g1094 ( 
.A1(n_930),
.A2(n_937),
.A3(n_883),
.B1(n_906),
.B2(n_943),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_903),
.B(n_883),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_912),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_858),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_SL g1098 ( 
.A1(n_862),
.A2(n_886),
.B1(n_904),
.B2(n_814),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_903),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_966),
.A2(n_918),
.B(n_968),
.Y(n_1100)
);

O2A1O1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_904),
.A2(n_909),
.B(n_878),
.C(n_910),
.Y(n_1101)
);

O2A1O1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_904),
.A2(n_878),
.B(n_910),
.C(n_870),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_960),
.B(n_936),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_903),
.B(n_878),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_903),
.Y(n_1105)
);

A2O1A1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_939),
.A2(n_936),
.B(n_970),
.C(n_935),
.Y(n_1106)
);

INVx1_ASAP7_75t_SL g1107 ( 
.A(n_840),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_840),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_840),
.Y(n_1109)
);

O2A1O1Ixp33_ASAP7_75t_SL g1110 ( 
.A1(n_859),
.A2(n_867),
.B(n_966),
.C(n_880),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_939),
.A2(n_970),
.B(n_925),
.C(n_932),
.Y(n_1111)
);

O2A1O1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_953),
.A2(n_952),
.B(n_934),
.C(n_947),
.Y(n_1112)
);

INVxp67_ASAP7_75t_SL g1113 ( 
.A(n_840),
.Y(n_1113)
);

NAND3xp33_ASAP7_75t_SL g1114 ( 
.A(n_958),
.B(n_947),
.C(n_963),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_982),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1036),
.A2(n_925),
.B(n_932),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1045),
.B(n_970),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1054),
.B(n_970),
.Y(n_1118)
);

INVx2_ASAP7_75t_SL g1119 ( 
.A(n_990),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_996),
.B(n_827),
.Y(n_1120)
);

OAI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1100),
.A2(n_965),
.B(n_975),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_1047),
.A2(n_953),
.B(n_934),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1035),
.B(n_952),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_980),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_1104),
.B(n_924),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_1077),
.A2(n_924),
.B(n_823),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1082),
.A2(n_924),
.B(n_978),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1037),
.Y(n_1128)
);

NOR2xp67_ASAP7_75t_SL g1129 ( 
.A(n_1031),
.B(n_924),
.Y(n_1129)
);

AND2x4_ASAP7_75t_L g1130 ( 
.A(n_1104),
.B(n_1069),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1035),
.B(n_1038),
.Y(n_1131)
);

INVx8_ASAP7_75t_L g1132 ( 
.A(n_1012),
.Y(n_1132)
);

OAI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1100),
.A2(n_1078),
.B(n_1086),
.Y(n_1133)
);

NOR2x1_ASAP7_75t_SL g1134 ( 
.A(n_994),
.B(n_1022),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_1001),
.B(n_1034),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1038),
.A2(n_1070),
.B1(n_1075),
.B2(n_1071),
.Y(n_1136)
);

AO31x2_ASAP7_75t_L g1137 ( 
.A1(n_988),
.A2(n_1091),
.A3(n_1092),
.B(n_1002),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_983),
.A2(n_986),
.B(n_984),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_1039),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_988),
.A2(n_1019),
.B(n_993),
.Y(n_1140)
);

AOI31xp67_ASAP7_75t_L g1141 ( 
.A1(n_1074),
.A2(n_1019),
.A3(n_1011),
.B(n_1005),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_993),
.A2(n_1110),
.B(n_992),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_1051),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_1055),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_1069),
.B(n_1046),
.Y(n_1145)
);

AO21x2_ASAP7_75t_L g1146 ( 
.A1(n_985),
.A2(n_1080),
.B(n_1106),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_SL g1147 ( 
.A1(n_1111),
.A2(n_1002),
.B(n_1058),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1056),
.B(n_1059),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_991),
.A2(n_1087),
.B(n_1059),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_SL g1150 ( 
.A1(n_1102),
.A2(n_1011),
.B(n_1039),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1087),
.A2(n_1093),
.B(n_1056),
.Y(n_1151)
);

AO21x2_ASAP7_75t_L g1152 ( 
.A1(n_1114),
.A2(n_1066),
.B(n_1103),
.Y(n_1152)
);

AO31x2_ASAP7_75t_L g1153 ( 
.A1(n_1066),
.A2(n_1004),
.A3(n_1094),
.B(n_1003),
.Y(n_1153)
);

AO21x2_ASAP7_75t_L g1154 ( 
.A1(n_1068),
.A2(n_1095),
.B(n_1016),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1109),
.A2(n_1090),
.B(n_979),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1030),
.B(n_1041),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_1044),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_1067),
.B(n_1026),
.Y(n_1158)
);

AO22x2_ASAP7_75t_L g1159 ( 
.A1(n_1031),
.A2(n_1043),
.B1(n_987),
.B2(n_1029),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_SL g1160 ( 
.A1(n_1033),
.A2(n_1007),
.B(n_997),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1028),
.A2(n_1021),
.B(n_1014),
.Y(n_1161)
);

INVxp67_ASAP7_75t_L g1162 ( 
.A(n_1052),
.Y(n_1162)
);

BUFx10_ASAP7_75t_L g1163 ( 
.A(n_1061),
.Y(n_1163)
);

BUFx2_ASAP7_75t_L g1164 ( 
.A(n_998),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1109),
.A2(n_979),
.B(n_1063),
.Y(n_1165)
);

AOI211x1_ASAP7_75t_L g1166 ( 
.A1(n_1079),
.A2(n_1084),
.B(n_1010),
.C(n_1006),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1018),
.A2(n_1094),
.B(n_1113),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_1063),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1018),
.A2(n_1094),
.B(n_1042),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1013),
.B(n_1020),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1107),
.A2(n_1105),
.B(n_1099),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1107),
.A2(n_1049),
.B(n_1040),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1009),
.A2(n_1073),
.B(n_1060),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1053),
.B(n_1083),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_1055),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_1064),
.B(n_1081),
.Y(n_1176)
);

OAI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1096),
.A2(n_1085),
.B(n_989),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1008),
.A2(n_977),
.B(n_999),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1015),
.A2(n_1062),
.B(n_1000),
.C(n_1108),
.Y(n_1179)
);

O2A1O1Ixp5_ASAP7_75t_L g1180 ( 
.A1(n_1029),
.A2(n_1098),
.B(n_1065),
.C(n_1017),
.Y(n_1180)
);

O2A1O1Ixp5_ASAP7_75t_L g1181 ( 
.A1(n_1029),
.A2(n_1065),
.B(n_1032),
.C(n_1024),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1012),
.A2(n_1050),
.B(n_1072),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1012),
.A2(n_1050),
.B1(n_1072),
.B2(n_1057),
.Y(n_1183)
);

OR2x2_ASAP7_75t_SL g1184 ( 
.A(n_1027),
.B(n_1025),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1050),
.A2(n_1057),
.B(n_1072),
.Y(n_1185)
);

INVxp67_ASAP7_75t_SL g1186 ( 
.A(n_1108),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_981),
.A2(n_995),
.B(n_1027),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_SL g1188 ( 
.A1(n_1036),
.A2(n_1111),
.B(n_1112),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1047),
.A2(n_1077),
.B(n_1088),
.Y(n_1189)
);

AO32x2_ASAP7_75t_L g1190 ( 
.A1(n_1066),
.A2(n_1002),
.A3(n_988),
.B1(n_743),
.B2(n_732),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_986),
.A2(n_865),
.B(n_671),
.C(n_805),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_1012),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_SL g1193 ( 
.A1(n_1036),
.A2(n_1111),
.B(n_1112),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1045),
.B(n_1054),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_SL g1195 ( 
.A1(n_1031),
.A2(n_865),
.B(n_671),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_1001),
.B(n_962),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1023),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_980),
.Y(n_1198)
);

A2O1A1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_986),
.A2(n_865),
.B(n_671),
.C(n_805),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1036),
.A2(n_1076),
.B(n_1082),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1047),
.A2(n_1077),
.B(n_1088),
.Y(n_1201)
);

NAND2xp33_ASAP7_75t_L g1202 ( 
.A(n_1068),
.B(n_865),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1045),
.B(n_1054),
.Y(n_1203)
);

AO31x2_ASAP7_75t_L g1204 ( 
.A1(n_1036),
.A2(n_946),
.A3(n_1048),
.B(n_1086),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_1051),
.Y(n_1205)
);

BUFx5_ASAP7_75t_L g1206 ( 
.A(n_1097),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_SL g1207 ( 
.A1(n_1089),
.A2(n_1101),
.B(n_1078),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1067),
.A2(n_671),
.B1(n_865),
.B2(n_805),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1047),
.A2(n_1077),
.B(n_1088),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_1012),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1047),
.A2(n_1077),
.B(n_1088),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_SL g1212 ( 
.A1(n_1031),
.A2(n_865),
.B(n_671),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1045),
.B(n_1054),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1047),
.A2(n_1077),
.B(n_1088),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1047),
.A2(n_1077),
.B(n_1088),
.Y(n_1215)
);

AO21x1_ASAP7_75t_L g1216 ( 
.A1(n_1078),
.A2(n_865),
.B(n_900),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1023),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_1001),
.B(n_962),
.Y(n_1218)
);

AO31x2_ASAP7_75t_L g1219 ( 
.A1(n_1036),
.A2(n_946),
.A3(n_1048),
.B(n_1086),
.Y(n_1219)
);

AOI31xp67_ASAP7_75t_L g1220 ( 
.A1(n_983),
.A2(n_865),
.A3(n_933),
.B(n_968),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1047),
.A2(n_1077),
.B(n_1088),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1036),
.A2(n_1076),
.B(n_1082),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1036),
.A2(n_1076),
.B(n_1082),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_SL g1224 ( 
.A1(n_1031),
.A2(n_865),
.B(n_671),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1047),
.A2(n_1077),
.B(n_1088),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1036),
.A2(n_1076),
.B(n_1082),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1012),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_998),
.Y(n_1228)
);

NOR4xp25_ASAP7_75t_L g1229 ( 
.A(n_997),
.B(n_1021),
.C(n_1028),
.D(n_1031),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1036),
.A2(n_1076),
.B(n_1082),
.Y(n_1230)
);

AOI21x1_ASAP7_75t_L g1231 ( 
.A1(n_978),
.A2(n_1047),
.B(n_1082),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_SL g1232 ( 
.A1(n_1036),
.A2(n_1111),
.B(n_1112),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1045),
.A2(n_865),
.B1(n_805),
.B2(n_900),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1036),
.A2(n_1076),
.B(n_1082),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1023),
.Y(n_1235)
);

AND2x4_ASAP7_75t_L g1236 ( 
.A(n_1104),
.B(n_1069),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1037),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1036),
.A2(n_1076),
.B(n_1082),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1045),
.B(n_1054),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1036),
.A2(n_1076),
.B(n_1082),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_R g1241 ( 
.A(n_998),
.B(n_512),
.Y(n_1241)
);

O2A1O1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_986),
.A2(n_805),
.B(n_671),
.C(n_900),
.Y(n_1242)
);

BUFx2_ASAP7_75t_L g1243 ( 
.A(n_982),
.Y(n_1243)
);

NAND3xp33_ASAP7_75t_L g1244 ( 
.A(n_1043),
.B(n_671),
.C(n_865),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1012),
.Y(n_1245)
);

O2A1O1Ixp5_ASAP7_75t_L g1246 ( 
.A1(n_1036),
.A2(n_805),
.B(n_900),
.C(n_671),
.Y(n_1246)
);

INVx2_ASAP7_75t_SL g1247 ( 
.A(n_990),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1054),
.B(n_805),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1045),
.B(n_1054),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1047),
.A2(n_1077),
.B(n_1088),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1045),
.B(n_1054),
.Y(n_1251)
);

BUFx3_ASAP7_75t_L g1252 ( 
.A(n_982),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1045),
.B(n_1054),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1047),
.A2(n_1077),
.B(n_1088),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1036),
.A2(n_865),
.B(n_805),
.Y(n_1255)
);

CKINVDCx16_ASAP7_75t_R g1256 ( 
.A(n_998),
.Y(n_1256)
);

INVx4_ASAP7_75t_L g1257 ( 
.A(n_994),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1047),
.A2(n_1077),
.B(n_1088),
.Y(n_1258)
);

XNOR2x2_ASAP7_75t_SL g1259 ( 
.A(n_1031),
.B(n_865),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_990),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1047),
.A2(n_1077),
.B(n_1088),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1047),
.A2(n_1077),
.B(n_1088),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_982),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1047),
.A2(n_1077),
.B(n_1088),
.Y(n_1264)
);

OAI222xp33_ASAP7_75t_L g1265 ( 
.A1(n_1208),
.A2(n_1129),
.B1(n_1233),
.B2(n_1259),
.C1(n_1135),
.C2(n_1242),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1191),
.A2(n_1199),
.B(n_1246),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1156),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1190),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1189),
.A2(n_1209),
.B(n_1201),
.Y(n_1269)
);

OAI221xp5_ASAP7_75t_L g1270 ( 
.A1(n_1195),
.A2(n_1224),
.B1(n_1212),
.B2(n_1244),
.C(n_1255),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1211),
.A2(n_1215),
.B(n_1214),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1156),
.Y(n_1272)
);

AOI221xp5_ASAP7_75t_L g1273 ( 
.A1(n_1195),
.A2(n_1212),
.B1(n_1224),
.B2(n_1229),
.C(n_1160),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1158),
.B(n_1248),
.Y(n_1274)
);

AOI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1127),
.A2(n_1222),
.B(n_1200),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1221),
.A2(n_1250),
.B(n_1225),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1252),
.Y(n_1277)
);

CKINVDCx6p67_ASAP7_75t_R g1278 ( 
.A(n_1228),
.Y(n_1278)
);

INVx8_ASAP7_75t_L g1279 ( 
.A(n_1132),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1263),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1194),
.B(n_1203),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1152),
.Y(n_1282)
);

BUFx10_ASAP7_75t_L g1283 ( 
.A(n_1143),
.Y(n_1283)
);

NAND2xp33_ASAP7_75t_SL g1284 ( 
.A(n_1131),
.B(n_1136),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1254),
.A2(n_1261),
.B(n_1258),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1159),
.B(n_1131),
.Y(n_1286)
);

NAND3xp33_ASAP7_75t_L g1287 ( 
.A(n_1202),
.B(n_1161),
.C(n_1160),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1262),
.A2(n_1264),
.B(n_1231),
.Y(n_1288)
);

BUFx8_ASAP7_75t_L g1289 ( 
.A(n_1164),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1159),
.B(n_1136),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1237),
.Y(n_1291)
);

INVx1_ASAP7_75t_SL g1292 ( 
.A(n_1115),
.Y(n_1292)
);

OAI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1161),
.A2(n_1233),
.B(n_1149),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1206),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1116),
.A2(n_1226),
.B(n_1240),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1243),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1223),
.A2(n_1238),
.B(n_1234),
.Y(n_1297)
);

AND2x4_ASAP7_75t_L g1298 ( 
.A(n_1125),
.B(n_1130),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1230),
.A2(n_1126),
.B(n_1142),
.Y(n_1299)
);

BUFx2_ASAP7_75t_L g1300 ( 
.A(n_1152),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_1157),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1206),
.Y(n_1302)
);

AOI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1167),
.A2(n_1169),
.B(n_1138),
.Y(n_1303)
);

OA21x2_ASAP7_75t_L g1304 ( 
.A1(n_1133),
.A2(n_1138),
.B(n_1140),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1142),
.A2(n_1140),
.B(n_1155),
.Y(n_1305)
);

OAI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1229),
.A2(n_1150),
.B(n_1151),
.Y(n_1306)
);

CKINVDCx20_ASAP7_75t_R g1307 ( 
.A(n_1241),
.Y(n_1307)
);

OA21x2_ASAP7_75t_L g1308 ( 
.A1(n_1133),
.A2(n_1121),
.B(n_1207),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1117),
.B(n_1148),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1206),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1172),
.A2(n_1188),
.B(n_1232),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1193),
.A2(n_1165),
.B(n_1171),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1213),
.B(n_1239),
.Y(n_1313)
);

AO21x2_ASAP7_75t_L g1314 ( 
.A1(n_1216),
.A2(n_1146),
.B(n_1147),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1190),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1196),
.A2(n_1218),
.B1(n_1120),
.B2(n_1145),
.Y(n_1316)
);

AOI221xp5_ASAP7_75t_L g1317 ( 
.A1(n_1181),
.A2(n_1180),
.B1(n_1166),
.B2(n_1251),
.C(n_1249),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1178),
.A2(n_1177),
.B(n_1117),
.Y(n_1318)
);

NAND2x1p5_ASAP7_75t_L g1319 ( 
.A(n_1125),
.B(n_1257),
.Y(n_1319)
);

OAI222xp33_ASAP7_75t_L g1320 ( 
.A1(n_1213),
.A2(n_1253),
.B1(n_1251),
.B2(n_1148),
.C1(n_1118),
.C2(n_1123),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1197),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1177),
.A2(n_1173),
.B(n_1183),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1141),
.A2(n_1253),
.B(n_1220),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1183),
.A2(n_1182),
.B(n_1185),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1217),
.Y(n_1325)
);

AO21x1_ASAP7_75t_L g1326 ( 
.A1(n_1123),
.A2(n_1190),
.B(n_1153),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1206),
.Y(n_1327)
);

INVx4_ASAP7_75t_SL g1328 ( 
.A(n_1137),
.Y(n_1328)
);

AO21x2_ASAP7_75t_L g1329 ( 
.A1(n_1146),
.A2(n_1154),
.B(n_1179),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1235),
.Y(n_1330)
);

AND2x4_ASAP7_75t_L g1331 ( 
.A(n_1130),
.B(n_1236),
.Y(n_1331)
);

OA21x2_ASAP7_75t_L g1332 ( 
.A1(n_1174),
.A2(n_1204),
.B(n_1219),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1170),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1256),
.B(n_1145),
.Y(n_1334)
);

CKINVDCx20_ASAP7_75t_R g1335 ( 
.A(n_1184),
.Y(n_1335)
);

OA21x2_ASAP7_75t_L g1336 ( 
.A1(n_1174),
.A2(n_1204),
.B(n_1219),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1176),
.B(n_1236),
.Y(n_1337)
);

OA21x2_ASAP7_75t_L g1338 ( 
.A1(n_1204),
.A2(n_1219),
.B(n_1137),
.Y(n_1338)
);

BUFx10_ASAP7_75t_L g1339 ( 
.A(n_1205),
.Y(n_1339)
);

OAI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1170),
.A2(n_1162),
.B(n_1186),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1176),
.B(n_1198),
.Y(n_1341)
);

AO21x2_ASAP7_75t_L g1342 ( 
.A1(n_1154),
.A2(n_1134),
.B(n_1153),
.Y(n_1342)
);

AND2x6_ASAP7_75t_L g1343 ( 
.A(n_1139),
.B(n_1168),
.Y(n_1343)
);

OAI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1187),
.A2(n_1257),
.B(n_1124),
.Y(n_1344)
);

CKINVDCx14_ASAP7_75t_R g1345 ( 
.A(n_1163),
.Y(n_1345)
);

OAI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1206),
.A2(n_1119),
.B(n_1247),
.Y(n_1346)
);

OA21x2_ASAP7_75t_L g1347 ( 
.A1(n_1137),
.A2(n_1153),
.B(n_1144),
.Y(n_1347)
);

AOI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1192),
.A2(n_1210),
.B(n_1227),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_L g1349 ( 
.A(n_1163),
.B(n_1260),
.Y(n_1349)
);

OR2x6_ASAP7_75t_L g1350 ( 
.A(n_1132),
.B(n_1175),
.Y(n_1350)
);

OA21x2_ASAP7_75t_L g1351 ( 
.A1(n_1192),
.A2(n_1210),
.B(n_1227),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1210),
.Y(n_1352)
);

AOI21xp33_ASAP7_75t_L g1353 ( 
.A1(n_1227),
.A2(n_1245),
.B(n_1132),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1245),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1245),
.B(n_1255),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_SL g1356 ( 
.A1(n_1244),
.A2(n_671),
.B1(n_962),
.B2(n_805),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1128),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1189),
.A2(n_1209),
.B(n_1201),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_1252),
.Y(n_1359)
);

AOI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1244),
.A2(n_671),
.B1(n_491),
.B2(n_486),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1156),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1248),
.B(n_1194),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1156),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1255),
.B(n_1159),
.Y(n_1364)
);

AND2x2_ASAP7_75t_SL g1365 ( 
.A(n_1229),
.B(n_1202),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1157),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1244),
.A2(n_671),
.B1(n_1202),
.B2(n_805),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1248),
.B(n_1194),
.Y(n_1368)
);

O2A1O1Ixp5_ASAP7_75t_L g1369 ( 
.A1(n_1161),
.A2(n_805),
.B(n_671),
.C(n_1191),
.Y(n_1369)
);

OAI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1191),
.A2(n_865),
.B(n_671),
.Y(n_1370)
);

HB1xp67_ASAP7_75t_L g1371 ( 
.A(n_1157),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1189),
.A2(n_1209),
.B(n_1201),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1248),
.B(n_1194),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1156),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1244),
.A2(n_671),
.B1(n_1202),
.B2(n_805),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1156),
.Y(n_1376)
);

OAI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1191),
.A2(n_865),
.B(n_671),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1156),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1156),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1189),
.A2(n_1209),
.B(n_1201),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1156),
.Y(n_1381)
);

AO21x2_ASAP7_75t_L g1382 ( 
.A1(n_1138),
.A2(n_1140),
.B(n_1142),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1128),
.Y(n_1383)
);

AO21x2_ASAP7_75t_L g1384 ( 
.A1(n_1138),
.A2(n_1140),
.B(n_1142),
.Y(n_1384)
);

AO21x2_ASAP7_75t_L g1385 ( 
.A1(n_1138),
.A2(n_1140),
.B(n_1142),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1157),
.Y(n_1386)
);

O2A1O1Ixp33_ASAP7_75t_L g1387 ( 
.A1(n_1195),
.A2(n_805),
.B(n_671),
.C(n_1212),
.Y(n_1387)
);

CKINVDCx16_ASAP7_75t_R g1388 ( 
.A(n_1241),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1208),
.A2(n_865),
.B1(n_671),
.B2(n_962),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1152),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1189),
.A2(n_1209),
.B(n_1201),
.Y(n_1391)
);

INVx2_ASAP7_75t_SL g1392 ( 
.A(n_1132),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1244),
.A2(n_671),
.B1(n_1202),
.B2(n_805),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1255),
.B(n_1159),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1189),
.A2(n_1209),
.B(n_1201),
.Y(n_1395)
);

OAI22x1_ASAP7_75t_L g1396 ( 
.A1(n_1244),
.A2(n_1208),
.B1(n_865),
.B2(n_962),
.Y(n_1396)
);

INVx2_ASAP7_75t_SL g1397 ( 
.A(n_1132),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1122),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1148),
.B(n_1152),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1128),
.Y(n_1400)
);

OAI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1191),
.A2(n_865),
.B(n_671),
.Y(n_1401)
);

OA21x2_ASAP7_75t_L g1402 ( 
.A1(n_1133),
.A2(n_1138),
.B(n_1140),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1189),
.A2(n_1209),
.B(n_1201),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1189),
.A2(n_1209),
.B(n_1201),
.Y(n_1404)
);

OAI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1191),
.A2(n_865),
.B(n_671),
.Y(n_1405)
);

AOI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1244),
.A2(n_671),
.B1(n_491),
.B2(n_486),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1128),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1270),
.B(n_1287),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1274),
.B(n_1396),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_SL g1410 ( 
.A1(n_1370),
.A2(n_1401),
.B(n_1377),
.Y(n_1410)
);

O2A1O1Ixp5_ASAP7_75t_L g1411 ( 
.A1(n_1405),
.A2(n_1369),
.B(n_1306),
.C(n_1293),
.Y(n_1411)
);

CKINVDCx16_ASAP7_75t_R g1412 ( 
.A(n_1388),
.Y(n_1412)
);

CKINVDCx16_ASAP7_75t_R g1413 ( 
.A(n_1307),
.Y(n_1413)
);

O2A1O1Ixp33_ASAP7_75t_L g1414 ( 
.A1(n_1389),
.A2(n_1387),
.B(n_1265),
.C(n_1367),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1281),
.B(n_1313),
.Y(n_1415)
);

OA22x2_ASAP7_75t_L g1416 ( 
.A1(n_1396),
.A2(n_1340),
.B1(n_1360),
.B2(n_1406),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1333),
.Y(n_1417)
);

INVx1_ASAP7_75t_SL g1418 ( 
.A(n_1292),
.Y(n_1418)
);

NAND3xp33_ASAP7_75t_L g1419 ( 
.A(n_1375),
.B(n_1393),
.C(n_1356),
.Y(n_1419)
);

AOI21x1_ASAP7_75t_SL g1420 ( 
.A1(n_1364),
.A2(n_1394),
.B(n_1290),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_SL g1421 ( 
.A1(n_1335),
.A2(n_1307),
.B1(n_1365),
.B2(n_1345),
.Y(n_1421)
);

AOI21xp5_ASAP7_75t_SL g1422 ( 
.A1(n_1362),
.A2(n_1373),
.B(n_1368),
.Y(n_1422)
);

AOI21x1_ASAP7_75t_SL g1423 ( 
.A1(n_1364),
.A2(n_1394),
.B(n_1290),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1365),
.A2(n_1273),
.B1(n_1267),
.B2(n_1363),
.Y(n_1424)
);

CKINVDCx11_ASAP7_75t_R g1425 ( 
.A(n_1283),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1272),
.A2(n_1361),
.B1(n_1374),
.B2(n_1381),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1376),
.A2(n_1379),
.B1(n_1378),
.B2(n_1402),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1277),
.Y(n_1428)
);

INVxp67_ASAP7_75t_L g1429 ( 
.A(n_1301),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1304),
.A2(n_1402),
.B1(n_1316),
.B2(n_1335),
.Y(n_1430)
);

INVx3_ASAP7_75t_SL g1431 ( 
.A(n_1278),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1309),
.B(n_1366),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1309),
.B(n_1341),
.Y(n_1433)
);

O2A1O1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1320),
.A2(n_1344),
.B(n_1371),
.C(n_1386),
.Y(n_1434)
);

NOR2xp67_ASAP7_75t_L g1435 ( 
.A(n_1349),
.B(n_1334),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1337),
.B(n_1278),
.Y(n_1436)
);

O2A1O1Ixp33_ASAP7_75t_L g1437 ( 
.A1(n_1382),
.A2(n_1385),
.B(n_1384),
.C(n_1317),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1331),
.B(n_1298),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1304),
.A2(n_1308),
.B1(n_1286),
.B2(n_1325),
.Y(n_1439)
);

AOI21xp5_ASAP7_75t_SL g1440 ( 
.A1(n_1346),
.A2(n_1350),
.B(n_1308),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1308),
.A2(n_1321),
.B1(n_1330),
.B2(n_1345),
.Y(n_1441)
);

A2O1A1Ixp33_ASAP7_75t_L g1442 ( 
.A1(n_1311),
.A2(n_1284),
.B(n_1297),
.C(n_1295),
.Y(n_1442)
);

AOI21x1_ASAP7_75t_SL g1443 ( 
.A1(n_1355),
.A2(n_1354),
.B(n_1329),
.Y(n_1443)
);

AOI221x1_ASAP7_75t_SL g1444 ( 
.A1(n_1291),
.A2(n_1407),
.B1(n_1400),
.B2(n_1383),
.C(n_1357),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1399),
.A2(n_1407),
.B1(n_1400),
.B2(n_1350),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_SL g1446 ( 
.A1(n_1350),
.A2(n_1384),
.B(n_1382),
.Y(n_1446)
);

AOI21x1_ASAP7_75t_SL g1447 ( 
.A1(n_1329),
.A2(n_1347),
.B(n_1326),
.Y(n_1447)
);

AOI21x1_ASAP7_75t_SL g1448 ( 
.A1(n_1329),
.A2(n_1347),
.B(n_1326),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1296),
.B(n_1382),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1352),
.B(n_1347),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1332),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1280),
.A2(n_1359),
.B1(n_1390),
.B2(n_1300),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1311),
.A2(n_1295),
.B(n_1385),
.Y(n_1453)
);

O2A1O1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1384),
.A2(n_1385),
.B(n_1323),
.C(n_1314),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1280),
.A2(n_1359),
.B1(n_1390),
.B2(n_1300),
.Y(n_1455)
);

AOI21xp5_ASAP7_75t_SL g1456 ( 
.A1(n_1319),
.A2(n_1397),
.B(n_1392),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1282),
.A2(n_1268),
.B1(n_1315),
.B2(n_1319),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_SL g1458 ( 
.A1(n_1319),
.A2(n_1397),
.B1(n_1392),
.B2(n_1351),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1338),
.B(n_1336),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1351),
.B(n_1328),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1282),
.A2(n_1268),
.B1(n_1315),
.B2(n_1338),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1338),
.A2(n_1332),
.B1(n_1336),
.B2(n_1303),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1336),
.A2(n_1303),
.B1(n_1327),
.B2(n_1294),
.Y(n_1463)
);

NOR2xp67_ASAP7_75t_L g1464 ( 
.A(n_1294),
.B(n_1327),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1302),
.A2(n_1310),
.B1(n_1275),
.B2(n_1279),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1318),
.Y(n_1466)
);

O2A1O1Ixp33_ASAP7_75t_L g1467 ( 
.A1(n_1314),
.A2(n_1353),
.B(n_1398),
.C(n_1310),
.Y(n_1467)
);

INVx1_ASAP7_75t_SL g1468 ( 
.A(n_1283),
.Y(n_1468)
);

AOI211xp5_ASAP7_75t_L g1469 ( 
.A1(n_1299),
.A2(n_1305),
.B(n_1312),
.C(n_1322),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1339),
.B(n_1289),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1289),
.B(n_1343),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1351),
.B(n_1342),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_SL g1473 ( 
.A1(n_1279),
.A2(n_1339),
.B(n_1343),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1348),
.Y(n_1474)
);

AOI21x1_ASAP7_75t_SL g1475 ( 
.A1(n_1342),
.A2(n_1324),
.B(n_1328),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1324),
.Y(n_1476)
);

INVx3_ASAP7_75t_SL g1477 ( 
.A(n_1279),
.Y(n_1477)
);

BUFx4f_ASAP7_75t_L g1478 ( 
.A(n_1343),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1288),
.A2(n_1269),
.B1(n_1271),
.B2(n_1276),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1288),
.B(n_1269),
.Y(n_1480)
);

AOI21x1_ASAP7_75t_SL g1481 ( 
.A1(n_1271),
.A2(n_1276),
.B(n_1285),
.Y(n_1481)
);

AOI21xp5_ASAP7_75t_SL g1482 ( 
.A1(n_1358),
.A2(n_1372),
.B(n_1380),
.Y(n_1482)
);

NOR2xp67_ASAP7_75t_L g1483 ( 
.A(n_1372),
.B(n_1380),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1391),
.B(n_1395),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1395),
.B(n_1403),
.Y(n_1485)
);

OA21x2_ASAP7_75t_L g1486 ( 
.A1(n_1404),
.A2(n_1306),
.B(n_1266),
.Y(n_1486)
);

O2A1O1Ixp5_ASAP7_75t_L g1487 ( 
.A1(n_1370),
.A2(n_1377),
.B(n_1405),
.C(n_1401),
.Y(n_1487)
);

AOI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1370),
.A2(n_1401),
.B(n_1377),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1370),
.A2(n_1401),
.B(n_1377),
.Y(n_1489)
);

A2O1A1Ixp33_ASAP7_75t_L g1490 ( 
.A1(n_1387),
.A2(n_865),
.B(n_671),
.C(n_1195),
.Y(n_1490)
);

AOI221xp5_ASAP7_75t_L g1491 ( 
.A1(n_1389),
.A2(n_671),
.B1(n_1244),
.B2(n_1377),
.C(n_1370),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1274),
.B(n_1396),
.Y(n_1492)
);

O2A1O1Ixp5_ASAP7_75t_L g1493 ( 
.A1(n_1370),
.A2(n_1377),
.B(n_1405),
.C(n_1401),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1281),
.B(n_1313),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1281),
.B(n_1313),
.Y(n_1495)
);

AOI221x1_ASAP7_75t_SL g1496 ( 
.A1(n_1389),
.A2(n_1244),
.B1(n_1287),
.B2(n_671),
.C(n_1031),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1451),
.Y(n_1497)
);

AOI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1479),
.A2(n_1483),
.B(n_1453),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1445),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1459),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1461),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1439),
.B(n_1457),
.Y(n_1502)
);

AO21x2_ASAP7_75t_L g1503 ( 
.A1(n_1488),
.A2(n_1489),
.B(n_1410),
.Y(n_1503)
);

INVx2_ASAP7_75t_SL g1504 ( 
.A(n_1484),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1417),
.B(n_1424),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1439),
.B(n_1457),
.Y(n_1506)
);

AO31x2_ASAP7_75t_L g1507 ( 
.A1(n_1462),
.A2(n_1461),
.A3(n_1463),
.B(n_1490),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1472),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1450),
.B(n_1486),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1466),
.Y(n_1510)
);

BUFx2_ASAP7_75t_L g1511 ( 
.A(n_1486),
.Y(n_1511)
);

OAI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1487),
.A2(n_1493),
.B(n_1491),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1462),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1427),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1463),
.B(n_1476),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1445),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1427),
.Y(n_1517)
);

AOI221xp5_ASAP7_75t_L g1518 ( 
.A1(n_1496),
.A2(n_1414),
.B1(n_1419),
.B2(n_1411),
.C(n_1424),
.Y(n_1518)
);

INVxp67_ASAP7_75t_L g1519 ( 
.A(n_1449),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1485),
.Y(n_1520)
);

CKINVDCx11_ASAP7_75t_R g1521 ( 
.A(n_1431),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1441),
.B(n_1452),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1454),
.B(n_1460),
.Y(n_1523)
);

AOI21xp33_ASAP7_75t_L g1524 ( 
.A1(n_1408),
.A2(n_1416),
.B(n_1437),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1480),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1469),
.B(n_1446),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1430),
.B(n_1442),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_L g1528 ( 
.A1(n_1475),
.A2(n_1481),
.B(n_1447),
.Y(n_1528)
);

INVx4_ASAP7_75t_L g1529 ( 
.A(n_1478),
.Y(n_1529)
);

AO21x2_ASAP7_75t_L g1530 ( 
.A1(n_1465),
.A2(n_1482),
.B(n_1430),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1474),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1409),
.B(n_1492),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1422),
.B(n_1426),
.Y(n_1533)
);

INVx3_ASAP7_75t_SL g1534 ( 
.A(n_1416),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1440),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_SL g1536 ( 
.A(n_1434),
.B(n_1426),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1467),
.Y(n_1537)
);

INVxp67_ASAP7_75t_L g1538 ( 
.A(n_1455),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1444),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1433),
.B(n_1432),
.Y(n_1540)
);

AO21x2_ASAP7_75t_L g1541 ( 
.A1(n_1464),
.A2(n_1448),
.B(n_1494),
.Y(n_1541)
);

INVx3_ASAP7_75t_L g1542 ( 
.A(n_1478),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1458),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1429),
.B(n_1418),
.Y(n_1544)
);

OA21x2_ASAP7_75t_L g1545 ( 
.A1(n_1415),
.A2(n_1495),
.B(n_1443),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1497),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1509),
.B(n_1438),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1510),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1531),
.Y(n_1549)
);

BUFx2_ASAP7_75t_L g1550 ( 
.A(n_1525),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1509),
.B(n_1435),
.Y(n_1551)
);

BUFx3_ASAP7_75t_L g1552 ( 
.A(n_1520),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1519),
.B(n_1436),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1519),
.B(n_1468),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1500),
.B(n_1456),
.Y(n_1555)
);

INVxp67_ASAP7_75t_SL g1556 ( 
.A(n_1531),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_1528),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1500),
.Y(n_1558)
);

NAND2x1_ASAP7_75t_L g1559 ( 
.A(n_1529),
.B(n_1473),
.Y(n_1559)
);

AND2x4_ASAP7_75t_L g1560 ( 
.A(n_1520),
.B(n_1471),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1534),
.A2(n_1421),
.B1(n_1412),
.B2(n_1470),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_SL g1562 ( 
.A1(n_1503),
.A2(n_1413),
.B1(n_1420),
.B2(n_1423),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1520),
.B(n_1428),
.Y(n_1563)
);

INVxp67_ASAP7_75t_L g1564 ( 
.A(n_1541),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1508),
.Y(n_1565)
);

INVx1_ASAP7_75t_SL g1566 ( 
.A(n_1511),
.Y(n_1566)
);

OAI221xp5_ASAP7_75t_L g1567 ( 
.A1(n_1518),
.A2(n_1425),
.B1(n_1477),
.B2(n_1512),
.C(n_1534),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1515),
.B(n_1507),
.Y(n_1568)
);

BUFx2_ASAP7_75t_L g1569 ( 
.A(n_1504),
.Y(n_1569)
);

INVx1_ASAP7_75t_SL g1570 ( 
.A(n_1508),
.Y(n_1570)
);

AO21x2_ASAP7_75t_L g1571 ( 
.A1(n_1564),
.A2(n_1524),
.B(n_1537),
.Y(n_1571)
);

BUFx2_ASAP7_75t_L g1572 ( 
.A(n_1569),
.Y(n_1572)
);

NAND3xp33_ASAP7_75t_SL g1573 ( 
.A(n_1567),
.B(n_1518),
.C(n_1512),
.Y(n_1573)
);

OAI221xp5_ASAP7_75t_L g1574 ( 
.A1(n_1567),
.A2(n_1534),
.B1(n_1524),
.B2(n_1533),
.C(n_1536),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1546),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1553),
.B(n_1554),
.Y(n_1576)
);

AOI221xp5_ASAP7_75t_L g1577 ( 
.A1(n_1568),
.A2(n_1534),
.B1(n_1536),
.B2(n_1537),
.C(n_1503),
.Y(n_1577)
);

INVx3_ASAP7_75t_L g1578 ( 
.A(n_1552),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1551),
.B(n_1532),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1562),
.A2(n_1534),
.B1(n_1503),
.B2(n_1532),
.Y(n_1580)
);

NAND4xp25_ASAP7_75t_L g1581 ( 
.A(n_1554),
.B(n_1533),
.C(n_1505),
.D(n_1537),
.Y(n_1581)
);

AOI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1561),
.A2(n_1503),
.B1(n_1532),
.B2(n_1527),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1562),
.A2(n_1503),
.B1(n_1527),
.B2(n_1543),
.Y(n_1583)
);

OR2x6_ASAP7_75t_L g1584 ( 
.A(n_1559),
.B(n_1535),
.Y(n_1584)
);

AOI31xp33_ASAP7_75t_L g1585 ( 
.A1(n_1561),
.A2(n_1543),
.A3(n_1505),
.B(n_1535),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1549),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1549),
.Y(n_1587)
);

OAI33xp33_ASAP7_75t_L g1588 ( 
.A1(n_1554),
.A2(n_1539),
.A3(n_1501),
.B1(n_1514),
.B2(n_1544),
.B3(n_1513),
.Y(n_1588)
);

NAND2xp33_ASAP7_75t_R g1589 ( 
.A(n_1563),
.B(n_1545),
.Y(n_1589)
);

AOI221xp5_ASAP7_75t_L g1590 ( 
.A1(n_1568),
.A2(n_1527),
.B1(n_1539),
.B2(n_1517),
.C(n_1501),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1553),
.B(n_1540),
.Y(n_1591)
);

BUFx12f_ASAP7_75t_L g1592 ( 
.A(n_1563),
.Y(n_1592)
);

AO21x2_ASAP7_75t_L g1593 ( 
.A1(n_1568),
.A2(n_1498),
.B(n_1526),
.Y(n_1593)
);

OAI33xp33_ASAP7_75t_L g1594 ( 
.A1(n_1553),
.A2(n_1539),
.A3(n_1501),
.B1(n_1514),
.B2(n_1544),
.B3(n_1513),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1565),
.Y(n_1595)
);

OAI221xp5_ASAP7_75t_L g1596 ( 
.A1(n_1561),
.A2(n_1535),
.B1(n_1543),
.B2(n_1555),
.C(n_1527),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1546),
.Y(n_1597)
);

AO21x2_ASAP7_75t_L g1598 ( 
.A1(n_1568),
.A2(n_1498),
.B(n_1526),
.Y(n_1598)
);

AOI221xp5_ASAP7_75t_L g1599 ( 
.A1(n_1555),
.A2(n_1517),
.B1(n_1538),
.B2(n_1499),
.C(n_1516),
.Y(n_1599)
);

BUFx2_ASAP7_75t_L g1600 ( 
.A(n_1569),
.Y(n_1600)
);

BUFx6f_ASAP7_75t_L g1601 ( 
.A(n_1559),
.Y(n_1601)
);

AOI221xp5_ASAP7_75t_L g1602 ( 
.A1(n_1555),
.A2(n_1538),
.B1(n_1499),
.B2(n_1516),
.C(n_1526),
.Y(n_1602)
);

OAI221xp5_ASAP7_75t_L g1603 ( 
.A1(n_1559),
.A2(n_1535),
.B1(n_1543),
.B2(n_1506),
.C(n_1502),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1565),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1570),
.B(n_1508),
.Y(n_1605)
);

INVxp67_ASAP7_75t_SL g1606 ( 
.A(n_1556),
.Y(n_1606)
);

OAI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1557),
.A2(n_1529),
.B1(n_1522),
.B2(n_1542),
.Y(n_1607)
);

INVx4_ASAP7_75t_SL g1608 ( 
.A(n_1601),
.Y(n_1608)
);

BUFx3_ASAP7_75t_L g1609 ( 
.A(n_1601),
.Y(n_1609)
);

OR2x6_ASAP7_75t_L g1610 ( 
.A(n_1584),
.B(n_1529),
.Y(n_1610)
);

BUFx2_ASAP7_75t_L g1611 ( 
.A(n_1584),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1575),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_SL g1613 ( 
.A(n_1577),
.B(n_1563),
.Y(n_1613)
);

OAI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1573),
.A2(n_1502),
.B(n_1506),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1595),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_SL g1616 ( 
.A(n_1585),
.B(n_1563),
.Y(n_1616)
);

AND2x6_ASAP7_75t_SL g1617 ( 
.A(n_1584),
.B(n_1521),
.Y(n_1617)
);

INVxp67_ASAP7_75t_L g1618 ( 
.A(n_1576),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1593),
.B(n_1550),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1586),
.B(n_1558),
.Y(n_1620)
);

HB1xp67_ASAP7_75t_L g1621 ( 
.A(n_1604),
.Y(n_1621)
);

BUFx3_ASAP7_75t_L g1622 ( 
.A(n_1601),
.Y(n_1622)
);

NAND3xp33_ASAP7_75t_L g1623 ( 
.A(n_1574),
.B(n_1602),
.C(n_1599),
.Y(n_1623)
);

BUFx8_ASAP7_75t_L g1624 ( 
.A(n_1601),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_1601),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1575),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1597),
.Y(n_1627)
);

BUFx3_ASAP7_75t_L g1628 ( 
.A(n_1571),
.Y(n_1628)
);

BUFx3_ASAP7_75t_L g1629 ( 
.A(n_1571),
.Y(n_1629)
);

AND4x1_ASAP7_75t_L g1630 ( 
.A(n_1583),
.B(n_1521),
.C(n_1514),
.D(n_1523),
.Y(n_1630)
);

INVxp67_ASAP7_75t_L g1631 ( 
.A(n_1571),
.Y(n_1631)
);

NOR2xp33_ASAP7_75t_L g1632 ( 
.A(n_1581),
.B(n_1544),
.Y(n_1632)
);

INVx2_ASAP7_75t_SL g1633 ( 
.A(n_1572),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1598),
.B(n_1579),
.Y(n_1634)
);

INVx1_ASAP7_75t_SL g1635 ( 
.A(n_1572),
.Y(n_1635)
);

OA21x2_ASAP7_75t_L g1636 ( 
.A1(n_1580),
.A2(n_1528),
.B(n_1548),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1618),
.B(n_1605),
.Y(n_1637)
);

AOI33xp33_ASAP7_75t_L g1638 ( 
.A1(n_1619),
.A2(n_1590),
.A3(n_1582),
.B1(n_1607),
.B2(n_1566),
.B3(n_1551),
.Y(n_1638)
);

INVxp67_ASAP7_75t_L g1639 ( 
.A(n_1632),
.Y(n_1639)
);

OAI21xp5_ASAP7_75t_SL g1640 ( 
.A1(n_1623),
.A2(n_1596),
.B(n_1603),
.Y(n_1640)
);

INVx3_ASAP7_75t_L g1641 ( 
.A(n_1617),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1608),
.B(n_1598),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1626),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1626),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1612),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1616),
.B(n_1579),
.Y(n_1646)
);

AOI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1623),
.A2(n_1594),
.B(n_1588),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1612),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1612),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1616),
.B(n_1598),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1627),
.Y(n_1651)
);

NAND2xp33_ASAP7_75t_SL g1652 ( 
.A(n_1613),
.B(n_1589),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1634),
.B(n_1578),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1632),
.B(n_1591),
.Y(n_1654)
);

BUFx2_ASAP7_75t_L g1655 ( 
.A(n_1617),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1618),
.B(n_1605),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1627),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1613),
.B(n_1587),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1627),
.Y(n_1659)
);

OR2x6_ASAP7_75t_L g1660 ( 
.A(n_1610),
.B(n_1529),
.Y(n_1660)
);

AOI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1614),
.A2(n_1530),
.B(n_1606),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1634),
.B(n_1551),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1634),
.B(n_1611),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1633),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1620),
.B(n_1570),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1614),
.A2(n_1530),
.B1(n_1592),
.B2(n_1560),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1633),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1615),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1634),
.B(n_1551),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1620),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1615),
.B(n_1570),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1611),
.B(n_1600),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1611),
.B(n_1600),
.Y(n_1673)
);

AND2x4_ASAP7_75t_SL g1674 ( 
.A(n_1610),
.B(n_1529),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1609),
.B(n_1547),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1621),
.B(n_1635),
.Y(n_1676)
);

BUFx2_ASAP7_75t_SL g1677 ( 
.A(n_1633),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1609),
.B(n_1547),
.Y(n_1678)
);

AND2x4_ASAP7_75t_L g1679 ( 
.A(n_1608),
.B(n_1609),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1668),
.Y(n_1680)
);

AOI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1652),
.A2(n_1636),
.B1(n_1610),
.B2(n_1530),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1645),
.Y(n_1682)
);

INVxp67_ASAP7_75t_L g1683 ( 
.A(n_1655),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1639),
.B(n_1654),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1647),
.B(n_1621),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1645),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1648),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1648),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1640),
.B(n_1630),
.Y(n_1689)
);

OAI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1655),
.A2(n_1502),
.B1(n_1506),
.B2(n_1636),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1664),
.Y(n_1691)
);

AOI211xp5_ASAP7_75t_L g1692 ( 
.A1(n_1641),
.A2(n_1661),
.B(n_1650),
.C(n_1658),
.Y(n_1692)
);

INVxp67_ASAP7_75t_L g1693 ( 
.A(n_1676),
.Y(n_1693)
);

AND2x4_ASAP7_75t_L g1694 ( 
.A(n_1679),
.B(n_1608),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1649),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1664),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1679),
.B(n_1608),
.Y(n_1697)
);

HB1xp67_ASAP7_75t_L g1698 ( 
.A(n_1676),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1649),
.Y(n_1699)
);

CKINVDCx16_ASAP7_75t_R g1700 ( 
.A(n_1679),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1638),
.B(n_1630),
.Y(n_1701)
);

INVxp67_ASAP7_75t_SL g1702 ( 
.A(n_1667),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1651),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1651),
.Y(n_1704)
);

INVx2_ASAP7_75t_SL g1705 ( 
.A(n_1667),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1672),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1641),
.B(n_1609),
.Y(n_1707)
);

AOI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1641),
.A2(n_1636),
.B1(n_1610),
.B2(n_1530),
.Y(n_1708)
);

AND2x4_ASAP7_75t_SL g1709 ( 
.A(n_1672),
.B(n_1673),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1658),
.B(n_1630),
.Y(n_1710)
);

INVx2_ASAP7_75t_SL g1711 ( 
.A(n_1673),
.Y(n_1711)
);

NOR2xp33_ASAP7_75t_SL g1712 ( 
.A(n_1650),
.B(n_1624),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1657),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1657),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1646),
.B(n_1617),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1698),
.Y(n_1716)
);

BUFx3_ASAP7_75t_L g1717 ( 
.A(n_1707),
.Y(n_1717)
);

INVxp67_ASAP7_75t_L g1718 ( 
.A(n_1698),
.Y(n_1718)
);

INVxp67_ASAP7_75t_L g1719 ( 
.A(n_1715),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1682),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1709),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1683),
.B(n_1646),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1683),
.B(n_1670),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1693),
.B(n_1684),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1709),
.B(n_1677),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1693),
.B(n_1670),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1711),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1700),
.B(n_1677),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1706),
.Y(n_1729)
);

INVx1_ASAP7_75t_SL g1730 ( 
.A(n_1694),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1694),
.B(n_1663),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1680),
.B(n_1675),
.Y(n_1732)
);

OAI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1701),
.A2(n_1666),
.B1(n_1636),
.B2(n_1660),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1689),
.B(n_1637),
.Y(n_1734)
);

AND2x2_ASAP7_75t_SL g1735 ( 
.A(n_1715),
.B(n_1642),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_SL g1736 ( 
.A(n_1692),
.B(n_1642),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1694),
.B(n_1663),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1685),
.B(n_1706),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1686),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1710),
.B(n_1675),
.Y(n_1740)
);

XNOR2xp5_ASAP7_75t_L g1741 ( 
.A(n_1681),
.B(n_1674),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1691),
.B(n_1637),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1722),
.B(n_1738),
.Y(n_1743)
);

A2O1A1Ixp33_ASAP7_75t_L g1744 ( 
.A1(n_1734),
.A2(n_1708),
.B(n_1712),
.C(n_1628),
.Y(n_1744)
);

AOI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1719),
.A2(n_1697),
.B1(n_1690),
.B2(n_1636),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1728),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1716),
.Y(n_1747)
);

OAI21xp33_ASAP7_75t_L g1748 ( 
.A1(n_1740),
.A2(n_1660),
.B(n_1697),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1728),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1716),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1729),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1729),
.Y(n_1752)
);

NOR3xp33_ASAP7_75t_L g1753 ( 
.A(n_1718),
.B(n_1702),
.C(n_1631),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1727),
.B(n_1705),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1729),
.Y(n_1755)
);

OAI21xp33_ASAP7_75t_L g1756 ( 
.A1(n_1717),
.A2(n_1660),
.B(n_1674),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1738),
.B(n_1656),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1731),
.B(n_1678),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1731),
.B(n_1678),
.Y(n_1759)
);

A2O1A1Ixp33_ASAP7_75t_L g1760 ( 
.A1(n_1736),
.A2(n_1629),
.B(n_1628),
.C(n_1642),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1725),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1727),
.B(n_1691),
.Y(n_1762)
);

OAI222xp33_ASAP7_75t_L g1763 ( 
.A1(n_1745),
.A2(n_1733),
.B1(n_1741),
.B2(n_1730),
.C1(n_1724),
.C2(n_1725),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1746),
.B(n_1737),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1746),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1751),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1749),
.B(n_1730),
.Y(n_1767)
);

INVxp67_ASAP7_75t_L g1768 ( 
.A(n_1749),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1747),
.B(n_1724),
.Y(n_1769)
);

OAI222xp33_ASAP7_75t_L g1770 ( 
.A1(n_1757),
.A2(n_1741),
.B1(n_1721),
.B2(n_1660),
.C1(n_1732),
.C2(n_1737),
.Y(n_1770)
);

NAND2x1_ASAP7_75t_L g1771 ( 
.A(n_1761),
.B(n_1721),
.Y(n_1771)
);

AND2x4_ASAP7_75t_SL g1772 ( 
.A(n_1761),
.B(n_1720),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1750),
.B(n_1723),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1770),
.B(n_1743),
.Y(n_1774)
);

OAI311xp33_ASAP7_75t_L g1775 ( 
.A1(n_1767),
.A2(n_1748),
.A3(n_1744),
.B1(n_1756),
.C1(n_1760),
.Y(n_1775)
);

OAI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1763),
.A2(n_1744),
.B(n_1760),
.Y(n_1776)
);

OAI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1771),
.A2(n_1735),
.B1(n_1717),
.B2(n_1754),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1768),
.Y(n_1778)
);

NAND4xp25_ASAP7_75t_L g1779 ( 
.A(n_1764),
.B(n_1717),
.C(n_1762),
.D(n_1753),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_SL g1780 ( 
.A(n_1769),
.B(n_1735),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1765),
.B(n_1758),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1772),
.Y(n_1782)
);

AOI211xp5_ASAP7_75t_L g1783 ( 
.A1(n_1769),
.A2(n_1753),
.B(n_1726),
.C(n_1755),
.Y(n_1783)
);

NOR2x1_ASAP7_75t_L g1784 ( 
.A(n_1782),
.B(n_1752),
.Y(n_1784)
);

AOI221xp5_ASAP7_75t_L g1785 ( 
.A1(n_1776),
.A2(n_1773),
.B1(n_1766),
.B2(n_1720),
.C(n_1739),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1778),
.Y(n_1786)
);

AOI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1774),
.A2(n_1735),
.B1(n_1759),
.B2(n_1773),
.Y(n_1787)
);

XOR2xp5_ASAP7_75t_L g1788 ( 
.A(n_1777),
.B(n_1742),
.Y(n_1788)
);

NAND3xp33_ASAP7_75t_L g1789 ( 
.A(n_1783),
.B(n_1742),
.C(n_1739),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1786),
.B(n_1781),
.Y(n_1790)
);

NOR3x1_ASAP7_75t_L g1791 ( 
.A(n_1789),
.B(n_1779),
.C(n_1780),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1784),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1787),
.B(n_1702),
.Y(n_1793)
);

INVx2_ASAP7_75t_SL g1794 ( 
.A(n_1788),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1785),
.B(n_1696),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1786),
.B(n_1696),
.Y(n_1796)
);

OAI321xp33_ASAP7_75t_L g1797 ( 
.A1(n_1793),
.A2(n_1775),
.A3(n_1631),
.B1(n_1713),
.B2(n_1704),
.C(n_1714),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1792),
.Y(n_1798)
);

NAND4xp25_ASAP7_75t_SL g1799 ( 
.A(n_1790),
.B(n_1703),
.C(n_1699),
.D(n_1695),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1796),
.Y(n_1800)
);

OAI21xp5_ASAP7_75t_SL g1801 ( 
.A1(n_1794),
.A2(n_1688),
.B(n_1687),
.Y(n_1801)
);

INVx1_ASAP7_75t_SL g1802 ( 
.A(n_1800),
.Y(n_1802)
);

AND2x4_ASAP7_75t_L g1803 ( 
.A(n_1798),
.B(n_1791),
.Y(n_1803)
);

NOR3xp33_ASAP7_75t_L g1804 ( 
.A(n_1797),
.B(n_1795),
.C(n_1629),
.Y(n_1804)
);

INVxp67_ASAP7_75t_SL g1805 ( 
.A(n_1803),
.Y(n_1805)
);

OAI322xp33_ASAP7_75t_L g1806 ( 
.A1(n_1805),
.A2(n_1802),
.A3(n_1804),
.B1(n_1801),
.B2(n_1799),
.C1(n_1643),
.C2(n_1644),
.Y(n_1806)
);

AOI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1806),
.A2(n_1643),
.B(n_1644),
.Y(n_1807)
);

OAI22x1_ASAP7_75t_L g1808 ( 
.A1(n_1806),
.A2(n_1633),
.B1(n_1635),
.B2(n_1659),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1807),
.A2(n_1656),
.B1(n_1629),
.B2(n_1628),
.Y(n_1809)
);

OAI22xp5_ASAP7_75t_SL g1810 ( 
.A1(n_1808),
.A2(n_1629),
.B1(n_1628),
.B2(n_1625),
.Y(n_1810)
);

AOI21xp33_ASAP7_75t_L g1811 ( 
.A1(n_1809),
.A2(n_1625),
.B(n_1622),
.Y(n_1811)
);

AOI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1810),
.A2(n_1653),
.B1(n_1622),
.B2(n_1625),
.Y(n_1812)
);

XNOR2xp5_ASAP7_75t_L g1813 ( 
.A(n_1812),
.B(n_1653),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1813),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1814),
.B(n_1811),
.Y(n_1815)
);

AOI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1815),
.A2(n_1622),
.B1(n_1625),
.B2(n_1659),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_SL g1817 ( 
.A1(n_1816),
.A2(n_1622),
.B1(n_1624),
.B2(n_1662),
.Y(n_1817)
);

AOI211xp5_ASAP7_75t_L g1818 ( 
.A1(n_1817),
.A2(n_1665),
.B(n_1671),
.C(n_1669),
.Y(n_1818)
);


endmodule