module fake_jpeg_14001_n_180 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_180);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_2),
.B(n_7),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx4f_ASAP7_75t_SL g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_40),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_29),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_30),
.Y(n_59)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_41),
.Y(n_52)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_44),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_5),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_45),
.B(n_25),
.Y(n_49)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_58),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_18),
.B1(n_21),
.B2(n_23),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_50),
.A2(n_68),
.B1(n_35),
.B2(n_42),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_23),
.B(n_21),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_22),
.Y(n_83)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_56),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_43),
.B(n_31),
.Y(n_58)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_30),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_65),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_17),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_17),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_40),
.A2(n_26),
.B1(n_20),
.B2(n_32),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_38),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_83),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_46),
.C(n_26),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_75),
.B(n_89),
.Y(n_103)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

BUFx24_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_92),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_56),
.A2(n_20),
.B1(n_22),
.B2(n_24),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_48),
.B(n_51),
.Y(n_98)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_53),
.B(n_22),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_53),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_50),
.A2(n_6),
.B(n_14),
.C(n_10),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_90),
.A2(n_71),
.B(n_88),
.C(n_78),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_70),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_95),
.A2(n_108),
.B(n_91),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_54),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_99),
.B(n_100),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_51),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_14),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_101),
.B(n_10),
.Y(n_123)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_71),
.B1(n_88),
.B2(n_85),
.Y(n_120)
);

AO22x1_ASAP7_75t_L g108 ( 
.A1(n_83),
.A2(n_68),
.B1(n_64),
.B2(n_69),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_109),
.C(n_103),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_118),
.C(n_108),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_109),
.A2(n_75),
.B1(n_89),
.B2(n_74),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_121),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_79),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_120),
.A2(n_124),
.B(n_127),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_79),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_93),
.Y(n_122)
);

AOI221xp5_ASAP7_75t_L g132 ( 
.A1(n_122),
.A2(n_105),
.B1(n_95),
.B2(n_102),
.C(n_106),
.Y(n_132)
);

NAND3xp33_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_127),
.C(n_94),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_73),
.B(n_90),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_91),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_125),
.B(n_94),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_94),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_104),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_57),
.B1(n_48),
.B2(n_81),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_129),
.A2(n_111),
.B1(n_120),
.B2(n_102),
.Y(n_137)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_132),
.B(n_136),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

AOI322xp5_ASAP7_75t_L g136 ( 
.A1(n_116),
.A2(n_108),
.A3(n_94),
.B1(n_110),
.B2(n_104),
.C1(n_111),
.C2(n_24),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_122),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_141),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_143),
.Y(n_153)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_115),
.C(n_118),
.Y(n_146)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_130),
.C(n_139),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_131),
.A2(n_117),
.B1(n_98),
.B2(n_119),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

NAND2x1_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_121),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_152),
.A2(n_142),
.B(n_130),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_155),
.A2(n_153),
.B(n_148),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_158),
.C(n_159),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_152),
.C(n_150),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_124),
.Y(n_159)
);

AOI321xp33_ASAP7_75t_L g160 ( 
.A1(n_154),
.A2(n_143),
.A3(n_141),
.B1(n_135),
.B2(n_128),
.C(n_129),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_145),
.Y(n_165)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_162),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_151),
.A2(n_128),
.B1(n_57),
.B2(n_3),
.Y(n_162)
);

OAI21x1_ASAP7_75t_L g163 ( 
.A1(n_158),
.A2(n_153),
.B(n_151),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_166),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_167),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_156),
.A2(n_144),
.B(n_81),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_164),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_169),
.B(n_170),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_168),
.B(n_156),
.Y(n_170)
);

NOR2xp67_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_5),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_172),
.A2(n_80),
.B(n_1),
.Y(n_176)
);

AOI322xp5_ASAP7_75t_L g175 ( 
.A1(n_173),
.A2(n_171),
.A3(n_172),
.B1(n_7),
.B2(n_24),
.C1(n_80),
.C2(n_69),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_176),
.A2(n_0),
.B(n_1),
.Y(n_178)
);

NOR3xp33_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_174),
.C(n_3),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_177),
.Y(n_180)
);


endmodule