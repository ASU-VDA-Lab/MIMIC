module real_aes_18404_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_1404;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_1011;
wire n_286;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1403;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1352;
wire n_1323;
wire n_1280;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_SL g1099 ( .A1(n_0), .A2(n_66), .B1(n_505), .B2(n_507), .Y(n_1099) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_0), .A2(n_226), .B1(n_607), .B2(n_952), .Y(n_1107) );
INVx1_ASAP7_75t_L g718 ( .A(n_1), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_1), .A2(n_97), .B1(n_607), .B2(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g1103 ( .A(n_2), .Y(n_1103) );
OAI211xp5_ASAP7_75t_L g465 ( .A1(n_3), .A2(n_466), .B(n_468), .C(n_478), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_3), .B(n_497), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_4), .A2(n_117), .B1(n_934), .B2(n_936), .Y(n_933) );
AOI22xp33_ASAP7_75t_SL g951 ( .A1(n_4), .A2(n_122), .B1(n_606), .B2(n_952), .Y(n_951) );
INVx1_ASAP7_75t_L g322 ( .A(n_5), .Y(n_322) );
AO22x1_ASAP7_75t_L g395 ( .A1(n_5), .A2(n_137), .B1(n_396), .B2(n_398), .Y(n_395) );
INVx1_ASAP7_75t_L g263 ( .A(n_6), .Y(n_263) );
AND2x2_ASAP7_75t_L g293 ( .A(n_6), .B(n_294), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_6), .B(n_273), .Y(n_389) );
AND2x2_ASAP7_75t_L g407 ( .A(n_6), .B(n_205), .Y(n_407) );
INVx1_ASAP7_75t_L g343 ( .A(n_7), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_7), .A2(n_94), .B1(n_391), .B2(n_393), .Y(n_390) );
INVx1_ASAP7_75t_L g987 ( .A(n_8), .Y(n_987) );
AOI221xp5_ASAP7_75t_L g1096 ( .A1(n_9), .A2(n_140), .B1(n_1093), .B2(n_1097), .C(n_1098), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_9), .A2(n_59), .B1(n_607), .B2(n_1111), .Y(n_1110) );
AOI22xp33_ASAP7_75t_SL g931 ( .A1(n_10), .A2(n_150), .B1(n_364), .B2(n_932), .Y(n_931) );
AOI221xp5_ASAP7_75t_L g948 ( .A1(n_10), .A2(n_16), .B1(n_597), .B2(n_603), .C(n_949), .Y(n_948) );
INVx1_ASAP7_75t_L g1323 ( .A(n_11), .Y(n_1323) );
AOI22xp5_ASAP7_75t_L g1347 ( .A1(n_11), .A2(n_35), .B1(n_900), .B2(n_1348), .Y(n_1347) );
AOI22xp33_ASAP7_75t_SL g559 ( .A1(n_12), .A2(n_127), .B1(n_502), .B2(n_560), .Y(n_559) );
INVxp67_ASAP7_75t_SL g627 ( .A(n_12), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_13), .A2(n_142), .B1(n_736), .B2(n_768), .Y(n_767) );
AOI22xp33_ASAP7_75t_SL g801 ( .A1(n_13), .A2(n_230), .B1(n_502), .B2(n_692), .Y(n_801) );
CKINVDCx5p33_ASAP7_75t_R g1090 ( .A(n_14), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_15), .B(n_1129), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1131 ( .A(n_15), .B(n_98), .Y(n_1131) );
INVx2_ASAP7_75t_L g1135 ( .A(n_15), .Y(n_1135) );
AOI22xp33_ASAP7_75t_SL g940 ( .A1(n_16), .A2(n_34), .B1(n_574), .B2(n_822), .Y(n_940) );
CKINVDCx5p33_ASAP7_75t_R g1388 ( .A(n_17), .Y(n_1388) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_18), .A2(n_216), .B1(n_560), .B2(n_572), .Y(n_571) );
AOI221xp5_ASAP7_75t_L g596 ( .A1(n_18), .A2(n_127), .B1(n_597), .B2(n_599), .C(n_602), .Y(n_596) );
INVx1_ASAP7_75t_L g929 ( .A(n_19), .Y(n_929) );
OAI22xp33_ASAP7_75t_L g941 ( .A1(n_20), .A2(n_196), .B1(n_576), .B2(n_580), .Y(n_941) );
INVx1_ASAP7_75t_L g955 ( .A(n_20), .Y(n_955) );
INVx1_ASAP7_75t_L g1392 ( .A(n_21), .Y(n_1392) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_22), .A2(n_211), .B1(n_440), .B2(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g740 ( .A(n_23), .Y(n_740) );
AOI22xp33_ASAP7_75t_SL g719 ( .A1(n_24), .A2(n_67), .B1(n_502), .B2(n_503), .Y(n_719) );
AOI221xp5_ASAP7_75t_L g733 ( .A1(n_24), .A2(n_245), .B1(n_598), .B2(n_603), .C(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g762 ( .A(n_25), .Y(n_762) );
OAI22xp5_ASAP7_75t_L g786 ( .A1(n_25), .A2(n_215), .B1(n_440), .B2(n_589), .Y(n_786) );
INVx1_ASAP7_75t_L g655 ( .A(n_26), .Y(n_655) );
OAI22xp33_ASAP7_75t_L g680 ( .A1(n_26), .A2(n_158), .B1(n_576), .B2(n_681), .Y(n_680) );
OAI221xp5_ASAP7_75t_L g665 ( .A1(n_27), .A2(n_53), .B1(n_617), .B2(n_666), .C(n_668), .Y(n_665) );
INVx1_ASAP7_75t_L g694 ( .A(n_27), .Y(n_694) );
OAI211xp5_ASAP7_75t_L g479 ( .A1(n_28), .A2(n_480), .B(n_482), .C(n_484), .Y(n_479) );
INVx1_ASAP7_75t_L g540 ( .A(n_28), .Y(n_540) );
INVx1_ASAP7_75t_L g739 ( .A(n_29), .Y(n_739) );
XOR2x2_ASAP7_75t_L g975 ( .A(n_30), .B(n_976), .Y(n_975) );
AOI22xp5_ASAP7_75t_L g1169 ( .A1(n_30), .A2(n_159), .B1(n_1130), .B2(n_1136), .Y(n_1169) );
CKINVDCx5p33_ASAP7_75t_R g809 ( .A(n_31), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g1191 ( .A1(n_32), .A2(n_185), .B1(n_1126), .B2(n_1133), .Y(n_1191) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_33), .A2(n_245), .B1(n_502), .B2(n_503), .Y(n_727) );
AOI22xp33_ASAP7_75t_SL g745 ( .A1(n_33), .A2(n_67), .B1(n_605), .B2(n_664), .Y(n_745) );
A2O1A1Ixp33_ASAP7_75t_L g958 ( .A1(n_34), .A2(n_959), .B(n_960), .C(n_969), .Y(n_958) );
INVx1_ASAP7_75t_L g1335 ( .A(n_35), .Y(n_1335) );
INVx1_ASAP7_75t_L g1329 ( .A(n_36), .Y(n_1329) );
AOI22xp33_ASAP7_75t_L g1352 ( .A1(n_36), .A2(n_163), .B1(n_778), .B2(n_1348), .Y(n_1352) );
INVx1_ASAP7_75t_L g1000 ( .A(n_37), .Y(n_1000) );
OAI22xp5_ASAP7_75t_L g944 ( .A1(n_38), .A2(n_55), .B1(n_497), .B2(n_589), .Y(n_944) );
OAI211xp5_ASAP7_75t_L g946 ( .A1(n_38), .A2(n_651), .B(n_947), .C(n_953), .Y(n_946) );
AOI22xp5_ASAP7_75t_L g1143 ( .A1(n_39), .A2(n_108), .B1(n_1126), .B2(n_1133), .Y(n_1143) );
AOI22xp5_ASAP7_75t_L g1158 ( .A1(n_40), .A2(n_194), .B1(n_1126), .B2(n_1136), .Y(n_1158) );
INVx1_ASAP7_75t_L g1355 ( .A(n_40), .Y(n_1355) );
AOI22xp33_ASAP7_75t_L g1362 ( .A1(n_40), .A2(n_1363), .B1(n_1365), .B2(n_1411), .Y(n_1362) );
AOI22xp5_ASAP7_75t_L g1168 ( .A1(n_41), .A2(n_89), .B1(n_1126), .B2(n_1133), .Y(n_1168) );
XOR2x2_ASAP7_75t_L g548 ( .A(n_42), .B(n_549), .Y(n_548) );
XNOR2x2_ASAP7_75t_L g922 ( .A(n_43), .B(n_923), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_44), .A2(n_63), .B1(n_432), .B2(n_470), .Y(n_469) );
AOI22xp33_ASAP7_75t_SL g501 ( .A1(n_44), .A2(n_242), .B1(n_502), .B2(n_503), .Y(n_501) );
INVx1_ASAP7_75t_L g835 ( .A(n_45), .Y(n_835) );
INVx1_ASAP7_75t_L g314 ( .A(n_46), .Y(n_314) );
INVx1_ASAP7_75t_L g327 ( .A(n_46), .Y(n_327) );
INVxp67_ASAP7_75t_SL g644 ( .A(n_47), .Y(n_644) );
AND4x1_ASAP7_75t_L g697 ( .A(n_47), .B(n_646), .C(n_649), .D(n_678), .Y(n_697) );
INVx1_ASAP7_75t_L g703 ( .A(n_48), .Y(n_703) );
OAI22xp33_ASAP7_75t_L g575 ( .A1(n_49), .A2(n_162), .B1(n_576), .B2(n_580), .Y(n_575) );
INVx1_ASAP7_75t_L g610 ( .A(n_49), .Y(n_610) );
OAI221xp5_ASAP7_75t_L g1312 ( .A1(n_50), .A2(n_101), .B1(n_306), .B2(n_869), .C(n_1313), .Y(n_1312) );
INVxp67_ASAP7_75t_SL g1342 ( .A(n_50), .Y(n_1342) );
INVxp67_ASAP7_75t_SL g776 ( .A(n_51), .Y(n_776) );
AOI22xp33_ASAP7_75t_SL g798 ( .A1(n_51), .A2(n_126), .B1(n_565), .B2(n_799), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_52), .A2(n_122), .B1(n_936), .B2(n_938), .Y(n_937) );
AOI221xp5_ASAP7_75t_L g961 ( .A1(n_52), .A2(n_117), .B1(n_962), .B2(n_965), .C(n_966), .Y(n_961) );
INVx1_ASAP7_75t_L g696 ( .A(n_53), .Y(n_696) );
INVx1_ASAP7_75t_L g256 ( .A(n_54), .Y(n_256) );
INVx2_ASAP7_75t_L g310 ( .A(n_56), .Y(n_310) );
INVx1_ASAP7_75t_L g449 ( .A(n_57), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g1159 ( .A1(n_58), .A2(n_75), .B1(n_1133), .B2(n_1146), .Y(n_1159) );
AOI221xp5_ASAP7_75t_L g1092 ( .A1(n_59), .A2(n_65), .B1(n_822), .B2(n_1093), .C(n_1094), .Y(n_1092) );
NOR2xp33_ASAP7_75t_L g779 ( .A(n_60), .B(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g791 ( .A(n_60), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_61), .A2(n_76), .B1(n_825), .B2(n_827), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_61), .A2(n_209), .B1(n_446), .B2(n_736), .Y(n_841) );
INVx1_ASAP7_75t_L g1086 ( .A(n_62), .Y(n_1086) );
AOI22xp33_ASAP7_75t_SL g510 ( .A1(n_63), .A2(n_93), .B1(n_367), .B2(n_502), .Y(n_510) );
INVx1_ASAP7_75t_L g1085 ( .A(n_64), .Y(n_1085) );
AOI221xp5_ASAP7_75t_L g1106 ( .A1(n_65), .A2(n_140), .B1(n_477), .B2(n_598), .C(n_600), .Y(n_1106) );
AOI221xp5_ASAP7_75t_L g1112 ( .A1(n_66), .A2(n_71), .B1(n_600), .B2(n_638), .C(n_900), .Y(n_1112) );
AOI22xp33_ASAP7_75t_SL g1378 ( .A1(n_68), .A2(n_170), .B1(n_560), .B2(n_1379), .Y(n_1378) );
AOI22xp33_ASAP7_75t_SL g1408 ( .A1(n_68), .A2(n_213), .B1(n_664), .B2(n_952), .Y(n_1408) );
AOI22xp5_ASAP7_75t_L g1154 ( .A1(n_69), .A2(n_121), .B1(n_1126), .B2(n_1133), .Y(n_1154) );
INVx1_ASAP7_75t_L g891 ( .A(n_70), .Y(n_891) );
AOI221xp5_ASAP7_75t_L g906 ( .A1(n_70), .A2(n_123), .B1(n_734), .B2(n_900), .C(n_907), .Y(n_906) );
AOI22xp33_ASAP7_75t_SL g1095 ( .A1(n_71), .A2(n_226), .B1(n_505), .B2(n_507), .Y(n_1095) );
INVx1_ASAP7_75t_L g1333 ( .A(n_72), .Y(n_1333) );
AOI22xp33_ASAP7_75t_L g1349 ( .A1(n_72), .A2(n_208), .B1(n_446), .B2(n_470), .Y(n_1349) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_73), .A2(n_193), .B1(n_440), .B2(n_589), .Y(n_648) );
OAI211xp5_ASAP7_75t_L g650 ( .A1(n_73), .A2(n_651), .B(n_652), .C(n_656), .Y(n_650) );
OAI222xp33_ASAP7_75t_L g362 ( .A1(n_74), .A2(n_190), .B1(n_363), .B2(n_371), .C1(n_373), .C2(n_377), .Y(n_362) );
INVx1_ASAP7_75t_L g408 ( .A(n_74), .Y(n_408) );
AOI21xp33_ASAP7_75t_L g850 ( .A1(n_76), .A2(n_472), .B(n_476), .Y(n_850) );
OAI211xp5_ASAP7_75t_L g1027 ( .A1(n_77), .A2(n_1011), .B(n_1028), .C(n_1030), .Y(n_1027) );
INVx1_ASAP7_75t_L g1073 ( .A(n_77), .Y(n_1073) );
INVx1_ASAP7_75t_L g556 ( .A(n_78), .Y(n_556) );
OAI221xp5_ASAP7_75t_L g616 ( .A1(n_78), .A2(n_87), .B1(n_617), .B2(n_621), .C(n_624), .Y(n_616) );
OAI22xp33_ASAP7_75t_L g836 ( .A1(n_79), .A2(n_83), .B1(n_580), .B2(n_803), .Y(n_836) );
INVx1_ASAP7_75t_L g843 ( .A(n_79), .Y(n_843) );
AOI22xp33_ASAP7_75t_SL g831 ( .A1(n_80), .A2(n_235), .B1(n_819), .B2(n_822), .Y(n_831) );
AOI22xp33_ASAP7_75t_SL g851 ( .A1(n_80), .A2(n_161), .B1(n_852), .B2(n_853), .Y(n_851) );
CKINVDCx5p33_ASAP7_75t_R g1319 ( .A(n_81), .Y(n_1319) );
AOI22xp5_ASAP7_75t_L g1163 ( .A1(n_82), .A2(n_120), .B1(n_1126), .B2(n_1133), .Y(n_1163) );
INVx1_ASAP7_75t_L g844 ( .A(n_83), .Y(n_844) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_84), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_85), .A2(n_238), .B1(n_396), .B2(n_664), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_85), .A2(n_110), .B1(n_565), .B2(n_686), .Y(n_688) );
AOI22xp5_ASAP7_75t_SL g1162 ( .A1(n_86), .A2(n_232), .B1(n_1136), .B2(n_1146), .Y(n_1162) );
INVx1_ASAP7_75t_L g553 ( .A(n_87), .Y(n_553) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_88), .Y(n_258) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_88), .B(n_256), .Y(n_1127) );
AOI22xp33_ASAP7_75t_SL g1381 ( .A1(n_90), .A2(n_248), .B1(n_799), .B2(n_1382), .Y(n_1381) );
AOI21xp33_ASAP7_75t_L g1405 ( .A1(n_90), .A2(n_638), .B(n_1406), .Y(n_1405) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_91), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g1089 ( .A(n_92), .Y(n_1089) );
AOI221xp5_ASAP7_75t_SL g475 ( .A1(n_93), .A2(n_242), .B1(n_393), .B2(n_476), .C(n_477), .Y(n_475) );
INVx1_ASAP7_75t_L g337 ( .A(n_94), .Y(n_337) );
OAI22xp5_ASAP7_75t_L g1393 ( .A1(n_95), .A2(n_236), .B1(n_580), .B2(n_803), .Y(n_1393) );
INVx1_ASAP7_75t_L g1400 ( .A(n_95), .Y(n_1400) );
CKINVDCx5p33_ASAP7_75t_R g724 ( .A(n_96), .Y(n_724) );
INVx1_ASAP7_75t_L g726 ( .A(n_97), .Y(n_726) );
INVx1_ASAP7_75t_L g1129 ( .A(n_98), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_98), .B(n_1135), .Y(n_1137) );
AOI22xp33_ASAP7_75t_SL g1142 ( .A1(n_99), .A2(n_109), .B1(n_1130), .B2(n_1136), .Y(n_1142) );
INVxp67_ASAP7_75t_SL g674 ( .A(n_100), .Y(n_674) );
AOI22xp33_ASAP7_75t_SL g690 ( .A1(n_100), .A2(n_195), .B1(n_691), .B2(n_692), .Y(n_690) );
INVx1_ASAP7_75t_L g1354 ( .A(n_101), .Y(n_1354) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_102), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_103), .A2(n_243), .B1(n_1126), .B2(n_1130), .Y(n_1125) );
CKINVDCx5p33_ASAP7_75t_R g647 ( .A(n_104), .Y(n_647) );
INVx1_ASAP7_75t_L g1036 ( .A(n_105), .Y(n_1036) );
OAI211xp5_ASAP7_75t_L g1066 ( .A1(n_105), .A2(n_984), .B(n_1067), .C(n_1070), .Y(n_1066) );
INVxp67_ASAP7_75t_SL g773 ( .A(n_106), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_106), .A2(n_228), .B1(n_795), .B2(n_796), .Y(n_794) );
OAI211xp5_ASAP7_75t_SL g763 ( .A1(n_107), .A2(n_621), .B(n_764), .C(n_771), .Y(n_763) );
INVx1_ASAP7_75t_L g790 ( .A(n_107), .Y(n_790) );
AOI221xp5_ASAP7_75t_L g675 ( .A1(n_110), .A2(n_203), .B1(n_391), .B2(n_638), .C(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g713 ( .A(n_111), .Y(n_713) );
AOI21xp33_ASAP7_75t_L g744 ( .A1(n_111), .A2(n_638), .B(n_734), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_112), .B(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g340 ( .A(n_112), .Y(n_340) );
INVx1_ASAP7_75t_L g356 ( .A(n_112), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_113), .A2(n_144), .B1(n_352), .B2(n_457), .Y(n_894) );
INVx1_ASAP7_75t_L g908 ( .A(n_113), .Y(n_908) );
AOI22xp5_ASAP7_75t_L g1147 ( .A1(n_114), .A2(n_212), .B1(n_1126), .B2(n_1133), .Y(n_1147) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_115), .A2(n_134), .B1(n_480), .B2(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g519 ( .A(n_115), .Y(n_519) );
INVx1_ASAP7_75t_L g350 ( .A(n_116), .Y(n_350) );
NAND2xp33_ASAP7_75t_SL g433 ( .A(n_116), .B(n_393), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_118), .A2(n_207), .B1(n_440), .B2(n_705), .Y(n_704) );
OAI211xp5_ASAP7_75t_L g731 ( .A1(n_118), .A2(n_593), .B(n_732), .C(n_738), .Y(n_731) );
INVx1_ASAP7_75t_L g761 ( .A(n_119), .Y(n_761) );
OAI22xp33_ASAP7_75t_L g802 ( .A1(n_119), .A2(n_241), .B1(n_681), .B2(n_803), .Y(n_802) );
AOI221xp5_ASAP7_75t_L g881 ( .A1(n_123), .A2(n_221), .B1(n_369), .B2(n_882), .C(n_883), .Y(n_881) );
XNOR2xp5_ASAP7_75t_L g860 ( .A(n_124), .B(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g1336 ( .A(n_125), .Y(n_1336) );
AOI22xp33_ASAP7_75t_L g1353 ( .A1(n_125), .A2(n_175), .B1(n_605), .B2(n_607), .Y(n_1353) );
INVxp67_ASAP7_75t_SL g765 ( .A(n_126), .Y(n_765) );
INVx1_ASAP7_75t_L g980 ( .A(n_128), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_129), .A2(n_209), .B1(n_827), .B2(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g847 ( .A(n_129), .Y(n_847) );
INVx1_ASAP7_75t_L g999 ( .A(n_130), .Y(n_999) );
OAI22xp5_ASAP7_75t_L g1366 ( .A1(n_131), .A2(n_1367), .B1(n_1409), .B2(n_1410), .Y(n_1366) );
CKINVDCx5p33_ASAP7_75t_R g1409 ( .A(n_131), .Y(n_1409) );
INVxp67_ASAP7_75t_SL g1376 ( .A(n_132), .Y(n_1376) );
OAI211xp5_ASAP7_75t_L g1395 ( .A1(n_132), .A2(n_593), .B(n_1396), .C(n_1399), .Y(n_1395) );
AOI22xp33_ASAP7_75t_SL g1383 ( .A1(n_133), .A2(n_227), .B1(n_799), .B2(n_1382), .Y(n_1383) );
AOI22xp33_ASAP7_75t_L g1398 ( .A1(n_133), .A2(n_248), .B1(n_607), .B2(n_852), .Y(n_1398) );
INVx1_ASAP7_75t_L g536 ( .A(n_134), .Y(n_536) );
CKINVDCx16_ASAP7_75t_R g366 ( .A(n_135), .Y(n_366) );
OAI22xp33_ASAP7_75t_L g868 ( .A1(n_136), .A2(n_240), .B1(n_306), .B2(n_869), .Y(n_868) );
INVxp33_ASAP7_75t_SL g920 ( .A(n_136), .Y(n_920) );
AOI21xp5_ASAP7_75t_L g351 ( .A1(n_137), .A2(n_352), .B(n_355), .Y(n_351) );
NAND5xp2_ASAP7_75t_L g463 ( .A(n_138), .B(n_464), .C(n_498), .D(n_522), .E(n_531), .Y(n_463) );
INVx1_ASAP7_75t_L g544 ( .A(n_138), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g1152 ( .A1(n_138), .A2(n_224), .B1(n_1136), .B2(n_1153), .Y(n_1152) );
INVx1_ASAP7_75t_L g438 ( .A(n_139), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_141), .A2(n_237), .B1(n_562), .B2(n_565), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_141), .A2(n_176), .B1(n_605), .B2(n_606), .Y(n_604) );
AOI22xp33_ASAP7_75t_SL g793 ( .A1(n_142), .A2(n_165), .B1(n_502), .B2(n_684), .Y(n_793) );
BUFx3_ASAP7_75t_L g316 ( .A(n_143), .Y(n_316) );
INVx1_ASAP7_75t_L g902 ( .A(n_144), .Y(n_902) );
INVx1_ASAP7_75t_L g1373 ( .A(n_145), .Y(n_1373) );
OAI221xp5_ASAP7_75t_L g1402 ( .A1(n_145), .A2(n_146), .B1(n_667), .B2(n_780), .C(n_1403), .Y(n_1402) );
INVx1_ASAP7_75t_L g1374 ( .A(n_146), .Y(n_1374) );
CKINVDCx5p33_ASAP7_75t_R g874 ( .A(n_147), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g1384 ( .A1(n_148), .A2(n_213), .B1(n_560), .B2(n_1385), .Y(n_1384) );
AOI221xp5_ASAP7_75t_L g1397 ( .A1(n_148), .A2(n_170), .B1(n_598), .B2(n_603), .C(n_734), .Y(n_1397) );
INVx1_ASAP7_75t_L g878 ( .A(n_149), .Y(n_878) );
AOI221xp5_ASAP7_75t_L g899 ( .A1(n_149), .A2(n_184), .B1(n_734), .B2(n_900), .C(n_901), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g967 ( .A(n_150), .B(n_968), .Y(n_967) );
INVxp67_ASAP7_75t_L g807 ( .A(n_151), .Y(n_807) );
AOI22xp33_ASAP7_75t_SL g818 ( .A1(n_152), .A2(n_161), .B1(n_819), .B2(n_820), .Y(n_818) );
AOI221xp5_ASAP7_75t_L g840 ( .A1(n_152), .A2(n_235), .B1(n_391), .B2(n_603), .C(n_778), .Y(n_840) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_153), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_154), .A2(n_189), .B1(n_396), .B2(n_432), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_154), .A2(n_181), .B1(n_507), .B2(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g863 ( .A(n_155), .Y(n_863) );
INVx1_ASAP7_75t_L g1104 ( .A(n_156), .Y(n_1104) );
CKINVDCx5p33_ASAP7_75t_R g875 ( .A(n_157), .Y(n_875) );
INVx1_ASAP7_75t_L g653 ( .A(n_158), .Y(n_653) );
OAI21xp5_ASAP7_75t_SL g1114 ( .A1(n_160), .A2(n_705), .B(n_1115), .Y(n_1114) );
INVx1_ASAP7_75t_L g613 ( .A(n_162), .Y(n_613) );
INVx1_ASAP7_75t_L g1322 ( .A(n_163), .Y(n_1322) );
INVx1_ASAP7_75t_L g888 ( .A(n_164), .Y(n_888) );
AOI221xp5_ASAP7_75t_L g777 ( .A1(n_165), .A2(n_230), .B1(n_603), .B2(n_660), .C(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g812 ( .A(n_166), .Y(n_812) );
OAI221xp5_ASAP7_75t_SL g845 ( .A1(n_166), .A2(n_233), .B1(n_617), .B2(n_666), .C(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g298 ( .A(n_167), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_167), .B(n_306), .Y(n_305) );
XOR2x2_ASAP7_75t_L g754 ( .A(n_168), .B(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g993 ( .A(n_169), .Y(n_993) );
OAI22xp33_ASAP7_75t_L g1040 ( .A1(n_171), .A2(n_192), .B1(n_1041), .B2(n_1044), .Y(n_1040) );
OAI22xp33_ASAP7_75t_L g1052 ( .A1(n_171), .A2(n_192), .B1(n_1053), .B2(n_1054), .Y(n_1052) );
INVx1_ASAP7_75t_L g982 ( .A(n_172), .Y(n_982) );
AOI22xp5_ASAP7_75t_L g1145 ( .A1(n_173), .A2(n_246), .B1(n_1136), .B2(n_1146), .Y(n_1145) );
AOI22xp33_ASAP7_75t_L g1190 ( .A1(n_174), .A2(n_178), .B1(n_1130), .B2(n_1136), .Y(n_1190) );
INVx1_ASAP7_75t_L g1327 ( .A(n_175), .Y(n_1327) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_176), .A2(n_244), .B1(n_562), .B2(n_565), .Y(n_561) );
INVx1_ASAP7_75t_L g530 ( .A(n_177), .Y(n_530) );
INVxp67_ASAP7_75t_SL g672 ( .A(n_179), .Y(n_672) );
AOI22xp33_ASAP7_75t_SL g683 ( .A1(n_179), .A2(n_202), .B1(n_574), .B2(n_684), .Y(n_683) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_180), .Y(n_269) );
AOI221xp5_ASAP7_75t_L g471 ( .A1(n_181), .A2(n_219), .B1(n_391), .B2(n_393), .C(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g1031 ( .A(n_182), .Y(n_1031) );
INVx1_ASAP7_75t_L g1315 ( .A(n_183), .Y(n_1315) );
OAI22xp5_ASAP7_75t_L g1345 ( .A1(n_183), .A2(n_186), .B1(n_410), .B2(n_590), .Y(n_1345) );
AOI21xp33_ASAP7_75t_L g892 ( .A1(n_184), .A2(n_336), .B(n_893), .Y(n_892) );
INVx1_ASAP7_75t_L g1318 ( .A(n_186), .Y(n_1318) );
INVx1_ASAP7_75t_L g785 ( .A(n_187), .Y(n_785) );
CKINVDCx5p33_ASAP7_75t_R g943 ( .A(n_188), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_189), .A2(n_219), .B1(n_505), .B2(n_507), .Y(n_504) );
NOR2xp33_ASAP7_75t_R g416 ( .A(n_190), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g988 ( .A(n_191), .Y(n_988) );
AOI221xp5_ASAP7_75t_L g657 ( .A1(n_195), .A2(n_202), .B1(n_658), .B2(n_660), .C(n_662), .Y(n_657) );
INVx1_ASAP7_75t_L g954 ( .A(n_196), .Y(n_954) );
INVx1_ASAP7_75t_L g994 ( .A(n_197), .Y(n_994) );
OAI22xp5_ASAP7_75t_L g1019 ( .A1(n_198), .A2(n_206), .B1(n_1020), .B2(n_1024), .Y(n_1019) );
OAI22xp5_ASAP7_75t_L g1057 ( .A1(n_198), .A2(n_206), .B1(n_1058), .B2(n_1060), .Y(n_1057) );
INVx1_ASAP7_75t_L g282 ( .A(n_199), .Y(n_282) );
INVx1_ASAP7_75t_L g927 ( .A(n_200), .Y(n_927) );
OAI211xp5_ASAP7_75t_L g1316 ( .A1(n_201), .A2(n_358), .B(n_441), .C(n_1317), .Y(n_1316) );
INVxp33_ASAP7_75t_SL g1344 ( .A(n_201), .Y(n_1344) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_203), .A2(n_238), .B1(n_565), .B2(n_686), .Y(n_685) );
OAI211xp5_ASAP7_75t_SL g870 ( .A1(n_204), .A2(n_358), .B(n_871), .C(n_873), .Y(n_870) );
INVx1_ASAP7_75t_L g913 ( .A(n_204), .Y(n_913) );
BUFx3_ASAP7_75t_L g273 ( .A(n_205), .Y(n_273) );
INVx1_ASAP7_75t_L g294 ( .A(n_205), .Y(n_294) );
INVx1_ASAP7_75t_L g1325 ( .A(n_208), .Y(n_1325) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_210), .Y(n_486) );
OAI211xp5_ASAP7_75t_L g592 ( .A1(n_211), .A2(n_593), .B(n_595), .C(n_609), .Y(n_592) );
INVx1_ASAP7_75t_L g291 ( .A(n_214), .Y(n_291) );
INVx2_ASAP7_75t_L g382 ( .A(n_214), .Y(n_382) );
INVx1_ASAP7_75t_L g421 ( .A(n_214), .Y(n_421) );
INVxp67_ASAP7_75t_SL g633 ( .A(n_216), .Y(n_633) );
CKINVDCx5p33_ASAP7_75t_R g587 ( .A(n_217), .Y(n_587) );
XNOR2x1_ASAP7_75t_L g1081 ( .A(n_218), .B(n_1082), .Y(n_1081) );
INVx1_ASAP7_75t_L g328 ( .A(n_220), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_220), .A2(n_247), .B1(n_396), .B2(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g903 ( .A(n_221), .Y(n_903) );
INVxp67_ASAP7_75t_SL g815 ( .A(n_222), .Y(n_815) );
OAI211xp5_ASAP7_75t_SL g838 ( .A1(n_222), .A2(n_651), .B(n_839), .C(n_842), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g1132 ( .A1(n_223), .A2(n_225), .B1(n_1133), .B2(n_1136), .Y(n_1132) );
INVx1_ASAP7_75t_L g1404 ( .A(n_227), .Y(n_1404) );
AOI21xp5_ASAP7_75t_L g769 ( .A1(n_228), .A2(n_472), .B(n_770), .Y(n_769) );
OAI22xp33_ASAP7_75t_SL g728 ( .A1(n_229), .A2(n_239), .B1(n_555), .B2(n_729), .Y(n_728) );
OAI221xp5_ASAP7_75t_L g741 ( .A1(n_229), .A2(n_239), .B1(n_617), .B2(n_667), .C(n_742), .Y(n_741) );
OAI21xp33_ASAP7_75t_SL g1309 ( .A1(n_231), .A2(n_1310), .B(n_1311), .Y(n_1309) );
INVx1_ASAP7_75t_L g1314 ( .A(n_231), .Y(n_1314) );
XNOR2xp5_ASAP7_75t_L g700 ( .A(n_232), .B(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g813 ( .A(n_233), .Y(n_813) );
CKINVDCx5p33_ASAP7_75t_R g880 ( .A(n_234), .Y(n_880) );
INVx1_ASAP7_75t_L g1401 ( .A(n_236), .Y(n_1401) );
AOI221xp5_ASAP7_75t_L g634 ( .A1(n_237), .A2(n_244), .B1(n_635), .B2(n_636), .C(n_638), .Y(n_634) );
INVxp67_ASAP7_75t_SL g866 ( .A(n_240), .Y(n_866) );
INVx1_ASAP7_75t_L g759 ( .A(n_241), .Y(n_759) );
INVx1_ASAP7_75t_L g345 ( .A(n_247), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_274), .B(n_1119), .Y(n_249) );
BUFx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx3_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_259), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g1361 ( .A(n_253), .B(n_262), .Y(n_1361) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_255), .B(n_257), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g1364 ( .A(n_255), .B(n_258), .Y(n_1364) );
INVx1_ASAP7_75t_L g1415 ( .A(n_255), .Y(n_1415) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g1417 ( .A(n_258), .B(n_1415), .Y(n_1417) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_264), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x4_ASAP7_75t_L g1078 ( .A(n_262), .B(n_1079), .Y(n_1078) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x4_ASAP7_75t_L g425 ( .A(n_263), .B(n_273), .Y(n_425) );
AND2x4_ASAP7_75t_L g473 ( .A(n_263), .B(n_272), .Y(n_473) );
INVx1_ASAP7_75t_L g1053 ( .A(n_264), .Y(n_1053) );
AND2x4_ASAP7_75t_SL g1360 ( .A(n_264), .B(n_1361), .Y(n_1360) );
INVx3_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OR2x6_ASAP7_75t_L g265 ( .A(n_266), .B(n_271), .Y(n_265) );
INVxp67_ASAP7_75t_L g968 ( .A(n_266), .Y(n_968) );
OR2x6_ASAP7_75t_L g1059 ( .A(n_266), .B(n_1056), .Y(n_1059) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
BUFx4f_ASAP7_75t_L g481 ( .A(n_267), .Y(n_481) );
INVx3_ASAP7_75t_L g671 ( .A(n_267), .Y(n_671) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx2_ASAP7_75t_L g296 ( .A(n_269), .Y(n_296) );
AND2x2_ASAP7_75t_L g302 ( .A(n_269), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g394 ( .A(n_269), .B(n_270), .Y(n_394) );
INVx2_ASAP7_75t_L g400 ( .A(n_269), .Y(n_400) );
INVx1_ASAP7_75t_L g406 ( .A(n_269), .Y(n_406) );
NAND2x1_ASAP7_75t_L g419 ( .A(n_269), .B(n_270), .Y(n_419) );
INVx1_ASAP7_75t_L g297 ( .A(n_270), .Y(n_297) );
INVx2_ASAP7_75t_L g303 ( .A(n_270), .Y(n_303) );
AND2x2_ASAP7_75t_L g399 ( .A(n_270), .B(n_400), .Y(n_399) );
BUFx2_ASAP7_75t_L g415 ( .A(n_270), .Y(n_415) );
OR2x2_ASAP7_75t_L g430 ( .A(n_270), .B(n_296), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_270), .B(n_400), .Y(n_632) );
INVxp67_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g1069 ( .A(n_272), .Y(n_1069) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
BUFx2_ASAP7_75t_L g1065 ( .A(n_273), .Y(n_1065) );
AND2x4_ASAP7_75t_L g1076 ( .A(n_273), .B(n_405), .Y(n_1076) );
OAI22xp33_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_276), .B1(n_752), .B2(n_1118), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
XNOR2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_640), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
XNOR2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_458), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
XNOR2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
NOR2x1_ASAP7_75t_L g283 ( .A(n_284), .B(n_383), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_304), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_287), .B1(n_298), .B2(n_299), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_286), .A2(n_364), .B1(n_366), .B2(n_367), .Y(n_363) );
HB1xp67_ASAP7_75t_L g862 ( .A(n_287), .Y(n_862) );
INVx3_ASAP7_75t_L g1310 ( .A(n_287), .Y(n_1310) );
AND2x4_ASAP7_75t_L g287 ( .A(n_288), .B(n_292), .Y(n_287) );
AND2x4_ASAP7_75t_L g299 ( .A(n_288), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g403 ( .A(n_289), .B(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g442 ( .A(n_289), .Y(n_442) );
OR2x2_ASAP7_75t_L g590 ( .A(n_289), .B(n_404), .Y(n_590) );
INVx1_ASAP7_75t_L g1079 ( .A(n_289), .Y(n_1079) );
BUFx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g426 ( .A(n_290), .Y(n_426) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g612 ( .A(n_292), .Y(n_612) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_292), .Y(n_654) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
AND2x2_ASAP7_75t_L g300 ( .A(n_293), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_293), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g467 ( .A(n_293), .B(n_446), .Y(n_467) );
BUFx2_ASAP7_75t_L g492 ( .A(n_293), .Y(n_492) );
AND2x4_ASAP7_75t_L g594 ( .A(n_293), .B(n_398), .Y(n_594) );
AND2x4_ASAP7_75t_L g615 ( .A(n_293), .B(n_301), .Y(n_615) );
AND2x4_ASAP7_75t_SL g620 ( .A(n_293), .B(n_393), .Y(n_620) );
HB1xp67_ASAP7_75t_L g1056 ( .A(n_294), .Y(n_1056) );
INVx3_ASAP7_75t_L g397 ( .A(n_295), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_295), .B(n_407), .Y(n_453) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_295), .Y(n_470) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_296), .Y(n_488) );
INVx2_ASAP7_75t_L g529 ( .A(n_299), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_299), .B(n_866), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g1341 ( .A(n_299), .B(n_1342), .Y(n_1341) );
INVx2_ASAP7_75t_L g601 ( .A(n_301), .Y(n_601) );
BUFx6f_ASAP7_75t_L g1348 ( .A(n_301), .Y(n_1348) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g392 ( .A(n_302), .Y(n_392) );
BUFx3_ASAP7_75t_L g734 ( .A(n_302), .Y(n_734) );
AND2x4_ASAP7_75t_L g1055 ( .A(n_302), .B(n_1056), .Y(n_1055) );
OAI31xp33_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_317), .A3(n_362), .B(n_381), .Y(n_304) );
OR2x6_ASAP7_75t_SL g306 ( .A(n_307), .B(n_311), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_308), .Y(n_372) );
AND2x4_ASAP7_75t_L g456 ( .A(n_308), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g528 ( .A(n_309), .B(n_426), .Y(n_528) );
INVx1_ASAP7_75t_L g887 ( .A(n_309), .Y(n_887) );
BUFx3_ASAP7_75t_L g339 ( .A(n_310), .Y(n_339) );
INVx3_ASAP7_75t_L g357 ( .A(n_310), .Y(n_357) );
NAND2xp33_ASAP7_75t_SL g711 ( .A(n_310), .B(n_340), .Y(n_711) );
INVx3_ASAP7_75t_L g526 ( .A(n_311), .Y(n_526) );
OAI221xp5_ASAP7_75t_L g712 ( .A1(n_311), .A2(n_713), .B1(n_714), .B2(n_718), .C(n_719), .Y(n_712) );
BUFx2_ASAP7_75t_L g826 ( .A(n_311), .Y(n_826) );
BUFx2_ASAP7_75t_L g935 ( .A(n_311), .Y(n_935) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_312), .Y(n_336) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_312), .Y(n_506) );
BUFx8_ASAP7_75t_L g564 ( .A(n_312), .Y(n_564) );
AND2x4_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
INVxp67_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g321 ( .A(n_314), .Y(n_321) );
AND2x4_ASAP7_75t_L g353 ( .A(n_315), .B(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g320 ( .A(n_316), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_316), .B(n_327), .Y(n_326) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_316), .Y(n_333) );
AND2x4_ASAP7_75t_L g369 ( .A(n_316), .B(n_370), .Y(n_369) );
OAI221xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_329), .B1(n_341), .B2(n_346), .C(n_358), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_322), .B1(n_323), .B2(n_328), .Y(n_318) );
HB1xp67_ASAP7_75t_L g1004 ( .A(n_319), .Y(n_1004) );
INVx1_ASAP7_75t_L g1016 ( .A(n_319), .Y(n_1016) );
BUFx4f_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g578 ( .A(n_320), .Y(n_578) );
OR2x4_ASAP7_75t_L g1022 ( .A(n_320), .B(n_1023), .Y(n_1022) );
OR2x4_ASAP7_75t_L g1043 ( .A(n_320), .B(n_357), .Y(n_1043) );
BUFx3_ASAP7_75t_L g1332 ( .A(n_320), .Y(n_1332) );
INVx1_ASAP7_75t_L g354 ( .A(n_321), .Y(n_354) );
INVx3_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx3_ASAP7_75t_L g344 ( .A(n_324), .Y(n_344) );
CKINVDCx8_ASAP7_75t_R g725 ( .A(n_324), .Y(n_725) );
INVx3_ASAP7_75t_L g1017 ( .A(n_324), .Y(n_1017) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g539 ( .A(n_325), .Y(n_539) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx2_ASAP7_75t_L g717 ( .A(n_326), .Y(n_717) );
INVx1_ASAP7_75t_L g332 ( .A(n_327), .Y(n_332) );
INVx2_ASAP7_75t_L g370 ( .A(n_327), .Y(n_370) );
OAI221xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_334), .B1(n_335), .B2(n_337), .C(n_338), .Y(n_329) );
OR2x6_ASAP7_75t_L g358 ( .A(n_330), .B(n_359), .Y(n_358) );
BUFx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_331), .Y(n_349) );
BUFx3_ASAP7_75t_L g1012 ( .A(n_331), .Y(n_1012) );
NAND2x1p5_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
BUFx2_ASAP7_75t_L g1039 ( .A(n_332), .Y(n_1039) );
INVx2_ASAP7_75t_L g376 ( .A(n_333), .Y(n_376) );
AND2x4_ASAP7_75t_L g457 ( .A(n_333), .B(n_380), .Y(n_457) );
BUFx2_ASAP7_75t_L g1035 ( .A(n_333), .Y(n_1035) );
OAI211xp5_ASAP7_75t_L g427 ( .A1(n_334), .A2(n_428), .B(n_431), .C(n_433), .Y(n_427) );
OAI221xp5_ASAP7_75t_L g877 ( .A1(n_335), .A2(n_878), .B1(n_879), .B2(n_880), .C(n_881), .Y(n_877) );
INVx3_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_SL g342 ( .A(n_336), .Y(n_342) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_336), .Y(n_795) );
INVx2_ASAP7_75t_SL g800 ( .A(n_336), .Y(n_800) );
INVx5_ASAP7_75t_L g939 ( .A(n_336), .Y(n_939) );
OAI221xp5_ASAP7_75t_L g1321 ( .A1(n_338), .A2(n_563), .B1(n_1007), .B2(n_1322), .C(n_1323), .Y(n_1321) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
AND3x4_ASAP7_75t_L g500 ( .A(n_339), .B(n_340), .C(n_381), .Y(n_500) );
INVx3_ASAP7_75t_L g1034 ( .A(n_339), .Y(n_1034) );
INVx1_ASAP7_75t_L g361 ( .A(n_340), .Y(n_361) );
HB1xp67_ASAP7_75t_L g1048 ( .A(n_340), .Y(n_1048) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_343), .B1(n_344), .B2(n_345), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g1008 ( .A1(n_344), .A2(n_687), .B1(n_980), .B2(n_993), .Y(n_1008) );
OAI21xp5_ASAP7_75t_SL g346 ( .A1(n_347), .A2(n_350), .B(n_351), .Y(n_346) );
OAI211xp5_ASAP7_75t_L g890 ( .A1(n_347), .A2(n_891), .B(n_892), .C(n_894), .Y(n_890) );
INVx3_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx3_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g533 ( .A(n_349), .B(n_528), .Y(n_533) );
BUFx6f_ASAP7_75t_L g1007 ( .A(n_349), .Y(n_1007) );
INVx4_ASAP7_75t_L g1331 ( .A(n_349), .Y(n_1331) );
BUFx2_ASAP7_75t_L g691 ( .A(n_352), .Y(n_691) );
BUFx3_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx8_ASAP7_75t_L g365 ( .A(n_353), .Y(n_365) );
NAND2x1p5_ASAP7_75t_L g441 ( .A(n_353), .B(n_360), .Y(n_441) );
BUFx3_ASAP7_75t_L g574 ( .A(n_353), .Y(n_574) );
AND2x2_ASAP7_75t_L g886 ( .A(n_353), .B(n_887), .Y(n_886) );
OR2x6_ASAP7_75t_L g512 ( .A(n_355), .B(n_388), .Y(n_512) );
INVx3_ASAP7_75t_L g884 ( .A(n_355), .Y(n_884) );
OR2x2_ASAP7_75t_L g1094 ( .A(n_355), .B(n_388), .Y(n_1094) );
NAND2x1p5_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
NAND3x1_ASAP7_75t_L g569 ( .A(n_356), .B(n_357), .C(n_570), .Y(n_569) );
AND2x4_ASAP7_75t_L g360 ( .A(n_357), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g1023 ( .A(n_357), .Y(n_1023) );
OR2x6_ASAP7_75t_L g1026 ( .A(n_357), .B(n_717), .Y(n_1026) );
AND2x4_ASAP7_75t_L g1029 ( .A(n_357), .B(n_369), .Y(n_1029) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x6_ASAP7_75t_L g374 ( .A(n_360), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g378 ( .A(n_360), .B(n_379), .Y(n_378) );
AND2x4_ASAP7_75t_L g515 ( .A(n_360), .B(n_452), .Y(n_515) );
AND2x4_ASAP7_75t_L g534 ( .A(n_364), .B(n_535), .Y(n_534) );
AND2x4_ASAP7_75t_L g749 ( .A(n_364), .B(n_535), .Y(n_749) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx8_ASAP7_75t_L g502 ( .A(n_365), .Y(n_502) );
CKINVDCx5p33_ASAP7_75t_R g882 ( .A(n_365), .Y(n_882) );
INVx2_ASAP7_75t_L g1093 ( .A(n_365), .Y(n_1093) );
INVx3_ASAP7_75t_L g1385 ( .A(n_365), .Y(n_1385) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_366), .A2(n_402), .B1(n_408), .B2(n_409), .Y(n_401) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g692 ( .A(n_368), .Y(n_692) );
INVx2_ASAP7_75t_L g1097 ( .A(n_368), .Y(n_1097) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx2_ASAP7_75t_L g503 ( .A(n_369), .Y(n_503) );
BUFx2_ASAP7_75t_L g521 ( .A(n_369), .Y(n_521) );
BUFx3_ASAP7_75t_L g560 ( .A(n_369), .Y(n_560) );
BUFx2_ASAP7_75t_L g684 ( .A(n_369), .Y(n_684) );
BUFx2_ASAP7_75t_L g822 ( .A(n_369), .Y(n_822) );
AND2x2_ASAP7_75t_L g889 ( .A(n_369), .B(n_887), .Y(n_889) );
INVx1_ASAP7_75t_L g380 ( .A(n_370), .Y(n_380) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx4_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_374), .A2(n_378), .B1(n_874), .B2(n_875), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g1317 ( .A1(n_374), .A2(n_378), .B1(n_1318), .B2(n_1319), .Y(n_1317) );
AND2x4_ASAP7_75t_SL g514 ( .A(n_375), .B(n_515), .Y(n_514) );
NAND2x1_ASAP7_75t_L g555 ( .A(n_375), .B(n_515), .Y(n_555) );
AND2x2_ASAP7_75t_L g695 ( .A(n_375), .B(n_515), .Y(n_695) );
AND2x2_ASAP7_75t_L g928 ( .A(n_375), .B(n_515), .Y(n_928) );
INVx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g518 ( .A(n_379), .Y(n_518) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g495 ( .A(n_381), .Y(n_495) );
INVx2_ASAP7_75t_SL g639 ( .A(n_381), .Y(n_639) );
OAI31xp33_ASAP7_75t_SL g867 ( .A1(n_381), .A2(n_868), .A3(n_870), .B(n_876), .Y(n_867) );
OAI31xp33_ASAP7_75t_SL g1311 ( .A1(n_381), .A2(n_1312), .A3(n_1316), .B(n_1320), .Y(n_1311) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx2_ASAP7_75t_L g388 ( .A(n_382), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_382), .B(n_407), .Y(n_412) );
NAND3xp33_ASAP7_75t_L g383 ( .A(n_384), .B(n_437), .C(n_448), .Y(n_383) );
NOR3xp33_ASAP7_75t_SL g384 ( .A(n_385), .B(n_416), .C(n_422), .Y(n_384) );
OAI21xp5_ASAP7_75t_SL g385 ( .A1(n_386), .A2(n_395), .B(n_401), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_390), .Y(n_386) );
HB1xp67_ASAP7_75t_L g905 ( .A(n_387), .Y(n_905) );
INVx2_ASAP7_75t_L g985 ( .A(n_387), .Y(n_985) );
INVx4_ASAP7_75t_L g1351 ( .A(n_387), .Y(n_1351) );
AND2x4_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVx1_ASAP7_75t_L g455 ( .A(n_388), .Y(n_455) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g476 ( .A(n_392), .Y(n_476) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_393), .Y(n_598) );
AND2x6_ASAP7_75t_L g608 ( .A(n_393), .B(n_407), .Y(n_608) );
BUFx3_ASAP7_75t_L g635 ( .A(n_393), .Y(n_635) );
INVx1_ASAP7_75t_L g659 ( .A(n_393), .Y(n_659) );
BUFx3_ASAP7_75t_L g778 ( .A(n_393), .Y(n_778) );
BUFx3_ASAP7_75t_L g900 ( .A(n_393), .Y(n_900) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_393), .B(n_1069), .Y(n_1068) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g964 ( .A(n_394), .Y(n_964) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_SL g605 ( .A(n_397), .Y(n_605) );
INVx2_ASAP7_75t_L g952 ( .A(n_397), .Y(n_952) );
INVx1_ASAP7_75t_L g1111 ( .A(n_397), .Y(n_1111) );
BUFx2_ASAP7_75t_L g768 ( .A(n_398), .Y(n_768) );
INVx1_ASAP7_75t_L g854 ( .A(n_398), .Y(n_854) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx3_ASAP7_75t_L g432 ( .A(n_399), .Y(n_432) );
INVx2_ASAP7_75t_L g447 ( .A(n_399), .Y(n_447) );
BUFx3_ASAP7_75t_L g607 ( .A(n_399), .Y(n_607) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_405), .B(n_407), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g491 ( .A(n_407), .Y(n_491) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_407), .B(n_485), .Y(n_1113) );
INVx2_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g914 ( .A(n_410), .Y(n_914) );
NAND2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_413), .Y(n_410) );
INVx1_ASAP7_75t_L g436 ( .A(n_411), .Y(n_436) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx2_ASAP7_75t_L g485 ( .A(n_415), .Y(n_485) );
INVx1_ASAP7_75t_L g623 ( .A(n_415), .Y(n_623) );
AND2x4_ASAP7_75t_L g1072 ( .A(n_415), .B(n_1065), .Y(n_1072) );
OR2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_420), .Y(n_417) );
INVx2_ASAP7_75t_SL g849 ( .A(n_418), .Y(n_849) );
OR2x2_ASAP7_75t_L g898 ( .A(n_418), .B(n_420), .Y(n_898) );
BUFx3_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_419), .Y(n_435) );
INVx1_ASAP7_75t_L g445 ( .A(n_420), .Y(n_445) );
INVx1_ASAP7_75t_L g452 ( .A(n_421), .Y(n_452) );
INVx1_ASAP7_75t_L g570 ( .A(n_421), .Y(n_570) );
OAI21xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_427), .B(n_434), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_SL g424 ( .A(n_425), .B(n_426), .Y(n_424) );
INVx4_ASAP7_75t_L g477 ( .A(n_425), .Y(n_477) );
INVx4_ASAP7_75t_L g603 ( .A(n_425), .Y(n_603) );
INVx1_ASAP7_75t_SL g662 ( .A(n_425), .Y(n_662) );
AND2x4_ASAP7_75t_L g909 ( .A(n_425), .B(n_910), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_425), .B(n_910), .Y(n_997) );
OR2x2_ASAP7_75t_L g710 ( .A(n_426), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g911 ( .A(n_426), .Y(n_911) );
HB1xp67_ASAP7_75t_L g1050 ( .A(n_426), .Y(n_1050) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx2_ASAP7_75t_L g981 ( .A(n_430), .Y(n_981) );
CKINVDCx5p33_ASAP7_75t_R g921 ( .A(n_434), .Y(n_921) );
OR2x6_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVx4_ASAP7_75t_L g483 ( .A(n_435), .Y(n_483) );
BUFx4f_ASAP7_75t_L g494 ( .A(n_435), .Y(n_494) );
BUFx4f_ASAP7_75t_L g766 ( .A(n_435), .Y(n_766) );
BUFx6f_ASAP7_75t_L g984 ( .A(n_435), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_440), .B(n_443), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
OR2x6_ASAP7_75t_L g497 ( .A(n_441), .B(n_442), .Y(n_497) );
INVx2_ASAP7_75t_L g872 ( .A(n_441), .Y(n_872) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AOI222xp33_ASAP7_75t_L g912 ( .A1(n_444), .A2(n_874), .B1(n_888), .B2(n_913), .C1(n_914), .C2(n_915), .Y(n_912) );
AOI21xp33_ASAP7_75t_L g1343 ( .A1(n_444), .A2(n_1344), .B(n_1345), .Y(n_1343) );
AND2x4_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
INVx3_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g664 ( .A(n_447), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_454), .Y(n_450) );
AND2x4_ASAP7_75t_L g586 ( .A(n_451), .B(n_538), .Y(n_586) );
OR2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
INVx1_ASAP7_75t_L g918 ( .A(n_452), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_453), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
INVx1_ASAP7_75t_L g677 ( .A(n_455), .Y(n_677) );
BUFx2_ASAP7_75t_L g747 ( .A(n_455), .Y(n_747) );
INVx3_ASAP7_75t_L g869 ( .A(n_456), .Y(n_869) );
BUFx12f_ASAP7_75t_L g507 ( .A(n_457), .Y(n_507) );
BUFx3_ASAP7_75t_L g565 ( .A(n_457), .Y(n_565) );
INVx5_ASAP7_75t_L g797 ( .A(n_457), .Y(n_797) );
BUFx3_ASAP7_75t_L g936 ( .A(n_457), .Y(n_936) );
BUFx2_ASAP7_75t_L g1382 ( .A(n_457), .Y(n_1382) );
XNOR2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_548), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND3xp33_ASAP7_75t_L g462 ( .A(n_463), .B(n_541), .C(n_545), .Y(n_462) );
INVx1_ASAP7_75t_L g542 ( .A(n_464), .Y(n_542) );
AOI21x1_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_495), .B(n_496), .Y(n_464) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AOI221xp5_ASAP7_75t_L g1105 ( .A1(n_467), .A2(n_608), .B1(n_1085), .B2(n_1106), .C(n_1107), .Y(n_1105) );
AOI22xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_471), .B1(n_474), .B2(n_475), .Y(n_468) );
INVx3_ASAP7_75t_L g737 ( .A(n_470), .Y(n_737) );
BUFx6f_ASAP7_75t_L g852 ( .A(n_470), .Y(n_852) );
INVx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g638 ( .A(n_473), .Y(n_638) );
INVx2_ASAP7_75t_L g966 ( .A(n_473), .Y(n_966) );
INVx2_ASAP7_75t_L g637 ( .A(n_476), .Y(n_637) );
INVx1_ASAP7_75t_L g661 ( .A(n_476), .Y(n_661) );
HB1xp67_ASAP7_75t_L g965 ( .A(n_476), .Y(n_965) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_490), .B1(n_492), .B2(n_493), .Y(n_478) );
INVx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_481), .Y(n_626) );
OAI211xp5_ASAP7_75t_L g1403 ( .A1(n_482), .A2(n_1404), .B(n_1405), .C(n_1408), .Y(n_1403) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g743 ( .A(n_483), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B1(n_487), .B2(n_489), .Y(n_484) );
AOI221xp5_ASAP7_75t_L g513 ( .A1(n_486), .A2(n_514), .B1(n_516), .B2(n_519), .C(n_520), .Y(n_513) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AOI222xp33_ASAP7_75t_L g531 ( .A1(n_489), .A2(n_532), .B1(n_534), .B2(n_536), .C1(n_537), .C2(n_540), .Y(n_531) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NOR2x1_ASAP7_75t_L g622 ( .A(n_491), .B(n_623), .Y(n_622) );
BUFx2_ASAP7_75t_L g783 ( .A(n_495), .Y(n_783) );
INVx5_ASAP7_75t_L g816 ( .A(n_497), .Y(n_816) );
INVx3_ASAP7_75t_L g1084 ( .A(n_497), .Y(n_1084) );
INVx1_ASAP7_75t_L g543 ( .A(n_498), .Y(n_543) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_513), .Y(n_498) );
AOI33xp33_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_501), .A3(n_504), .B1(n_508), .B2(n_510), .B3(n_511), .Y(n_499) );
AOI33xp33_ASAP7_75t_L g558 ( .A1(n_500), .A2(n_559), .A3(n_561), .B1(n_566), .B2(n_567), .B3(n_571), .Y(n_558) );
AOI33xp33_ASAP7_75t_L g682 ( .A1(n_500), .A2(n_683), .A3(n_685), .B1(n_688), .B2(n_689), .B3(n_690), .Y(n_682) );
AOI33xp33_ASAP7_75t_L g792 ( .A1(n_500), .A2(n_567), .A3(n_793), .B1(n_794), .B2(n_798), .B3(n_801), .Y(n_792) );
BUFx3_ASAP7_75t_L g823 ( .A(n_500), .Y(n_823) );
INVx1_ASAP7_75t_L g1098 ( .A(n_500), .Y(n_1098) );
AOI33xp33_ASAP7_75t_L g1377 ( .A1(n_500), .A2(n_1378), .A3(n_1381), .B1(n_1383), .B2(n_1384), .B3(n_1386), .Y(n_1377) );
BUFx2_ASAP7_75t_L g819 ( .A(n_502), .Y(n_819) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_506), .Y(n_509) );
INVx2_ASAP7_75t_L g687 ( .A(n_506), .Y(n_687) );
INVx2_ASAP7_75t_L g723 ( .A(n_506), .Y(n_723) );
AND2x4_ASAP7_75t_L g1045 ( .A(n_506), .B(n_1023), .Y(n_1045) );
INVx1_ASAP7_75t_L g1010 ( .A(n_509), .Y(n_1010) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g1088 ( .A1(n_514), .A2(n_516), .B1(n_1089), .B2(n_1090), .Y(n_1088) );
AND2x4_ASAP7_75t_SL g516 ( .A(n_515), .B(n_517), .Y(n_516) );
AND2x4_ASAP7_75t_L g520 ( .A(n_515), .B(n_521), .Y(n_520) );
AND2x4_ASAP7_75t_L g557 ( .A(n_515), .B(n_517), .Y(n_557) );
INVx1_ASAP7_75t_L g729 ( .A(n_516), .Y(n_729) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx3_ASAP7_75t_L g583 ( .A(n_520), .Y(n_583) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_520), .Y(n_707) );
INVx3_ASAP7_75t_L g805 ( .A(n_520), .Y(n_805) );
BUFx2_ASAP7_75t_L g932 ( .A(n_521), .Y(n_932) );
INVx1_ASAP7_75t_L g547 ( .A(n_522), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_530), .Y(n_522) );
NAND2x1_ASAP7_75t_L g523 ( .A(n_524), .B(n_529), .Y(n_523) );
INVx2_ASAP7_75t_SL g524 ( .A(n_525), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_525), .A2(n_534), .B1(n_1103), .B2(n_1104), .Y(n_1115) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
INVxp67_ASAP7_75t_L g579 ( .A(n_527), .Y(n_579) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g535 ( .A(n_528), .Y(n_535) );
OR2x2_ASAP7_75t_L g538 ( .A(n_528), .B(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g546 ( .A(n_531), .Y(n_546) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x4_ASAP7_75t_L g589 ( .A(n_533), .B(n_590), .Y(n_589) );
AND2x4_ASAP7_75t_L g705 ( .A(n_533), .B(n_590), .Y(n_705) );
AND2x4_ASAP7_75t_L g581 ( .A(n_535), .B(n_564), .Y(n_581) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
BUFx3_ASAP7_75t_L g879 ( .A(n_539), .Y(n_879) );
INVx1_ASAP7_75t_L g1338 ( .A(n_539), .Y(n_1338) );
OAI21xp5_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_543), .B(n_544), .Y(n_541) );
OAI21xp33_ASAP7_75t_L g545 ( .A1(n_544), .A2(n_546), .B(n_547), .Y(n_545) );
NAND3xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_584), .C(n_591), .Y(n_549) );
NOR3xp33_ASAP7_75t_L g550 ( .A(n_551), .B(n_575), .C(n_582), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_558), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_554), .B1(n_556), .B2(n_557), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g1372 ( .A1(n_554), .A2(n_557), .B1(n_1373), .B2(n_1374), .Y(n_1372) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_557), .A2(n_694), .B1(n_695), .B2(n_696), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_557), .A2(n_695), .B1(n_790), .B2(n_791), .Y(n_789) );
AOI22xp5_ASAP7_75t_L g811 ( .A1(n_557), .A2(n_695), .B1(n_812), .B2(n_813), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_557), .A2(n_927), .B1(n_928), .B2(n_929), .Y(n_926) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g1334 ( .A1(n_563), .A2(n_1335), .B1(n_1336), .B2(n_1337), .Y(n_1334) );
INVx3_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx3_ASAP7_75t_L g830 ( .A(n_564), .Y(n_830) );
AOI33xp33_ASAP7_75t_L g930 ( .A1(n_567), .A2(n_823), .A3(n_931), .B1(n_933), .B2(n_937), .B3(n_940), .Y(n_930) );
BUFx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
BUFx2_ASAP7_75t_L g689 ( .A(n_568), .Y(n_689) );
BUFx2_ASAP7_75t_L g1386 ( .A(n_568), .Y(n_1386) );
INVx3_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx3_ASAP7_75t_L g721 ( .A(n_569), .Y(n_721) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx2_ASAP7_75t_SL g1380 ( .A(n_574), .Y(n_1380) );
OR2x6_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .Y(n_576) );
OR2x2_ASAP7_75t_L g803 ( .A(n_577), .B(n_579), .Y(n_803) );
INVx2_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
INVx3_ASAP7_75t_L g1326 ( .A(n_578), .Y(n_1326) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g681 ( .A(n_581), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_581), .A2(n_739), .B1(n_740), .B2(n_749), .Y(n_748) );
INVx2_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
AND4x1_ASAP7_75t_L g678 ( .A(n_583), .B(n_679), .C(n_682), .D(n_693), .Y(n_678) );
NAND3xp33_ASAP7_75t_SL g1087 ( .A(n_583), .B(n_1088), .C(n_1091), .Y(n_1087) );
AOI21xp33_ASAP7_75t_SL g584 ( .A1(n_585), .A2(n_587), .B(n_588), .Y(n_584) );
AOI21xp33_ASAP7_75t_L g646 ( .A1(n_585), .A2(n_647), .B(n_648), .Y(n_646) );
AOI21xp5_ASAP7_75t_L g702 ( .A1(n_585), .A2(n_703), .B(n_704), .Y(n_702) );
AOI21xp33_ASAP7_75t_SL g784 ( .A1(n_585), .A2(n_785), .B(n_786), .Y(n_784) );
AOI211x1_ASAP7_75t_L g808 ( .A1(n_585), .A2(n_809), .B(n_810), .C(n_832), .Y(n_808) );
AOI21xp5_ASAP7_75t_L g942 ( .A1(n_585), .A2(n_943), .B(n_944), .Y(n_942) );
AOI221xp5_ASAP7_75t_L g1083 ( .A1(n_585), .A2(n_1084), .B1(n_1085), .B2(n_1086), .C(n_1087), .Y(n_1083) );
NAND2xp33_ASAP7_75t_L g1387 ( .A(n_585), .B(n_1388), .Y(n_1387) );
INVx8_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g834 ( .A(n_589), .Y(n_834) );
INVx2_ASAP7_75t_SL g915 ( .A(n_590), .Y(n_915) );
OAI21xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_616), .B(n_639), .Y(n_591) );
INVx2_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
INVx3_ASAP7_75t_L g651 ( .A(n_594), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_594), .A2(n_654), .B1(n_761), .B2(n_762), .Y(n_760) );
AOI21xp5_ASAP7_75t_SL g595 ( .A1(n_596), .A2(n_604), .B(n_608), .Y(n_595) );
BUFx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g950 ( .A(n_600), .Y(n_950) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
HB1xp67_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
BUFx3_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AOI21xp5_ASAP7_75t_L g656 ( .A1(n_608), .A2(n_657), .B(n_663), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g732 ( .A1(n_608), .A2(n_733), .B(n_735), .Y(n_732) );
AOI21xp5_ASAP7_75t_L g758 ( .A1(n_608), .A2(n_614), .B(n_759), .Y(n_758) );
AOI21xp5_ASAP7_75t_L g839 ( .A1(n_608), .A2(n_840), .B(n_841), .Y(n_839) );
AOI21xp5_ASAP7_75t_L g947 ( .A1(n_608), .A2(n_948), .B(n_951), .Y(n_947) );
AOI21xp5_ASAP7_75t_L g1396 ( .A1(n_608), .A2(n_1397), .B(n_1398), .Y(n_1396) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_611), .B1(n_613), .B2(n_614), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_611), .A2(n_954), .B1(n_955), .B2(n_956), .Y(n_953) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_614), .A2(n_653), .B1(n_654), .B2(n_655), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_614), .A2(n_654), .B1(n_843), .B2(n_844), .Y(n_842) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_615), .A2(n_654), .B1(n_739), .B2(n_740), .Y(n_738) );
INVx1_ASAP7_75t_L g957 ( .A(n_615), .Y(n_957) );
AOI22xp5_ASAP7_75t_L g1102 ( .A1(n_615), .A2(n_654), .B1(n_1103), .B2(n_1104), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g1399 ( .A1(n_615), .A2(n_654), .B1(n_1400), .B2(n_1401), .Y(n_1399) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g780 ( .A(n_618), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_618), .A2(n_622), .B1(n_927), .B2(n_929), .Y(n_969) );
INVx4_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
BUFx3_ASAP7_75t_L g1109 ( .A(n_620), .Y(n_1109) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g667 ( .A(n_622), .Y(n_667) );
OAI221xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_627), .B1(n_628), .B2(n_633), .C(n_634), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
BUFx2_ASAP7_75t_L g673 ( .A(n_628), .Y(n_673) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_SL g775 ( .A(n_630), .Y(n_775) );
INVx2_ASAP7_75t_L g904 ( .A(n_630), .Y(n_904) );
BUFx6f_ASAP7_75t_L g959 ( .A(n_630), .Y(n_959) );
INVx4_ASAP7_75t_L g991 ( .A(n_630), .Y(n_991) );
INVx8_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g1064 ( .A(n_631), .B(n_1065), .Y(n_1064) );
BUFx6f_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g770 ( .A(n_637), .Y(n_770) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B1(n_698), .B2(n_750), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AO21x2_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_645), .B(n_697), .Y(n_643) );
NAND3xp33_ASAP7_75t_SL g645 ( .A(n_646), .B(n_649), .C(n_678), .Y(n_645) );
OAI21xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_665), .B(n_677), .Y(n_649) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g676 ( .A(n_659), .Y(n_676) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
BUFx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
OAI221xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_672), .B1(n_673), .B2(n_674), .C(n_675), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g986 ( .A1(n_669), .A2(n_987), .B1(n_988), .B2(n_989), .Y(n_986) );
OAI22xp33_ASAP7_75t_L g992 ( .A1(n_669), .A2(n_984), .B1(n_993), .B2(n_994), .Y(n_992) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx2_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
BUFx6f_ASAP7_75t_L g772 ( .A(n_671), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g901 ( .A1(n_671), .A2(n_902), .B1(n_903), .B2(n_904), .Y(n_901) );
OAI22x1_ASAP7_75t_SL g907 ( .A1(n_671), .A2(n_880), .B1(n_904), .B2(n_908), .Y(n_907) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g1013 ( .A(n_689), .Y(n_1013) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g751 ( .A(n_699), .Y(n_751) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AND4x1_ASAP7_75t_L g701 ( .A(n_702), .B(n_706), .C(n_730), .D(n_748), .Y(n_701) );
NOR3xp33_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .C(n_728), .Y(n_706) );
NOR3xp33_ASAP7_75t_L g924 ( .A(n_707), .B(n_925), .C(n_941), .Y(n_924) );
OAI22xp5_ASAP7_75t_SL g708 ( .A1(n_709), .A2(n_712), .B1(n_720), .B2(n_722), .Y(n_708) );
BUFx3_ASAP7_75t_L g1002 ( .A(n_709), .Y(n_1002) );
BUFx4f_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
BUFx2_ASAP7_75t_L g893 ( .A(n_711), .Y(n_893) );
INVx3_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
BUFx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AOI33xp33_ASAP7_75t_L g817 ( .A1(n_721), .A2(n_818), .A3(n_823), .B1(n_824), .B2(n_828), .B3(n_831), .Y(n_817) );
OAI221xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_724), .B1(n_725), .B2(n_726), .C(n_727), .Y(n_722) );
OAI211xp5_ASAP7_75t_L g742 ( .A1(n_724), .A2(n_743), .B(n_744), .C(n_745), .Y(n_742) );
OAI21xp5_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_741), .B(n_746), .Y(n_730) );
INVx1_ASAP7_75t_L g1407 ( .A(n_734), .Y(n_1407) );
INVx2_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
AOI21xp5_ASAP7_75t_L g1100 ( .A1(n_746), .A2(n_1101), .B(n_1114), .Y(n_1100) );
OAI21xp5_ASAP7_75t_L g1394 ( .A1(n_746), .A2(n_1395), .B(n_1402), .Y(n_1394) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g855 ( .A(n_747), .Y(n_855) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g1118 ( .A(n_752), .Y(n_1118) );
XNOR2xp5_ASAP7_75t_L g752 ( .A(n_753), .B(n_856), .Y(n_752) );
XNOR2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_806), .Y(n_753) );
NAND3xp33_ASAP7_75t_L g755 ( .A(n_756), .B(n_784), .C(n_787), .Y(n_755) );
OAI31xp33_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_763), .A3(n_779), .B(n_781), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_758), .B(n_760), .Y(n_757) );
OAI211xp5_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_766), .B(n_767), .C(n_769), .Y(n_764) );
OAI221xp5_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_773), .B1(n_774), .B2(n_776), .C(n_777), .Y(n_771) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g971 ( .A(n_783), .Y(n_971) );
NOR3xp33_ASAP7_75t_L g787 ( .A(n_788), .B(n_802), .C(n_804), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_789), .B(n_792), .Y(n_788) );
INVx2_ASAP7_75t_R g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g827 ( .A(n_797), .Y(n_827) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
NAND4xp25_ASAP7_75t_SL g810 ( .A(n_805), .B(n_811), .C(n_814), .D(n_817), .Y(n_810) );
NAND4xp25_ASAP7_75t_SL g1371 ( .A(n_805), .B(n_1372), .C(n_1375), .D(n_1377), .Y(n_1371) );
XNOR2x2_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g1375 ( .A(n_816), .B(n_1376), .Y(n_1375) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_833), .B(n_837), .Y(n_832) );
AOI21xp5_ASAP7_75t_L g833 ( .A1(n_834), .A2(n_835), .B(n_836), .Y(n_833) );
AOI21xp5_ASAP7_75t_L g1391 ( .A1(n_834), .A2(n_1392), .B(n_1393), .Y(n_1391) );
OAI21xp33_ASAP7_75t_L g837 ( .A1(n_838), .A2(n_845), .B(n_855), .Y(n_837) );
OAI211xp5_ASAP7_75t_L g846 ( .A1(n_847), .A2(n_848), .B(n_850), .C(n_851), .Y(n_846) );
INVx5_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
AOI22xp5_ASAP7_75t_SL g856 ( .A1(n_857), .A2(n_858), .B1(n_974), .B2(n_1117), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
OAI22xp5_ASAP7_75t_L g858 ( .A1(n_859), .A2(n_922), .B1(n_972), .B2(n_973), .Y(n_858) );
INVx1_ASAP7_75t_L g973 ( .A(n_859), .Y(n_973) );
HB1xp67_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
AOI211x1_ASAP7_75t_L g861 ( .A1(n_862), .A2(n_863), .B(n_864), .C(n_895), .Y(n_861) );
AOI22xp5_ASAP7_75t_L g885 ( .A1(n_863), .A2(n_886), .B1(n_888), .B2(n_889), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_865), .B(n_867), .Y(n_864) );
INVx2_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
AOI222xp33_ASAP7_75t_L g896 ( .A1(n_875), .A2(n_897), .B1(n_899), .B2(n_905), .C1(n_906), .C2(n_909), .Y(n_896) );
NAND3xp33_ASAP7_75t_L g876 ( .A(n_877), .B(n_885), .C(n_890), .Y(n_876) );
INVx3_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
OAI221xp5_ASAP7_75t_L g1328 ( .A1(n_884), .A2(n_1329), .B1(n_1330), .B2(n_1332), .C(n_1333), .Y(n_1328) );
AOI22xp5_ASAP7_75t_L g1313 ( .A1(n_886), .A2(n_889), .B1(n_1314), .B2(n_1315), .Y(n_1313) );
NAND3xp33_ASAP7_75t_L g895 ( .A(n_896), .B(n_912), .C(n_916), .Y(n_895) );
AOI21xp5_ASAP7_75t_L g1340 ( .A1(n_897), .A2(n_921), .B(n_1319), .Y(n_1340) );
INVx2_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
AOI332xp33_ASAP7_75t_L g1346 ( .A1(n_909), .A2(n_917), .A3(n_1347), .B1(n_1349), .B2(n_1350), .B3(n_1352), .C1(n_1353), .C2(n_1354), .Y(n_1346) );
INVx1_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
AOI21xp33_ASAP7_75t_SL g916 ( .A1(n_917), .A2(n_920), .B(n_921), .Y(n_916) );
AND2x4_ASAP7_75t_L g917 ( .A(n_918), .B(n_919), .Y(n_917) );
INVx1_ASAP7_75t_L g972 ( .A(n_922), .Y(n_972) );
NAND3xp33_ASAP7_75t_L g923 ( .A(n_924), .B(n_942), .C(n_945), .Y(n_923) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_926), .B(n_930), .Y(n_925) );
INVx2_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx8_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
OAI21xp5_ASAP7_75t_L g945 ( .A1(n_946), .A2(n_958), .B(n_970), .Y(n_945) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
INVx1_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g960 ( .A(n_961), .B(n_967), .Y(n_960) );
INVx2_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
BUFx2_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
INVx2_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
INVx1_ASAP7_75t_L g1117 ( .A(n_974), .Y(n_1117) );
AO22x1_ASAP7_75t_L g974 ( .A1(n_975), .A2(n_1080), .B1(n_1081), .B2(n_1116), .Y(n_974) );
INVx1_ASAP7_75t_L g1116 ( .A(n_975), .Y(n_1116) );
NAND3xp33_ASAP7_75t_L g976 ( .A(n_977), .B(n_1018), .C(n_1051), .Y(n_976) );
NOR2xp33_ASAP7_75t_L g977 ( .A(n_978), .B(n_1001), .Y(n_977) );
OAI33xp33_ASAP7_75t_L g978 ( .A1(n_979), .A2(n_985), .A3(n_986), .B1(n_992), .B2(n_995), .B3(n_998), .Y(n_978) );
OAI22xp5_ASAP7_75t_L g979 ( .A1(n_980), .A2(n_981), .B1(n_982), .B2(n_983), .Y(n_979) );
OAI22xp5_ASAP7_75t_L g998 ( .A1(n_981), .A2(n_989), .B1(n_999), .B2(n_1000), .Y(n_998) );
OAI22xp5_ASAP7_75t_L g1009 ( .A1(n_982), .A2(n_994), .B1(n_1010), .B2(n_1011), .Y(n_1009) );
HB1xp67_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
OAI22xp33_ASAP7_75t_L g1003 ( .A1(n_987), .A2(n_999), .B1(n_1004), .B2(n_1005), .Y(n_1003) );
OAI22xp5_ASAP7_75t_L g1014 ( .A1(n_988), .A2(n_1000), .B1(n_1015), .B2(n_1017), .Y(n_1014) );
INVx2_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
INVx2_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
INVx2_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
INVx1_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
OAI33xp33_ASAP7_75t_L g1001 ( .A1(n_1002), .A2(n_1003), .A3(n_1008), .B1(n_1009), .B2(n_1013), .B3(n_1014), .Y(n_1001) );
INVx2_ASAP7_75t_SL g1005 ( .A(n_1006), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
BUFx6f_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
INVx2_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
OAI22xp5_ASAP7_75t_L g1324 ( .A1(n_1017), .A2(n_1325), .B1(n_1326), .B2(n_1327), .Y(n_1324) );
OAI31xp33_ASAP7_75t_L g1018 ( .A1(n_1019), .A2(n_1027), .A3(n_1040), .B(n_1046), .Y(n_1018) );
INVx1_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
INVx2_ASAP7_75t_SL g1021 ( .A(n_1022), .Y(n_1021) );
INVx2_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
INVx2_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
CKINVDCx8_ASAP7_75t_R g1028 ( .A(n_1029), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g1030 ( .A1(n_1031), .A2(n_1032), .B1(n_1036), .B2(n_1037), .Y(n_1030) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_1031), .A2(n_1071), .B1(n_1073), .B2(n_1074), .Y(n_1070) );
BUFx3_ASAP7_75t_L g1032 ( .A(n_1033), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1035), .Y(n_1033) );
AND2x4_ASAP7_75t_L g1038 ( .A(n_1034), .B(n_1039), .Y(n_1038) );
BUFx6f_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
INVx1_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
INVx1_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
AND2x2_ASAP7_75t_SL g1046 ( .A(n_1047), .B(n_1049), .Y(n_1046) );
INVx1_ASAP7_75t_SL g1047 ( .A(n_1048), .Y(n_1047) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
OAI31xp33_ASAP7_75t_SL g1051 ( .A1(n_1052), .A2(n_1057), .A3(n_1066), .B(n_1077), .Y(n_1051) );
INVx3_ASAP7_75t_SL g1054 ( .A(n_1055), .Y(n_1054) );
HB1xp67_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
INVx2_ASAP7_75t_L g1060 ( .A(n_1061), .Y(n_1060) );
INVx2_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
INVx2_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
INVx3_ASAP7_75t_L g1067 ( .A(n_1068), .Y(n_1067) );
BUFx3_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
INVx2_ASAP7_75t_L g1074 ( .A(n_1075), .Y(n_1074) );
INVx2_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
BUFx3_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1081), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1100), .Y(n_1082) );
AOI222xp33_ASAP7_75t_L g1108 ( .A1(n_1089), .A2(n_1090), .B1(n_1109), .B2(n_1110), .C1(n_1112), .C2(n_1113), .Y(n_1108) );
AOI22xp5_ASAP7_75t_L g1091 ( .A1(n_1092), .A2(n_1095), .B1(n_1096), .B2(n_1099), .Y(n_1091) );
NAND3xp33_ASAP7_75t_L g1101 ( .A(n_1102), .B(n_1105), .C(n_1108), .Y(n_1101) );
OAI221xp5_ASAP7_75t_L g1119 ( .A1(n_1120), .A2(n_1304), .B1(n_1307), .B2(n_1356), .C(n_1362), .Y(n_1119) );
NOR3xp33_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1243), .C(n_1280), .Y(n_1120) );
AOI32xp33_ASAP7_75t_L g1121 ( .A1(n_1122), .A2(n_1209), .A3(n_1228), .B1(n_1232), .B2(n_1242), .Y(n_1121) );
AOI211xp5_ASAP7_75t_L g1122 ( .A1(n_1123), .A2(n_1138), .B(n_1173), .C(n_1197), .Y(n_1122) );
OAI311xp33_ASAP7_75t_L g1173 ( .A1(n_1123), .A2(n_1174), .A3(n_1179), .B1(n_1180), .C1(n_1192), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1241 ( .A(n_1123), .B(n_1144), .Y(n_1241) );
AOI21xp33_ASAP7_75t_L g1276 ( .A1(n_1123), .A2(n_1277), .B(n_1279), .Y(n_1276) );
OR2x2_ASAP7_75t_L g1288 ( .A(n_1123), .B(n_1140), .Y(n_1288) );
AND2x2_ASAP7_75t_L g1302 ( .A(n_1123), .B(n_1167), .Y(n_1302) );
INVx3_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
NOR2xp33_ASAP7_75t_L g1181 ( .A(n_1124), .B(n_1182), .Y(n_1181) );
OR2x2_ASAP7_75t_L g1186 ( .A(n_1124), .B(n_1144), .Y(n_1186) );
OR2x2_ASAP7_75t_L g1211 ( .A(n_1124), .B(n_1212), .Y(n_1211) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1124), .B(n_1178), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1124), .B(n_1193), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1124), .B(n_1208), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1263 ( .A(n_1124), .B(n_1264), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1273 ( .A(n_1124), .B(n_1242), .Y(n_1273) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1124), .B(n_1144), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_1124), .B(n_1164), .Y(n_1293) );
AND2x4_ASAP7_75t_SL g1124 ( .A(n_1125), .B(n_1132), .Y(n_1124) );
INVx2_ASAP7_75t_L g1306 ( .A(n_1126), .Y(n_1306) );
AND2x6_ASAP7_75t_L g1126 ( .A(n_1127), .B(n_1128), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_1127), .B(n_1131), .Y(n_1130) );
AND2x4_ASAP7_75t_L g1133 ( .A(n_1127), .B(n_1134), .Y(n_1133) );
AND2x6_ASAP7_75t_L g1136 ( .A(n_1127), .B(n_1137), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_1127), .B(n_1131), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_1127), .B(n_1131), .Y(n_1153) );
HB1xp67_ASAP7_75t_L g1414 ( .A(n_1128), .Y(n_1414) );
AND2x2_ASAP7_75t_L g1134 ( .A(n_1129), .B(n_1135), .Y(n_1134) );
OAI22xp5_ASAP7_75t_L g1138 ( .A1(n_1139), .A2(n_1148), .B1(n_1164), .B2(n_1166), .Y(n_1138) );
A2O1A1Ixp33_ASAP7_75t_L g1224 ( .A1(n_1139), .A2(n_1167), .B(n_1225), .C(n_1226), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1139), .B(n_1199), .Y(n_1252) );
NAND2xp5_ASAP7_75t_L g1301 ( .A(n_1139), .B(n_1302), .Y(n_1301) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
OR2x2_ASAP7_75t_L g1140 ( .A(n_1141), .B(n_1144), .Y(n_1140) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1141), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1141), .B(n_1144), .Y(n_1178) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1141), .Y(n_1183) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1141), .Y(n_1193) );
NAND2xp5_ASAP7_75t_L g1141 ( .A(n_1142), .B(n_1143), .Y(n_1141) );
OR2x2_ASAP7_75t_L g1212 ( .A(n_1144), .B(n_1183), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g1299 ( .A(n_1144), .B(n_1236), .Y(n_1299) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_1145), .B(n_1147), .Y(n_1144) );
AND2x4_ASAP7_75t_L g1200 ( .A(n_1145), .B(n_1147), .Y(n_1200) );
AOI31xp33_ASAP7_75t_L g1250 ( .A1(n_1148), .A2(n_1246), .A3(n_1248), .B(n_1251), .Y(n_1250) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
OAI21xp5_ASAP7_75t_L g1257 ( .A1(n_1149), .A2(n_1258), .B(n_1260), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1150), .B(n_1155), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1150), .B(n_1195), .Y(n_1194) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1150), .B(n_1172), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1150), .B(n_1219), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1226 ( .A(n_1150), .B(n_1227), .Y(n_1226) );
OR2x2_ASAP7_75t_L g1248 ( .A(n_1150), .B(n_1249), .Y(n_1248) );
CKINVDCx5p33_ASAP7_75t_R g1150 ( .A(n_1151), .Y(n_1150) );
NAND2xp5_ASAP7_75t_L g1171 ( .A(n_1151), .B(n_1172), .Y(n_1171) );
NOR2xp33_ASAP7_75t_L g1184 ( .A(n_1151), .B(n_1157), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1151), .B(n_1156), .Y(n_1187) );
NOR2xp33_ASAP7_75t_L g1234 ( .A(n_1151), .B(n_1167), .Y(n_1234) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_1151), .B(n_1227), .Y(n_1240) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1151), .B(n_1167), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_1152), .B(n_1154), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1152), .B(n_1154), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1155), .B(n_1176), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1155), .B(n_1213), .Y(n_1238) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1155), .Y(n_1297) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1156), .B(n_1160), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
OR2x2_ASAP7_75t_L g1196 ( .A(n_1157), .B(n_1160), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1207 ( .A(n_1157), .B(n_1160), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1157), .B(n_1161), .Y(n_1227) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1157), .Y(n_1274) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1158), .B(n_1159), .Y(n_1157) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1160), .Y(n_1172) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1161), .Y(n_1179) );
NAND2xp5_ASAP7_75t_L g1161 ( .A(n_1162), .B(n_1163), .Y(n_1161) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1164), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_1164), .B(n_1268), .Y(n_1278) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
NAND2xp5_ASAP7_75t_L g1166 ( .A(n_1167), .B(n_1170), .Y(n_1166) );
INVx3_ASAP7_75t_L g1177 ( .A(n_1167), .Y(n_1177) );
OR2x2_ASAP7_75t_L g1182 ( .A(n_1167), .B(n_1183), .Y(n_1182) );
INVx2_ASAP7_75t_L g1199 ( .A(n_1167), .Y(n_1199) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1168), .B(n_1169), .Y(n_1167) );
OAI332xp33_ASAP7_75t_L g1295 ( .A1(n_1170), .A2(n_1211), .A3(n_1274), .B1(n_1296), .B2(n_1299), .B3(n_1300), .C1(n_1301), .C2(n_1303), .Y(n_1295) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
OR2x2_ASAP7_75t_L g1259 ( .A(n_1171), .B(n_1176), .Y(n_1259) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1176), .B(n_1178), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1176), .B(n_1206), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1176), .B(n_1184), .Y(n_1282) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1177), .Y(n_1176) );
NOR2xp33_ASAP7_75t_L g1195 ( .A(n_1177), .B(n_1196), .Y(n_1195) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_1177), .B(n_1207), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1177), .B(n_1238), .Y(n_1294) );
CKINVDCx14_ASAP7_75t_R g1203 ( .A(n_1178), .Y(n_1203) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1179), .Y(n_1225) );
AOI221xp5_ASAP7_75t_L g1180 ( .A1(n_1181), .A2(n_1184), .B1(n_1185), .B2(n_1187), .C(n_1188), .Y(n_1180) );
CKINVDCx14_ASAP7_75t_R g1262 ( .A(n_1182), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1183), .B(n_1200), .Y(n_1272) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
OAI221xp5_ASAP7_75t_L g1270 ( .A1(n_1186), .A2(n_1198), .B1(n_1271), .B2(n_1274), .C(n_1275), .Y(n_1270) );
NAND2xp5_ASAP7_75t_L g1198 ( .A(n_1187), .B(n_1199), .Y(n_1198) );
CKINVDCx14_ASAP7_75t_R g1303 ( .A(n_1187), .Y(n_1303) );
OAI31xp33_ASAP7_75t_L g1244 ( .A1(n_1188), .A2(n_1245), .A3(n_1250), .B(n_1253), .Y(n_1244) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1189), .Y(n_1188) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1189), .Y(n_1242) );
AOI21xp33_ASAP7_75t_SL g1290 ( .A1(n_1189), .A2(n_1291), .B(n_1292), .Y(n_1290) );
AND2x2_ASAP7_75t_L g1189 ( .A(n_1190), .B(n_1191), .Y(n_1189) );
NAND2xp5_ASAP7_75t_L g1192 ( .A(n_1193), .B(n_1194), .Y(n_1192) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1193), .Y(n_1206) );
A2O1A1Ixp33_ASAP7_75t_SL g1232 ( .A1(n_1193), .A2(n_1233), .B(n_1235), .C(n_1241), .Y(n_1232) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1194), .Y(n_1279) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1196), .Y(n_1219) );
OAI221xp5_ASAP7_75t_L g1197 ( .A1(n_1198), .A2(n_1200), .B1(n_1201), .B2(n_1203), .C(n_1204), .Y(n_1197) );
OR2x2_ASAP7_75t_L g1230 ( .A(n_1199), .B(n_1231), .Y(n_1230) );
AOI22xp33_ASAP7_75t_L g1235 ( .A1(n_1199), .A2(n_1236), .B1(n_1237), .B2(n_1239), .Y(n_1235) );
INVx2_ASAP7_75t_L g1236 ( .A(n_1199), .Y(n_1236) );
INVx2_ASAP7_75t_L g1208 ( .A(n_1200), .Y(n_1208) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1202), .Y(n_1201) );
AOI21xp33_ASAP7_75t_L g1245 ( .A1(n_1203), .A2(n_1246), .B(n_1248), .Y(n_1245) );
A2O1A1Ixp33_ASAP7_75t_L g1266 ( .A1(n_1203), .A2(n_1255), .B(n_1267), .C(n_1269), .Y(n_1266) );
NAND3xp33_ASAP7_75t_L g1204 ( .A(n_1205), .B(n_1207), .C(n_1208), .Y(n_1204) );
NAND2xp5_ASAP7_75t_L g1228 ( .A(n_1206), .B(n_1229), .Y(n_1228) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1207), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_1207), .B(n_1234), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1207), .B(n_1247), .Y(n_1268) );
AOI221xp5_ASAP7_75t_L g1209 ( .A1(n_1210), .A2(n_1213), .B1(n_1214), .B2(n_1215), .C(n_1216), .Y(n_1209) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
INVx2_ASAP7_75t_SL g1264 ( .A(n_1212), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1213), .B(n_1221), .Y(n_1284) );
NAND2xp5_ASAP7_75t_L g1269 ( .A(n_1214), .B(n_1218), .Y(n_1269) );
AOI321xp33_ASAP7_75t_L g1289 ( .A1(n_1215), .A2(n_1236), .A3(n_1285), .B1(n_1290), .B2(n_1294), .C(n_1295), .Y(n_1289) );
A2O1A1Ixp33_ASAP7_75t_L g1216 ( .A1(n_1217), .A2(n_1220), .B(n_1222), .C(n_1224), .Y(n_1216) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1219), .B(n_1234), .Y(n_1233) );
NAND2xp5_ASAP7_75t_L g1246 ( .A(n_1219), .B(n_1247), .Y(n_1246) );
A2O1A1Ixp33_ASAP7_75t_L g1280 ( .A1(n_1220), .A2(n_1281), .B(n_1283), .C(n_1289), .Y(n_1280) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1226), .Y(n_1231) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1227), .Y(n_1298) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
NAND3xp33_ASAP7_75t_L g1271 ( .A(n_1236), .B(n_1272), .C(n_1273), .Y(n_1271) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
OAI21xp5_ASAP7_75t_L g1275 ( .A1(n_1238), .A2(n_1258), .B(n_1264), .Y(n_1275) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
OAI21xp33_ASAP7_75t_L g1261 ( .A1(n_1240), .A2(n_1262), .B(n_1263), .Y(n_1261) );
NAND2xp5_ASAP7_75t_L g1243 ( .A(n_1244), .B(n_1265), .Y(n_1243) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
OAI211xp5_ASAP7_75t_L g1253 ( .A1(n_1254), .A2(n_1255), .B(n_1257), .C(n_1261), .Y(n_1253) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1259), .Y(n_1258) );
NOR3xp33_ASAP7_75t_L g1265 ( .A(n_1266), .B(n_1270), .C(n_1276), .Y(n_1265) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1268), .Y(n_1267) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1272), .Y(n_1291) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1273), .Y(n_1300) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
CKINVDCx14_ASAP7_75t_R g1281 ( .A(n_1282), .Y(n_1281) );
AOI21xp5_ASAP7_75t_L g1283 ( .A1(n_1284), .A2(n_1285), .B(n_1287), .Y(n_1283) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1288), .Y(n_1287) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1293), .Y(n_1292) );
NAND2xp5_ASAP7_75t_L g1296 ( .A(n_1297), .B(n_1298), .Y(n_1296) );
CKINVDCx20_ASAP7_75t_R g1304 ( .A(n_1305), .Y(n_1304) );
CKINVDCx20_ASAP7_75t_R g1305 ( .A(n_1306), .Y(n_1305) );
XOR2x2_ASAP7_75t_L g1307 ( .A(n_1308), .B(n_1355), .Y(n_1307) );
NOR2xp33_ASAP7_75t_L g1308 ( .A(n_1309), .B(n_1339), .Y(n_1308) );
OAI22xp5_ASAP7_75t_L g1320 ( .A1(n_1321), .A2(n_1324), .B1(n_1328), .B2(n_1334), .Y(n_1320) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1331), .Y(n_1330) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
NAND4xp25_ASAP7_75t_SL g1339 ( .A(n_1340), .B(n_1341), .C(n_1343), .D(n_1346), .Y(n_1339) );
INVx2_ASAP7_75t_SL g1350 ( .A(n_1351), .Y(n_1350) );
CKINVDCx20_ASAP7_75t_R g1356 ( .A(n_1357), .Y(n_1356) );
CKINVDCx20_ASAP7_75t_R g1357 ( .A(n_1358), .Y(n_1357) );
INVx3_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
BUFx3_ASAP7_75t_L g1359 ( .A(n_1360), .Y(n_1359) );
HB1xp67_ASAP7_75t_SL g1363 ( .A(n_1364), .Y(n_1363) );
INVxp33_ASAP7_75t_SL g1365 ( .A(n_1366), .Y(n_1365) );
INVx1_ASAP7_75t_L g1410 ( .A(n_1367), .Y(n_1410) );
NAND2xp5_ASAP7_75t_L g1367 ( .A(n_1368), .B(n_1389), .Y(n_1367) );
INVxp67_ASAP7_75t_L g1368 ( .A(n_1369), .Y(n_1368) );
NAND2xp5_ASAP7_75t_L g1369 ( .A(n_1370), .B(n_1387), .Y(n_1369) );
INVxp67_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
INVx2_ASAP7_75t_L g1379 ( .A(n_1380), .Y(n_1379) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
NAND2xp5_ASAP7_75t_L g1390 ( .A(n_1391), .B(n_1394), .Y(n_1390) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1407), .Y(n_1406) );
INVx2_ASAP7_75t_SL g1411 ( .A(n_1412), .Y(n_1411) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1413), .Y(n_1412) );
OAI21xp5_ASAP7_75t_L g1413 ( .A1(n_1414), .A2(n_1415), .B(n_1416), .Y(n_1413) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
endmodule