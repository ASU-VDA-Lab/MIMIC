module real_jpeg_983_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx2_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_1),
.A2(n_59),
.B1(n_60),
.B2(n_71),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_1),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_1),
.A2(n_34),
.B1(n_35),
.B2(n_71),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_71),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_1),
.A2(n_49),
.B1(n_50),
.B2(n_71),
.Y(n_180)
);

BUFx4f_ASAP7_75t_L g87 ( 
.A(n_2),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_3),
.A2(n_59),
.B1(n_60),
.B2(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_3),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_136),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_3),
.A2(n_34),
.B1(n_35),
.B2(n_136),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_3),
.A2(n_49),
.B1(n_50),
.B2(n_136),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_4),
.B(n_165),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_4),
.B(n_28),
.C(n_30),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_4),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_4),
.B(n_27),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_4),
.B(n_46),
.C(n_49),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_200),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_4),
.B(n_87),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_4),
.B(n_52),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_200),
.Y(n_265)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_6),
.A2(n_59),
.B1(n_60),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_6),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_6),
.A2(n_34),
.B1(n_35),
.B2(n_97),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_97),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_6),
.A2(n_49),
.B1(n_50),
.B2(n_97),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_7),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_38),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_7),
.A2(n_38),
.B1(n_59),
.B2(n_60),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_7),
.A2(n_38),
.B1(n_49),
.B2(n_50),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_12),
.A2(n_59),
.B1(n_60),
.B2(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_12),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_12),
.A2(n_34),
.B1(n_35),
.B2(n_164),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_164),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_12),
.A2(n_49),
.B1(n_50),
.B2(n_164),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_14),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_14),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_14),
.A2(n_34),
.B1(n_35),
.B2(n_62),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_62),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_14),
.A2(n_49),
.B1(n_50),
.B2(n_62),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_15),
.A2(n_49),
.B1(n_50),
.B2(n_55),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_15),
.A2(n_34),
.B1(n_35),
.B2(n_55),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_16),
.A2(n_34),
.B1(n_35),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_16),
.A2(n_29),
.B1(n_30),
.B2(n_41),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_16),
.A2(n_41),
.B1(n_49),
.B2(n_50),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_111),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_109),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_98),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_20),
.B(n_98),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_73),
.C(n_79),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_21),
.B(n_73),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_56),
.B1(n_57),
.B2(n_72),
.Y(n_21)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_42),
.B2(n_43),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_SL g108 ( 
.A(n_23),
.B(n_43),
.C(n_57),
.Y(n_108)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_25),
.A2(n_37),
.B1(n_39),
.B2(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_25),
.A2(n_39),
.B1(n_40),
.B2(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_25),
.A2(n_39),
.B1(n_75),
.B2(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_25),
.A2(n_39),
.B1(n_173),
.B2(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_25),
.A2(n_265),
.B(n_266),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_25),
.A2(n_204),
.B(n_266),
.Y(n_284)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_26),
.B(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_33),
.Y(n_26)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_27),
.B(n_161),
.Y(n_266)
);

AO22x2_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_27)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_L g45 ( 
.A1(n_29),
.A2(n_30),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_30),
.B(n_239),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_34),
.A2(n_35),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_34),
.B(n_190),
.Y(n_189)
);

NAND2xp33_ASAP7_75t_SL g214 ( 
.A(n_34),
.B(n_67),
.Y(n_214)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI32xp33_ASAP7_75t_L g212 ( 
.A1(n_35),
.A2(n_60),
.A3(n_66),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_39),
.A2(n_132),
.B(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_39),
.A2(n_160),
.B(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_42),
.A2(n_43),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_52),
.B(n_53),
.Y(n_43)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_44),
.A2(n_52),
.B1(n_92),
.B2(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_44),
.A2(n_52),
.B1(n_130),
.B2(n_155),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_44),
.A2(n_182),
.B(n_184),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_44),
.B(n_186),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_48),
.Y(n_44)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_48),
.A2(n_54),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_48),
.A2(n_77),
.B1(n_78),
.B2(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_48),
.A2(n_206),
.B(n_207),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_48),
.A2(n_207),
.B(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_48),
.A2(n_77),
.B1(n_183),
.B2(n_233),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_49),
.B(n_246),
.Y(n_245)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_52),
.B(n_186),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_56),
.A2(n_57),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_63),
.B1(n_65),
.B2(n_70),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_58),
.A2(n_65),
.B(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_59),
.A2(n_60),
.B1(n_66),
.B2(n_67),
.Y(n_69)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_60),
.A2(n_63),
.B(n_200),
.C(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_60),
.B(n_200),
.Y(n_201)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_63),
.A2(n_65),
.B1(n_70),
.B2(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_63),
.A2(n_134),
.B(n_137),
.Y(n_133)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_64),
.A2(n_135),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_69),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_65),
.B(n_96),
.Y(n_138)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_65),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_65),
.A2(n_94),
.B(n_286),
.Y(n_285)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_73),
.A2(n_74),
.B(n_76),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_76),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_77),
.A2(n_185),
.B(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_83),
.B(n_93),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_80),
.A2(n_81),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_90),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_82),
.A2(n_83),
.B1(n_93),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_82),
.A2(n_83),
.B1(n_90),
.B2(n_150),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_87),
.B(n_88),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_84),
.A2(n_87),
.B1(n_127),
.B2(n_157),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_84),
.A2(n_200),
.B(n_227),
.Y(n_247)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_85),
.A2(n_86),
.B1(n_89),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_85),
.A2(n_86),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_85),
.B(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_85),
.A2(n_86),
.B1(n_180),
.B2(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_85),
.A2(n_225),
.B(n_226),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_85),
.A2(n_86),
.B1(n_225),
.B2(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_86),
.A2(n_179),
.B(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_86),
.B(n_194),
.Y(n_227)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_87),
.A2(n_193),
.B(n_250),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_90),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_93),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_108),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_139),
.B(n_314),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_113),
.B(n_115),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_121),
.C(n_122),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_117),
.B1(n_121),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_131),
.C(n_133),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_124),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_125),
.A2(n_128),
.B1(n_129),
.B2(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_125),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_131),
.B(n_133),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_138),
.B(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

AO21x1_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_166),
.B(n_313),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_145),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_142),
.B(n_145),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_149),
.C(n_151),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_146),
.B(n_149),
.Y(n_311)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_151),
.B(n_311),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_158),
.C(n_162),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_152),
.A2(n_153),
.B1(n_301),
.B2(n_303),
.Y(n_300)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_154),
.B(n_156),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_155),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_157),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_158),
.A2(n_159),
.B1(n_162),
.B2(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_162),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_163),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_308),
.B(n_312),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_277),
.B(n_305),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_219),
.B(n_276),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_195),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_170),
.B(n_195),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_181),
.C(n_187),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_171),
.B(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_172),
.B(n_175),
.C(n_178),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_181),
.B(n_187),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_188),
.A2(n_189),
.B1(n_191),
.B2(n_269),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_191),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_209),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_196),
.B(n_210),
.C(n_218),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_202),
.B2(n_208),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_197),
.B(n_203),
.C(n_205),
.Y(n_290)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_201),
.Y(n_213)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_202),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_218),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_215),
.B2(n_216),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_211),
.B(n_216),
.Y(n_281)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_271),
.B(n_275),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_260),
.B(n_270),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_242),
.B(n_259),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_236),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_223),
.B(n_236),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_228),
.B1(n_234),
.B2(n_235),
.Y(n_223)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_224),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_228),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_231),
.C(n_234),
.Y(n_261)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_240),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_237),
.A2(n_238),
.B1(n_240),
.B2(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_253),
.B(n_258),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_248),
.B(n_252),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_251),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_250),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_256),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_262),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_268),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_267),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_267),
.C(n_268),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_272),
.B(n_274),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_292),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_291),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_279),
.B(n_291),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_288),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_289),
.C(n_290),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_283),
.C(n_287),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_285),
.B2(n_287),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_285),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_292),
.A2(n_306),
.B(n_307),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_304),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_304),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_296),
.B2(n_297),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_298),
.C(n_300),
.Y(n_309)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_300),
.Y(n_297)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_301),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_309),
.B(n_310),
.Y(n_312)
);


endmodule