module fake_jpeg_10991_n_67 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_67);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_67;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_32;
wire n_66;

INVx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_15),
.B(n_4),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_35),
.Y(n_44)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_32),
.A2(n_27),
.B1(n_29),
.B2(n_23),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_40),
.B1(n_0),
.B2(n_1),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_27),
.B(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_25),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_23),
.B1(n_25),
.B2(n_28),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_47),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_10),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_50),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_1),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_2),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_58),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_46),
.A2(n_42),
.B1(n_5),
.B2(n_3),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_57),
.Y(n_61)
);

MAJx2_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_49),
.C(n_9),
.Y(n_57)
);

FAx1_ASAP7_75t_SL g58 ( 
.A(n_47),
.B(n_8),
.CI(n_12),
.CON(n_58),
.SN(n_58)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_14),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_62),
.C(n_57),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_52),
.A2(n_42),
.B(n_18),
.Y(n_62)
);

NAND5xp2_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_59),
.C(n_58),
.D(n_61),
.E(n_53),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_64),
.A2(n_59),
.B(n_54),
.Y(n_65)
);

AOI211xp5_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_16),
.B(n_19),
.C(n_21),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_22),
.Y(n_67)
);


endmodule