module fake_aes_399_n_13 (n_1, n_2, n_0, n_13);
input n_1;
input n_2;
input n_0;
output n_13;
wire n_11;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx2_ASAP7_75t_L g3 ( .A(n_2), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_0), .Y(n_4) );
INVx2_ASAP7_75t_L g5 ( .A(n_1), .Y(n_5) );
OAI21xp5_ASAP7_75t_L g6 ( .A1(n_4), .A2(n_0), .B(n_2), .Y(n_6) );
CKINVDCx5p33_ASAP7_75t_R g7 ( .A(n_3), .Y(n_7) );
NAND2xp5_ASAP7_75t_L g8 ( .A(n_7), .B(n_5), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_8), .Y(n_9) );
NAND3xp33_ASAP7_75t_SL g10 ( .A(n_9), .B(n_6), .C(n_0), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_10), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_11), .Y(n_12) );
INVxp67_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
endmodule