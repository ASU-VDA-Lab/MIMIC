module fake_jpeg_4726_n_93 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_93);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_93;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_8),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_20),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_23),
.Y(n_28)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_23),
.A2(n_12),
.B1(n_16),
.B2(n_15),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

NAND2xp33_ASAP7_75t_SL g29 ( 
.A(n_19),
.B(n_13),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_28),
.Y(n_40)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_34),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_21),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_33),
.B(n_28),
.Y(n_43)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_30),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_40),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_22),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_26),
.Y(n_45)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

OAI22x1_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_29),
.B1(n_28),
.B2(n_30),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_49),
.B1(n_22),
.B2(n_23),
.Y(n_57)
);

OAI32xp33_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_31),
.A3(n_28),
.B1(n_19),
.B2(n_21),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_19),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_19),
.B(n_39),
.C(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_51),
.B(n_23),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_52),
.B(n_50),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_58),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_57),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_54),
.B(n_14),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_70)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_9),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_47),
.C(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_25),
.Y(n_64)
);

AOI322xp5_ASAP7_75t_L g72 ( 
.A1(n_64),
.A2(n_18),
.A3(n_17),
.B1(n_11),
.B2(n_16),
.C1(n_15),
.C2(n_13),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_71),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_25),
.C(n_20),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_10),
.C(n_1),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_63),
.A2(n_20),
.B1(n_18),
.B2(n_17),
.Y(n_71)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_67),
.A2(n_55),
.B1(n_20),
.B2(n_11),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_69),
.B1(n_71),
.B2(n_70),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_10),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_10),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_66),
.C(n_1),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_78),
.A2(n_76),
.B1(n_77),
.B2(n_73),
.Y(n_82)
);

MAJx2_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_74),
.C(n_68),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_79),
.A2(n_8),
.B1(n_7),
.B2(n_6),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_0),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_0),
.C(n_2),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_82),
.B(n_85),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_84),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_84),
.A2(n_79),
.B(n_3),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_2),
.Y(n_90)
);

AO21x1_ASAP7_75t_L g89 ( 
.A1(n_88),
.A2(n_2),
.B(n_3),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_89),
.A2(n_90),
.B(n_3),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_87),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_4),
.Y(n_93)
);


endmodule