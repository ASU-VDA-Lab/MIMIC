module fake_aes_6895_n_28 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_28);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_28;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_7), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_9), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_3), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_11), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_0), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_1), .Y(n_17) );
OAI22xp5_ASAP7_75t_L g18 ( .A1(n_16), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_18) );
AOI22xp33_ASAP7_75t_L g19 ( .A1(n_13), .A2(n_2), .B1(n_4), .B2(n_5), .Y(n_19) );
HB1xp67_ASAP7_75t_L g20 ( .A(n_18), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_20), .B(n_17), .Y(n_21) );
INVx1_ASAP7_75t_SL g22 ( .A(n_21), .Y(n_22) );
NOR4xp25_ASAP7_75t_L g23 ( .A(n_22), .B(n_19), .C(n_13), .D(n_12), .Y(n_23) );
INVx1_ASAP7_75t_SL g24 ( .A(n_23), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
OAI22xp5_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_14), .B1(n_15), .B2(n_10), .Y(n_26) );
NAND2x1_ASAP7_75t_L g27 ( .A(n_25), .B(n_6), .Y(n_27) );
AOI22xp33_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_24), .B1(n_27), .B2(n_8), .Y(n_28) );
endmodule