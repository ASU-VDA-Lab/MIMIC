module fake_aes_12476_n_30 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_30);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_2), .Y(n_13) );
BUFx2_ASAP7_75t_L g14 ( .A(n_1), .Y(n_14) );
NAND2xp33_ASAP7_75t_R g15 ( .A(n_1), .B(n_3), .Y(n_15) );
NAND2xp5_ASAP7_75t_SL g16 ( .A(n_4), .B(n_8), .Y(n_16) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_9), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_7), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_14), .Y(n_19) );
NOR3xp33_ASAP7_75t_SL g20 ( .A(n_15), .B(n_0), .C(n_2), .Y(n_20) );
AOI22xp33_ASAP7_75t_L g21 ( .A1(n_19), .A2(n_14), .B1(n_13), .B2(n_16), .Y(n_21) );
INVx5_ASAP7_75t_L g22 ( .A(n_20), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_22), .B(n_18), .Y(n_23) );
INVx4_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
AOI31xp33_ASAP7_75t_SL g25 ( .A1(n_24), .A2(n_15), .A3(n_21), .B(n_17), .Y(n_25) );
AOI221xp5_ASAP7_75t_SL g26 ( .A1(n_25), .A2(n_22), .B1(n_24), .B2(n_4), .C(n_5), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
AOI22xp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_22), .B1(n_3), .B2(n_5), .Y(n_28) );
NOR3x2_ASAP7_75t_L g29 ( .A(n_28), .B(n_26), .C(n_27), .Y(n_29) );
AOI322xp5_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_0), .A3(n_6), .B1(n_10), .B2(n_11), .C1(n_12), .C2(n_27), .Y(n_30) );
endmodule