module fake_netlist_5_1633_n_1668 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1668);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1668;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1538;
wire n_272;
wire n_1162;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_72),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_88),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_100),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_13),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_14),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_5),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_86),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_31),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_81),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_55),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_71),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_102),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_27),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_47),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_31),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_155),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_60),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_123),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_25),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_121),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_110),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_34),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_61),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_14),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_120),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_136),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_51),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_85),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_39),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_10),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_51),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_91),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_132),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_153),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_2),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_39),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_145),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_64),
.Y(n_195)
);

INVx4_ASAP7_75t_R g196 ( 
.A(n_130),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_83),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_108),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_7),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_80),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_26),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_45),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_3),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_139),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_131),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_79),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_97),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_4),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_76),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_33),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_10),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_89),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_128),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_96),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_129),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_48),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_45),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_54),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_113),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_66),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_65),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_68),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_11),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_23),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_47),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_105),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_32),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_92),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_41),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_119),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_107),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_134),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_34),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_82),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_122),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_50),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_117),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_30),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_150),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_74),
.Y(n_240)
);

BUFx5_ASAP7_75t_L g241 ( 
.A(n_26),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_1),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_78),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_0),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_125),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_138),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_149),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_103),
.Y(n_248)
);

BUFx4f_ASAP7_75t_SL g249 ( 
.A(n_152),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_21),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_75),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_142),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_8),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_106),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_50),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_126),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_3),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_9),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_7),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_57),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_15),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_6),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_147),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_151),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_146),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_19),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_143),
.Y(n_267)
);

BUFx8_ASAP7_75t_SL g268 ( 
.A(n_17),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_133),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_99),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_109),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_84),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_11),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_154),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_90),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_44),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_32),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_29),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_41),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_93),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_17),
.Y(n_281)
);

BUFx2_ASAP7_75t_SL g282 ( 
.A(n_104),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_16),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_2),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_59),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_53),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_42),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_25),
.Y(n_288)
);

BUFx10_ASAP7_75t_L g289 ( 
.A(n_48),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_67),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_111),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_21),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_112),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_15),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_49),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_98),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_5),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_8),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_114),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_29),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_94),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_37),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_135),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_12),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_141),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_101),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_241),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_180),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_268),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_241),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_241),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_241),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_191),
.B(n_4),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_158),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_241),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_241),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_162),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_171),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_280),
.B(n_6),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_180),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_165),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_168),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_190),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_194),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_198),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_191),
.B(n_9),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_168),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_168),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_168),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_189),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_212),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_214),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_213),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_187),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_200),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_187),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_218),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_219),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_221),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_167),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_222),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_214),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_187),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_230),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_187),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_171),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_223),
.B(n_12),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_224),
.Y(n_348)
);

NOR2xp67_ASAP7_75t_L g349 ( 
.A(n_226),
.B(n_13),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_224),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_231),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_235),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_224),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_239),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_252),
.B(n_18),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_224),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_225),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_225),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_225),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_246),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_247),
.Y(n_361)
);

NOR2xp67_ASAP7_75t_L g362 ( 
.A(n_226),
.B(n_18),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_254),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_226),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_252),
.B(n_19),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_232),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_225),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_163),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_205),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_200),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_223),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_163),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_292),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_289),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_260),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_250),
.B(n_20),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_206),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_274),
.B(n_20),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_206),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_274),
.B(n_22),
.Y(n_380)
);

NOR2xp67_ASAP7_75t_L g381 ( 
.A(n_217),
.B(n_22),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_243),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_217),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_227),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_256),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_314),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_340),
.B(n_209),
.Y(n_387)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_307),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_318),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_317),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_346),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_371),
.B(n_292),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_322),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_374),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_321),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_322),
.Y(n_396)
);

OAI21x1_ASAP7_75t_L g397 ( 
.A1(n_307),
.A2(n_204),
.B(n_195),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_327),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_327),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_328),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_328),
.Y(n_401)
);

INVx4_ASAP7_75t_L g402 ( 
.A(n_382),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_329),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_382),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_323),
.B(n_195),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_334),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_382),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_334),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_324),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_308),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_320),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_336),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_336),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_343),
.Y(n_414)
);

BUFx8_ASAP7_75t_L g415 ( 
.A(n_347),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_343),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_345),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_325),
.B(n_204),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_382),
.Y(n_419)
);

AND3x2_ASAP7_75t_L g420 ( 
.A(n_319),
.B(n_283),
.C(n_227),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_331),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_364),
.B(n_207),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_310),
.Y(n_423)
);

BUFx6f_ASAP7_75t_SL g424 ( 
.A(n_345),
.Y(n_424)
);

AND2x6_ASAP7_75t_L g425 ( 
.A(n_347),
.B(n_243),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_333),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_348),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_337),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_349),
.B(n_207),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_348),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_310),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_350),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_330),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_338),
.B(n_290),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_311),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_350),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_353),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_353),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_356),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_311),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_312),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_356),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_357),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_339),
.B(n_237),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_357),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_312),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_358),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_358),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_341),
.B(n_290),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_344),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_315),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_359),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_359),
.Y(n_453)
);

CKINVDCx8_ASAP7_75t_R g454 ( 
.A(n_340),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_351),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_352),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_354),
.Y(n_457)
);

BUFx12f_ASAP7_75t_L g458 ( 
.A(n_309),
.Y(n_458)
);

OR2x6_ASAP7_75t_L g459 ( 
.A(n_450),
.B(n_458),
.Y(n_459)
);

AND2x6_ASAP7_75t_L g460 ( 
.A(n_422),
.B(n_293),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_422),
.B(n_373),
.Y(n_461)
);

AND2x2_ASAP7_75t_SL g462 ( 
.A(n_429),
.B(n_313),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_444),
.B(n_360),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_388),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_405),
.B(n_361),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_389),
.B(n_366),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_392),
.B(n_332),
.Y(n_467)
);

OR2x6_ASAP7_75t_L g468 ( 
.A(n_450),
.B(n_282),
.Y(n_468)
);

AND2x6_ASAP7_75t_L g469 ( 
.A(n_422),
.B(n_293),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_392),
.B(n_342),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_422),
.B(n_368),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_418),
.B(n_434),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_431),
.Y(n_473)
);

NAND2xp33_ASAP7_75t_L g474 ( 
.A(n_425),
.B(n_200),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_449),
.B(n_363),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_410),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_388),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_388),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_411),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_423),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_391),
.B(n_385),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_435),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g483 ( 
.A1(n_429),
.A2(n_326),
.B1(n_355),
.B2(n_380),
.Y(n_483)
);

BUFx10_ASAP7_75t_L g484 ( 
.A(n_386),
.Y(n_484)
);

OR2x6_ASAP7_75t_L g485 ( 
.A(n_458),
.B(n_362),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_435),
.Y(n_486)
);

AND2x4_ASAP7_75t_L g487 ( 
.A(n_429),
.B(n_367),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_390),
.B(n_366),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_431),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_395),
.B(n_375),
.Y(n_490)
);

AND2x6_ASAP7_75t_L g491 ( 
.A(n_429),
.B(n_243),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_435),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_431),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g494 ( 
.A(n_394),
.B(n_375),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_394),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_435),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_L g497 ( 
.A1(n_425),
.A2(n_365),
.B1(n_378),
.B2(n_381),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_402),
.B(n_367),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_440),
.Y(n_499)
);

INVx4_ASAP7_75t_L g500 ( 
.A(n_431),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_393),
.B(n_368),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_425),
.A2(n_381),
.B1(n_193),
.B2(n_253),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_388),
.Y(n_503)
);

BUFx8_ASAP7_75t_SL g504 ( 
.A(n_433),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_427),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_427),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_440),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_440),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_420),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_441),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_431),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_387),
.B(n_376),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_441),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_425),
.A2(n_176),
.B1(n_181),
.B2(n_169),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_442),
.Y(n_515)
);

AO22x2_ASAP7_75t_L g516 ( 
.A1(n_441),
.A2(n_259),
.B1(n_199),
.B2(n_201),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_431),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_446),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_446),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_442),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_397),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_446),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_451),
.Y(n_523)
);

INVxp33_ASAP7_75t_L g524 ( 
.A(n_421),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_454),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_407),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_425),
.A2(n_261),
.B1(n_202),
.B2(n_203),
.Y(n_527)
);

OAI22xp33_ASAP7_75t_L g528 ( 
.A1(n_409),
.A2(n_186),
.B1(n_188),
.B2(n_184),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_407),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_415),
.Y(n_530)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_457),
.B(n_376),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_397),
.B(n_372),
.Y(n_532)
);

AND2x2_ASAP7_75t_SL g533 ( 
.A(n_402),
.B(n_243),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_451),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_419),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_451),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_415),
.B(n_303),
.Y(n_537)
);

INVx6_ASAP7_75t_L g538 ( 
.A(n_415),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_415),
.B(n_303),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_451),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_451),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_402),
.B(n_315),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_425),
.B(n_316),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_393),
.B(n_372),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_425),
.B(n_316),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_451),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_404),
.Y(n_547)
);

INVxp67_ASAP7_75t_SL g548 ( 
.A(n_404),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_419),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_404),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_396),
.Y(n_551)
);

AND2x6_ASAP7_75t_L g552 ( 
.A(n_404),
.B(n_303),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_398),
.Y(n_553)
);

NAND3x1_ASAP7_75t_L g554 ( 
.A(n_454),
.B(n_208),
.C(n_161),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_399),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_399),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_400),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_400),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_401),
.B(n_267),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_401),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_426),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_424),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_428),
.B(n_303),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_403),
.B(n_285),
.Y(n_564)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_424),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_403),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_406),
.B(n_383),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_408),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_408),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_412),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_412),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_413),
.Y(n_572)
);

OR2x6_ASAP7_75t_L g573 ( 
.A(n_413),
.B(n_210),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_414),
.Y(n_574)
);

OR2x6_ASAP7_75t_L g575 ( 
.A(n_414),
.B(n_233),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_416),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_455),
.B(n_164),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_416),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_417),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_417),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_430),
.B(n_301),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_456),
.B(n_166),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_430),
.B(n_264),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_432),
.B(n_170),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_432),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_424),
.A2(n_270),
.B1(n_220),
.B2(n_215),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_436),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_436),
.B(n_269),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_437),
.B(n_369),
.Y(n_589)
);

BUFx6f_ASAP7_75t_SL g590 ( 
.A(n_437),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_438),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_438),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_439),
.B(n_271),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_443),
.B(n_172),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_443),
.B(n_272),
.Y(n_595)
);

OAI22xp33_ASAP7_75t_L g596 ( 
.A1(n_445),
.A2(n_216),
.B1(n_262),
.B2(n_244),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_445),
.B(n_377),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_471),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g599 ( 
.A1(n_483),
.A2(n_234),
.B1(n_209),
.B2(n_215),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_465),
.B(n_447),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_463),
.B(n_448),
.Y(n_601)
);

AO22x1_ASAP7_75t_L g602 ( 
.A1(n_509),
.A2(n_179),
.B1(n_300),
.B2(n_304),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_462),
.A2(n_220),
.B1(n_234),
.B2(n_305),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_533),
.B(n_200),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_461),
.B(n_452),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_461),
.B(n_452),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_471),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_467),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_460),
.A2(n_469),
.B1(n_462),
.B2(n_532),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_467),
.B(n_379),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_532),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_487),
.B(n_185),
.Y(n_612)
);

NAND2xp33_ASAP7_75t_L g613 ( 
.A(n_460),
.B(n_200),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_501),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_460),
.A2(n_469),
.B1(n_532),
.B2(n_470),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_470),
.B(n_453),
.Y(n_616)
);

OR2x6_ASAP7_75t_L g617 ( 
.A(n_538),
.B(n_197),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_475),
.B(n_248),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_533),
.B(n_548),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_547),
.B(n_200),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_481),
.B(n_577),
.Y(n_621)
);

AND2x2_ASAP7_75t_SL g622 ( 
.A(n_474),
.B(n_240),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_501),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_556),
.B(n_453),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_547),
.B(n_200),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_577),
.B(n_248),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_556),
.B(n_245),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_555),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_547),
.B(n_251),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_582),
.B(n_270),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_504),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_556),
.B(n_263),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_543),
.B(n_265),
.Y(n_633)
);

INVxp67_ASAP7_75t_SL g634 ( 
.A(n_489),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_495),
.B(n_289),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_570),
.B(n_275),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_551),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_460),
.A2(n_296),
.B1(n_306),
.B2(n_424),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_555),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_551),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_544),
.B(n_567),
.Y(n_641)
);

NOR3xp33_ASAP7_75t_L g642 ( 
.A(n_586),
.B(n_597),
.C(n_589),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_566),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_566),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_545),
.B(n_299),
.Y(n_645)
);

INVxp67_ASAP7_75t_L g646 ( 
.A(n_494),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_571),
.B(n_291),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_487),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_576),
.B(n_156),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_460),
.A2(n_335),
.B1(n_370),
.B2(n_257),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_572),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_572),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_582),
.B(n_299),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_489),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_542),
.B(n_305),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_576),
.B(n_156),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_544),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_553),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_567),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_576),
.B(n_157),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_574),
.B(n_157),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_574),
.B(n_550),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_580),
.B(n_173),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_580),
.B(n_173),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_580),
.B(n_174),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_574),
.B(n_174),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_573),
.B(n_383),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_487),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_560),
.B(n_175),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_553),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_574),
.B(n_175),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_557),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_578),
.B(n_177),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_587),
.B(n_178),
.Y(n_674)
);

NAND2xp33_ASAP7_75t_L g675 ( 
.A(n_460),
.B(n_178),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_591),
.B(n_182),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_592),
.B(n_182),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_480),
.B(n_183),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_573),
.B(n_384),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_482),
.B(n_486),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_466),
.B(n_304),
.Y(n_681)
);

NOR3xp33_ASAP7_75t_L g682 ( 
.A(n_528),
.B(n_531),
.C(n_509),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_469),
.A2(n_497),
.B1(n_516),
.B2(n_521),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_573),
.B(n_255),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_573),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_492),
.B(n_183),
.Y(n_686)
);

NAND3xp33_ASAP7_75t_L g687 ( 
.A(n_563),
.B(n_160),
.C(n_159),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_496),
.B(n_469),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_558),
.Y(n_689)
);

NAND2xp33_ASAP7_75t_L g690 ( 
.A(n_469),
.B(n_228),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_558),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_575),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_469),
.B(n_249),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_512),
.B(n_179),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_521),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_478),
.B(n_192),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_575),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_498),
.B(n_211),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_568),
.B(n_569),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_569),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_538),
.Y(n_701)
);

AND2x2_ASAP7_75t_SL g702 ( 
.A(n_474),
.B(n_302),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_562),
.B(n_242),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_579),
.B(n_229),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_579),
.B(n_236),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_585),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_505),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_583),
.B(n_238),
.Y(n_708)
);

BUFx12f_ASAP7_75t_L g709 ( 
.A(n_484),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_505),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_588),
.B(n_281),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_562),
.B(n_565),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_593),
.B(n_284),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_506),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_595),
.B(n_258),
.Y(n_715)
);

A2O1A1Ixp33_ASAP7_75t_L g716 ( 
.A1(n_537),
.A2(n_288),
.B(n_298),
.C(n_278),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_511),
.B(n_266),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_563),
.B(n_297),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_506),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_515),
.Y(n_720)
);

INVx4_ASAP7_75t_L g721 ( 
.A(n_489),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_511),
.B(n_273),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_562),
.B(n_287),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_516),
.A2(n_279),
.B1(n_295),
.B2(n_300),
.Y(n_724)
);

OAI221xp5_ASAP7_75t_L g725 ( 
.A1(n_575),
.A2(n_294),
.B1(n_277),
.B2(n_276),
.C(n_196),
.Y(n_725)
);

AND2x2_ASAP7_75t_SL g726 ( 
.A(n_502),
.B(n_250),
.Y(n_726)
);

NOR2xp67_ASAP7_75t_L g727 ( 
.A(n_561),
.B(n_58),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_565),
.B(n_289),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_515),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_524),
.B(n_488),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_489),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_520),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_511),
.B(n_56),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_565),
.B(n_286),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_523),
.B(n_140),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_537),
.B(n_539),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_L g737 ( 
.A1(n_468),
.A2(n_137),
.B1(n_127),
.B2(n_124),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_526),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_523),
.B(n_534),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_575),
.B(n_118),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_524),
.B(n_23),
.Y(n_741)
);

NOR2x1p5_ASAP7_75t_L g742 ( 
.A(n_559),
.B(n_24),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_523),
.B(n_116),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_709),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_600),
.B(n_564),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_611),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_SL g747 ( 
.A(n_709),
.B(n_484),
.Y(n_747)
);

A2O1A1Ixp33_ASAP7_75t_L g748 ( 
.A1(n_621),
.A2(n_530),
.B(n_490),
.C(n_581),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_631),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_601),
.B(n_534),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_611),
.A2(n_473),
.B(n_500),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_648),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_626),
.A2(n_468),
.B1(n_590),
.B2(n_530),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_648),
.Y(n_754)
);

OAI21xp5_ASAP7_75t_L g755 ( 
.A1(n_619),
.A2(n_536),
.B(n_540),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_630),
.A2(n_468),
.B1(n_590),
.B2(n_538),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_613),
.A2(n_609),
.B(n_615),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_618),
.B(n_476),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_653),
.A2(n_468),
.B1(n_590),
.B2(n_525),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_599),
.B(n_484),
.Y(n_760)
);

HB1xp67_ASAP7_75t_L g761 ( 
.A(n_610),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_613),
.A2(n_473),
.B(n_500),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_608),
.A2(n_554),
.B1(n_546),
.B2(n_541),
.Y(n_763)
);

O2A1O1Ixp5_ASAP7_75t_L g764 ( 
.A1(n_736),
.A2(n_594),
.B(n_584),
.C(n_541),
.Y(n_764)
);

OAI21xp5_ASAP7_75t_L g765 ( 
.A1(n_604),
.A2(n_508),
.B(n_518),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_646),
.B(n_479),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_641),
.B(n_596),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_730),
.B(n_479),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_616),
.B(n_513),
.Y(n_769)
);

O2A1O1Ixp33_ASAP7_75t_SL g770 ( 
.A1(n_604),
.A2(n_510),
.B(n_507),
.C(n_519),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_637),
.Y(n_771)
);

BUFx12f_ASAP7_75t_L g772 ( 
.A(n_742),
.Y(n_772)
);

OAI21xp5_ASAP7_75t_L g773 ( 
.A1(n_688),
.A2(n_522),
.B(n_499),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_605),
.A2(n_493),
.B(n_517),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_606),
.A2(n_493),
.B(n_517),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_603),
.B(n_485),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_699),
.A2(n_503),
.B(n_464),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_683),
.A2(n_503),
.B(n_464),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_637),
.Y(n_779)
);

AND2x2_ASAP7_75t_SL g780 ( 
.A(n_726),
.B(n_514),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_719),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_641),
.B(n_517),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_598),
.B(n_516),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_607),
.B(n_614),
.Y(n_784)
);

AOI21x1_ASAP7_75t_L g785 ( 
.A1(n_662),
.A2(n_477),
.B(n_549),
.Y(n_785)
);

OAI22xp5_ASAP7_75t_L g786 ( 
.A1(n_702),
.A2(n_527),
.B1(n_554),
.B2(n_485),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_623),
.B(n_477),
.Y(n_787)
);

OAI21x1_ASAP7_75t_L g788 ( 
.A1(n_739),
.A2(n_526),
.B(n_549),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_640),
.Y(n_789)
);

O2A1O1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_645),
.A2(n_529),
.B(n_535),
.C(n_485),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_622),
.A2(n_517),
.B(n_493),
.Y(n_791)
);

O2A1O1Ixp33_ASAP7_75t_L g792 ( 
.A1(n_645),
.A2(n_529),
.B(n_459),
.C(n_491),
.Y(n_792)
);

OAI21xp5_ASAP7_75t_L g793 ( 
.A1(n_622),
.A2(n_491),
.B(n_552),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_702),
.A2(n_493),
.B(n_491),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_620),
.A2(n_491),
.B(n_459),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_658),
.Y(n_796)
);

BUFx4f_ASAP7_75t_L g797 ( 
.A(n_617),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_698),
.B(n_552),
.Y(n_798)
);

A2O1A1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_718),
.A2(n_27),
.B(n_28),
.C(n_33),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_635),
.B(n_35),
.Y(n_800)
);

BUFx2_ASAP7_75t_L g801 ( 
.A(n_740),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_729),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_657),
.B(n_35),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_670),
.Y(n_804)
);

OAI21xp5_ASAP7_75t_L g805 ( 
.A1(n_680),
.A2(n_115),
.B(n_95),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_659),
.B(n_36),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_727),
.B(n_87),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_L g808 ( 
.A1(n_695),
.A2(n_77),
.B1(n_73),
.B2(n_70),
.Y(n_808)
);

AOI22xp5_ASAP7_75t_L g809 ( 
.A1(n_682),
.A2(n_69),
.B1(n_63),
.B2(n_62),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_708),
.B(n_37),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_734),
.B(n_38),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_734),
.B(n_38),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_711),
.B(n_40),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_672),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_667),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_713),
.B(n_43),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_715),
.B(n_628),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_625),
.A2(n_46),
.B(n_49),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_695),
.A2(n_52),
.B1(n_53),
.B2(n_726),
.Y(n_819)
);

HB1xp67_ASAP7_75t_L g820 ( 
.A(n_667),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_650),
.A2(n_52),
.B(n_633),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_633),
.A2(n_624),
.B(n_647),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_639),
.B(n_643),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_627),
.A2(n_636),
.B(n_632),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_684),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_679),
.B(n_684),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_675),
.A2(n_690),
.B(n_717),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_679),
.B(n_681),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_644),
.B(n_651),
.Y(n_829)
);

INVxp67_ASAP7_75t_L g830 ( 
.A(n_741),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_675),
.A2(n_690),
.B(n_722),
.Y(n_831)
);

BUFx4f_ASAP7_75t_L g832 ( 
.A(n_617),
.Y(n_832)
);

A2O1A1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_668),
.A2(n_697),
.B(n_685),
.C(n_692),
.Y(n_833)
);

AOI21xp33_ASAP7_75t_L g834 ( 
.A1(n_669),
.A2(n_674),
.B(n_673),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_649),
.A2(n_665),
.B(n_664),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_SL g836 ( 
.A1(n_740),
.A2(n_725),
.B1(n_692),
.B2(n_685),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_695),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_656),
.A2(n_663),
.B(n_660),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_689),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_691),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_629),
.A2(n_696),
.B(n_634),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_652),
.B(n_700),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_701),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_706),
.B(n_612),
.Y(n_844)
);

A2O1A1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_697),
.A2(n_687),
.B(n_612),
.C(n_716),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_612),
.Y(n_846)
);

NAND3xp33_ASAP7_75t_L g847 ( 
.A(n_724),
.B(n_678),
.C(n_677),
.Y(n_847)
);

NOR3xp33_ASAP7_75t_L g848 ( 
.A(n_728),
.B(n_602),
.C(n_723),
.Y(n_848)
);

NAND3xp33_ASAP7_75t_SL g849 ( 
.A(n_728),
.B(n_716),
.C(n_723),
.Y(n_849)
);

AOI21xp33_ASAP7_75t_L g850 ( 
.A1(n_676),
.A2(n_704),
.B(n_705),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_686),
.A2(n_661),
.B(n_671),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_707),
.A2(n_710),
.B1(n_720),
.B2(n_714),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_703),
.B(n_671),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_661),
.A2(n_666),
.B(n_721),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_654),
.A2(n_721),
.B(n_712),
.Y(n_855)
);

AND2x6_ASAP7_75t_L g856 ( 
.A(n_701),
.B(n_743),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_732),
.Y(n_857)
);

AOI21x1_ASAP7_75t_L g858 ( 
.A1(n_738),
.A2(n_733),
.B(n_735),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_731),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_617),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_703),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_654),
.A2(n_721),
.B(n_712),
.Y(n_862)
);

BUFx4f_ASAP7_75t_L g863 ( 
.A(n_617),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_693),
.A2(n_638),
.B(n_731),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_731),
.B(n_737),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_610),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_648),
.Y(n_867)
);

AO21x1_ASAP7_75t_L g868 ( 
.A1(n_736),
.A2(n_621),
.B(n_604),
.Y(n_868)
);

A2O1A1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_621),
.A2(n_626),
.B(n_653),
.C(n_630),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_611),
.Y(n_870)
);

O2A1O1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_621),
.A2(n_608),
.B(n_645),
.C(n_655),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_621),
.B(n_618),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_600),
.B(n_472),
.Y(n_873)
);

INVx1_ASAP7_75t_SL g874 ( 
.A(n_610),
.Y(n_874)
);

OAI21x1_ASAP7_75t_L g875 ( 
.A1(n_688),
.A2(n_739),
.B(n_680),
.Y(n_875)
);

O2A1O1Ixp5_ASAP7_75t_L g876 ( 
.A1(n_736),
.A2(n_621),
.B(n_604),
.C(n_696),
.Y(n_876)
);

A2O1A1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_621),
.A2(n_626),
.B(n_653),
.C(n_630),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_600),
.B(n_472),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_641),
.B(n_648),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_621),
.A2(n_626),
.B1(n_653),
.B2(n_630),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_611),
.A2(n_619),
.B(n_613),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_621),
.B(n_618),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_648),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_600),
.B(n_472),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_611),
.Y(n_885)
);

NOR2xp67_ASAP7_75t_L g886 ( 
.A(n_709),
.B(n_561),
.Y(n_886)
);

BUFx3_ASAP7_75t_L g887 ( 
.A(n_709),
.Y(n_887)
);

OR2x2_ASAP7_75t_L g888 ( 
.A(n_694),
.B(n_610),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_600),
.B(n_472),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_611),
.A2(n_619),
.B(n_604),
.Y(n_890)
);

A2O1A1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_621),
.A2(n_626),
.B(n_653),
.C(n_630),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_600),
.B(n_472),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_611),
.A2(n_619),
.B(n_613),
.Y(n_893)
);

OAI22xp5_ASAP7_75t_L g894 ( 
.A1(n_621),
.A2(n_615),
.B1(n_683),
.B2(n_609),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_611),
.A2(n_619),
.B(n_613),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_610),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_746),
.Y(n_897)
);

INVx2_ASAP7_75t_SL g898 ( 
.A(n_888),
.Y(n_898)
);

AOI21x1_ASAP7_75t_L g899 ( 
.A1(n_827),
.A2(n_831),
.B(n_841),
.Y(n_899)
);

OAI21xp33_ASAP7_75t_L g900 ( 
.A1(n_872),
.A2(n_882),
.B(n_880),
.Y(n_900)
);

AOI221xp5_ASAP7_75t_SL g901 ( 
.A1(n_869),
.A2(n_877),
.B1(n_891),
.B2(n_892),
.C(n_884),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_873),
.B(n_878),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_885),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_L g904 ( 
.A1(n_889),
.A2(n_894),
.B1(n_780),
.B2(n_757),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_760),
.A2(n_853),
.B1(n_826),
.B2(n_776),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_757),
.A2(n_876),
.B(n_778),
.Y(n_906)
);

OR2x2_ASAP7_75t_L g907 ( 
.A(n_874),
.B(n_896),
.Y(n_907)
);

NAND2x1p5_ASAP7_75t_L g908 ( 
.A(n_837),
.B(n_752),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_762),
.A2(n_824),
.B(n_864),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_745),
.B(n_769),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_761),
.B(n_866),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_850),
.B(n_817),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_870),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_881),
.A2(n_895),
.B(n_893),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_893),
.A2(n_895),
.B(n_890),
.Y(n_915)
);

OAI21x1_ASAP7_75t_L g916 ( 
.A1(n_777),
.A2(n_751),
.B(n_858),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_879),
.B(n_754),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_871),
.A2(n_847),
.B(n_812),
.C(n_811),
.Y(n_918)
);

AOI21x1_ASAP7_75t_L g919 ( 
.A1(n_835),
.A2(n_838),
.B(n_791),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_830),
.B(n_758),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_773),
.A2(n_862),
.B(n_855),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_SL g922 ( 
.A1(n_845),
.A2(n_799),
.B(n_833),
.C(n_748),
.Y(n_922)
);

AND2x6_ASAP7_75t_L g923 ( 
.A(n_809),
.B(n_837),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_784),
.B(n_834),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_815),
.Y(n_925)
);

AO31x2_ASAP7_75t_L g926 ( 
.A1(n_868),
.A2(n_851),
.A3(n_822),
.B(n_854),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_828),
.B(n_750),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_837),
.Y(n_928)
);

OAI21x1_ASAP7_75t_L g929 ( 
.A1(n_751),
.A2(n_775),
.B(n_774),
.Y(n_929)
);

OAI22xp5_ASAP7_75t_L g930 ( 
.A1(n_801),
.A2(n_819),
.B1(n_865),
.B2(n_783),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_861),
.B(n_810),
.Y(n_931)
);

AO31x2_ASAP7_75t_L g932 ( 
.A1(n_794),
.A2(n_786),
.A3(n_813),
.B(n_816),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_768),
.B(n_820),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_825),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_848),
.A2(n_879),
.B1(n_849),
.B2(n_767),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_766),
.B(n_759),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_752),
.B(n_800),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_771),
.B(n_779),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_823),
.B(n_829),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_839),
.B(n_840),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_859),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_842),
.B(n_846),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_764),
.A2(n_765),
.B(n_798),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_844),
.A2(n_790),
.B(n_793),
.Y(n_944)
);

AOI21xp33_ASAP7_75t_L g945 ( 
.A1(n_792),
.A2(n_803),
.B(n_806),
.Y(n_945)
);

NAND2x1_ASAP7_75t_L g946 ( 
.A(n_859),
.B(n_802),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_857),
.B(n_787),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_782),
.A2(n_770),
.B(n_807),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_795),
.A2(n_805),
.B(n_763),
.C(n_756),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_789),
.B(n_814),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_796),
.B(n_804),
.Y(n_951)
);

NAND2x1p5_ASAP7_75t_L g952 ( 
.A(n_859),
.B(n_754),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_781),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_836),
.A2(n_821),
.B(n_852),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_797),
.A2(n_863),
.B1(n_832),
.B2(n_753),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_754),
.B(n_867),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_867),
.B(n_883),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_867),
.B(n_883),
.Y(n_958)
);

OAI21x1_ASAP7_75t_L g959 ( 
.A1(n_821),
.A2(n_808),
.B(n_818),
.Y(n_959)
);

OR2x2_ASAP7_75t_L g960 ( 
.A(n_843),
.B(n_860),
.Y(n_960)
);

OAI21x1_ASAP7_75t_L g961 ( 
.A1(n_856),
.A2(n_886),
.B(n_747),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_856),
.Y(n_962)
);

OAI21x1_ASAP7_75t_L g963 ( 
.A1(n_856),
.A2(n_744),
.B(n_887),
.Y(n_963)
);

OAI21x1_ASAP7_75t_L g964 ( 
.A1(n_856),
.A2(n_749),
.B(n_788),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_873),
.B(n_878),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_837),
.Y(n_966)
);

BUFx3_ASAP7_75t_L g967 ( 
.A(n_744),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_826),
.B(n_610),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_885),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_873),
.B(n_878),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_872),
.B(n_882),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_880),
.A2(n_869),
.B1(n_891),
.B2(n_877),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_896),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_757),
.A2(n_877),
.B(n_869),
.Y(n_974)
);

NOR2xp67_ASAP7_75t_L g975 ( 
.A(n_861),
.B(n_709),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_872),
.A2(n_882),
.B(n_869),
.C(n_877),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_872),
.A2(n_882),
.B(n_869),
.C(n_877),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_873),
.B(n_878),
.Y(n_978)
);

AOI21xp33_ASAP7_75t_L g979 ( 
.A1(n_872),
.A2(n_882),
.B(n_880),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_746),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_757),
.A2(n_877),
.B(n_869),
.Y(n_981)
);

OAI21x1_ASAP7_75t_SL g982 ( 
.A1(n_868),
.A2(n_757),
.B(n_795),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_825),
.B(n_879),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_872),
.A2(n_882),
.B(n_869),
.C(n_877),
.Y(n_984)
);

BUFx12f_ASAP7_75t_L g985 ( 
.A(n_772),
.Y(n_985)
);

AND3x4_ASAP7_75t_L g986 ( 
.A(n_749),
.B(n_682),
.C(n_642),
.Y(n_986)
);

AND2x2_ASAP7_75t_SL g987 ( 
.A(n_872),
.B(n_882),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_757),
.A2(n_877),
.B(n_869),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_SL g989 ( 
.A1(n_757),
.A2(n_894),
.B(n_877),
.Y(n_989)
);

INVx5_ASAP7_75t_L g990 ( 
.A(n_837),
.Y(n_990)
);

AOI211x1_ASAP7_75t_L g991 ( 
.A1(n_873),
.A2(n_878),
.B(n_889),
.C(n_884),
.Y(n_991)
);

OAI21x1_ASAP7_75t_L g992 ( 
.A1(n_788),
.A2(n_785),
.B(n_875),
.Y(n_992)
);

AO21x2_ASAP7_75t_L g993 ( 
.A1(n_755),
.A2(n_831),
.B(n_827),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_873),
.B(n_878),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_873),
.B(n_878),
.Y(n_995)
);

OAI21x1_ASAP7_75t_L g996 ( 
.A1(n_788),
.A2(n_785),
.B(n_875),
.Y(n_996)
);

OAI21x1_ASAP7_75t_SL g997 ( 
.A1(n_868),
.A2(n_757),
.B(n_795),
.Y(n_997)
);

INVx2_ASAP7_75t_SL g998 ( 
.A(n_888),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_826),
.B(n_610),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_873),
.B(n_878),
.Y(n_1000)
);

AO31x2_ASAP7_75t_L g1001 ( 
.A1(n_868),
.A2(n_877),
.A3(n_891),
.B(n_869),
.Y(n_1001)
);

OAI21x1_ASAP7_75t_L g1002 ( 
.A1(n_788),
.A2(n_785),
.B(n_875),
.Y(n_1002)
);

OAI21x1_ASAP7_75t_L g1003 ( 
.A1(n_788),
.A2(n_785),
.B(n_875),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_885),
.Y(n_1004)
);

INVx3_ASAP7_75t_L g1005 ( 
.A(n_837),
.Y(n_1005)
);

AOI21x1_ASAP7_75t_L g1006 ( 
.A1(n_827),
.A2(n_831),
.B(n_841),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_SL g1007 ( 
.A1(n_757),
.A2(n_894),
.B(n_877),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_872),
.A2(n_882),
.B(n_869),
.C(n_877),
.Y(n_1008)
);

OAI22x1_ASAP7_75t_L g1009 ( 
.A1(n_880),
.A2(n_760),
.B1(n_882),
.B2(n_872),
.Y(n_1009)
);

OA21x2_ASAP7_75t_L g1010 ( 
.A1(n_755),
.A2(n_773),
.B(n_876),
.Y(n_1010)
);

INVx4_ASAP7_75t_L g1011 ( 
.A(n_837),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_815),
.Y(n_1012)
);

AO221x2_ASAP7_75t_L g1013 ( 
.A1(n_819),
.A2(n_599),
.B1(n_786),
.B2(n_602),
.C(n_528),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_873),
.B(n_878),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_837),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_837),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_788),
.A2(n_785),
.B(n_875),
.Y(n_1017)
);

INVx2_ASAP7_75t_SL g1018 ( 
.A(n_888),
.Y(n_1018)
);

AOI21xp33_ASAP7_75t_L g1019 ( 
.A1(n_872),
.A2(n_882),
.B(n_880),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_921),
.A2(n_970),
.B(n_902),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_941),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_971),
.A2(n_978),
.B1(n_1014),
.B2(n_994),
.Y(n_1022)
);

HB1xp67_ASAP7_75t_L g1023 ( 
.A(n_973),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_965),
.A2(n_1000),
.B(n_995),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_940),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_965),
.A2(n_995),
.B1(n_1000),
.B2(n_910),
.Y(n_1026)
);

A2O1A1Ixp33_ASAP7_75t_SL g1027 ( 
.A1(n_974),
.A2(n_988),
.B(n_981),
.C(n_945),
.Y(n_1027)
);

INVx2_ASAP7_75t_SL g1028 ( 
.A(n_960),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_900),
.B(n_910),
.Y(n_1029)
);

INVx2_ASAP7_75t_SL g1030 ( 
.A(n_967),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_985),
.Y(n_1031)
);

INVx5_ASAP7_75t_L g1032 ( 
.A(n_966),
.Y(n_1032)
);

OR2x2_ASAP7_75t_L g1033 ( 
.A(n_907),
.B(n_911),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_903),
.Y(n_1034)
);

A2O1A1Ixp33_ASAP7_75t_SL g1035 ( 
.A1(n_974),
.A2(n_988),
.B(n_981),
.C(n_945),
.Y(n_1035)
);

BUFx10_ASAP7_75t_L g1036 ( 
.A(n_933),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_979),
.B(n_1019),
.Y(n_1037)
);

CKINVDCx20_ASAP7_75t_R g1038 ( 
.A(n_898),
.Y(n_1038)
);

INVx1_ASAP7_75t_SL g1039 ( 
.A(n_968),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_925),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_SL g1041 ( 
.A1(n_987),
.A2(n_936),
.B1(n_986),
.B2(n_1009),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_969),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_998),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1004),
.Y(n_1044)
);

BUFx3_ASAP7_75t_L g1045 ( 
.A(n_1018),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_979),
.B(n_1019),
.Y(n_1046)
);

NOR2xp67_ASAP7_75t_L g1047 ( 
.A(n_931),
.B(n_1012),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_941),
.Y(n_1048)
);

OAI22xp33_ASAP7_75t_L g1049 ( 
.A1(n_905),
.A2(n_920),
.B1(n_924),
.B2(n_912),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_976),
.A2(n_984),
.B(n_1008),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_983),
.B(n_917),
.Y(n_1051)
);

INVxp67_ASAP7_75t_L g1052 ( 
.A(n_999),
.Y(n_1052)
);

INVx2_ASAP7_75t_SL g1053 ( 
.A(n_934),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_977),
.A2(n_904),
.B1(n_972),
.B2(n_991),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_983),
.B(n_956),
.Y(n_1055)
);

OR2x6_ASAP7_75t_L g1056 ( 
.A(n_955),
.B(n_975),
.Y(n_1056)
);

INVx2_ASAP7_75t_SL g1057 ( 
.A(n_956),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_897),
.Y(n_1058)
);

INVx2_ASAP7_75t_SL g1059 ( 
.A(n_957),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_957),
.B(n_958),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_958),
.B(n_942),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_912),
.B(n_1013),
.Y(n_1062)
);

OAI21xp33_ASAP7_75t_L g1063 ( 
.A1(n_918),
.A2(n_972),
.B(n_939),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_944),
.A2(n_989),
.B(n_1007),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_927),
.B(n_937),
.Y(n_1065)
);

OAI22x1_ASAP7_75t_L g1066 ( 
.A1(n_935),
.A2(n_962),
.B1(n_908),
.B2(n_952),
.Y(n_1066)
);

INVx6_ASAP7_75t_L g1067 ( 
.A(n_990),
.Y(n_1067)
);

INVx2_ASAP7_75t_SL g1068 ( 
.A(n_966),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_904),
.A2(n_930),
.B1(n_954),
.B2(n_955),
.Y(n_1069)
);

INVx1_ASAP7_75t_SL g1070 ( 
.A(n_966),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_1015),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_938),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_947),
.B(n_930),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_901),
.B(n_1001),
.Y(n_1074)
);

OR2x6_ASAP7_75t_SL g1075 ( 
.A(n_913),
.B(n_980),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_1015),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_901),
.B(n_1001),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1001),
.B(n_951),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_915),
.A2(n_914),
.B(n_949),
.Y(n_1079)
);

NOR2x1_ASAP7_75t_SL g1080 ( 
.A(n_990),
.B(n_1016),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_953),
.B(n_932),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_941),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_993),
.A2(n_943),
.B(n_922),
.Y(n_1083)
);

AOI22xp33_ASAP7_75t_L g1084 ( 
.A1(n_954),
.A2(n_923),
.B1(n_982),
.B2(n_997),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_1015),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_SL g1086 ( 
.A1(n_906),
.A2(n_943),
.B(n_948),
.C(n_928),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_932),
.B(n_951),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_950),
.A2(n_990),
.B1(n_908),
.B2(n_952),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_946),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_1016),
.Y(n_1090)
);

BUFx3_ASAP7_75t_L g1091 ( 
.A(n_1016),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_932),
.B(n_1005),
.Y(n_1092)
);

INVxp67_ASAP7_75t_SL g1093 ( 
.A(n_928),
.Y(n_1093)
);

OR2x2_ASAP7_75t_L g1094 ( 
.A(n_1005),
.B(n_1011),
.Y(n_1094)
);

BUFx10_ASAP7_75t_L g1095 ( 
.A(n_923),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_963),
.B(n_990),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_926),
.Y(n_1097)
);

AOI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_923),
.A2(n_959),
.B1(n_1010),
.B2(n_961),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_923),
.B(n_964),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1010),
.B(n_926),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_916),
.A2(n_929),
.B(n_1017),
.Y(n_1101)
);

INVx4_ASAP7_75t_L g1102 ( 
.A(n_899),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_1006),
.Y(n_1103)
);

AND2x2_ASAP7_75t_SL g1104 ( 
.A(n_992),
.B(n_996),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1002),
.A2(n_921),
.B(n_902),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_SL g1106 ( 
.A(n_1003),
.B(n_599),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_985),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_903),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_971),
.A2(n_902),
.B1(n_978),
.B2(n_970),
.Y(n_1109)
);

OAI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_971),
.A2(n_880),
.B1(n_599),
.B2(n_603),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_940),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_921),
.A2(n_970),
.B(n_902),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_902),
.B(n_970),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_983),
.B(n_826),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_973),
.Y(n_1115)
);

OA21x2_ASAP7_75t_L g1116 ( 
.A1(n_906),
.A2(n_915),
.B(n_974),
.Y(n_1116)
);

OR2x6_ASAP7_75t_L g1117 ( 
.A(n_955),
.B(n_709),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_902),
.B(n_970),
.Y(n_1118)
);

BUFx3_ASAP7_75t_L g1119 ( 
.A(n_973),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_SL g1120 ( 
.A(n_971),
.B(n_599),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_973),
.Y(n_1121)
);

AOI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_1013),
.A2(n_882),
.B1(n_872),
.B2(n_971),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_908),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_908),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_971),
.B(n_987),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_971),
.A2(n_902),
.B1(n_978),
.B2(n_970),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_908),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_971),
.A2(n_882),
.B(n_872),
.C(n_877),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_940),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_908),
.Y(n_1130)
);

AOI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_971),
.A2(n_882),
.B1(n_872),
.B2(n_880),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_987),
.B(n_880),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_902),
.B(n_970),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_941),
.Y(n_1134)
);

CKINVDCx11_ASAP7_75t_R g1135 ( 
.A(n_985),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_908),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_902),
.B(n_970),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_987),
.B(n_968),
.Y(n_1138)
);

CKINVDCx8_ASAP7_75t_R g1139 ( 
.A(n_973),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_941),
.Y(n_1140)
);

OR2x6_ASAP7_75t_L g1141 ( 
.A(n_955),
.B(n_709),
.Y(n_1141)
);

AND2x4_ASAP7_75t_L g1142 ( 
.A(n_983),
.B(n_826),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_987),
.B(n_880),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_902),
.B(n_970),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_971),
.A2(n_882),
.B(n_872),
.C(n_877),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_902),
.B(n_970),
.Y(n_1146)
);

INVx1_ASAP7_75t_SL g1147 ( 
.A(n_907),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_940),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_971),
.B(n_987),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_940),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_902),
.B(n_970),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_973),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_987),
.B(n_968),
.Y(n_1153)
);

CKINVDCx8_ASAP7_75t_R g1154 ( 
.A(n_973),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_1120),
.A2(n_1110),
.B1(n_1041),
.B2(n_1122),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1062),
.B(n_1037),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_1023),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_1120),
.A2(n_1041),
.B1(n_1132),
.B2(n_1143),
.Y(n_1158)
);

INVx3_ASAP7_75t_L g1159 ( 
.A(n_1095),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_1060),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_1135),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_1067),
.Y(n_1162)
);

AOI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1131),
.A2(n_1149),
.B1(n_1125),
.B2(n_1022),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_SL g1164 ( 
.A1(n_1050),
.A2(n_1126),
.B1(n_1109),
.B2(n_1022),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_1131),
.B(n_1138),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1046),
.A2(n_1037),
.B1(n_1069),
.B2(n_1063),
.Y(n_1166)
);

NAND2x1p5_ASAP7_75t_L g1167 ( 
.A(n_1099),
.B(n_1096),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_1095),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1034),
.Y(n_1169)
);

HB1xp67_ASAP7_75t_L g1170 ( 
.A(n_1040),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1118),
.A2(n_1133),
.B1(n_1151),
.B2(n_1146),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1042),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1065),
.B(n_1128),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1108),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_SL g1175 ( 
.A1(n_1145),
.A2(n_1050),
.B(n_1064),
.Y(n_1175)
);

AOI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1063),
.A2(n_1153),
.B1(n_1073),
.B2(n_1049),
.Y(n_1176)
);

INVx5_ASAP7_75t_L g1177 ( 
.A(n_1096),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1060),
.B(n_1026),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1026),
.B(n_1029),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1044),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1081),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1078),
.Y(n_1182)
);

INVx1_ASAP7_75t_SL g1183 ( 
.A(n_1121),
.Y(n_1183)
);

INVx6_ASAP7_75t_L g1184 ( 
.A(n_1032),
.Y(n_1184)
);

AO21x2_ASAP7_75t_L g1185 ( 
.A1(n_1083),
.A2(n_1079),
.B(n_1105),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1039),
.A2(n_1029),
.B1(n_1056),
.B2(n_1142),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1087),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1092),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_1123),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_1039),
.A2(n_1056),
.B1(n_1114),
.B2(n_1142),
.Y(n_1190)
);

NAND2x1p5_ASAP7_75t_L g1191 ( 
.A(n_1098),
.B(n_1116),
.Y(n_1191)
);

BUFx12f_ASAP7_75t_L g1192 ( 
.A(n_1031),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_1067),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1056),
.A2(n_1114),
.B1(n_1052),
.B2(n_1054),
.Y(n_1194)
);

AND2x4_ASAP7_75t_L g1195 ( 
.A(n_1055),
.B(n_1051),
.Y(n_1195)
);

NAND2x1p5_ASAP7_75t_L g1196 ( 
.A(n_1098),
.B(n_1116),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1054),
.A2(n_1117),
.B1(n_1141),
.B2(n_1106),
.Y(n_1197)
);

INVxp33_ASAP7_75t_L g1198 ( 
.A(n_1033),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1058),
.Y(n_1199)
);

OAI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1113),
.A2(n_1137),
.B1(n_1144),
.B2(n_1146),
.Y(n_1200)
);

AO21x2_ASAP7_75t_L g1201 ( 
.A1(n_1027),
.A2(n_1035),
.B(n_1086),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1074),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1113),
.B(n_1137),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1072),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1025),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1144),
.B(n_1024),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1111),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1129),
.Y(n_1208)
);

OR2x2_ASAP7_75t_L g1209 ( 
.A(n_1077),
.B(n_1147),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1148),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1150),
.Y(n_1211)
);

CKINVDCx20_ASAP7_75t_R g1212 ( 
.A(n_1038),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1061),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1075),
.A2(n_1047),
.B1(n_1084),
.B2(n_1154),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_SL g1215 ( 
.A(n_1115),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1117),
.A2(n_1141),
.B1(n_1106),
.B2(n_1036),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1061),
.Y(n_1217)
);

CKINVDCx20_ASAP7_75t_R g1218 ( 
.A(n_1107),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1057),
.Y(n_1219)
);

BUFx2_ASAP7_75t_R g1220 ( 
.A(n_1139),
.Y(n_1220)
);

INVx1_ASAP7_75t_SL g1221 ( 
.A(n_1147),
.Y(n_1221)
);

OA21x2_ASAP7_75t_L g1222 ( 
.A1(n_1100),
.A2(n_1020),
.B(n_1112),
.Y(n_1222)
);

BUFx8_ASAP7_75t_SL g1223 ( 
.A(n_1076),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1103),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1100),
.Y(n_1225)
);

NOR2x1_ASAP7_75t_R g1226 ( 
.A(n_1119),
.B(n_1152),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1028),
.A2(n_1053),
.B1(n_1043),
.B2(n_1045),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_SL g1228 ( 
.A(n_1030),
.B(n_1036),
.Y(n_1228)
);

INVxp67_ASAP7_75t_SL g1229 ( 
.A(n_1059),
.Y(n_1229)
);

BUFx2_ASAP7_75t_L g1230 ( 
.A(n_1055),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1102),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1093),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_L g1233 ( 
.A(n_1071),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1088),
.A2(n_1089),
.B(n_1136),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1051),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1066),
.Y(n_1236)
);

NAND2x1p5_ASAP7_75t_L g1237 ( 
.A(n_1104),
.B(n_1136),
.Y(n_1237)
);

INVx3_ASAP7_75t_L g1238 ( 
.A(n_1124),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1124),
.A2(n_1127),
.B(n_1130),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1094),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1091),
.A2(n_1021),
.B1(n_1134),
.B2(n_1048),
.Y(n_1241)
);

CKINVDCx12_ASAP7_75t_R g1242 ( 
.A(n_1032),
.Y(n_1242)
);

OR2x2_ASAP7_75t_L g1243 ( 
.A(n_1070),
.B(n_1068),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1070),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1080),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1021),
.Y(n_1246)
);

INVx2_ASAP7_75t_SL g1247 ( 
.A(n_1032),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1021),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1048),
.A2(n_1082),
.B(n_1085),
.Y(n_1249)
);

INVxp67_ASAP7_75t_L g1250 ( 
.A(n_1048),
.Y(n_1250)
);

INVx6_ASAP7_75t_L g1251 ( 
.A(n_1082),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1082),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1085),
.A2(n_1090),
.B1(n_1134),
.B2(n_1140),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1085),
.B(n_1090),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1090),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1134),
.B(n_1140),
.Y(n_1256)
);

INVx2_ASAP7_75t_SL g1257 ( 
.A(n_1140),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1095),
.Y(n_1258)
);

INVxp33_ASAP7_75t_L g1259 ( 
.A(n_1023),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1120),
.A2(n_872),
.B1(n_882),
.B2(n_1013),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1034),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_SL g1262 ( 
.A1(n_1120),
.A2(n_1041),
.B1(n_760),
.B2(n_987),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1120),
.A2(n_872),
.B1(n_882),
.B2(n_1013),
.Y(n_1263)
);

INVx3_ASAP7_75t_L g1264 ( 
.A(n_1095),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1131),
.A2(n_971),
.B1(n_880),
.B2(n_1122),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1120),
.A2(n_872),
.B1(n_882),
.B2(n_1013),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_1038),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_1060),
.Y(n_1268)
);

BUFx10_ASAP7_75t_L g1269 ( 
.A(n_1067),
.Y(n_1269)
);

AOI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1101),
.A2(n_919),
.B(n_909),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1097),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1179),
.B(n_1200),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1181),
.B(n_1188),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_1177),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1181),
.B(n_1188),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1265),
.A2(n_1155),
.B1(n_1263),
.B2(n_1260),
.Y(n_1276)
);

INVxp67_ASAP7_75t_L g1277 ( 
.A(n_1209),
.Y(n_1277)
);

INVx2_ASAP7_75t_SL g1278 ( 
.A(n_1237),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1271),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1182),
.B(n_1187),
.Y(n_1280)
);

OAI21xp33_ASAP7_75t_SL g1281 ( 
.A1(n_1206),
.A2(n_1266),
.B(n_1203),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1262),
.A2(n_1163),
.B1(n_1158),
.B2(n_1176),
.Y(n_1282)
);

OR2x2_ASAP7_75t_L g1283 ( 
.A(n_1209),
.B(n_1225),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1231),
.B(n_1236),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1156),
.B(n_1179),
.Y(n_1285)
);

OA21x2_ASAP7_75t_L g1286 ( 
.A1(n_1175),
.A2(n_1270),
.B(n_1202),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_L g1287 ( 
.A(n_1198),
.B(n_1165),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1236),
.Y(n_1288)
);

OR2x2_ASAP7_75t_L g1289 ( 
.A(n_1156),
.B(n_1178),
.Y(n_1289)
);

OR2x2_ASAP7_75t_L g1290 ( 
.A(n_1178),
.B(n_1191),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1191),
.B(n_1196),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1231),
.Y(n_1292)
);

INVx4_ASAP7_75t_L g1293 ( 
.A(n_1177),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1191),
.B(n_1196),
.Y(n_1294)
);

INVxp67_ASAP7_75t_SL g1295 ( 
.A(n_1196),
.Y(n_1295)
);

INVxp67_ASAP7_75t_SL g1296 ( 
.A(n_1204),
.Y(n_1296)
);

OR2x2_ASAP7_75t_L g1297 ( 
.A(n_1201),
.B(n_1185),
.Y(n_1297)
);

AND2x4_ASAP7_75t_L g1298 ( 
.A(n_1234),
.B(n_1224),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1222),
.Y(n_1299)
);

INVx1_ASAP7_75t_SL g1300 ( 
.A(n_1221),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1222),
.Y(n_1301)
);

BUFx2_ASAP7_75t_L g1302 ( 
.A(n_1237),
.Y(n_1302)
);

BUFx2_ASAP7_75t_L g1303 ( 
.A(n_1237),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1201),
.B(n_1173),
.Y(n_1304)
);

INVx2_ASAP7_75t_SL g1305 ( 
.A(n_1234),
.Y(n_1305)
);

INVx3_ASAP7_75t_L g1306 ( 
.A(n_1167),
.Y(n_1306)
);

BUFx2_ASAP7_75t_L g1307 ( 
.A(n_1167),
.Y(n_1307)
);

INVxp33_ASAP7_75t_L g1308 ( 
.A(n_1226),
.Y(n_1308)
);

AO21x2_ASAP7_75t_L g1309 ( 
.A1(n_1180),
.A2(n_1217),
.B(n_1213),
.Y(n_1309)
);

OA21x2_ASAP7_75t_L g1310 ( 
.A1(n_1197),
.A2(n_1166),
.B(n_1180),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1164),
.B(n_1167),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1216),
.B(n_1160),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1160),
.B(n_1268),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1205),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1207),
.Y(n_1315)
);

OA21x2_ASAP7_75t_L g1316 ( 
.A1(n_1186),
.A2(n_1194),
.B(n_1208),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1210),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1268),
.B(n_1211),
.Y(n_1318)
);

AO31x2_ASAP7_75t_L g1319 ( 
.A1(n_1171),
.A2(n_1174),
.A3(n_1172),
.B(n_1169),
.Y(n_1319)
);

INVx3_ASAP7_75t_L g1320 ( 
.A(n_1239),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1261),
.B(n_1240),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1235),
.B(n_1195),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1199),
.Y(n_1323)
);

AOI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1232),
.A2(n_1214),
.B(n_1230),
.Y(n_1324)
);

INVxp67_ASAP7_75t_SL g1325 ( 
.A(n_1170),
.Y(n_1325)
);

INVx3_ASAP7_75t_L g1326 ( 
.A(n_1159),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1277),
.B(n_1229),
.Y(n_1327)
);

AND2x4_ASAP7_75t_L g1328 ( 
.A(n_1298),
.B(n_1258),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1277),
.B(n_1157),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1276),
.A2(n_1190),
.B1(n_1195),
.B2(n_1267),
.Y(n_1330)
);

INVx3_ASAP7_75t_L g1331 ( 
.A(n_1298),
.Y(n_1331)
);

INVx2_ASAP7_75t_SL g1332 ( 
.A(n_1298),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1304),
.B(n_1195),
.Y(n_1333)
);

INVxp67_ASAP7_75t_L g1334 ( 
.A(n_1288),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1304),
.B(n_1219),
.Y(n_1335)
);

BUFx2_ASAP7_75t_L g1336 ( 
.A(n_1298),
.Y(n_1336)
);

BUFx2_ASAP7_75t_L g1337 ( 
.A(n_1284),
.Y(n_1337)
);

OR2x2_ASAP7_75t_L g1338 ( 
.A(n_1290),
.B(n_1289),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1291),
.B(n_1244),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1291),
.B(n_1294),
.Y(n_1340)
);

OR2x2_ASAP7_75t_L g1341 ( 
.A(n_1290),
.B(n_1183),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1294),
.B(n_1279),
.Y(n_1342)
);

NOR2x1_ASAP7_75t_L g1343 ( 
.A(n_1293),
.B(n_1159),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1287),
.B(n_1267),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1285),
.B(n_1189),
.Y(n_1345)
);

AND2x4_ASAP7_75t_L g1346 ( 
.A(n_1320),
.B(n_1305),
.Y(n_1346)
);

CKINVDCx6p67_ASAP7_75t_R g1347 ( 
.A(n_1274),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1272),
.B(n_1285),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1289),
.B(n_1233),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1285),
.B(n_1238),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_1284),
.Y(n_1351)
);

NAND2x1p5_ASAP7_75t_L g1352 ( 
.A(n_1293),
.B(n_1168),
.Y(n_1352)
);

INVx1_ASAP7_75t_SL g1353 ( 
.A(n_1300),
.Y(n_1353)
);

INVx3_ASAP7_75t_L g1354 ( 
.A(n_1284),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1286),
.B(n_1168),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1272),
.B(n_1168),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1309),
.Y(n_1357)
);

INVxp67_ASAP7_75t_L g1358 ( 
.A(n_1288),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1286),
.B(n_1264),
.Y(n_1359)
);

INVx2_ASAP7_75t_SL g1360 ( 
.A(n_1284),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1286),
.B(n_1264),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1283),
.B(n_1258),
.Y(n_1362)
);

INVxp67_ASAP7_75t_L g1363 ( 
.A(n_1325),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1283),
.B(n_1319),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1340),
.B(n_1342),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1356),
.B(n_1325),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1330),
.A2(n_1276),
.B1(n_1282),
.B2(n_1312),
.Y(n_1367)
);

OAI21xp33_ASAP7_75t_SL g1368 ( 
.A1(n_1360),
.A2(n_1296),
.B(n_1282),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1356),
.B(n_1281),
.Y(n_1369)
);

NAND3xp33_ASAP7_75t_L g1370 ( 
.A(n_1344),
.B(n_1281),
.C(n_1312),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1353),
.B(n_1318),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1353),
.B(n_1318),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1348),
.B(n_1318),
.Y(n_1373)
);

NAND3xp33_ASAP7_75t_L g1374 ( 
.A(n_1327),
.B(n_1312),
.C(n_1311),
.Y(n_1374)
);

OAI21xp33_ASAP7_75t_L g1375 ( 
.A1(n_1348),
.A2(n_1311),
.B(n_1324),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1335),
.B(n_1313),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1341),
.A2(n_1311),
.B1(n_1300),
.B2(n_1308),
.Y(n_1377)
);

NAND4xp25_ASAP7_75t_L g1378 ( 
.A(n_1329),
.B(n_1228),
.C(n_1321),
.D(n_1314),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1335),
.B(n_1313),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1335),
.B(n_1313),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1327),
.B(n_1315),
.Y(n_1381)
);

NOR2xp33_ASAP7_75t_L g1382 ( 
.A(n_1341),
.B(n_1324),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1329),
.B(n_1362),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1342),
.B(n_1295),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1362),
.B(n_1315),
.Y(n_1385)
);

OA21x2_ASAP7_75t_L g1386 ( 
.A1(n_1355),
.A2(n_1301),
.B(n_1299),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1349),
.B(n_1315),
.Y(n_1387)
);

NAND3xp33_ASAP7_75t_L g1388 ( 
.A(n_1363),
.B(n_1316),
.C(n_1310),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1342),
.B(n_1273),
.Y(n_1389)
);

OAI21xp33_ASAP7_75t_L g1390 ( 
.A1(n_1364),
.A2(n_1259),
.B(n_1275),
.Y(n_1390)
);

OAI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1343),
.A2(n_1278),
.B(n_1297),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1349),
.B(n_1317),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1347),
.A2(n_1220),
.B1(n_1302),
.B2(n_1303),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1337),
.B(n_1273),
.Y(n_1394)
);

NOR3xp33_ASAP7_75t_L g1395 ( 
.A(n_1343),
.B(n_1258),
.C(n_1227),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1363),
.B(n_1345),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1345),
.B(n_1317),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1351),
.B(n_1275),
.Y(n_1398)
);

AOI221xp5_ASAP7_75t_L g1399 ( 
.A1(n_1334),
.A2(n_1321),
.B1(n_1314),
.B2(n_1323),
.C(n_1292),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1347),
.A2(n_1303),
.B1(n_1302),
.B2(n_1316),
.Y(n_1400)
);

NOR3xp33_ASAP7_75t_L g1401 ( 
.A(n_1355),
.B(n_1326),
.C(n_1306),
.Y(n_1401)
);

NAND3xp33_ASAP7_75t_L g1402 ( 
.A(n_1355),
.B(n_1316),
.C(n_1310),
.Y(n_1402)
);

AOI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1339),
.A2(n_1316),
.B1(n_1310),
.B2(n_1322),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1345),
.B(n_1317),
.Y(n_1404)
);

OAI221xp5_ASAP7_75t_L g1405 ( 
.A1(n_1352),
.A2(n_1278),
.B1(n_1307),
.B2(n_1306),
.C(n_1161),
.Y(n_1405)
);

OAI221xp5_ASAP7_75t_L g1406 ( 
.A1(n_1352),
.A2(n_1278),
.B1(n_1307),
.B2(n_1306),
.C(n_1161),
.Y(n_1406)
);

OA21x2_ASAP7_75t_L g1407 ( 
.A1(n_1359),
.A2(n_1301),
.B(n_1299),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1350),
.B(n_1292),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_SL g1409 ( 
.A(n_1328),
.B(n_1322),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1350),
.B(n_1280),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1350),
.B(n_1280),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_SL g1412 ( 
.A1(n_1352),
.A2(n_1212),
.B1(n_1218),
.B2(n_1242),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1338),
.B(n_1280),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1386),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1389),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1386),
.Y(n_1416)
);

BUFx2_ASAP7_75t_L g1417 ( 
.A(n_1386),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1369),
.B(n_1364),
.Y(n_1418)
);

INVx1_ASAP7_75t_SL g1419 ( 
.A(n_1387),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1407),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1389),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1397),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1407),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1407),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1382),
.B(n_1334),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1365),
.Y(n_1426)
);

INVxp67_ASAP7_75t_SL g1427 ( 
.A(n_1382),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1402),
.B(n_1338),
.Y(n_1428)
);

AND2x4_ASAP7_75t_SL g1429 ( 
.A(n_1401),
.B(n_1347),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1404),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1383),
.B(n_1358),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1384),
.Y(n_1432)
);

AND2x4_ASAP7_75t_SL g1433 ( 
.A(n_1395),
.B(n_1293),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1403),
.B(n_1336),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1403),
.B(n_1331),
.Y(n_1435)
);

OR2x2_ASAP7_75t_L g1436 ( 
.A(n_1388),
.B(n_1332),
.Y(n_1436)
);

AND2x4_ASAP7_75t_L g1437 ( 
.A(n_1409),
.B(n_1346),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1366),
.B(n_1332),
.Y(n_1438)
);

INVx2_ASAP7_75t_SL g1439 ( 
.A(n_1409),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1396),
.B(n_1332),
.Y(n_1440)
);

INVx2_ASAP7_75t_SL g1441 ( 
.A(n_1394),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1385),
.B(n_1357),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1398),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_L g1444 ( 
.A(n_1378),
.B(n_1333),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1410),
.B(n_1361),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1411),
.B(n_1361),
.Y(n_1446)
);

AND2x4_ASAP7_75t_SL g1447 ( 
.A(n_1368),
.B(n_1293),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1413),
.B(n_1361),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1444),
.B(n_1412),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1428),
.B(n_1392),
.Y(n_1450)
);

INVxp67_ASAP7_75t_L g1451 ( 
.A(n_1444),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1415),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1428),
.B(n_1408),
.Y(n_1453)
);

AOI221xp5_ASAP7_75t_L g1454 ( 
.A1(n_1427),
.A2(n_1370),
.B1(n_1375),
.B2(n_1367),
.C(n_1377),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1427),
.B(n_1373),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1419),
.B(n_1371),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1433),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1426),
.B(n_1354),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1417),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1419),
.B(n_1372),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1417),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1438),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1415),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1421),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1421),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1432),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1418),
.A2(n_1405),
.B(n_1406),
.Y(n_1467)
);

OAI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1418),
.A2(n_1374),
.B1(n_1393),
.B2(n_1400),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1426),
.B(n_1354),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1432),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1428),
.B(n_1376),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1426),
.B(n_1437),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1417),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1432),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1432),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1414),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1425),
.B(n_1379),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1426),
.B(n_1354),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1438),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1425),
.B(n_1380),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1414),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1414),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1442),
.B(n_1436),
.Y(n_1483)
);

OR2x6_ASAP7_75t_L g1484 ( 
.A(n_1436),
.B(n_1391),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1438),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1433),
.A2(n_1390),
.B1(n_1399),
.B2(n_1352),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1431),
.B(n_1381),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1483),
.B(n_1436),
.Y(n_1488)
);

OR2x6_ASAP7_75t_L g1489 ( 
.A(n_1484),
.B(n_1274),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1484),
.B(n_1457),
.Y(n_1490)
);

NOR2x1_ASAP7_75t_L g1491 ( 
.A(n_1468),
.B(n_1431),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1451),
.B(n_1422),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_SL g1493 ( 
.A(n_1449),
.B(n_1368),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1483),
.B(n_1442),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1462),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1452),
.Y(n_1496)
);

INVxp33_ASAP7_75t_L g1497 ( 
.A(n_1454),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1484),
.B(n_1457),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1485),
.B(n_1429),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1452),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1467),
.B(n_1422),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_1479),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1463),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1459),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1484),
.B(n_1439),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1484),
.B(n_1439),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1485),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1487),
.B(n_1430),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_L g1509 ( 
.A(n_1477),
.B(n_1192),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1459),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1463),
.Y(n_1511)
);

NOR2xp67_ASAP7_75t_L g1512 ( 
.A(n_1471),
.B(n_1439),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1472),
.B(n_1434),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1464),
.Y(n_1514)
);

AOI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1486),
.A2(n_1433),
.B1(n_1434),
.B2(n_1447),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1461),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1477),
.B(n_1480),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1453),
.B(n_1450),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1472),
.B(n_1429),
.Y(n_1519)
);

NAND3xp33_ASAP7_75t_L g1520 ( 
.A(n_1450),
.B(n_1434),
.C(n_1435),
.Y(n_1520)
);

OR2x2_ASAP7_75t_SL g1521 ( 
.A(n_1471),
.B(n_1416),
.Y(n_1521)
);

INVx2_ASAP7_75t_SL g1522 ( 
.A(n_1461),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1473),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1480),
.B(n_1430),
.Y(n_1524)
);

INVx1_ASAP7_75t_SL g1525 ( 
.A(n_1456),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1473),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1476),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1458),
.B(n_1469),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1464),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1455),
.B(n_1448),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1497),
.A2(n_1435),
.B1(n_1433),
.B2(n_1322),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1490),
.B(n_1458),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1490),
.B(n_1469),
.Y(n_1533)
);

CKINVDCx16_ASAP7_75t_R g1534 ( 
.A(n_1493),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1517),
.B(n_1453),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1491),
.B(n_1465),
.Y(n_1536)
);

OR2x6_ASAP7_75t_L g1537 ( 
.A(n_1489),
.B(n_1192),
.Y(n_1537)
);

NOR2x1_ASAP7_75t_L g1538 ( 
.A(n_1501),
.B(n_1218),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1497),
.B(n_1465),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1496),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1522),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1496),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1509),
.A2(n_1520),
.B1(n_1525),
.B2(n_1495),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1500),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1502),
.B(n_1445),
.Y(n_1545)
);

AND2x2_ASAP7_75t_SL g1546 ( 
.A(n_1498),
.B(n_1447),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_L g1547 ( 
.A(n_1492),
.B(n_1223),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1516),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1500),
.Y(n_1549)
);

INVxp67_ASAP7_75t_L g1550 ( 
.A(n_1512),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1503),
.Y(n_1551)
);

INVx1_ASAP7_75t_SL g1552 ( 
.A(n_1498),
.Y(n_1552)
);

INVx3_ASAP7_75t_SL g1553 ( 
.A(n_1521),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1503),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1523),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1511),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1508),
.B(n_1445),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1524),
.B(n_1445),
.Y(n_1558)
);

INVx6_ASAP7_75t_L g1559 ( 
.A(n_1499),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1511),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1529),
.Y(n_1561)
);

INVxp67_ASAP7_75t_L g1562 ( 
.A(n_1505),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_1499),
.Y(n_1563)
);

INVx3_ASAP7_75t_SL g1564 ( 
.A(n_1521),
.Y(n_1564)
);

INVxp67_ASAP7_75t_L g1565 ( 
.A(n_1505),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1515),
.A2(n_1435),
.B1(n_1322),
.B2(n_1310),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1552),
.B(n_1507),
.Y(n_1567)
);

OA21x2_ASAP7_75t_SL g1568 ( 
.A1(n_1536),
.A2(n_1499),
.B(n_1519),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1548),
.Y(n_1569)
);

AOI33xp33_ASAP7_75t_L g1570 ( 
.A1(n_1543),
.A2(n_1506),
.A3(n_1522),
.B1(n_1504),
.B2(n_1510),
.B3(n_1526),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1563),
.B(n_1519),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1548),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1553),
.A2(n_1519),
.B1(n_1489),
.B2(n_1518),
.Y(n_1573)
);

OAI221xp5_ASAP7_75t_L g1574 ( 
.A1(n_1553),
.A2(n_1564),
.B1(n_1538),
.B2(n_1543),
.C(n_1539),
.Y(n_1574)
);

AOI221xp5_ASAP7_75t_SL g1575 ( 
.A1(n_1562),
.A2(n_1506),
.B1(n_1513),
.B2(n_1488),
.C(n_1529),
.Y(n_1575)
);

INVx2_ASAP7_75t_SL g1576 ( 
.A(n_1559),
.Y(n_1576)
);

AOI221xp5_ASAP7_75t_L g1577 ( 
.A1(n_1564),
.A2(n_1526),
.B1(n_1504),
.B2(n_1510),
.C(n_1488),
.Y(n_1577)
);

AOI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1534),
.A2(n_1489),
.B1(n_1447),
.B2(n_1429),
.Y(n_1578)
);

OAI33xp33_ASAP7_75t_L g1579 ( 
.A1(n_1565),
.A2(n_1494),
.A3(n_1514),
.B1(n_1518),
.B2(n_1527),
.B3(n_1530),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1550),
.B(n_1513),
.Y(n_1580)
);

AOI211xp5_ASAP7_75t_L g1581 ( 
.A1(n_1547),
.A2(n_1494),
.B(n_1527),
.C(n_1420),
.Y(n_1581)
);

INVx1_ASAP7_75t_SL g1582 ( 
.A(n_1559),
.Y(n_1582)
);

AOI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1555),
.A2(n_1489),
.B(n_1420),
.Y(n_1583)
);

INVx2_ASAP7_75t_SL g1584 ( 
.A(n_1559),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1537),
.A2(n_1447),
.B1(n_1429),
.B2(n_1528),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1541),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1555),
.Y(n_1587)
);

AOI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1546),
.A2(n_1437),
.B1(n_1460),
.B2(n_1328),
.Y(n_1588)
);

OAI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1537),
.A2(n_1441),
.B1(n_1440),
.B2(n_1443),
.Y(n_1589)
);

AOI211xp5_ASAP7_75t_L g1590 ( 
.A1(n_1547),
.A2(n_1416),
.B(n_1528),
.C(n_1481),
.Y(n_1590)
);

AOI222xp33_ASAP7_75t_L g1591 ( 
.A1(n_1566),
.A2(n_1474),
.B1(n_1466),
.B2(n_1470),
.C1(n_1475),
.C2(n_1424),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1540),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_SL g1593 ( 
.A(n_1574),
.B(n_1546),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1569),
.Y(n_1594)
);

INVxp67_ASAP7_75t_L g1595 ( 
.A(n_1574),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1572),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1580),
.B(n_1535),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1587),
.Y(n_1598)
);

AND2x4_ASAP7_75t_SL g1599 ( 
.A(n_1571),
.B(n_1212),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1592),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1567),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1582),
.B(n_1545),
.Y(n_1602)
);

INVxp67_ASAP7_75t_SL g1603 ( 
.A(n_1576),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1584),
.B(n_1541),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1586),
.Y(n_1605)
);

CKINVDCx16_ASAP7_75t_R g1606 ( 
.A(n_1573),
.Y(n_1606)
);

NOR2x1_ASAP7_75t_L g1607 ( 
.A(n_1583),
.B(n_1537),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1570),
.B(n_1532),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1575),
.B(n_1533),
.Y(n_1609)
);

A2O1A1Ixp33_ASAP7_75t_L g1610 ( 
.A1(n_1581),
.A2(n_1577),
.B(n_1590),
.C(n_1583),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1579),
.B(n_1558),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1577),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1591),
.B(n_1542),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1594),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_SL g1615 ( 
.A1(n_1595),
.A2(n_1568),
.B1(n_1544),
.B2(n_1551),
.Y(n_1615)
);

O2A1O1Ixp33_ASAP7_75t_SL g1616 ( 
.A1(n_1610),
.A2(n_1612),
.B(n_1613),
.C(n_1609),
.Y(n_1616)
);

AND5x1_ASAP7_75t_L g1617 ( 
.A(n_1593),
.B(n_1578),
.C(n_1588),
.D(n_1585),
.E(n_1589),
.Y(n_1617)
);

NAND3xp33_ASAP7_75t_SL g1618 ( 
.A(n_1593),
.B(n_1566),
.C(n_1531),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1599),
.B(n_1531),
.Y(n_1619)
);

OAI211xp5_ASAP7_75t_L g1620 ( 
.A1(n_1607),
.A2(n_1561),
.B(n_1560),
.C(n_1556),
.Y(n_1620)
);

AOI21xp33_ASAP7_75t_L g1621 ( 
.A1(n_1603),
.A2(n_1554),
.B(n_1549),
.Y(n_1621)
);

NAND3xp33_ASAP7_75t_SL g1622 ( 
.A(n_1611),
.B(n_1557),
.C(n_1223),
.Y(n_1622)
);

A2O1A1Ixp33_ASAP7_75t_L g1623 ( 
.A1(n_1613),
.A2(n_1414),
.B(n_1424),
.C(n_1423),
.Y(n_1623)
);

AOI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1606),
.A2(n_1437),
.B1(n_1215),
.B2(n_1470),
.Y(n_1624)
);

OAI21xp33_ASAP7_75t_L g1625 ( 
.A1(n_1608),
.A2(n_1481),
.B(n_1476),
.Y(n_1625)
);

NAND4xp25_ASAP7_75t_SL g1626 ( 
.A(n_1620),
.B(n_1604),
.C(n_1602),
.D(n_1597),
.Y(n_1626)
);

NAND5xp2_ASAP7_75t_L g1627 ( 
.A(n_1616),
.B(n_1601),
.C(n_1598),
.D(n_1596),
.E(n_1605),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_1614),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1622),
.B(n_1600),
.Y(n_1629)
);

AOI211xp5_ASAP7_75t_SL g1630 ( 
.A1(n_1618),
.A2(n_1253),
.B(n_1250),
.C(n_1242),
.Y(n_1630)
);

NOR2xp67_ASAP7_75t_L g1631 ( 
.A(n_1624),
.B(n_1482),
.Y(n_1631)
);

AOI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1618),
.A2(n_1215),
.B1(n_1437),
.B2(n_1482),
.Y(n_1632)
);

NOR3xp33_ASAP7_75t_L g1633 ( 
.A(n_1621),
.B(n_1193),
.C(n_1162),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1615),
.B(n_1466),
.Y(n_1634)
);

NOR2x1_ASAP7_75t_L g1635 ( 
.A(n_1619),
.B(n_1248),
.Y(n_1635)
);

NAND4xp25_ASAP7_75t_L g1636 ( 
.A(n_1627),
.B(n_1625),
.C(n_1617),
.D(n_1623),
.Y(n_1636)
);

OAI221xp5_ASAP7_75t_L g1637 ( 
.A1(n_1632),
.A2(n_1475),
.B1(n_1474),
.B2(n_1441),
.C(n_1442),
.Y(n_1637)
);

NAND3xp33_ASAP7_75t_SL g1638 ( 
.A(n_1630),
.B(n_1215),
.C(n_1241),
.Y(n_1638)
);

OAI211xp5_ASAP7_75t_L g1639 ( 
.A1(n_1629),
.A2(n_1162),
.B(n_1193),
.C(n_1247),
.Y(n_1639)
);

AOI211x1_ASAP7_75t_SL g1640 ( 
.A1(n_1631),
.A2(n_1424),
.B(n_1423),
.C(n_1252),
.Y(n_1640)
);

NOR4xp25_ASAP7_75t_L g1641 ( 
.A(n_1626),
.B(n_1246),
.C(n_1255),
.D(n_1424),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1641),
.B(n_1628),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1639),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1636),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1640),
.Y(n_1645)
);

BUFx2_ASAP7_75t_L g1646 ( 
.A(n_1638),
.Y(n_1646)
);

INVxp67_ASAP7_75t_SL g1647 ( 
.A(n_1637),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1639),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1644),
.B(n_1647),
.Y(n_1649)
);

NOR3xp33_ASAP7_75t_L g1650 ( 
.A(n_1646),
.B(n_1635),
.C(n_1633),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1643),
.Y(n_1651)
);

NOR3xp33_ASAP7_75t_L g1652 ( 
.A(n_1642),
.B(n_1634),
.C(n_1247),
.Y(n_1652)
);

INVx1_ASAP7_75t_SL g1653 ( 
.A(n_1648),
.Y(n_1653)
);

XOR2x1_ASAP7_75t_L g1654 ( 
.A(n_1649),
.B(n_1645),
.Y(n_1654)
);

NAND3x1_ASAP7_75t_L g1655 ( 
.A(n_1652),
.B(n_1647),
.C(n_1256),
.Y(n_1655)
);

AOI22x1_ASAP7_75t_L g1656 ( 
.A1(n_1653),
.A2(n_1423),
.B1(n_1257),
.B2(n_1441),
.Y(n_1656)
);

OAI22xp5_ASAP7_75t_SL g1657 ( 
.A1(n_1654),
.A2(n_1651),
.B1(n_1650),
.B2(n_1184),
.Y(n_1657)
);

AOI21xp33_ASAP7_75t_L g1658 ( 
.A1(n_1657),
.A2(n_1655),
.B(n_1656),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1658),
.Y(n_1659)
);

AO21x2_ASAP7_75t_L g1660 ( 
.A1(n_1658),
.A2(n_1423),
.B(n_1249),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1659),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1660),
.B(n_1478),
.Y(n_1662)
);

AOI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1661),
.A2(n_1660),
.B(n_1257),
.Y(n_1663)
);

AOI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1662),
.A2(n_1184),
.B1(n_1478),
.B2(n_1269),
.Y(n_1664)
);

OA21x2_ASAP7_75t_L g1665 ( 
.A1(n_1663),
.A2(n_1664),
.B(n_1249),
.Y(n_1665)
);

AOI222xp33_ASAP7_75t_L g1666 ( 
.A1(n_1665),
.A2(n_1269),
.B1(n_1184),
.B2(n_1248),
.C1(n_1251),
.C2(n_1446),
.Y(n_1666)
);

OAI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1666),
.A2(n_1184),
.B1(n_1251),
.B2(n_1243),
.C(n_1245),
.Y(n_1667)
);

AOI211xp5_ASAP7_75t_L g1668 ( 
.A1(n_1667),
.A2(n_1256),
.B(n_1254),
.C(n_1243),
.Y(n_1668)
);


endmodule