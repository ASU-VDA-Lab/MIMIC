module fake_netlist_5_874_n_89 (n_16, n_0, n_12, n_9, n_18, n_1, n_8, n_10, n_4, n_11, n_17, n_19, n_7, n_15, n_20, n_5, n_14, n_2, n_13, n_3, n_6, n_89);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_1;
input n_8;
input n_10;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_20;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_89;

wire n_82;
wire n_24;
wire n_86;
wire n_83;
wire n_61;
wire n_75;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_37;
wire n_31;
wire n_66;
wire n_60;
wire n_43;
wire n_58;
wire n_69;
wire n_42;
wire n_22;
wire n_45;
wire n_46;
wire n_21;
wire n_38;
wire n_80;
wire n_35;
wire n_73;
wire n_30;
wire n_33;
wire n_84;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_62;
wire n_71;
wire n_85;
wire n_59;
wire n_26;
wire n_55;
wire n_49;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_87;
wire n_27;
wire n_64;
wire n_77;
wire n_81;
wire n_28;
wire n_70;
wire n_68;
wire n_72;
wire n_32;
wire n_41;
wire n_56;
wire n_51;
wire n_63;
wire n_48;
wire n_50;
wire n_52;
wire n_88;

INVx5_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

AND2x4_ASAP7_75t_L g25 ( 
.A(n_0),
.B(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_9),
.B(n_20),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_1),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

AND2x6_ASAP7_75t_SL g41 ( 
.A(n_25),
.B(n_5),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_13),
.B(n_14),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_32),
.B(n_25),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_29),
.A2(n_34),
.B1(n_36),
.B2(n_31),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

OAI21x1_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_33),
.B(n_27),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

AOI21x1_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_28),
.B(n_23),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_45),
.A2(n_26),
.B(n_30),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_21),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

OA21x2_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_43),
.B(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_49),
.Y(n_61)
);

NOR2xp67_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_47),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVxp67_ASAP7_75t_SL g65 ( 
.A(n_57),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVxp67_ASAP7_75t_SL g67 ( 
.A(n_58),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

NAND2x1p5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_60),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_59),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_46),
.B(n_67),
.C(n_49),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_69),
.A2(n_63),
.B(n_21),
.C(n_24),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_61),
.B(n_63),
.Y(n_76)
);

AND3x4_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_70),
.C(n_71),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_63),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_SL g80 ( 
.A(n_77),
.B(n_74),
.C(n_22),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_77),
.Y(n_82)
);

AO22x2_ASAP7_75t_L g83 ( 
.A1(n_80),
.A2(n_78),
.B1(n_21),
.B2(n_24),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_81),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

OA21x2_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_84),
.B(n_85),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_83),
.Y(n_89)
);


endmodule