module fake_jpeg_661_n_539 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_539);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_539;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_3),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_58),
.Y(n_202)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_59),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_60),
.B(n_61),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_19),
.B(n_18),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_62),
.B(n_66),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_19),
.B(n_52),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_64),
.B(n_65),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_47),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g162 ( 
.A(n_67),
.Y(n_162)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_33),
.B(n_16),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_69),
.B(n_76),
.Y(n_169)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_70),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_33),
.A2(n_16),
.B1(n_1),
.B2(n_2),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_72),
.B(n_101),
.C(n_2),
.Y(n_179)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_73),
.Y(n_166)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_33),
.B(n_0),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_37),
.B(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_77),
.B(n_88),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_24),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_78),
.B(n_79),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_24),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_37),
.B(n_36),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_80),
.B(n_82),
.Y(n_172)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_81),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_24),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_85),
.B(n_91),
.Y(n_175)
);

BUFx8_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g200 ( 
.A(n_86),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_20),
.B(n_0),
.Y(n_88)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_89),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_39),
.Y(n_90)
);

NAND2xp33_ASAP7_75t_SL g142 ( 
.A(n_90),
.B(n_121),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_48),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_92),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_21),
.B(n_1),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_93),
.B(n_112),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_38),
.B(n_1),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_94),
.B(n_124),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_95),
.Y(n_157)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_96),
.Y(n_150)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_97),
.Y(n_156)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_99),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_100),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_56),
.B(n_51),
.C(n_31),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_102),
.Y(n_194)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_22),
.Y(n_103)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_104),
.Y(n_209)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_26),
.Y(n_105)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_105),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_109),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_29),
.Y(n_110)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_46),
.Y(n_111)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_111),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_23),
.B(n_32),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_46),
.Y(n_113)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_113),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_51),
.Y(n_114)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_114),
.Y(n_193)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_46),
.Y(n_115)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_115),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_23),
.B(n_2),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_116),
.B(n_125),
.Y(n_201)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_46),
.Y(n_117)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_117),
.Y(n_173)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_49),
.Y(n_118)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_118),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_119),
.Y(n_189)
);

INVx4_ASAP7_75t_SL g120 ( 
.A(n_49),
.Y(n_120)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_120),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_31),
.Y(n_121)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_49),
.Y(n_122)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_122),
.Y(n_208)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_49),
.Y(n_123)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_123),
.Y(n_196)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_49),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_54),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_72),
.A2(n_55),
.B1(n_38),
.B2(n_41),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_127),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_120),
.A2(n_31),
.B1(n_54),
.B2(n_53),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_86),
.A2(n_54),
.B1(n_28),
.B2(n_53),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_86),
.A2(n_54),
.B1(n_28),
.B2(n_44),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_101),
.A2(n_55),
.B1(n_41),
.B2(n_27),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_140),
.A2(n_144),
.B1(n_154),
.B2(n_158),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_80),
.A2(n_35),
.B1(n_44),
.B2(n_42),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_141),
.A2(n_205),
.B1(n_211),
.B2(n_130),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_90),
.A2(n_54),
.B1(n_42),
.B2(n_35),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_109),
.A2(n_34),
.B1(n_32),
.B2(n_40),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_57),
.A2(n_34),
.B1(n_40),
.B2(n_29),
.Y(n_158)
);

AND2x2_ASAP7_75t_SL g160 ( 
.A(n_68),
.B(n_40),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_160),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_74),
.A2(n_40),
.B1(n_29),
.B2(n_5),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_161),
.A2(n_167),
.B1(n_177),
.B2(n_180),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_103),
.B(n_2),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_165),
.B(n_181),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_70),
.A2(n_40),
.B1(n_4),
.B2(n_5),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_75),
.A2(n_105),
.B1(n_121),
.B2(n_115),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_179),
.B(n_164),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_63),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_83),
.B(n_4),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_113),
.B(n_117),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_182),
.B(n_183),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_58),
.B(n_4),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_119),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_186),
.A2(n_187),
.B1(n_190),
.B2(n_195),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_99),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_98),
.A2(n_124),
.B1(n_114),
.B2(n_123),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_125),
.B(n_11),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_191),
.B(n_204),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_71),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_73),
.A2(n_13),
.B1(n_15),
.B2(n_84),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_198),
.A2(n_200),
.B1(n_143),
.B2(n_135),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_89),
.B(n_13),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_87),
.A2(n_13),
.B1(n_106),
.B2(n_92),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_104),
.A2(n_108),
.B1(n_95),
.B2(n_100),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_206),
.A2(n_210),
.B1(n_192),
.B2(n_170),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_102),
.B(n_107),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_207),
.B(n_212),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_122),
.A2(n_67),
.B1(n_111),
.B2(n_118),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_67),
.A2(n_110),
.B1(n_60),
.B2(n_61),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_62),
.B(n_66),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_126),
.Y(n_213)
);

INVx6_ASAP7_75t_L g303 ( 
.A(n_213),
.Y(n_303)
);

BUFx12f_ASAP7_75t_L g214 ( 
.A(n_148),
.Y(n_214)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_214),
.Y(n_312)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_166),
.Y(n_215)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_215),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_201),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_216),
.B(n_248),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_138),
.B(n_185),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_217),
.B(n_221),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_168),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_218),
.B(n_225),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_219),
.A2(n_259),
.B1(n_237),
.B2(n_220),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_169),
.B(n_176),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_126),
.Y(n_222)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_222),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_151),
.B(n_178),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_223),
.B(n_231),
.Y(n_294)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_163),
.Y(n_224)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_224),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_175),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_172),
.A2(n_142),
.B(n_141),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_227),
.A2(n_232),
.B(n_267),
.Y(n_288)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_166),
.Y(n_229)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_229),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_202),
.Y(n_230)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_230),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_147),
.B(n_149),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_150),
.A2(n_156),
.B1(n_170),
.B2(n_193),
.Y(n_232)
);

INVx8_ASAP7_75t_L g233 ( 
.A(n_200),
.Y(n_233)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_233),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_129),
.B(n_139),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_234),
.B(n_235),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_142),
.B(n_164),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_155),
.Y(n_236)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_236),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_238),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_131),
.B(n_137),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_240),
.B(n_245),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_197),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_242),
.B(n_247),
.Y(n_335)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_171),
.Y(n_243)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_243),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_134),
.B(n_135),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_200),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_160),
.B(n_159),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_160),
.B(n_173),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_249),
.B(n_250),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_155),
.B(n_189),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_251),
.B(n_258),
.Y(n_309)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_202),
.Y(n_252)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_252),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_143),
.B(n_196),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_253),
.B(n_255),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_136),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_254),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_128),
.B(n_208),
.Y(n_255)
);

AND2x6_ASAP7_75t_L g256 ( 
.A(n_132),
.B(n_133),
.Y(n_256)
);

AND2x6_ASAP7_75t_L g291 ( 
.A(n_256),
.B(n_271),
.Y(n_291)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_148),
.Y(n_257)
);

INVx6_ASAP7_75t_SL g310 ( 
.A(n_257),
.Y(n_310)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_128),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_259),
.B(n_260),
.Y(n_314)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_188),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_136),
.A2(n_157),
.B1(n_145),
.B2(n_194),
.Y(n_261)
);

OAI22x1_ASAP7_75t_L g322 ( 
.A1(n_261),
.A2(n_262),
.B1(n_280),
.B2(n_232),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_174),
.B(n_209),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_262),
.B(n_274),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_146),
.B(n_199),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_263),
.B(n_268),
.Y(n_337)
);

INVx13_ASAP7_75t_L g264 ( 
.A(n_162),
.Y(n_264)
);

INVx13_ASAP7_75t_L g290 ( 
.A(n_264),
.Y(n_290)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_171),
.Y(n_266)
);

INVx13_ASAP7_75t_L g304 ( 
.A(n_266),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_193),
.A2(n_199),
.B1(n_161),
.B2(n_190),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_146),
.B(n_203),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_203),
.Y(n_269)
);

INVx13_ASAP7_75t_L g307 ( 
.A(n_269),
.Y(n_307)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_197),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_270),
.B(n_272),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_177),
.B(n_144),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_246),
.C(n_239),
.Y(n_297)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_209),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_198),
.A2(n_180),
.B1(n_194),
.B2(n_157),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_273),
.A2(n_275),
.B1(n_282),
.B2(n_279),
.Y(n_323)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_174),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_145),
.A2(n_184),
.B1(n_162),
.B2(n_153),
.Y(n_275)
);

BUFx12f_ASAP7_75t_L g276 ( 
.A(n_162),
.Y(n_276)
);

INVx13_ASAP7_75t_L g320 ( 
.A(n_276),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_152),
.B(n_153),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_277),
.Y(n_289)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_152),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_278),
.B(n_283),
.Y(n_327)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_184),
.Y(n_279)
);

BUFx16f_ASAP7_75t_L g302 ( 
.A(n_279),
.Y(n_302)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_126),
.Y(n_280)
);

BUFx12_ASAP7_75t_L g295 ( 
.A(n_280),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_142),
.Y(n_281)
);

BUFx12_ASAP7_75t_L g333 ( 
.A(n_281),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_142),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_163),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_168),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_284),
.B(n_241),
.Y(n_334)
);

AO22x2_ASAP7_75t_L g285 ( 
.A1(n_140),
.A2(n_158),
.B1(n_167),
.B2(n_127),
.Y(n_285)
);

NOR2x1p5_ASAP7_75t_L g321 ( 
.A(n_285),
.B(n_283),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_291),
.B(n_233),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_216),
.B(n_251),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_293),
.B(n_297),
.C(n_306),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_281),
.A2(n_282),
.B(n_235),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_299),
.A2(n_332),
.B(n_215),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_226),
.A2(n_285),
.B1(n_251),
.B2(n_219),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_300),
.A2(n_301),
.B1(n_317),
.B2(n_321),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_227),
.B(n_226),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_285),
.A2(n_248),
.B1(n_249),
.B2(n_267),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_322),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_323),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_285),
.A2(n_256),
.B1(n_228),
.B2(n_250),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_326),
.A2(n_339),
.B1(n_314),
.B2(n_293),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_224),
.B(n_284),
.C(n_218),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_331),
.B(n_264),
.C(n_214),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_243),
.A2(n_266),
.B(n_244),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_334),
.B(n_260),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_242),
.A2(n_278),
.B1(n_274),
.B2(n_270),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_308),
.B(n_265),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_340),
.B(n_345),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_341),
.B(n_350),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_299),
.B(n_229),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_342),
.A2(n_336),
.B(n_313),
.Y(n_394)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_324),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_343),
.Y(n_407)
);

CKINVDCx14_ASAP7_75t_R g344 ( 
.A(n_288),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_344),
.B(n_353),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_321),
.B(n_236),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_321),
.B(n_272),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_346),
.B(n_351),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_296),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_347),
.B(n_349),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_348),
.A2(n_380),
.B(n_295),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_334),
.B(n_257),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_308),
.B(n_258),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_327),
.Y(n_352)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_352),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_327),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_301),
.A2(n_213),
.B1(n_254),
.B2(n_222),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_354),
.A2(n_366),
.B1(n_375),
.B2(n_376),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_328),
.A2(n_230),
.B(n_269),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_355),
.A2(n_379),
.B(n_320),
.Y(n_409)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_324),
.Y(n_356)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_356),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_331),
.B(n_214),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_358),
.B(n_363),
.Y(n_408)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_338),
.Y(n_359)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_359),
.Y(n_396)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_319),
.Y(n_360)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_360),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_361),
.B(n_325),
.C(n_312),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_326),
.B(n_252),
.Y(n_363)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_319),
.Y(n_365)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_365),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_314),
.A2(n_276),
.B1(n_317),
.B2(n_300),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_339),
.Y(n_368)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_368),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_286),
.B(n_276),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_369),
.B(n_372),
.Y(n_411)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_287),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_370),
.B(n_371),
.Y(n_390)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_310),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_305),
.B(n_337),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_294),
.B(n_292),
.Y(n_373)
);

OR2x2_ASAP7_75t_L g389 ( 
.A(n_373),
.B(n_298),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_288),
.A2(n_315),
.B(n_291),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_374),
.A2(n_333),
.B(n_313),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_314),
.A2(n_297),
.B1(n_316),
.B2(n_309),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_289),
.B(n_332),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_377),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_316),
.A2(n_309),
.B1(n_323),
.B2(n_315),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_378),
.A2(n_329),
.B1(n_330),
.B2(n_325),
.Y(n_395)
);

XNOR2x2_ASAP7_75t_SL g379 ( 
.A(n_306),
.B(n_309),
.Y(n_379)
);

A2O1A1O1Ixp25_ASAP7_75t_L g380 ( 
.A1(n_333),
.A2(n_335),
.B(n_310),
.C(n_311),
.D(n_322),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_383),
.A2(n_394),
.B(n_409),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_374),
.A2(n_333),
.B(n_336),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_387),
.A2(n_342),
.B(n_348),
.Y(n_428)
);

MAJx2_ASAP7_75t_L g388 ( 
.A(n_357),
.B(n_318),
.C(n_298),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_388),
.B(n_403),
.Y(n_429)
);

NAND3xp33_ASAP7_75t_L g430 ( 
.A(n_389),
.B(n_385),
.C(n_399),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_395),
.A2(n_400),
.B1(n_401),
.B2(n_402),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_397),
.B(n_404),
.C(n_413),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_367),
.A2(n_330),
.B1(n_302),
.B2(n_312),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_367),
.A2(n_302),
.B1(n_304),
.B2(n_303),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_366),
.A2(n_302),
.B1(n_304),
.B2(n_303),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_357),
.B(n_290),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_358),
.B(n_290),
.C(n_307),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_346),
.A2(n_295),
.B1(n_307),
.B2(n_320),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_405),
.A2(n_364),
.B1(n_368),
.B2(n_371),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_412),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_375),
.B(n_295),
.C(n_361),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_391),
.B(n_353),
.Y(n_414)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_414),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_415),
.B(n_426),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_399),
.B(n_373),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_419),
.B(n_431),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_403),
.B(n_379),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_420),
.B(n_408),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_392),
.A2(n_363),
.B1(n_345),
.B2(n_378),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_421),
.A2(n_433),
.B1(n_406),
.B2(n_384),
.Y(n_448)
);

A2O1A1Ixp33_ASAP7_75t_SL g422 ( 
.A1(n_412),
.A2(n_349),
.B(n_342),
.C(n_362),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_422),
.A2(n_430),
.B(n_387),
.Y(n_462)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_386),
.Y(n_423)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_423),
.Y(n_452)
);

OAI21x1_ASAP7_75t_L g424 ( 
.A1(n_381),
.A2(n_377),
.B(n_350),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_424),
.B(n_438),
.Y(n_467)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_386),
.Y(n_425)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_425),
.Y(n_456)
);

INVx4_ASAP7_75t_SL g426 ( 
.A(n_389),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_391),
.B(n_398),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_427),
.B(n_437),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_428),
.A2(n_409),
.B(n_383),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_396),
.B(n_372),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_390),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_432),
.B(n_435),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_392),
.A2(n_376),
.B1(n_362),
.B2(n_354),
.Y(n_433)
);

FAx1_ASAP7_75t_SL g434 ( 
.A(n_388),
.B(n_379),
.CI(n_340),
.CON(n_434),
.SN(n_434)
);

BUFx24_ASAP7_75t_SL g453 ( 
.A(n_434),
.Y(n_453)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_410),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_398),
.B(n_352),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_396),
.B(n_369),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_411),
.B(n_359),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_439),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_411),
.B(n_341),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_440),
.A2(n_382),
.B1(n_385),
.B2(n_365),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_413),
.B(n_349),
.C(n_360),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_441),
.B(n_429),
.C(n_420),
.Y(n_461)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_410),
.Y(n_442)
);

INVx13_ASAP7_75t_L g455 ( 
.A(n_442),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_443),
.B(n_390),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_433),
.A2(n_406),
.B1(n_384),
.B2(n_393),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_445),
.A2(n_466),
.B1(n_400),
.B2(n_401),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_448),
.A2(n_437),
.B1(n_432),
.B2(n_418),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_450),
.A2(n_462),
.B(n_464),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_436),
.B(n_388),
.C(n_397),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_451),
.B(n_459),
.C(n_460),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_457),
.B(n_434),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_436),
.B(n_408),
.C(n_404),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_441),
.B(n_381),
.C(n_382),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_461),
.B(n_463),
.C(n_428),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_429),
.B(n_351),
.C(n_355),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_417),
.A2(n_394),
.B(n_380),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_417),
.A2(n_389),
.B(n_395),
.Y(n_465)
);

CKINVDCx14_ASAP7_75t_R g477 ( 
.A(n_465),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_421),
.A2(n_426),
.B1(n_414),
.B2(n_427),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_468),
.A2(n_470),
.B1(n_485),
.B2(n_464),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_469),
.B(n_478),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_SL g470 ( 
.A1(n_447),
.A2(n_416),
.B1(n_364),
.B2(n_422),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_458),
.B(n_454),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_472),
.B(n_479),
.Y(n_488)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_452),
.Y(n_473)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_473),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_461),
.B(n_416),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_474),
.B(n_483),
.C(n_461),
.Y(n_495)
);

FAx1_ASAP7_75t_SL g475 ( 
.A(n_462),
.B(n_434),
.CI(n_422),
.CON(n_475),
.SN(n_475)
);

O2A1O1Ixp33_ASAP7_75t_L g498 ( 
.A1(n_475),
.A2(n_486),
.B(n_446),
.C(n_463),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_444),
.B(n_442),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_454),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_480),
.B(n_481),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_444),
.B(n_435),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_450),
.A2(n_422),
.B(n_415),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_482),
.B(n_484),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_451),
.B(n_425),
.C(n_423),
.Y(n_483)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_466),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_486),
.B(n_445),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_472),
.B(n_458),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_487),
.B(n_499),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_489),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_493),
.B(n_496),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_495),
.B(n_500),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_471),
.B(n_483),
.C(n_478),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_468),
.A2(n_447),
.B1(n_446),
.B2(n_467),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_497),
.A2(n_484),
.B1(n_485),
.B2(n_481),
.Y(n_510)
);

A2O1A1Ixp33_ASAP7_75t_L g503 ( 
.A1(n_498),
.A2(n_422),
.B(n_476),
.C(n_475),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_471),
.B(n_459),
.C(n_460),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_471),
.B(n_457),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_488),
.B(n_467),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_502),
.B(n_508),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_503),
.A2(n_504),
.B(n_505),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_498),
.A2(n_477),
.B(n_476),
.Y(n_504)
);

AOI21x1_ASAP7_75t_L g505 ( 
.A1(n_494),
.A2(n_470),
.B(n_482),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_499),
.B(n_443),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_493),
.A2(n_477),
.B(n_465),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_509),
.B(n_512),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_510),
.B(n_490),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_490),
.A2(n_479),
.B(n_453),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_506),
.B(n_496),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_513),
.B(n_515),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_502),
.B(n_497),
.Y(n_514)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_514),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_507),
.B(n_495),
.C(n_500),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_507),
.B(n_492),
.C(n_489),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_517),
.B(n_501),
.C(n_504),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_518),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_511),
.B(n_448),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_521),
.B(n_501),
.Y(n_523)
);

O2A1O1Ixp33_ASAP7_75t_SL g530 ( 
.A1(n_523),
.A2(n_519),
.B(n_456),
.C(n_452),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_516),
.Y(n_524)
);

AOI322xp5_ASAP7_75t_L g532 ( 
.A1(n_524),
.A2(n_527),
.A3(n_455),
.B1(n_449),
.B2(n_456),
.C1(n_475),
.C2(n_407),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_525),
.B(n_518),
.C(n_520),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_514),
.Y(n_527)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_529),
.Y(n_535)
);

AOI322xp5_ASAP7_75t_L g533 ( 
.A1(n_530),
.A2(n_531),
.A3(n_532),
.B1(n_522),
.B2(n_455),
.C1(n_527),
.C2(n_526),
.Y(n_533)
);

A2O1A1O1Ixp25_ASAP7_75t_L g531 ( 
.A1(n_528),
.A2(n_503),
.B(n_509),
.C(n_492),
.D(n_474),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_533),
.B(n_534),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_529),
.Y(n_534)
);

BUFx24_ASAP7_75t_SL g536 ( 
.A(n_535),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_536),
.A2(n_449),
.B(n_491),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_538),
.B(n_537),
.Y(n_539)
);


endmodule