module real_aes_4003_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_673;
wire n_905;
wire n_518;
wire n_254;
wire n_792;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_955;
wire n_889;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_961;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_478;
wire n_356;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_962;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_860;
wire n_748;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_960;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_142;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_957;
wire n_296;
wire n_954;
wire n_702;
wire n_969;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_965;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_720;
wire n_354;
wire n_265;
wire n_972;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_922;
wire n_149;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_959;
wire n_715;
wire n_134;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_166;
wire n_224;
wire n_839;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_967;
wire n_566;
wire n_719;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_968;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
OAI22xp5_ASAP7_75t_SL g543 ( .A1(n_0), .A2(n_17), .B1(n_544), .B2(n_545), .Y(n_543) );
CKINVDCx16_ASAP7_75t_R g545 ( .A(n_0), .Y(n_545) );
INVx1_ASAP7_75t_L g612 ( .A(n_1), .Y(n_612) );
INVx1_ASAP7_75t_L g308 ( .A(n_2), .Y(n_308) );
AOI22xp5_ASAP7_75t_L g278 ( .A1(n_3), .A2(n_22), .B1(n_215), .B2(n_258), .Y(n_278) );
AOI22x1_ASAP7_75t_SL g559 ( .A1(n_4), .A2(n_55), .B1(n_560), .B2(n_561), .Y(n_559) );
INVx1_ASAP7_75t_L g561 ( .A(n_4), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_5), .A2(n_558), .B1(n_562), .B2(n_563), .Y(n_557) );
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_5), .Y(n_562) );
INVx2_ASAP7_75t_L g165 ( .A(n_6), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_7), .B(n_625), .Y(n_723) );
INVx1_ASAP7_75t_SL g227 ( .A(n_8), .Y(n_227) );
INVxp67_ASAP7_75t_L g116 ( .A(n_9), .Y(n_116) );
BUFx2_ASAP7_75t_L g569 ( .A(n_9), .Y(n_569) );
INVx1_ASAP7_75t_L g959 ( .A(n_9), .Y(n_959) );
NAND2xp5_ASAP7_75t_SL g724 ( .A(n_10), .B(n_204), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_11), .A2(n_44), .B1(n_624), .B2(n_675), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_12), .A2(n_50), .B1(n_256), .B2(n_604), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_13), .A2(n_74), .B1(n_587), .B2(n_588), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_14), .B(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_15), .B(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g607 ( .A(n_16), .Y(n_607) );
INVx1_ASAP7_75t_L g544 ( .A(n_17), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_18), .A2(n_60), .B1(n_203), .B2(n_204), .Y(n_202) );
INVx1_ASAP7_75t_L g610 ( .A(n_19), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_20), .A2(n_542), .B1(n_543), .B2(n_546), .Y(n_541) );
CKINVDCx14_ASAP7_75t_R g546 ( .A(n_20), .Y(n_546) );
OA21x2_ASAP7_75t_L g144 ( .A1(n_21), .A2(n_78), .B(n_145), .Y(n_144) );
OA21x2_ASAP7_75t_L g197 ( .A1(n_21), .A2(n_78), .B(n_145), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_23), .A2(n_76), .B1(n_587), .B2(n_588), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_24), .B(n_161), .Y(n_268) );
AOI22xp5_ASAP7_75t_L g147 ( .A1(n_25), .A2(n_88), .B1(n_148), .B2(n_151), .Y(n_147) );
INVx2_ASAP7_75t_L g262 ( .A(n_26), .Y(n_262) );
INVx1_ASAP7_75t_L g603 ( .A(n_27), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g279 ( .A1(n_28), .A2(n_32), .B1(n_187), .B2(n_226), .Y(n_279) );
BUFx3_ASAP7_75t_L g111 ( .A(n_29), .Y(n_111) );
O2A1O1Ixp5_ASAP7_75t_L g255 ( .A1(n_30), .A2(n_185), .B(n_256), .C(n_257), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g157 ( .A1(n_31), .A2(n_71), .B1(n_158), .B2(n_160), .Y(n_157) );
OAI22xp5_ASAP7_75t_L g123 ( .A1(n_33), .A2(n_66), .B1(n_124), .B2(n_125), .Y(n_123) );
INVx1_ASAP7_75t_L g125 ( .A(n_33), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_34), .Y(n_189) );
AO22x1_ASAP7_75t_L g720 ( .A1(n_35), .A2(n_86), .B1(n_232), .B2(n_721), .Y(n_720) );
CKINVDCx5p33_ASAP7_75t_R g628 ( .A(n_36), .Y(n_628) );
AND2x2_ASAP7_75t_L g638 ( .A(n_37), .B(n_604), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_38), .B(n_232), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_39), .A2(n_89), .B1(n_212), .B2(n_214), .Y(n_211) );
INVx1_ASAP7_75t_L g121 ( .A(n_40), .Y(n_121) );
INVx1_ASAP7_75t_L g251 ( .A(n_41), .Y(n_251) );
AOI22x1_ASAP7_75t_L g660 ( .A1(n_42), .A2(n_102), .B1(n_587), .B2(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_43), .B(n_663), .Y(n_676) );
AND2x2_ASAP7_75t_L g967 ( .A(n_45), .B(n_968), .Y(n_967) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_46), .B(n_247), .Y(n_303) );
INVx2_ASAP7_75t_L g259 ( .A(n_47), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_48), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g646 ( .A(n_49), .B(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g267 ( .A(n_51), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_52), .B(n_301), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g551 ( .A(n_53), .Y(n_551) );
INVx1_ASAP7_75t_SL g231 ( .A(n_54), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_55), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_56), .B(n_226), .Y(n_692) );
INVx1_ASAP7_75t_L g181 ( .A(n_57), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_58), .B(n_253), .Y(n_631) );
INVx1_ASAP7_75t_L g145 ( .A(n_59), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g956 ( .A(n_61), .Y(n_956) );
AOI22xp5_ASAP7_75t_L g105 ( .A1(n_62), .A2(n_106), .B1(n_961), .B2(n_970), .Y(n_105) );
AND2x4_ASAP7_75t_L g139 ( .A(n_63), .B(n_140), .Y(n_139) );
AND2x4_ASAP7_75t_L g176 ( .A(n_63), .B(n_140), .Y(n_176) );
INVx1_ASAP7_75t_L g236 ( .A(n_64), .Y(n_236) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_65), .Y(n_156) );
INVx2_ASAP7_75t_L g124 ( .A(n_66), .Y(n_124) );
XOR2xp5_ASAP7_75t_SL g558 ( .A(n_67), .B(n_559), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_68), .A2(n_81), .B1(n_624), .B2(n_661), .Y(n_671) );
CKINVDCx14_ASAP7_75t_R g726 ( .A(n_69), .Y(n_726) );
AND2x2_ASAP7_75t_L g644 ( .A(n_70), .B(n_232), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_72), .B(n_229), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_73), .B(n_301), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_75), .B(n_295), .Y(n_686) );
NAND2x1p5_ASAP7_75t_L g648 ( .A(n_77), .B(n_591), .Y(n_648) );
CKINVDCx14_ASAP7_75t_R g665 ( .A(n_79), .Y(n_665) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_80), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_82), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_83), .B(n_625), .Y(n_690) );
OR2x6_ASAP7_75t_L g118 ( .A(n_84), .B(n_119), .Y(n_118) );
NAND3xp33_ASAP7_75t_L g966 ( .A(n_84), .B(n_116), .C(n_967), .Y(n_966) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_85), .B(n_152), .Y(n_233) );
INVx1_ASAP7_75t_L g120 ( .A(n_87), .Y(n_120) );
INVx1_ASAP7_75t_L g968 ( .A(n_90), .Y(n_968) );
INVx1_ASAP7_75t_L g150 ( .A(n_91), .Y(n_150) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_91), .Y(n_153) );
BUFx5_ASAP7_75t_L g188 ( .A(n_91), .Y(n_188) );
INVx2_ASAP7_75t_L g614 ( .A(n_92), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_93), .B(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g270 ( .A(n_94), .Y(n_270) );
INVx1_ASAP7_75t_L g274 ( .A(n_95), .Y(n_274) );
NAND2xp33_ASAP7_75t_L g640 ( .A(n_96), .B(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g195 ( .A(n_97), .Y(n_195) );
INVx2_ASAP7_75t_SL g140 ( .A(n_98), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_99), .B(n_178), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_100), .B(n_647), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_101), .B(n_295), .Y(n_294) );
AO32x2_ASAP7_75t_L g276 ( .A1(n_103), .A2(n_260), .A3(n_277), .B1(n_281), .B2(n_282), .Y(n_276) );
AO22x2_ASAP7_75t_L g313 ( .A1(n_103), .A2(n_277), .B1(n_314), .B2(n_316), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_104), .B(n_635), .Y(n_634) );
AO21x2_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_112), .B(n_554), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
BUFx3_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_111), .Y(n_565) );
OAI21x1_ASAP7_75t_SL g112 ( .A1(n_113), .A2(n_122), .B(n_549), .Y(n_112) );
INVx3_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
BUFx12f_ASAP7_75t_L g553 ( .A(n_114), .Y(n_553) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_117), .B(n_565), .Y(n_564) );
INVx8_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OR2x6_ASAP7_75t_L g958 ( .A(n_118), .B(n_959), .Y(n_958) );
HB1xp67_ASAP7_75t_L g969 ( .A(n_119), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
OAI22xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_126), .B1(n_127), .B2(n_548), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g548 ( .A(n_123), .Y(n_548) );
OR2x2_ASAP7_75t_L g589 ( .A(n_124), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AOI22xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_129), .B1(n_541), .B2(n_547), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
XNOR2x1_ASAP7_75t_L g570 ( .A(n_129), .B(n_545), .Y(n_570) );
AND2x4_ASAP7_75t_L g129 ( .A(n_130), .B(n_465), .Y(n_129) );
NOR2xp67_ASAP7_75t_L g130 ( .A(n_131), .B(n_387), .Y(n_130) );
NAND3xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_329), .C(n_366), .Y(n_131) );
AOI21xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_237), .B(n_283), .Y(n_132) );
OAI31xp33_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_167), .A3(n_198), .B(n_218), .Y(n_133) );
INVx1_ASAP7_75t_L g524 ( .A(n_134), .Y(n_524) );
BUFx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OR2x2_ASAP7_75t_L g361 ( .A(n_135), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g393 ( .A(n_135), .B(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_135), .B(n_320), .Y(n_407) );
AND2x2_ASAP7_75t_L g511 ( .A(n_135), .B(n_497), .Y(n_511) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g385 ( .A(n_136), .B(n_341), .Y(n_385) );
AND2x2_ASAP7_75t_L g424 ( .A(n_136), .B(n_321), .Y(n_424) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_136), .Y(n_458) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g338 ( .A(n_137), .Y(n_338) );
INVx1_ASAP7_75t_L g357 ( .A(n_137), .Y(n_357) );
AOI21x1_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_146), .B(n_164), .Y(n_137) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_141), .Y(n_138) );
INVx3_ASAP7_75t_L g207 ( .A(n_139), .Y(n_207) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_139), .Y(n_281) );
AND2x2_ASAP7_75t_L g314 ( .A(n_139), .B(n_315), .Y(n_314) );
INVx3_ASAP7_75t_L g585 ( .A(n_139), .Y(n_585) );
INVx1_ASAP7_75t_L g599 ( .A(n_139), .Y(n_599) );
AOI21xp33_ASAP7_75t_SL g651 ( .A1(n_141), .A2(n_584), .B(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_142), .B(n_207), .Y(n_223) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx3_ASAP7_75t_L g591 ( .A(n_143), .Y(n_591) );
INVx4_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g166 ( .A(n_144), .Y(n_166) );
BUFx3_ASAP7_75t_L g193 ( .A(n_144), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_154), .B1(n_157), .B2(n_162), .Y(n_146) );
INVx2_ASAP7_75t_L g721 ( .A(n_148), .Y(n_721) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g173 ( .A(n_149), .Y(n_173) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g159 ( .A(n_150), .Y(n_159) );
INVx1_ASAP7_75t_L g588 ( .A(n_151), .Y(n_588) );
INVx1_ASAP7_75t_L g675 ( .A(n_151), .Y(n_675) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g204 ( .A(n_152), .Y(n_204) );
INVx2_ASAP7_75t_L g226 ( .A(n_152), .Y(n_226) );
INVx1_ASAP7_75t_L g299 ( .A(n_152), .Y(n_299) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx6_ASAP7_75t_L g161 ( .A(n_153), .Y(n_161) );
INVx2_ASAP7_75t_L g179 ( .A(n_153), .Y(n_179) );
INVx2_ASAP7_75t_L g215 ( .A(n_153), .Y(n_215) );
AOI21x1_ASAP7_75t_L g719 ( .A1(n_154), .A2(n_720), .B(n_722), .Y(n_719) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_155), .B(n_206), .Y(n_205) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_155), .A2(n_225), .B(n_227), .C(n_228), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g269 ( .A1(n_155), .A2(n_173), .B(n_270), .C(n_271), .Y(n_269) );
INVx1_ASAP7_75t_L g280 ( .A(n_155), .Y(n_280) );
INVxp67_ASAP7_75t_L g633 ( .A(n_155), .Y(n_633) );
INVx2_ASAP7_75t_SL g650 ( .A(n_155), .Y(n_650) );
INVx1_ASAP7_75t_L g694 ( .A(n_155), .Y(n_694) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx3_ASAP7_75t_L g163 ( .A(n_156), .Y(n_163) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_156), .Y(n_185) );
INVx1_ASAP7_75t_L g217 ( .A(n_156), .Y(n_217) );
INVx4_ASAP7_75t_L g248 ( .A(n_156), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_156), .B(n_603), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_156), .B(n_607), .Y(n_606) );
INVxp67_ASAP7_75t_L g642 ( .A(n_156), .Y(n_642) );
INVx3_ASAP7_75t_L g256 ( .A(n_158), .Y(n_256) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g229 ( .A(n_159), .Y(n_229) );
INVx1_ASAP7_75t_L g266 ( .A(n_160), .Y(n_266) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g190 ( .A(n_161), .Y(n_190) );
INVx2_ASAP7_75t_L g245 ( .A(n_161), .Y(n_245) );
INVx2_ASAP7_75t_SL g258 ( .A(n_161), .Y(n_258) );
INVx1_ASAP7_75t_L g641 ( .A(n_161), .Y(n_641) );
INVx1_ASAP7_75t_L g647 ( .A(n_161), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_162), .B(n_175), .Y(n_174) );
NOR3xp33_ASAP7_75t_L g180 ( .A(n_162), .B(n_175), .C(n_181), .Y(n_180) );
NAND3xp33_ASAP7_75t_L g593 ( .A(n_162), .B(n_583), .C(n_584), .Y(n_593) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_163), .A2(n_231), .B(n_232), .C(n_233), .Y(n_230) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_163), .A2(n_266), .B(n_267), .C(n_268), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_165), .B(n_166), .Y(n_164) );
BUFx3_ASAP7_75t_L g260 ( .A(n_166), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_166), .B(n_262), .Y(n_261) );
INVx3_ASAP7_75t_L g295 ( .A(n_166), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_166), .B(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g348 ( .A(n_167), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_167), .B(n_349), .Y(n_441) );
BUFx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
OR2x2_ASAP7_75t_L g221 ( .A(n_168), .B(n_222), .Y(n_221) );
INVx2_ASAP7_75t_L g326 ( .A(n_168), .Y(n_326) );
AND2x2_ASAP7_75t_L g459 ( .A(n_168), .B(n_362), .Y(n_459) );
AO21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_192), .B(n_194), .Y(n_168) );
AO21x2_ASAP7_75t_L g289 ( .A1(n_169), .A2(n_194), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_170), .B(n_182), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_174), .B1(n_177), .B2(n_180), .Y(n_170) );
NOR2xp67_ASAP7_75t_L g171 ( .A(n_172), .B(n_173), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_175), .B(n_184), .Y(n_183) );
AOI221x1_ASAP7_75t_L g242 ( .A1(n_175), .A2(n_243), .B1(n_246), .B2(n_250), .C(n_252), .Y(n_242) );
INVx4_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g213 ( .A(n_179), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_183), .B(n_186), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_184), .B(n_627), .Y(n_626) );
OAI22x1_ASAP7_75t_L g657 ( .A1(n_184), .A2(n_658), .B1(n_659), .B2(n_660), .Y(n_657) );
INVx4_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
OAI22xp5_ASAP7_75t_L g277 ( .A1(n_185), .A2(n_278), .B1(n_279), .B2(n_280), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_185), .A2(n_298), .B(n_300), .Y(n_297) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_185), .A2(n_624), .B1(n_626), .B2(n_629), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_185), .B(n_670), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_185), .A2(n_689), .B(n_690), .Y(n_688) );
OAI22xp33_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_189), .B1(n_190), .B2(n_191), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g203 ( .A(n_188), .Y(n_203) );
INVx2_ASAP7_75t_L g232 ( .A(n_188), .Y(n_232) );
INVx2_ASAP7_75t_L g301 ( .A(n_188), .Y(n_301) );
INVx1_ASAP7_75t_L g305 ( .A(n_188), .Y(n_305) );
INVx2_ASAP7_75t_L g625 ( .A(n_188), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_190), .B(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g604 ( .A(n_190), .Y(n_604) );
NOR2xp67_ASAP7_75t_SL g664 ( .A(n_192), .B(n_665), .Y(n_664) );
OR2x2_ASAP7_75t_L g725 ( .A(n_192), .B(n_726), .Y(n_725) );
INVx3_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
OA21x2_ASAP7_75t_L g621 ( .A1(n_193), .A2(n_622), .B(n_634), .Y(n_621) );
OA21x2_ASAP7_75t_L g712 ( .A1(n_193), .A2(n_622), .B(n_634), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
INVx1_ASAP7_75t_L g282 ( .A(n_196), .Y(n_282) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NOR2xp67_ASAP7_75t_L g206 ( .A(n_197), .B(n_207), .Y(n_206) );
BUFx3_ASAP7_75t_L g209 ( .A(n_197), .Y(n_209) );
INVx1_ASAP7_75t_L g235 ( .A(n_197), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_197), .B(n_207), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_197), .B(n_207), .Y(n_309) );
INVx1_ASAP7_75t_L g315 ( .A(n_197), .Y(n_315) );
INVx2_ASAP7_75t_L g583 ( .A(n_197), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_197), .B(n_207), .Y(n_670) );
BUFx3_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g489 ( .A(n_199), .B(n_400), .Y(n_489) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g220 ( .A(n_200), .Y(n_220) );
INVx2_ASAP7_75t_L g325 ( .A(n_200), .Y(n_325) );
AND2x2_ASAP7_75t_L g344 ( .A(n_200), .B(n_293), .Y(n_344) );
AND2x2_ASAP7_75t_L g349 ( .A(n_200), .B(n_350), .Y(n_349) );
NAND2x1p5_ASAP7_75t_L g200 ( .A(n_201), .B(n_210), .Y(n_200) );
AND2x2_ASAP7_75t_SL g288 ( .A(n_201), .B(n_210), .Y(n_288) );
OA21x2_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_205), .B(n_208), .Y(n_201) );
INVx2_ASAP7_75t_L g587 ( .A(n_203), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_206), .B(n_217), .Y(n_216) );
OR2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_216), .Y(n_210) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVxp67_ASAP7_75t_SL g214 ( .A(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g253 ( .A(n_215), .Y(n_253) );
INVx1_ASAP7_75t_L g659 ( .A(n_217), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_217), .B(n_670), .Y(n_673) );
INVx2_ASAP7_75t_L g503 ( .A(n_218), .Y(n_503) );
OR2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_221), .Y(n_218) );
AND2x4_ASAP7_75t_L g428 ( .A(n_219), .B(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g443 ( .A(n_220), .B(n_327), .Y(n_443) );
INVx2_ASAP7_75t_L g405 ( .A(n_221), .Y(n_405) );
INVx1_ASAP7_75t_L g310 ( .A(n_222), .Y(n_310) );
INVx2_ASAP7_75t_L g328 ( .A(n_222), .Y(n_328) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_222), .Y(n_343) );
INVx2_ASAP7_75t_L g362 ( .A(n_222), .Y(n_362) );
AND2x2_ASAP7_75t_L g376 ( .A(n_222), .B(n_289), .Y(n_376) );
INVx1_ASAP7_75t_L g401 ( .A(n_222), .Y(n_401) );
AO31x2_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .A3(n_230), .B(n_234), .Y(n_222) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_232), .A2(n_253), .B1(n_609), .B2(n_611), .Y(n_608) );
NOR2xp33_ASAP7_75t_SL g234 ( .A(n_235), .B(n_236), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_235), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g663 ( .A(n_235), .Y(n_663) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_239), .B(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_275), .Y(n_239) );
AND2x2_ASAP7_75t_L g332 ( .A(n_240), .B(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g360 ( .A(n_240), .Y(n_360) );
INVx2_ASAP7_75t_L g418 ( .A(n_240), .Y(n_418) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_263), .Y(n_240) );
INVx2_ASAP7_75t_L g321 ( .A(n_241), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_241), .B(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g392 ( .A(n_241), .B(n_338), .Y(n_392) );
INVx1_ASAP7_75t_L g433 ( .A(n_241), .Y(n_433) );
AND2x2_ASAP7_75t_L g497 ( .A(n_241), .B(n_341), .Y(n_497) );
AO31x2_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_254), .A3(n_260), .B(n_261), .Y(n_241) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_249), .Y(n_246) );
AND2x2_ASAP7_75t_L g250 ( .A(n_247), .B(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_248), .B(n_308), .Y(n_307) );
NAND3xp33_ASAP7_75t_SL g582 ( .A(n_248), .B(n_583), .C(n_584), .Y(n_582) );
NOR2xp33_ASAP7_75t_SL g609 ( .A(n_248), .B(n_610), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_248), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_253), .B(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
INVx2_ASAP7_75t_L g316 ( .A(n_260), .Y(n_316) );
BUFx3_ASAP7_75t_L g317 ( .A(n_263), .Y(n_317) );
INVx2_ASAP7_75t_L g341 ( .A(n_263), .Y(n_341) );
AND2x4_ASAP7_75t_L g353 ( .A(n_263), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g395 ( .A(n_263), .Y(n_395) );
AND2x4_ASAP7_75t_L g432 ( .A(n_263), .B(n_433), .Y(n_432) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AO31x2_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_269), .A3(n_272), .B(n_273), .Y(n_264) );
INVx1_ASAP7_75t_L g408 ( .A(n_275), .Y(n_408) );
INVx2_ASAP7_75t_L g410 ( .A(n_275), .Y(n_410) );
AND2x4_ASAP7_75t_L g439 ( .A(n_275), .B(n_424), .Y(n_439) );
AND2x2_ASAP7_75t_L g505 ( .A(n_275), .B(n_506), .Y(n_505) );
BUFx8_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g354 ( .A(n_276), .Y(n_354) );
AND2x2_ASAP7_75t_L g369 ( .A(n_276), .B(n_370), .Y(n_369) );
OAI21x1_ASAP7_75t_L g622 ( .A1(n_281), .A2(n_623), .B(n_630), .Y(n_622) );
AO31x2_ASAP7_75t_L g656 ( .A1(n_281), .A2(n_657), .A3(n_662), .B(n_664), .Y(n_656) );
AO31x2_ASAP7_75t_L g700 ( .A1(n_281), .A2(n_657), .A3(n_662), .B(n_664), .Y(n_700) );
INVxp67_ASAP7_75t_L g290 ( .A(n_282), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_311), .B1(n_318), .B2(n_322), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_284), .B(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AOI211xp5_ASAP7_75t_L g484 ( .A1(n_285), .A2(n_367), .B(n_485), .C(n_491), .Y(n_484) );
AND2x4_ASAP7_75t_L g285 ( .A(n_286), .B(n_291), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
NOR2xp67_ASAP7_75t_SL g478 ( .A(n_287), .B(n_380), .Y(n_478) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g413 ( .A(n_288), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g420 ( .A(n_288), .B(n_414), .Y(n_420) );
INVx1_ASAP7_75t_L g526 ( .A(n_288), .Y(n_526) );
OR2x2_ASAP7_75t_L g365 ( .A(n_289), .B(n_350), .Y(n_365) );
AND2x2_ASAP7_75t_L g372 ( .A(n_289), .B(n_325), .Y(n_372) );
AND2x2_ASAP7_75t_L g490 ( .A(n_289), .B(n_292), .Y(n_490) );
AND2x2_ASAP7_75t_L g449 ( .A(n_291), .B(n_372), .Y(n_449) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_310), .Y(n_291) );
OR2x2_ASAP7_75t_L g380 ( .A(n_292), .B(n_326), .Y(n_380) );
INVx1_ASAP7_75t_L g474 ( .A(n_292), .Y(n_474) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g327 ( .A(n_293), .B(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g350 ( .A(n_293), .Y(n_350) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_293), .Y(n_402) );
INVx1_ASAP7_75t_L g414 ( .A(n_293), .Y(n_414) );
AND2x4_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
NOR2x1_ASAP7_75t_L g695 ( .A(n_295), .B(n_585), .Y(n_695) );
OAI21xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_302), .B(n_309), .Y(n_296) );
OAI21xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_304), .B(n_306), .Y(n_302) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVxp67_ASAP7_75t_L g386 ( .A(n_310), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_310), .B(n_500), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_311), .A2(n_406), .B(n_539), .C(n_540), .Y(n_538) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x4_ASAP7_75t_L g312 ( .A(n_313), .B(n_317), .Y(n_312) );
INVx1_ASAP7_75t_L g333 ( .A(n_313), .Y(n_333) );
AND2x4_ASAP7_75t_L g340 ( .A(n_313), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g396 ( .A(n_313), .Y(n_396) );
AND2x2_ASAP7_75t_L g514 ( .A(n_313), .B(n_338), .Y(n_514) );
INVx2_ASAP7_75t_SL g390 ( .A(n_317), .Y(n_390) );
INVxp67_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_319), .B(n_390), .Y(n_462) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g381 ( .A(n_320), .B(n_354), .Y(n_381) );
INVx2_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g368 ( .A(n_321), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_321), .B(n_354), .Y(n_383) );
BUFx3_ASAP7_75t_L g481 ( .A(n_321), .Y(n_481) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_327), .Y(n_323) );
AOI22xp33_ASAP7_75t_SL g378 ( .A1(n_324), .A2(n_379), .B1(n_381), .B2(n_382), .Y(n_378) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_325), .Y(n_453) );
BUFx2_ASAP7_75t_L g500 ( .A(n_325), .Y(n_500) );
AND2x4_ASAP7_75t_L g437 ( .A(n_326), .B(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g371 ( .A(n_327), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g438 ( .A(n_328), .Y(n_438) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_342), .B(n_345), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_331), .B(n_334), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_332), .B(n_524), .Y(n_529) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_339), .Y(n_335) );
OAI21xp33_ASAP7_75t_SL g373 ( .A1(n_336), .A2(n_339), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g469 ( .A(n_336), .Y(n_469) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g506 ( .A(n_337), .Y(n_506) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_338), .Y(n_537) );
INVx4_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_340), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
AND2x2_ASAP7_75t_L g375 ( .A(n_344), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g456 ( .A(n_344), .Y(n_456) );
AND2x2_ASAP7_75t_L g504 ( .A(n_344), .B(n_459), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_351), .B1(n_358), .B2(n_363), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_348), .B(n_531), .Y(n_530) );
NAND2xp67_ASAP7_75t_L g404 ( .A(n_349), .B(n_405), .Y(n_404) );
BUFx3_ASAP7_75t_L g426 ( .A(n_349), .Y(n_426) );
AND2x2_ASAP7_75t_L g534 ( .A(n_349), .B(n_437), .Y(n_534) );
AND2x2_ASAP7_75t_L g540 ( .A(n_349), .B(n_376), .Y(n_540) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_353), .B(n_356), .Y(n_374) );
INVx2_ASAP7_75t_L g486 ( .A(n_353), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_354), .B(n_370), .Y(n_448) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
HB1xp67_ASAP7_75t_SL g421 ( .A(n_356), .Y(n_421) );
AND2x2_ASAP7_75t_L g522 ( .A(n_356), .B(n_432), .Y(n_522) );
BUFx3_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g370 ( .A(n_357), .Y(n_370) );
INVxp67_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
NOR2xp67_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVxp67_ASAP7_75t_SL g464 ( .A(n_362), .Y(n_464) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g509 ( .A(n_364), .B(n_489), .Y(n_509) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVxp67_ASAP7_75t_L g429 ( .A(n_365), .Y(n_429) );
OR2x6_ASAP7_75t_L g463 ( .A(n_365), .B(n_464), .Y(n_463) );
INVxp67_ASAP7_75t_SL g483 ( .A(n_365), .Y(n_483) );
AOI221xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_371), .B1(n_373), .B2(n_375), .C(n_377), .Y(n_366) );
AND2x4_ASAP7_75t_SL g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx1_ASAP7_75t_L g493 ( .A(n_369), .Y(n_493) );
AND2x4_ASAP7_75t_L g398 ( .A(n_372), .B(n_399), .Y(n_398) );
NOR3xp33_ASAP7_75t_L g377 ( .A(n_378), .B(n_384), .C(n_386), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVxp67_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g536 ( .A(n_383), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g480 ( .A(n_385), .B(n_481), .Y(n_480) );
NAND4xp25_ASAP7_75t_L g387 ( .A(n_388), .B(n_415), .C(n_431), .D(n_444), .Y(n_387) );
O2A1O1Ixp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_393), .B(n_397), .C(n_403), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g455 ( .A(n_390), .Y(n_455) );
OAI32xp33_ASAP7_75t_L g523 ( .A1(n_390), .A2(n_411), .A3(n_492), .B1(n_524), .B2(n_525), .Y(n_523) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OR2x2_ASAP7_75t_L g409 ( .A(n_392), .B(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g518 ( .A(n_392), .Y(n_518) );
INVx1_ASAP7_75t_L g454 ( .A(n_394), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_394), .B(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g539 ( .A(n_394), .B(n_481), .Y(n_539) );
AND2x4_ASAP7_75t_SL g394 ( .A(n_395), .B(n_396), .Y(n_394) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_402), .Y(n_399) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_400), .Y(n_412) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OAI32xp33_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_406), .A3(n_408), .B1(n_409), .B2(n_411), .Y(n_403) );
AND2x2_ASAP7_75t_L g419 ( .A(n_405), .B(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g470 ( .A(n_409), .Y(n_470) );
AND2x2_ASAP7_75t_L g496 ( .A(n_410), .B(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
INVx1_ASAP7_75t_L g531 ( .A(n_413), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_421), .B(n_422), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_419), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_418), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_418), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g436 ( .A(n_420), .B(n_437), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_425), .B1(n_427), .B2(n_430), .Y(n_422) );
NOR2xp33_ASAP7_75t_SL g461 ( .A(n_424), .B(n_447), .Y(n_461) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx3_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AOI21xp33_ASAP7_75t_L g485 ( .A1(n_430), .A2(n_486), .B(n_487), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_434), .B1(n_439), .B2(n_440), .Y(n_431) );
INVx2_ASAP7_75t_L g494 ( .A(n_432), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_432), .B(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AND2x4_ASAP7_75t_L g473 ( .A(n_437), .B(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g499 ( .A(n_437), .B(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AOI221xp5_ASAP7_75t_SL g444 ( .A1(n_445), .A2(n_449), .B1(n_450), .B2(n_457), .C(n_460), .Y(n_444) );
INVxp67_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_454), .B1(n_455), .B2(n_456), .Y(n_450) );
INVxp67_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_452), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AND2x4_ASAP7_75t_L g482 ( .A(n_453), .B(n_483), .Y(n_482) );
AND2x4_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
INVx2_ASAP7_75t_L g521 ( .A(n_459), .Y(n_521) );
NAND2x1p5_ASAP7_75t_L g525 ( .A(n_459), .B(n_526), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_462), .B(n_463), .Y(n_460) );
NOR2x1_ASAP7_75t_L g465 ( .A(n_466), .B(n_501), .Y(n_465) );
NAND3xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_475), .C(n_484), .Y(n_466) );
OAI21xp33_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_470), .B(n_471), .Y(n_467) );
CKINVDCx5p33_ASAP7_75t_R g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVxp67_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_479), .Y(n_476) );
AOI221xp5_ASAP7_75t_L g515 ( .A1(n_478), .A2(n_516), .B1(n_519), .B2(n_522), .C(n_523), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_482), .Y(n_479) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x4_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_495), .B(n_498), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g520 ( .A(n_500), .Y(n_520) );
NAND3xp33_ASAP7_75t_SL g501 ( .A(n_502), .B(n_515), .C(n_527), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_504), .B(n_505), .C(n_507), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_510), .B1(n_512), .B2(n_513), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
NOR2x1p5_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_530), .B(n_532), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_535), .B(n_538), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVxp33_ASAP7_75t_SL g547 ( .A(n_541), .Y(n_547) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVxp67_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
OAI21xp33_ASAP7_75t_L g954 ( .A1(n_550), .A2(n_955), .B(n_960), .Y(n_954) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
BUFx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OAI221xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_566), .B1(n_951), .B2(n_952), .C(n_953), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_564), .Y(n_555) );
INVxp33_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_R g952 ( .A(n_557), .B(n_564), .Y(n_952) );
INVxp33_ASAP7_75t_SL g563 ( .A(n_558), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g960 ( .A(n_565), .Y(n_960) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_571), .Y(n_566) );
HB1xp67_ASAP7_75t_L g951 ( .A(n_567), .Y(n_951) );
OR2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
BUFx8_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_569), .Y(n_572) );
OA21x2_ASAP7_75t_L g953 ( .A1(n_571), .A2(n_952), .B(n_954), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2x1p5_ASAP7_75t_L g574 ( .A(n_575), .B(n_825), .Y(n_574) );
NOR4xp75_ASAP7_75t_L g575 ( .A(n_576), .B(n_738), .C(n_756), .D(n_782), .Y(n_575) );
AO21x1_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_615), .B(n_706), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_579), .B(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g746 ( .A(n_579), .B(n_716), .Y(n_746) );
INVx2_ASAP7_75t_L g808 ( .A(n_579), .Y(n_808) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_595), .Y(n_579) );
INVx1_ASAP7_75t_L g680 ( .A(n_580), .Y(n_680) );
INVx1_ASAP7_75t_L g705 ( .A(n_580), .Y(n_705) );
AND2x2_ASAP7_75t_L g728 ( .A(n_580), .B(n_596), .Y(n_728) );
INVx1_ASAP7_75t_L g759 ( .A(n_580), .Y(n_759) );
INVx2_ASAP7_75t_L g791 ( .A(n_580), .Y(n_791) );
NOR2x1_ASAP7_75t_L g833 ( .A(n_580), .B(n_834), .Y(n_833) );
HB1xp67_ASAP7_75t_L g848 ( .A(n_580), .Y(n_848) );
AND2x2_ASAP7_75t_L g897 ( .A(n_580), .B(n_684), .Y(n_897) );
OR2x6_ASAP7_75t_L g580 ( .A(n_581), .B(n_592), .Y(n_580) );
OAI21x1_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_586), .B(n_589), .Y(n_581) );
INVx1_ASAP7_75t_L g598 ( .A(n_583), .Y(n_598) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g635 ( .A(n_590), .Y(n_635) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NOR2xp67_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
AND2x2_ASAP7_75t_L g790 ( .A(n_595), .B(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g795 ( .A(n_596), .B(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g815 ( .A(n_596), .Y(n_815) );
INVx1_ASAP7_75t_L g834 ( .A(n_596), .Y(n_834) );
AND2x2_ASAP7_75t_L g896 ( .A(n_596), .B(n_761), .Y(n_896) );
INVxp67_ASAP7_75t_L g926 ( .A(n_596), .Y(n_926) );
AO21x2_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_600), .B(n_613), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
OR2x2_ASAP7_75t_L g718 ( .A(n_599), .B(n_635), .Y(n_718) );
NAND3xp33_ASAP7_75t_SL g600 ( .A(n_601), .B(n_605), .C(n_608), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_677), .B1(n_696), .B2(n_703), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AND2x4_ASAP7_75t_L g617 ( .A(n_618), .B(n_653), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g867 ( .A(n_619), .Y(n_867) );
OR2x2_ASAP7_75t_L g949 ( .A(n_619), .B(n_781), .Y(n_949) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g780 ( .A(n_620), .B(n_781), .Y(n_780) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_636), .Y(n_620) );
AND2x2_ASAP7_75t_L g697 ( .A(n_621), .B(n_698), .Y(n_697) );
NAND2x1_ASAP7_75t_L g742 ( .A(n_621), .B(n_655), .Y(n_742) );
AND2x2_ASAP7_75t_L g877 ( .A(n_621), .B(n_667), .Y(n_877) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_632), .B(n_633), .Y(n_630) );
AND2x2_ASAP7_75t_L g707 ( .A(n_636), .B(n_700), .Y(n_707) );
AND2x4_ASAP7_75t_L g731 ( .A(n_636), .B(n_732), .Y(n_731) );
OR2x2_ASAP7_75t_L g850 ( .A(n_636), .B(n_700), .Y(n_850) );
AO21x2_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_643), .B(n_651), .Y(n_636) );
AO21x2_ASAP7_75t_L g702 ( .A1(n_637), .A2(n_643), .B(n_651), .Y(n_702) );
OAI21x1_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_639), .B(n_642), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g661 ( .A(n_641), .Y(n_661) );
OAI21x1_ASAP7_75t_SL g643 ( .A1(n_644), .A2(n_645), .B(n_649), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_648), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_648), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g652 ( .A(n_648), .Y(n_652) );
AOI21x1_ASAP7_75t_L g722 ( .A1(n_650), .A2(n_723), .B(n_724), .Y(n_722) );
AND2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_666), .Y(n_653) );
INVx2_ASAP7_75t_L g733 ( .A(n_654), .Y(n_733) );
INVx1_ASAP7_75t_L g765 ( .A(n_654), .Y(n_765) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g755 ( .A(n_655), .B(n_702), .Y(n_755) );
INVx1_ASAP7_75t_L g769 ( .A(n_655), .Y(n_769) );
AND2x2_ASAP7_75t_L g909 ( .A(n_655), .B(n_713), .Y(n_909) );
INVx3_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g781 ( .A(n_666), .Y(n_781) );
OR2x2_ASAP7_75t_L g893 ( .A(n_666), .B(n_742), .Y(n_893) );
INVx2_ASAP7_75t_L g901 ( .A(n_666), .Y(n_901) );
INVx2_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_672), .Y(n_667) );
NAND2x1p5_ASAP7_75t_L g698 ( .A(n_668), .B(n_672), .Y(n_698) );
OR2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_671), .Y(n_668) );
OA21x2_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_674), .B(n_676), .Y(n_672) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_681), .Y(n_678) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g816 ( .A(n_680), .B(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g841 ( .A(n_682), .B(n_801), .Y(n_841) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OR2x2_ASAP7_75t_L g775 ( .A(n_683), .B(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g716 ( .A(n_684), .B(n_717), .Y(n_716) );
INVx3_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx2_ASAP7_75t_L g737 ( .A(n_685), .Y(n_737) );
AND2x2_ASAP7_75t_L g760 ( .A(n_685), .B(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g772 ( .A(n_685), .B(n_717), .Y(n_772) );
AND2x4_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
OAI21x1_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_691), .B(n_695), .Y(n_687) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_693), .B(n_694), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_697), .B(n_699), .Y(n_696) );
AND2x2_ASAP7_75t_L g797 ( .A(n_697), .B(n_741), .Y(n_797) );
INVx1_ASAP7_75t_L g910 ( .A(n_697), .Y(n_910) );
AND2x2_ASAP7_75t_L g942 ( .A(n_697), .B(n_769), .Y(n_942) );
INVx2_ASAP7_75t_L g713 ( .A(n_698), .Y(n_713) );
AND2x2_ASAP7_75t_L g752 ( .A(n_698), .B(n_711), .Y(n_752) );
INVx1_ASAP7_75t_L g802 ( .A(n_698), .Y(n_802) );
INVx1_ASAP7_75t_L g854 ( .A(n_698), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_698), .B(n_821), .Y(n_862) );
BUFx3_ASAP7_75t_L g749 ( .A(n_699), .Y(n_749) );
NOR2xp67_ASAP7_75t_L g869 ( .A(n_699), .B(n_751), .Y(n_869) );
AND2x4_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
INVx1_ASAP7_75t_L g779 ( .A(n_700), .Y(n_779) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVxp67_ASAP7_75t_L g741 ( .A(n_702), .Y(n_741) );
INVx1_ASAP7_75t_L g821 ( .A(n_702), .Y(n_821) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g771 ( .A(n_704), .B(n_772), .Y(n_771) );
OR2x2_ASAP7_75t_L g774 ( .A(n_704), .B(n_775), .Y(n_774) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_704), .Y(n_803) );
OR2x2_ASAP7_75t_L g930 ( .A(n_704), .B(n_807), .Y(n_930) );
INVx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g793 ( .A(n_705), .B(n_794), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_705), .B(n_859), .Y(n_858) );
OAI32xp33_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_708), .A3(n_714), .B1(n_729), .B2(n_734), .Y(n_706) );
INVx2_ASAP7_75t_L g865 ( .A(n_707), .Y(n_865) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g892 ( .A(n_709), .Y(n_892) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVxp67_ASAP7_75t_L g812 ( .A(n_710), .Y(n_812) );
OR2x2_ASAP7_75t_L g819 ( .A(n_710), .B(n_820), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_711), .B(n_713), .Y(n_710) );
INVx1_ASAP7_75t_L g904 ( .A(n_711), .Y(n_904) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g732 ( .A(n_712), .Y(n_732) );
HB1xp67_ASAP7_75t_L g860 ( .A(n_712), .Y(n_860) );
INVx1_ASAP7_75t_L g754 ( .A(n_713), .Y(n_754) );
INVx2_ASAP7_75t_L g744 ( .A(n_714), .Y(n_744) );
OR2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_727), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AND2x4_ASAP7_75t_L g832 ( .A(n_716), .B(n_833), .Y(n_832) );
AND2x2_ASAP7_75t_L g919 ( .A(n_716), .B(n_790), .Y(n_919) );
INVx2_ASAP7_75t_SL g761 ( .A(n_717), .Y(n_761) );
OAI21x1_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_719), .B(n_725), .Y(n_717) );
OAI21xp5_ASAP7_75t_L g796 ( .A1(n_718), .A2(n_719), .B(n_725), .Y(n_796) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g868 ( .A(n_728), .B(n_772), .Y(n_868) );
NAND2x1_ASAP7_75t_SL g890 ( .A(n_728), .B(n_760), .Y(n_890) );
AND2x2_ASAP7_75t_L g899 ( .A(n_728), .B(n_788), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_728), .B(n_941), .Y(n_940) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_L g943 ( .A(n_730), .B(n_801), .Y(n_943) );
AND2x2_ASAP7_75t_L g730 ( .A(n_731), .B(n_733), .Y(n_730) );
AND2x4_ASAP7_75t_SL g768 ( .A(n_731), .B(n_769), .Y(n_768) );
BUFx3_ASAP7_75t_L g844 ( .A(n_731), .Y(n_844) );
INVxp67_ASAP7_75t_SL g837 ( .A(n_732), .Y(n_837) );
INVx1_ASAP7_75t_L g870 ( .A(n_734), .Y(n_870) );
AOI211xp5_ASAP7_75t_SL g857 ( .A1(n_735), .A2(n_769), .B(n_858), .C(n_860), .Y(n_857) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g814 ( .A(n_736), .B(n_815), .Y(n_814) );
OR2x2_ASAP7_75t_L g872 ( .A(n_736), .B(n_873), .Y(n_872) );
AND2x2_ASAP7_75t_L g939 ( .A(n_736), .B(n_790), .Y(n_939) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g823 ( .A(n_737), .B(n_759), .Y(n_823) );
OR2x2_ASAP7_75t_L g838 ( .A(n_737), .B(n_795), .Y(n_838) );
NOR2xp33_ASAP7_75t_L g925 ( .A(n_737), .B(n_926), .Y(n_925) );
OAI22xp5_ASAP7_75t_SL g738 ( .A1(n_739), .A2(n_743), .B1(n_745), .B2(n_747), .Y(n_738) );
OR2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_742), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
HB1xp67_ASAP7_75t_L g836 ( .A(n_741), .Y(n_836) );
AND3x2_ASAP7_75t_L g916 ( .A(n_741), .B(n_901), .C(n_904), .Y(n_916) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
OA21x2_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_750), .B(n_753), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g935 ( .A(n_750), .Y(n_935) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g766 ( .A(n_752), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
BUFx3_ASAP7_75t_L g830 ( .A(n_755), .Y(n_830) );
AND2x2_ASAP7_75t_L g900 ( .A(n_755), .B(n_901), .Y(n_900) );
OAI21xp5_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_762), .B(n_770), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
AND2x2_ASAP7_75t_L g880 ( .A(n_760), .B(n_790), .Y(n_880) );
INVx2_ASAP7_75t_L g888 ( .A(n_760), .Y(n_888) );
INVx1_ASAP7_75t_L g776 ( .A(n_761), .Y(n_776) );
INVx1_ASAP7_75t_L g805 ( .A(n_761), .Y(n_805) );
INVxp67_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
NAND2xp5_ASAP7_75t_SL g763 ( .A(n_764), .B(n_767), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g799 ( .A1(n_764), .A2(n_785), .B1(n_800), .B2(n_806), .Y(n_799) );
OR2x2_ASAP7_75t_L g764 ( .A(n_765), .B(n_766), .Y(n_764) );
OR2x2_ASAP7_75t_L g875 ( .A(n_765), .B(n_876), .Y(n_875) );
INVx2_ASAP7_75t_SL g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g785 ( .A(n_768), .Y(n_785) );
OAI21xp5_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_773), .B(n_777), .Y(n_770) );
INVx2_ASAP7_75t_L g807 ( .A(n_772), .Y(n_807) );
AND2x2_ASAP7_75t_L g852 ( .A(n_772), .B(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
OAI22xp5_ASAP7_75t_L g902 ( .A1(n_774), .A2(n_875), .B1(n_903), .B2(n_905), .Y(n_902) );
INVxp67_ASAP7_75t_SL g788 ( .A(n_776), .Y(n_788) );
AND2x2_ASAP7_75t_L g777 ( .A(n_778), .B(n_780), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_778), .B(n_812), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_778), .B(n_892), .Y(n_891) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
NAND3x1_ASAP7_75t_L g782 ( .A(n_783), .B(n_798), .C(n_809), .Y(n_782) );
AOI21x1_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_786), .B(n_792), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
OAI22xp5_ASAP7_75t_L g948 ( .A1(n_787), .A2(n_872), .B1(n_949), .B2(n_950), .Y(n_948) );
OR2x2_ASAP7_75t_L g787 ( .A(n_788), .B(n_789), .Y(n_787) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
AND2x2_ASAP7_75t_L g792 ( .A(n_793), .B(n_797), .Y(n_792) );
INVx1_ASAP7_75t_L g842 ( .A(n_794), .Y(n_842) );
AND2x2_ASAP7_75t_L g922 ( .A(n_794), .B(n_848), .Y(n_922) );
INVx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g824 ( .A(n_795), .Y(n_824) );
BUFx2_ASAP7_75t_L g817 ( .A(n_796), .Y(n_817) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
NAND3xp33_ASAP7_75t_L g800 ( .A(n_801), .B(n_803), .C(n_804), .Y(n_800) );
INVx2_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
AND2x2_ASAP7_75t_L g856 ( .A(n_805), .B(n_815), .Y(n_856) );
OR2x2_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
INVxp67_ASAP7_75t_L g846 ( .A(n_808), .Y(n_846) );
AOI22xp5_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_813), .B1(n_818), .B2(n_822), .Y(n_809) );
INVx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
NAND3xp33_ASAP7_75t_SL g864 ( .A(n_811), .B(n_865), .C(n_866), .Y(n_864) );
AND2x2_ASAP7_75t_L g813 ( .A(n_814), .B(n_816), .Y(n_813) );
AND2x2_ASAP7_75t_L g924 ( .A(n_816), .B(n_925), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g945 ( .A(n_816), .B(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g859 ( .A(n_817), .Y(n_859) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_820), .B(n_854), .Y(n_950) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g845 ( .A1(n_821), .A2(n_846), .B1(n_847), .B2(n_849), .Y(n_845) );
AND2x2_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .Y(n_822) );
NAND2x2_ASAP7_75t_L g933 ( .A(n_823), .B(n_934), .Y(n_933) );
NOR2x1_ASAP7_75t_L g825 ( .A(n_826), .B(n_911), .Y(n_825) );
NAND4xp25_ASAP7_75t_L g826 ( .A(n_827), .B(n_863), .C(n_878), .D(n_898), .Y(n_826) );
NOR2xp67_ASAP7_75t_L g827 ( .A(n_828), .B(n_839), .Y(n_827) );
OAI22xp5_ASAP7_75t_L g828 ( .A1(n_829), .A2(n_831), .B1(n_835), .B2(n_838), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
AOI21xp33_ASAP7_75t_L g920 ( .A1(n_831), .A2(n_843), .B(n_921), .Y(n_920) );
INVx2_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx2_ASAP7_75t_L g873 ( .A(n_833), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_836), .B(n_837), .Y(n_835) );
OAI211xp5_ASAP7_75t_SL g855 ( .A1(n_837), .A2(n_856), .B(n_857), .C(n_861), .Y(n_855) );
INVx1_ASAP7_75t_L g882 ( .A(n_837), .Y(n_882) );
AOI21xp33_ASAP7_75t_L g907 ( .A1(n_838), .A2(n_908), .B(n_910), .Y(n_907) );
OAI321xp33_ASAP7_75t_L g839 ( .A1(n_840), .A2(n_842), .A3(n_843), .B1(n_845), .B2(n_851), .C(n_855), .Y(n_839) );
INVx2_ASAP7_75t_SL g840 ( .A(n_841), .Y(n_840) );
OR2x2_ASAP7_75t_L g905 ( .A(n_842), .B(n_906), .Y(n_905) );
INVx2_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_844), .B(n_885), .Y(n_884) );
NOR2x1_ASAP7_75t_R g927 ( .A(n_844), .B(n_908), .Y(n_927) );
HB1xp67_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
AND2x2_ASAP7_75t_L g928 ( .A(n_849), .B(n_877), .Y(n_928) );
INVx2_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
OR2x2_ASAP7_75t_L g903 ( .A(n_850), .B(n_904), .Y(n_903) );
INVx2_ASAP7_75t_L g915 ( .A(n_850), .Y(n_915) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g885 ( .A(n_854), .Y(n_885) );
INVxp67_ASAP7_75t_L g941 ( .A(n_859), .Y(n_941) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
AOI222xp33_ASAP7_75t_L g863 ( .A1(n_864), .A2(n_868), .B1(n_869), .B2(n_870), .C1(n_871), .C2(n_874), .Y(n_863) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g932 ( .A(n_867), .Y(n_932) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
OR2x2_ASAP7_75t_L g887 ( .A(n_873), .B(n_888), .Y(n_887) );
INVx2_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
AOI221x1_ASAP7_75t_L g878 ( .A1(n_879), .A2(n_881), .B1(n_883), .B2(n_886), .C(n_889), .Y(n_878) );
HB1xp67_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
OAI22xp33_ASAP7_75t_SL g889 ( .A1(n_890), .A2(n_891), .B1(n_893), .B2(n_894), .Y(n_889) );
INVx2_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
AND2x4_ASAP7_75t_L g895 ( .A(n_896), .B(n_897), .Y(n_895) );
BUFx3_ASAP7_75t_L g934 ( .A(n_896), .Y(n_934) );
INVx2_ASAP7_75t_L g906 ( .A(n_897), .Y(n_906) );
AOI211xp5_ASAP7_75t_L g898 ( .A1(n_899), .A2(n_900), .B(n_902), .C(n_907), .Y(n_898) );
NAND2x1_ASAP7_75t_L g914 ( .A(n_901), .B(n_915), .Y(n_914) );
OAI22xp5_ASAP7_75t_SL g931 ( .A1(n_905), .A2(n_932), .B1(n_933), .B2(n_935), .Y(n_931) );
INVx2_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
NAND3xp33_ASAP7_75t_SL g911 ( .A(n_912), .B(n_923), .C(n_936), .Y(n_911) );
O2A1O1Ixp33_ASAP7_75t_L g912 ( .A1(n_913), .A2(n_916), .B(n_917), .C(n_920), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
INVx2_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
INVx2_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
AOI221xp5_ASAP7_75t_L g923 ( .A1(n_924), .A2(n_927), .B1(n_928), .B2(n_929), .C(n_931), .Y(n_923) );
HB1xp67_ASAP7_75t_L g947 ( .A(n_926), .Y(n_947) );
INVxp67_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
AOI221xp5_ASAP7_75t_L g936 ( .A1(n_937), .A2(n_942), .B1(n_943), .B2(n_944), .C(n_948), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g937 ( .A(n_938), .B(n_940), .Y(n_937) );
INVx2_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
INVxp67_ASAP7_75t_SL g944 ( .A(n_945), .Y(n_944) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
NOR2xp33_ASAP7_75t_L g955 ( .A(n_956), .B(n_957), .Y(n_955) );
HB1xp67_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
CKINVDCx5p33_ASAP7_75t_R g961 ( .A(n_962), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
INVx1_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
BUFx5_ASAP7_75t_L g972 ( .A(n_964), .Y(n_972) );
BUFx3_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
OR2x2_ASAP7_75t_L g965 ( .A(n_966), .B(n_969), .Y(n_965) );
CKINVDCx5p33_ASAP7_75t_R g970 ( .A(n_971), .Y(n_970) );
CKINVDCx5p33_ASAP7_75t_R g971 ( .A(n_972), .Y(n_971) );
endmodule