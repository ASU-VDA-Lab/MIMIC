module fake_jpeg_24359_n_58 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_58);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_58;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_16;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_56;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx16f_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_6),
.B(n_2),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx11_ASAP7_75t_SL g16 ( 
.A(n_7),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_0),
.C(n_1),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_23),
.C(n_15),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_2),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_19),
.B(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_22),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_9),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_14),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_26),
.B(n_29),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_23),
.B(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_19),
.B(n_10),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_8),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_12),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_37),
.C(n_29),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_36),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_9),
.Y(n_37)
);

OA21x2_ASAP7_75t_L g39 ( 
.A1(n_28),
.A2(n_20),
.B(n_21),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_20),
.B(n_21),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_43),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_SL g43 ( 
.A(n_39),
.B(n_5),
.C(n_7),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_32),
.B1(n_38),
.B2(n_33),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_49),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_47),
.B(n_24),
.Y(n_52)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_45),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_48),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_53),
.B(n_51),
.Y(n_55)
);

OAI311xp33_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_50),
.A3(n_54),
.B1(n_40),
.C1(n_42),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_25),
.B(n_16),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_25),
.Y(n_58)
);


endmodule