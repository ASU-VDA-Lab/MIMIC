module fake_jpeg_17667_n_231 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_231);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_22),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_39),
.Y(n_48)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_25),
.Y(n_33)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_38),
.A2(n_15),
.B1(n_16),
.B2(n_20),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_42),
.A2(n_44),
.B1(n_45),
.B2(n_54),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_32),
.A2(n_20),
.B1(n_15),
.B2(n_21),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_36),
.A2(n_15),
.B1(n_23),
.B2(n_21),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_16),
.B1(n_23),
.B2(n_21),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_46),
.A2(n_50),
.B1(n_51),
.B2(n_55),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_0),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_49),
.A2(n_57),
.B1(n_29),
.B2(n_26),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_16),
.B1(n_23),
.B2(n_20),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_34),
.A2(n_30),
.B1(n_19),
.B2(n_17),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_35),
.A2(n_30),
.B1(n_19),
.B2(n_17),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_34),
.A2(n_30),
.B1(n_19),
.B2(n_17),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_1),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_35),
.A2(n_29),
.B1(n_26),
.B2(n_22),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_61),
.A2(n_29),
.B1(n_26),
.B2(n_33),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_61),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_76),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_22),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_64),
.B(n_73),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_71),
.Y(n_102)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_27),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_80),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_55),
.B1(n_60),
.B2(n_53),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_69),
.A2(n_42),
.B1(n_41),
.B2(n_57),
.Y(n_90)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_40),
.C(n_33),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_40),
.C(n_58),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_33),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_56),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_56),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_83),
.Y(n_98)
);

OAI32xp33_ASAP7_75t_L g80 ( 
.A1(n_49),
.A2(n_18),
.A3(n_28),
.B1(n_40),
.B2(n_41),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_57),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_57),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_52),
.Y(n_83)
);

NAND3xp33_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_9),
.C(n_12),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_84),
.A2(n_47),
.B1(n_10),
.B2(n_3),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_59),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_85),
.B(n_83),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_88),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_90),
.A2(n_94),
.B1(n_78),
.B2(n_84),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_75),
.A2(n_47),
.B1(n_11),
.B2(n_4),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_66),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_97),
.B(n_79),
.Y(n_120)
);

CKINVDCx10_ASAP7_75t_R g100 ( 
.A(n_67),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_107),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_64),
.B(n_58),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_108),
.Y(n_119)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_47),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_68),
.B(n_1),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_106),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_89),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_118),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_95),
.B(n_71),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_113),
.B(n_132),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_72),
.C(n_63),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_117),
.C(n_95),
.Y(n_137)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

AND2x4_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_80),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_116),
.A2(n_120),
.B(n_131),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_76),
.C(n_73),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_92),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_97),
.A2(n_86),
.B1(n_91),
.B2(n_90),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_126),
.B1(n_102),
.B2(n_74),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_99),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_124),
.Y(n_151)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_79),
.B1(n_85),
.B2(n_81),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_92),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_127),
.B(n_77),
.Y(n_146)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

XNOR2x1_ASAP7_75t_L g131 ( 
.A(n_86),
.B(n_40),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_88),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_137),
.C(n_141),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_112),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_136),
.A2(n_143),
.B(n_148),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_131),
.A2(n_98),
.B1(n_102),
.B2(n_109),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_138),
.A2(n_150),
.B1(n_129),
.B2(n_59),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_99),
.C(n_103),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_102),
.B(n_103),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_96),
.Y(n_145)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_125),
.A2(n_93),
.B1(n_107),
.B2(n_104),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_116),
.A2(n_59),
.B1(n_65),
.B2(n_105),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_111),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_134),
.A2(n_115),
.B1(n_126),
.B2(n_122),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_156),
.A2(n_169),
.B1(n_148),
.B2(n_143),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_126),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_152),
.Y(n_161)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_161),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_118),
.C(n_126),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_133),
.C(n_137),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_165),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_146),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_128),
.Y(n_166)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_153),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_167),
.A2(n_144),
.B1(n_151),
.B2(n_136),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_128),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_147),
.Y(n_178)
);

AOI322xp5_ASAP7_75t_SL g170 ( 
.A1(n_149),
.A2(n_9),
.A3(n_11),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_170),
.B(n_12),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_179),
.C(n_183),
.Y(n_192)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_162),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_174),
.A2(n_170),
.B(n_157),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_141),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_181),
.Y(n_188)
);

OAI22x1_ASAP7_75t_L g176 ( 
.A1(n_156),
.A2(n_142),
.B1(n_150),
.B2(n_135),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_176),
.A2(n_182),
.B1(n_165),
.B2(n_166),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_185),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_135),
.C(n_149),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_147),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_154),
.A2(n_151),
.B1(n_144),
.B2(n_18),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_105),
.C(n_62),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_155),
.C(n_157),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_180),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_186),
.A2(n_194),
.B1(n_195),
.B2(n_9),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_164),
.Y(n_187)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_174),
.Y(n_201)
);

OAI31xp33_ASAP7_75t_L g191 ( 
.A1(n_176),
.A2(n_160),
.A3(n_161),
.B(n_155),
.Y(n_191)
);

A2O1A1O1Ixp25_ASAP7_75t_L g196 ( 
.A1(n_179),
.A2(n_160),
.B(n_185),
.C(n_181),
.D(n_171),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_196),
.B(n_197),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_178),
.A2(n_168),
.B(n_169),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_175),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_200),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_184),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_201),
.B(n_204),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_177),
.C(n_164),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_186),
.Y(n_208)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_203),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_189),
.A2(n_8),
.B1(n_12),
.B2(n_4),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_193),
.A2(n_10),
.B1(n_11),
.B2(n_5),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_205),
.B(n_6),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_209),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_192),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_198),
.A2(n_194),
.B(n_196),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_211),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_191),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_203),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_217),
.Y(n_222)
);

INVx11_ASAP7_75t_L g216 ( 
.A(n_213),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_199),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_200),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_202),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_214),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_207),
.Y(n_221)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_221),
.Y(n_227)
);

AOI322xp5_ASAP7_75t_L g225 ( 
.A1(n_223),
.A2(n_218),
.A3(n_216),
.B1(n_215),
.B2(n_220),
.C1(n_217),
.C2(n_105),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_224),
.A2(n_1),
.B(n_2),
.Y(n_226)
);

OAI211xp5_ASAP7_75t_L g228 ( 
.A1(n_225),
.A2(n_226),
.B(n_222),
.C(n_2),
.Y(n_228)
);

BUFx24_ASAP7_75t_SL g229 ( 
.A(n_228),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_229),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_227),
.Y(n_231)
);


endmodule