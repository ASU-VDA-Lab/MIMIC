module real_jpeg_15842_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_466),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_0),
.B(n_467),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_1),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_67)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_1),
.A2(n_176),
.B1(n_179),
.B2(n_180),
.Y(n_175)
);

OAI32xp33_ASAP7_75t_L g190 ( 
.A1(n_1),
.A2(n_123),
.A3(n_191),
.B1(n_192),
.B2(n_195),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_1),
.A2(n_201),
.B1(n_202),
.B2(n_205),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_1),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_1),
.B(n_151),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_1),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_1),
.B(n_317),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_2),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_63)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_2),
.A2(n_66),
.B1(n_116),
.B2(n_221),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_L g231 ( 
.A1(n_2),
.A2(n_66),
.B1(n_232),
.B2(n_235),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_2),
.A2(n_66),
.B1(n_245),
.B2(n_248),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_3),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_3),
.Y(n_95)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_3),
.Y(n_267)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_3),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_4),
.Y(n_126)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_4),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_4),
.Y(n_135)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_5),
.A2(n_109),
.B1(n_110),
.B2(n_115),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g211 ( 
.A(n_6),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_6),
.Y(n_217)
);

BUFx5_ASAP7_75t_L g254 ( 
.A(n_6),
.Y(n_254)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_6),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_7),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_7),
.Y(n_97)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_7),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_7),
.Y(n_138)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_7),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_7),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_8),
.A2(n_55),
.B1(n_58),
.B2(n_59),
.Y(n_54)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_8),
.A2(n_59),
.B1(n_99),
.B2(n_102),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_8),
.A2(n_59),
.B1(n_143),
.B2(n_145),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g365 ( 
.A1(n_8),
.A2(n_59),
.B1(n_366),
.B2(n_370),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_9),
.Y(n_467)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_11),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_12),
.Y(n_80)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_12),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g204 ( 
.A(n_12),
.Y(n_204)
);

BUFx4f_ASAP7_75t_L g369 ( 
.A(n_12),
.Y(n_369)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_13),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_160),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_159),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_60),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_19),
.B(n_60),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_34),
.B1(n_42),
.B2(n_54),
.Y(n_19)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_20),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_21),
.A2(n_34),
.B1(n_63),
.B2(n_67),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g170 ( 
.A1(n_21),
.A2(n_34),
.B1(n_63),
.B2(n_67),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_21),
.B(n_34),
.Y(n_391)
);

OAI21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_29),
.B(n_34),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_22),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_26),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_31),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g349 ( 
.A(n_33),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_34),
.A2(n_42),
.B(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_34),
.Y(n_317)
);

OA22x2_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_40),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_47),
.B1(n_49),
.B2(n_53),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_47),
.A2(n_48),
.B1(n_360),
.B2(n_363),
.Y(n_359)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_53),
.A2(n_197),
.B1(n_381),
.B2(n_382),
.Y(n_380)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_152),
.C(n_156),
.Y(n_60)
);

FAx1_ASAP7_75t_SL g181 ( 
.A(n_61),
.B(n_152),
.CI(n_156),
.CON(n_181),
.SN(n_181)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_74),
.C(n_107),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_62),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_62),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_62),
.B(n_219),
.C(n_357),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_62),
.A2(n_166),
.B1(n_219),
.B2(n_237),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_62),
.B(n_312),
.C(n_419),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_62),
.A2(n_166),
.B1(n_312),
.B2(n_318),
.Y(n_427)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_67),
.Y(n_154)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_70),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_70),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_70),
.B(n_230),
.Y(n_229)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_74),
.B(n_107),
.Y(n_168)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_74),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_74),
.B(n_173),
.Y(n_451)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_98),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_85),
.Y(n_75)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_76),
.Y(n_296)
);

AOI21x1_ASAP7_75t_SL g328 ( 
.A1(n_76),
.A2(n_329),
.B(n_331),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_76),
.A2(n_380),
.B(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NOR2x1_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_87),
.Y(n_86)
);

AO22x2_ASAP7_75t_L g223 ( 
.A1(n_77),
.A2(n_86),
.B1(n_224),
.B2(n_231),
.Y(n_223)
);

AO22x1_ASAP7_75t_L g241 ( 
.A1(n_77),
.A2(n_86),
.B1(n_224),
.B2(n_231),
.Y(n_241)
);

AO22x2_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_81),
.B2(n_84),
.Y(n_77)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_79),
.Y(n_212)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_80),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_81),
.Y(n_364)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_83),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_85),
.Y(n_385)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_86),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_91),
.B1(n_93),
.B2(n_96),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_89),
.Y(n_236)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_90),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_96),
.Y(n_191)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_96),
.Y(n_197)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_98),
.A2(n_296),
.B1(n_379),
.B2(n_385),
.Y(n_378)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_106),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_120),
.B1(n_142),
.B2(n_151),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_108),
.A2(n_120),
.B1(n_151),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_109),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_110),
.A2(n_337),
.B1(n_346),
.B2(n_350),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_114),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g345 ( 
.A(n_114),
.Y(n_345)
);

BUFx2_ASAP7_75t_SL g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_118),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

OA22x2_ASAP7_75t_L g219 ( 
.A1(n_121),
.A2(n_133),
.B1(n_175),
.B2(n_220),
.Y(n_219)
);

OA22x2_ASAP7_75t_L g312 ( 
.A1(n_121),
.A2(n_133),
.B1(n_175),
.B2(n_220),
.Y(n_312)
);

AO21x1_ASAP7_75t_L g411 ( 
.A1(n_121),
.A2(n_133),
.B(n_175),
.Y(n_411)
);

NAND2x1p5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_133),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_128),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_127),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_132),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_133),
.B(n_158),
.Y(n_157)
);

OA22x2_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_136),
.B1(n_139),
.B2(n_140),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_138),
.Y(n_263)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_154),
.B(n_391),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_182),
.B(n_464),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_181),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_163),
.B(n_181),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_169),
.C(n_171),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_L g448 ( 
.A1(n_164),
.A2(n_165),
.B1(n_169),
.B2(n_170),
.Y(n_448)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_172),
.C(n_173),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_169),
.B(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_169),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_169),
.B(n_237),
.C(n_328),
.Y(n_433)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_170),
.B(n_411),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_170),
.B(n_451),
.Y(n_450)
);

XOR2x2_ASAP7_75t_L g447 ( 
.A(n_171),
.B(n_448),
.Y(n_447)
);

INVxp33_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_179),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_179),
.B(n_347),
.Y(n_346)
);

BUFx24_ASAP7_75t_SL g469 ( 
.A(n_181),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_445),
.B(n_461),
.Y(n_182)
);

AO221x1_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_352),
.B1(n_354),
.B2(n_438),
.C(n_444),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_322),
.B(n_351),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_305),
.B(n_321),
.Y(n_185)
);

OAI21x1_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_256),
.B(n_304),
.Y(n_186)
);

NOR2xp67_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_239),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_188),
.B(n_239),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_218),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_189),
.B(n_223),
.C(n_237),
.Y(n_320)
);

XOR2x2_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_198),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_190),
.B(n_198),
.Y(n_308)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_208),
.Y(n_198)
);

OA22x2_ASAP7_75t_L g242 ( 
.A1(n_199),
.A2(n_243),
.B1(n_244),
.B2(n_251),
.Y(n_242)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_200),
.B(n_209),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_201),
.A2(n_225),
.B(n_229),
.Y(n_224)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_204),
.Y(n_207)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_204),
.Y(n_247)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_204),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_204),
.Y(n_370)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g389 ( 
.A(n_208),
.B(n_365),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_213),
.Y(n_208)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_209),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI32xp33_ASAP7_75t_L g259 ( 
.A1(n_212),
.A2(n_229),
.A3(n_260),
.B1(n_264),
.B2(n_268),
.Y(n_259)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g288 ( 
.A(n_214),
.Y(n_288)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_223),
.B1(n_237),
.B2(n_238),
.Y(n_218)
);

INVx3_ASAP7_75t_SL g237 ( 
.A(n_219),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_219),
.A2(n_237),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_223),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_223),
.A2(n_238),
.B1(n_259),
.B2(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_223),
.B(n_405),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_223),
.A2(n_238),
.B1(n_405),
.B2(n_431),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_224),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_224),
.B(n_330),
.Y(n_396)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.C(n_255),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_240),
.A2(n_241),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_240),
.B(n_308),
.C(n_310),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_240),
.A2(n_241),
.B1(n_358),
.B2(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_241),
.B(n_255),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_241),
.B(n_358),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_242),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_242),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_242),
.B(n_294),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_242),
.B(n_294),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_242),
.A2(n_275),
.B1(n_335),
.B2(n_336),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_243),
.A2(n_359),
.B1(n_365),
.B2(n_371),
.Y(n_358)
);

OA21x2_ASAP7_75t_L g289 ( 
.A1(n_244),
.A2(n_290),
.B(n_292),
.Y(n_289)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_250),
.Y(n_362)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_254),
.Y(n_291)
);

AOI21x1_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_278),
.B(n_303),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_274),
.Y(n_257)
);

NOR2xp67_ASAP7_75t_SL g303 ( 
.A(n_258),
.B(n_274),
.Y(n_303)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_259),
.Y(n_301)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_271),
.Y(n_268)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_275),
.B(n_336),
.Y(n_419)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_298),
.B(n_302),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_293),
.B(n_297),
.Y(n_279)
);

NOR2x1_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_289),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_287),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_289),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_289),
.A2(n_299),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_289),
.B(n_312),
.C(n_316),
.Y(n_333)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_292),
.A2(n_359),
.B(n_406),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp33_ASAP7_75t_SL g302 ( 
.A(n_299),
.B(n_300),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_320),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_320),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_310),
.B1(n_311),
.B2(n_319),
.Y(n_306)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_307),
.Y(n_319)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_308),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_312),
.A2(n_313),
.B1(n_314),
.B2(n_318),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_312),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_312),
.A2(n_378),
.B(n_386),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_312),
.B(n_378),
.Y(n_386)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_323),
.B(n_324),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_332),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_325),
.B(n_333),
.C(n_334),
.Y(n_424)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_342),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_SL g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_422),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_412),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_355),
.B(n_397),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_R g444 ( 
.A(n_355),
.B(n_397),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_376),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_356),
.B(n_377),
.C(n_457),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_357),
.B(n_400),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_358),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_375),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_387),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_386),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_386),
.A2(n_450),
.B1(n_452),
.B2(n_460),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_387),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_394),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_389),
.A2(n_390),
.B1(n_392),
.B2(n_393),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_389),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_389),
.A2(n_392),
.B1(n_395),
.B2(n_402),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_389),
.A2(n_393),
.B(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_390),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_392),
.B(n_395),
.Y(n_394)
);

INVxp33_ASAP7_75t_L g454 ( 
.A(n_394),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_395),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_401),
.C(n_403),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_399),
.B(n_401),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_403),
.B(n_421),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_409),
.C(n_410),
.Y(n_403)
);

XNOR2x1_ASAP7_75t_L g414 ( 
.A(n_404),
.B(n_415),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_405),
.Y(n_431)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_412),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_420),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_413),
.B(n_420),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_416),
.C(n_418),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_414),
.B(n_416),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_418),
.B(n_436),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_419),
.B(n_427),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_434),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_425),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_424),
.B(n_425),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_428),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_426),
.B(n_430),
.C(n_432),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_429),
.A2(n_430),
.B1(n_432),
.B2(n_433),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_433),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_434),
.B(n_441),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_437),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_435),
.B(n_437),
.Y(n_439)
);

A2O1A1Ixp33_ASAP7_75t_L g438 ( 
.A1(n_439),
.A2(n_440),
.B(n_442),
.C(n_443),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_455),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_446),
.A2(n_462),
.B(n_463),
.Y(n_461)
);

NOR2xp67_ASAP7_75t_SL g446 ( 
.A(n_447),
.B(n_449),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_447),
.B(n_449),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_452),
.C(n_453),
.Y(n_449)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_450),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_453),
.B(n_459),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_458),
.Y(n_455)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_456),
.B(n_458),
.Y(n_462)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);


endmodule