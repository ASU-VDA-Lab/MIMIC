module real_jpeg_15456_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_516),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_0),
.B(n_517),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_1),
.A2(n_65),
.B1(n_68),
.B2(n_73),
.Y(n_64)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_1),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_1),
.A2(n_73),
.B1(n_160),
.B2(n_165),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_1),
.A2(n_73),
.B1(n_266),
.B2(n_269),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_SL g417 ( 
.A1(n_1),
.A2(n_73),
.B1(n_418),
.B2(n_419),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_2),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_2),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_2),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_2),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_3),
.Y(n_77)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_3),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_3),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_3),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_4),
.A2(n_183),
.B1(n_185),
.B2(n_186),
.Y(n_182)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_4),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_4),
.A2(n_185),
.B1(n_231),
.B2(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_4),
.A2(n_185),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_4),
.A2(n_185),
.B1(n_330),
.B2(n_333),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_5),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_6),
.Y(n_200)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_6),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_7),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_7),
.A2(n_22),
.B1(n_99),
.B2(n_101),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_7),
.B(n_133),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_7),
.A2(n_22),
.B1(n_202),
.B2(n_206),
.Y(n_201)
);

OAI32xp33_ASAP7_75t_L g303 ( 
.A1(n_7),
.A2(n_304),
.A3(n_307),
.B1(n_310),
.B2(n_314),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_7),
.B(n_123),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_7),
.B(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_7),
.B(n_75),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_8),
.Y(n_90)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_8),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_8),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_8),
.Y(n_104)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_8),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_8),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_8),
.Y(n_232)
);

BUFx5_ASAP7_75t_L g257 ( 
.A(n_8),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_9),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_9),
.A2(n_56),
.B1(n_108),
.B2(n_111),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_9),
.B(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_9),
.A2(n_56),
.B1(n_341),
.B2(n_344),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_10),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_11),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_12),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_12),
.Y(n_196)
);

BUFx4f_ASAP7_75t_L g205 ( 
.A(n_12),
.Y(n_205)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_12),
.Y(n_209)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_145),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_144),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_60),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_19),
.B(n_60),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_40),
.Y(n_19)
);

NAND2xp33_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_31),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_21),
.B(n_42),
.Y(n_155)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_21),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B(n_27),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_22),
.B(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_R g221 ( 
.A(n_22),
.B(n_32),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_22),
.B(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_22),
.B(n_311),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_26),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_27),
.A2(n_274),
.B1(n_277),
.B2(n_286),
.Y(n_273)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_31),
.B(n_54),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_31),
.B(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_43),
.Y(n_42)
);

OAI21xp33_ASAP7_75t_SL g63 ( 
.A1(n_32),
.A2(n_40),
.B(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_32),
.A2(n_137),
.B1(n_458),
.B2(n_459),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_32),
.A2(n_137),
.B(n_459),
.Y(n_480)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_32)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_33),
.Y(n_276)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_34),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_34),
.Y(n_122)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_34),
.Y(n_164)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_38),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_41),
.B(n_289),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_54),
.Y(n_41)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_42),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_42),
.B(n_290),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_45),
.B1(n_49),
.B2(n_53),
.Y(n_43)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_56),
.B(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g291 ( 
.A(n_59),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_136),
.C(n_139),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_61),
.B(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_74),
.C(n_105),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_62),
.A2(n_63),
.B1(n_150),
.B2(n_153),
.Y(n_149)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21x1_ASAP7_75t_R g136 ( 
.A1(n_64),
.A2(n_137),
.B(n_138),
.Y(n_136)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_67),
.Y(n_293)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_74),
.A2(n_105),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_74),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_R g157 ( 
.A(n_74),
.B(n_158),
.C(n_170),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_74),
.A2(n_152),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_74),
.A2(n_152),
.B1(n_158),
.B2(n_500),
.Y(n_499)
);

OA21x2_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_86),
.B(n_98),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_75),
.B(n_98),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_75),
.B(n_255),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_75),
.B(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_75),
.B(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_76),
.B(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_80),
.B2(n_84),
.Y(n_76)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_79),
.Y(n_269)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_79),
.Y(n_332)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_88),
.B1(n_91),
.B2(n_94),
.Y(n_87)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_86),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_86),
.B(n_98),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_86),
.B(n_340),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_86),
.Y(n_452)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_90),
.Y(n_343)
);

INVx6_ASAP7_75t_L g347 ( 
.A(n_90),
.Y(n_347)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_97),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g242 ( 
.A(n_104),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_105),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_130),
.Y(n_105)
);

AND2x4_ASAP7_75t_SL g296 ( 
.A(n_106),
.B(n_297),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_106),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_114),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_107),
.B(n_123),
.Y(n_169)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

INVx6_ASAP7_75t_L g286 ( 
.A(n_111),
.Y(n_286)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_112),
.A2(n_116),
.B1(n_118),
.B2(n_121),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_114),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_114),
.B(n_182),
.Y(n_181)
);

NOR2x1_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_123),
.Y(n_114)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_119),
.Y(n_236)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_119),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_121),
.Y(n_227)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_123),
.B(n_182),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_123),
.A2(n_473),
.B(n_474),
.Y(n_472)
);

AO22x2_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_126),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AND2x4_ASAP7_75t_SL g406 ( 
.A(n_130),
.B(n_181),
.Y(n_406)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

OAI32xp33_ASAP7_75t_L g223 ( 
.A1(n_134),
.A2(n_224),
.A3(n_228),
.B1(n_233),
.B2(n_237),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_136),
.A2(n_139),
.B1(n_140),
.B2(n_173),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_136),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_138),
.B(n_409),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_139),
.A2(n_140),
.B1(n_429),
.B2(n_430),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_139),
.B(n_424),
.C(n_430),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_140),
.Y(n_139)
);

AOI21x1_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_142),
.B(n_143),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_141),
.A2(n_159),
.B(n_169),
.Y(n_158)
);

NOR2x1_ASAP7_75t_L g388 ( 
.A(n_141),
.B(n_143),
.Y(n_388)
);

OAI21x1_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_174),
.B(n_514),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_171),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_148),
.B(n_171),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_154),
.C(n_156),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_149),
.A2(n_154),
.B1(n_170),
.B2(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_149),
.Y(n_509)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_150),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_152),
.B(n_288),
.C(n_296),
.Y(n_436)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_154),
.B(n_499),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_155),
.B(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_157),
.B(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_158),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_159),
.Y(n_473)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_169),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_493),
.B(n_511),
.Y(n_174)
);

AO221x1_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_400),
.B1(n_486),
.B2(n_491),
.C(n_492),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_298),
.B(n_399),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_258),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_178),
.B(n_258),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_222),
.C(n_250),
.Y(n_178)
);

XOR2x1_ASAP7_75t_L g394 ( 
.A(n_179),
.B(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_188),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_180),
.B(n_189),
.C(n_221),
.Y(n_261)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_220),
.B2(n_221),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_210),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_191),
.B(n_362),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_201),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_192),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_192),
.B(n_214),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_192),
.B(n_329),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_192),
.A2(n_265),
.B(n_427),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_197),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_195),
.Y(n_268)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_196),
.Y(n_309)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_197),
.Y(n_327)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_200),
.Y(n_365)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_201),
.Y(n_249)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_204),
.Y(n_313)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_205),
.Y(n_215)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_207),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_208),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_209),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_210),
.B(n_328),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_210),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_214),
.B(n_216),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_218),
.Y(n_270)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_222),
.A2(n_250),
.B1(n_251),
.B2(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_222),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_243),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_223),
.A2(n_243),
.B1(n_390),
.B2(n_391),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_223),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_231),
.Y(n_306)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_241),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_243),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_243),
.A2(n_390),
.B1(n_449),
.B2(n_450),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_243),
.A2(n_390),
.B1(n_480),
.B2(n_481),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_243),
.B(n_450),
.Y(n_482)
);

OA21x2_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_248),
.B(n_249),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_246),
.Y(n_360)
);

INVx4_ASAP7_75t_SL g414 ( 
.A(n_246),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

AO21x1_ASAP7_75t_L g325 ( 
.A1(n_249),
.A2(n_326),
.B(n_328),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_249),
.A2(n_272),
.B(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_253),
.B(n_384),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_254),
.B(n_339),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_287),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_260),
.B(n_263),
.C(n_287),
.Y(n_439)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_273),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_264),
.B(n_273),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_270),
.B(n_271),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_271),
.B(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_282),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_279),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_294),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_290),
.Y(n_458)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_297),
.B(n_387),
.Y(n_386)
);

AOI21x1_ASAP7_75t_SL g298 ( 
.A1(n_299),
.A2(n_393),
.B(n_398),
.Y(n_298)
);

OAI21x1_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_376),
.B(n_392),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_351),
.B(n_375),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_324),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_302),
.B(n_324),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_321),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_303),
.B(n_321),
.Y(n_373)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_318),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx5_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_322),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_323),
.B(n_339),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_337),
.Y(n_324)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_325),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_329),
.B(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_338),
.A2(n_348),
.B1(n_349),
.B2(n_350),
.Y(n_337)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_338),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_339),
.A2(n_451),
.B(n_452),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_342),
.Y(n_418)
);

INVx5_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_348),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_348),
.B(n_349),
.C(n_378),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_352),
.A2(n_370),
.B(n_374),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_353),
.A2(n_366),
.B(n_369),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_361),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_358),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_362),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_367),
.B(n_368),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_367),
.B(n_368),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_373),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_371),
.B(n_373),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_379),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_377),
.B(n_379),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_389),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_381),
.A2(n_382),
.B1(n_385),
.B2(n_386),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_381),
.B(n_386),
.C(n_389),
.Y(n_397)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_384),
.Y(n_422)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

NOR2xp67_ASAP7_75t_SL g455 ( 
.A(n_388),
.B(n_456),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_390),
.A2(n_483),
.B(n_503),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_394),
.B(n_397),
.Y(n_393)
);

NOR2xp67_ASAP7_75t_L g398 ( 
.A(n_394),
.B(n_397),
.Y(n_398)
);

NOR3xp33_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_442),
.C(n_463),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_402),
.B(n_438),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_402),
.B(n_489),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_431),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_403),
.B(n_431),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_410),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_404),
.B(n_411),
.C(n_444),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_406),
.C(n_407),
.Y(n_404)
);

XOR2x1_ASAP7_75t_SL g433 ( 
.A(n_405),
.B(n_434),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_406),
.A2(n_407),
.B1(n_408),
.B2(n_435),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_406),
.Y(n_435)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_423),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_415),
.Y(n_411)
);

AOI21x1_ASAP7_75t_SL g460 ( 
.A1(n_412),
.A2(n_416),
.B(n_422),
.Y(n_460)
);

INVx4_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_422),
.Y(n_415)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_417),
.Y(n_451)
);

INVx4_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_423),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_428),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_426),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_425),
.B(n_426),
.Y(n_437)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_429),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_436),
.C(n_437),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_433),
.B(n_441),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_436),
.B(n_437),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_440),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_439),
.B(n_440),
.Y(n_489)
);

A2O1A1Ixp33_ASAP7_75t_L g486 ( 
.A1(n_442),
.A2(n_487),
.B(n_488),
.C(n_490),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_445),
.Y(n_442)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_443),
.B(n_445),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_447),
.Y(n_445)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_446),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_448),
.A2(n_453),
.B1(n_461),
.B2(n_462),
.Y(n_447)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_448),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_448),
.B(n_461),
.C(n_465),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_453),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_460),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_457),
.Y(n_454)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_455),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_457),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_460),
.B(n_468),
.C(n_469),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_463),
.Y(n_491)
);

NOR2x1_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_466),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_464),
.B(n_466),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_470),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_467),
.B(n_471),
.C(n_505),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_471),
.A2(n_477),
.B1(n_484),
.B2(n_485),
.Y(n_470)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_471),
.Y(n_484)
);

OA21x2_ASAP7_75t_L g471 ( 
.A1(n_472),
.A2(n_475),
.B(n_476),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_472),
.B(n_475),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_476),
.A2(n_497),
.B1(n_498),
.B2(n_501),
.Y(n_496)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_476),
.Y(n_501)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_477),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_478),
.A2(n_479),
.B1(n_482),
.B2(n_483),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_480),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_480),
.Y(n_503)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_482),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_485),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_506),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_495),
.B(n_504),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_495),
.B(n_504),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_502),
.Y(n_495)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_498),
.B(n_501),
.C(n_502),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_506),
.A2(n_512),
.B(n_513),
.Y(n_511)
);

NOR2xp67_ASAP7_75t_SL g506 ( 
.A(n_507),
.B(n_510),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_507),
.B(n_510),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);


endmodule