module fake_jpeg_13308_n_173 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_173);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_13),
.B(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_21),
.B(n_8),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_38),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_14),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_18),
.Y(n_50)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

NAND3xp33_ASAP7_75t_L g97 ( 
.A(n_50),
.B(n_73),
.C(n_74),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_15),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_19),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_18),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_27),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_27),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_45),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_25),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_25),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_35),
.B(n_17),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_91),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_15),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_76),
.Y(n_100)
);

OAI22x1_ASAP7_75t_SL g79 ( 
.A1(n_69),
.A2(n_43),
.B1(n_24),
.B2(n_46),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_95),
.B1(n_55),
.B2(n_54),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_90),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_49),
.B1(n_44),
.B2(n_39),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_82),
.A2(n_83),
.B1(n_59),
.B2(n_54),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_58),
.A2(n_61),
.B1(n_64),
.B2(n_70),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_36),
.B(n_28),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_85),
.A2(n_86),
.B(n_87),
.Y(n_114)
);

AO22x1_ASAP7_75t_L g86 ( 
.A1(n_61),
.A2(n_34),
.B1(n_17),
.B2(n_22),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_55),
.A2(n_28),
.B(n_19),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_28),
.C(n_72),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_24),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_67),
.Y(n_92)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_22),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_96),
.Y(n_107)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_59),
.A2(n_29),
.B1(n_26),
.B2(n_31),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_106),
.C(n_91),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_82),
.B1(n_83),
.B2(n_93),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_78),
.B(n_12),
.Y(n_103)
);

NOR4xp25_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_115),
.C(n_10),
.D(n_86),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_70),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_109),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_105),
.A2(n_108),
.B1(n_79),
.B2(n_84),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_63),
.B(n_72),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_81),
.A2(n_29),
.B1(n_63),
.B2(n_62),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_0),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_0),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_104),
.Y(n_127)
);

NAND3xp33_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_11),
.C(n_12),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_85),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_126),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_118),
.A2(n_106),
.B1(n_99),
.B2(n_116),
.Y(n_133)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_122),
.B(n_125),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_123),
.A2(n_110),
.B(n_114),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_124),
.A2(n_130),
.B1(n_101),
.B2(n_102),
.Y(n_137)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_91),
.C(n_84),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_128),
.Y(n_134)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_107),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_129),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_94),
.B1(n_86),
.B2(n_75),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_131),
.Y(n_140)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_119),
.A2(n_102),
.B1(n_113),
.B2(n_114),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_117),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_138),
.C(n_92),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_123),
.B1(n_124),
.B2(n_130),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_99),
.Y(n_138)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_141),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_146),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_109),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_147),
.B(n_149),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_152),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_134),
.B(n_120),
.Y(n_149)
);

NOR3xp33_ASAP7_75t_SL g150 ( 
.A(n_140),
.B(n_120),
.C(n_126),
.Y(n_150)
);

NOR2xp67_ASAP7_75t_R g158 ( 
.A(n_150),
.B(n_132),
.Y(n_158)
);

OAI321xp33_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_113),
.A3(n_29),
.B1(n_3),
.B2(n_4),
.C(n_2),
.Y(n_151)
);

AOI311xp33_ASAP7_75t_L g156 ( 
.A1(n_151),
.A2(n_137),
.A3(n_143),
.B(n_3),
.C(n_4),
.Y(n_156)
);

AOI321xp33_ASAP7_75t_L g154 ( 
.A1(n_150),
.A2(n_132),
.A3(n_138),
.B1(n_143),
.B2(n_141),
.C(n_133),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_154),
.B(n_1),
.Y(n_162)
);

NOR3xp33_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_158),
.C(n_159),
.Y(n_164)
);

OAI21x1_ASAP7_75t_L g159 ( 
.A1(n_152),
.A2(n_142),
.B(n_31),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_145),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_162),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_155),
.A2(n_145),
.B(n_148),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_161),
.A2(n_163),
.B(n_3),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_1),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_164),
.A2(n_155),
.B1(n_157),
.B2(n_2),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_166),
.A2(n_168),
.B(n_31),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_62),
.Y(n_167)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_167),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_169),
.B(n_165),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_165),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_170),
.Y(n_173)
);


endmodule