module fake_jpeg_21809_n_111 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_111);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVxp67_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx4_ASAP7_75t_SL g27 ( 
.A(n_18),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_28),
.Y(n_38)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_31),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g32 ( 
.A(n_17),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_0),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_12),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_29),
.A2(n_13),
.B1(n_17),
.B2(n_21),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_43),
.B1(n_45),
.B2(n_37),
.Y(n_57)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_27),
.A2(n_28),
.B1(n_15),
.B2(n_23),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_47),
.Y(n_62)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_49),
.B(n_51),
.Y(n_65)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

NAND3xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_15),
.C(n_4),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_52),
.B(n_53),
.Y(n_64)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

AND2x6_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_2),
.Y(n_54)
);

AND2x6_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_10),
.Y(n_63)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_57),
.A2(n_58),
.B1(n_41),
.B2(n_24),
.Y(n_72)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_37),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_16),
.Y(n_67)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_70),
.B1(n_72),
.B2(n_16),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_67),
.B(n_56),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_32),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_49),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_37),
.B1(n_41),
.B2(n_12),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_77),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_69),
.A2(n_54),
.B(n_47),
.Y(n_75)
);

A2O1A1O1Ixp25_ASAP7_75t_L g85 ( 
.A1(n_75),
.A2(n_78),
.B(n_55),
.C(n_50),
.D(n_66),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_14),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_26),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_48),
.C(n_59),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_81),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_65),
.B(n_25),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_68),
.Y(n_90)
);

AOI22x1_ASAP7_75t_L g84 ( 
.A1(n_80),
.A2(n_72),
.B1(n_63),
.B2(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_89),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_78),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_77),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_87),
.B(n_90),
.Y(n_92)
);

AOI22x1_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_66),
.B1(n_71),
.B2(n_68),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_79),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_93),
.B(n_95),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_86),
.C(n_92),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_88),
.B(n_75),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_88),
.B(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_98),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_6),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_94),
.B(n_14),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_101),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_99),
.B(n_19),
.Y(n_101)
);

AO22x1_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_2),
.B1(n_20),
.B2(n_8),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_103),
.B(n_7),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_102),
.A2(n_7),
.B1(n_11),
.B2(n_2),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_104),
.A2(n_11),
.B(n_106),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_101),
.Y(n_107)
);

INVxp33_ASAP7_75t_L g109 ( 
.A(n_107),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_109),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_108),
.Y(n_111)
);


endmodule