module fake_jpeg_19206_n_213 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_213);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_213;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_45;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_4),
.B(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_33),
.Y(n_62)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_17),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_20),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_29),
.B(n_24),
.Y(n_44)
);

AOI21xp33_ASAP7_75t_L g69 ( 
.A1(n_44),
.A2(n_41),
.B(n_27),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_29),
.B1(n_30),
.B2(n_23),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_46),
.A2(n_54),
.B1(n_63),
.B2(n_38),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_31),
.B(n_18),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_47),
.B(n_16),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_29),
.B1(n_30),
.B2(n_18),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_58),
.B1(n_27),
.B2(n_19),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_49),
.A2(n_59),
.B(n_36),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_34),
.A2(n_15),
.B1(n_25),
.B2(n_24),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_32),
.A2(n_15),
.B1(n_25),
.B2(n_23),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_32),
.B(n_20),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_43),
.B1(n_39),
.B2(n_33),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_73),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_69),
.A2(n_91),
.B(n_21),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_76),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

AO22x1_ASAP7_75t_SL g72 ( 
.A1(n_62),
.A2(n_42),
.B1(n_37),
.B2(n_43),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_72),
.A2(n_95),
.B1(n_91),
.B2(n_73),
.Y(n_121)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_51),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_81),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_36),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_75),
.B(n_77),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_33),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_78),
.B(n_86),
.Y(n_111)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_82),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_26),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_26),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_26),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_88),
.Y(n_108)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_49),
.B(n_16),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_55),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_49),
.B(n_16),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_90),
.Y(n_112)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_62),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_37),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_20),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_93),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_20),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_55),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_98),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_59),
.A2(n_38),
.B1(n_22),
.B2(n_2),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_60),
.A2(n_21),
.B(n_28),
.C(n_4),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_95),
.Y(n_125)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_52),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_99),
.Y(n_106)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_109),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_64),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_124),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_121),
.A2(n_113),
.B1(n_125),
.B2(n_105),
.Y(n_128)
);

NAND3xp33_ASAP7_75t_L g122 ( 
.A(n_70),
.B(n_0),
.C(n_1),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_122),
.B(n_0),
.Y(n_141)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_76),
.Y(n_127)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_100),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_128),
.A2(n_131),
.B1(n_142),
.B2(n_145),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_67),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_130),
.B(n_139),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_113),
.A2(n_79),
.B1(n_77),
.B2(n_75),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_102),
.A2(n_90),
.B1(n_99),
.B2(n_72),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_132),
.A2(n_109),
.B(n_107),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_85),
.C(n_84),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_137),
.C(n_111),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_100),
.A2(n_98),
.B1(n_68),
.B2(n_72),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_135),
.A2(n_146),
.B1(n_132),
.B2(n_101),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_97),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_66),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_126),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_141),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_121),
.A2(n_45),
.B1(n_22),
.B2(n_28),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_144),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_100),
.A2(n_45),
.B1(n_28),
.B2(n_6),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_146),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_136),
.A2(n_124),
.B1(n_110),
.B2(n_102),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_148),
.A2(n_149),
.B1(n_157),
.B2(n_162),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_138),
.A2(n_110),
.B1(n_118),
.B2(n_104),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_153),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_11),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_155),
.A2(n_103),
.B1(n_138),
.B2(n_6),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_128),
.A2(n_142),
.B1(n_131),
.B2(n_137),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_109),
.B(n_114),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_159),
.A2(n_161),
.B(n_106),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_134),
.B(n_111),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_160),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_135),
.A2(n_129),
.B(n_145),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_132),
.A2(n_114),
.B1(n_143),
.B2(n_112),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_147),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_165),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_147),
.Y(n_165)
);

AOI322xp5_ASAP7_75t_L g166 ( 
.A1(n_160),
.A2(n_133),
.A3(n_132),
.B1(n_119),
.B2(n_116),
.C1(n_103),
.C2(n_106),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_170),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_119),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_169),
.C(n_175),
.Y(n_185)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_168),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_116),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_161),
.B1(n_151),
.B2(n_152),
.Y(n_183)
);

AOI322xp5_ASAP7_75t_L g174 ( 
.A1(n_150),
.A2(n_0),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_156),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_153),
.C(n_162),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_152),
.C(n_7),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_179),
.B(n_176),
.Y(n_190)
);

XNOR2x1_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_155),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_180),
.A2(n_183),
.B1(n_171),
.B2(n_169),
.Y(n_193)
);

INVxp33_ASAP7_75t_L g182 ( 
.A(n_164),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_173),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_168),
.B(n_151),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_186),
.Y(n_188)
);

BUFx12_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_187),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_195),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_180),
.A2(n_172),
.B1(n_171),
.B2(n_175),
.Y(n_191)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_191),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_192),
.A2(n_194),
.B(n_182),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_193),
.A2(n_177),
.B1(n_178),
.B2(n_185),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_181),
.A2(n_163),
.B(n_167),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_5),
.C(n_8),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_197),
.B(n_199),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_187),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_201),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_187),
.Y(n_201)
);

AOI322xp5_ASAP7_75t_L g202 ( 
.A1(n_198),
.A2(n_194),
.A3(n_192),
.B1(n_189),
.B2(n_195),
.C1(n_186),
.C2(n_9),
.Y(n_202)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g208 ( 
.A1(n_202),
.A2(n_196),
.B(n_11),
.C(n_9),
.D(n_197),
.Y(n_208)
);

NOR2x1_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_189),
.Y(n_203)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_203),
.Y(n_207)
);

INVxp33_ASAP7_75t_SL g206 ( 
.A(n_205),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_206),
.B(n_208),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_207),
.B(n_204),
.C(n_198),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_210),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_211),
.B(n_209),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_202),
.Y(n_213)
);


endmodule