module fake_jpeg_12388_n_390 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_390);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_390;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_25),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_52),
.Y(n_91)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_25),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_31),
.B(n_9),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_58),
.B(n_61),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVxp67_ASAP7_75t_SL g84 ( 
.A(n_59),
.Y(n_84)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_31),
.B(n_9),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_25),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_62),
.B(n_67),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_28),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_25),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_68),
.B(n_43),
.Y(n_115)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_71),
.Y(n_99)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_34),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_79),
.B(n_24),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_42),
.B1(n_41),
.B2(n_39),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_86),
.A2(n_78),
.B1(n_45),
.B2(n_37),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_53),
.A2(n_35),
.B1(n_26),
.B2(n_23),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_88),
.A2(n_97),
.B1(n_100),
.B2(n_103),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_57),
.A2(n_35),
.B1(n_39),
.B2(n_42),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_92),
.A2(n_102),
.B1(n_111),
.B2(n_59),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_53),
.A2(n_35),
.B1(n_26),
.B2(n_23),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_71),
.A2(n_26),
.B1(n_23),
.B2(n_41),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_48),
.A2(n_55),
.B1(n_73),
.B2(n_42),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_72),
.A2(n_22),
.B1(n_39),
.B2(n_41),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_48),
.A2(n_32),
.B1(n_27),
.B2(n_28),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_63),
.Y(n_124)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_60),
.A2(n_45),
.B1(n_44),
.B2(n_24),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_118),
.A2(n_76),
.B(n_32),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_143),
.Y(n_157)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_123),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_125),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_91),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_126),
.B(n_128),
.Y(n_169)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_58),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_79),
.B(n_51),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_133),
.Y(n_159)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_82),
.B(n_56),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_134),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_47),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_136),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_64),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_90),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_144),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_49),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_149),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_116),
.A2(n_73),
.B1(n_55),
.B2(n_50),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_139),
.A2(n_141),
.B1(n_142),
.B2(n_146),
.Y(n_160)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_86),
.A2(n_74),
.B1(n_70),
.B2(n_75),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_107),
.A2(n_62),
.B1(n_52),
.B2(n_68),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_93),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_95),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_107),
.A2(n_77),
.B1(n_76),
.B2(n_44),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_95),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_152),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_66),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_153),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_27),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_99),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_150),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_151),
.A2(n_126),
.B1(n_129),
.B2(n_149),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_37),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_87),
.B(n_33),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_87),
.B(n_33),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_85),
.Y(n_174)
);

INVx6_ASAP7_75t_SL g155 ( 
.A(n_84),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_155),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_156),
.A2(n_141),
.B1(n_130),
.B2(n_132),
.Y(n_193)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_104),
.B(n_29),
.C(n_112),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_161),
.B(n_150),
.Y(n_204)
);

FAx1_ASAP7_75t_SL g162 ( 
.A(n_136),
.B(n_105),
.CI(n_112),
.CON(n_162),
.SN(n_162)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_162),
.B(n_173),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_146),
.A2(n_104),
.B1(n_85),
.B2(n_106),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_164),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_106),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_148),
.C(n_153),
.Y(n_198)
);

FAx1_ASAP7_75t_SL g173 ( 
.A(n_128),
.B(n_125),
.CI(n_138),
.CON(n_173),
.SN(n_173)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_174),
.B(n_148),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_131),
.A2(n_83),
.B1(n_113),
.B2(n_66),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_185),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_121),
.A2(n_89),
.B1(n_80),
.B2(n_96),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_183),
.A2(n_80),
.B1(n_89),
.B2(n_109),
.Y(n_206)
);

FAx1_ASAP7_75t_SL g185 ( 
.A(n_123),
.B(n_83),
.CI(n_29),
.CON(n_185),
.SN(n_185)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_172),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_187),
.B(n_190),
.Y(n_229)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_188),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_184),
.Y(n_189)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_158),
.Y(n_190)
);

BUFx16f_ASAP7_75t_L g191 ( 
.A(n_182),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_194),
.Y(n_226)
);

MAJx2_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_124),
.C(n_134),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_196),
.C(n_169),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_193),
.B(n_201),
.Y(n_225)
);

INVxp33_ASAP7_75t_L g194 ( 
.A(n_186),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_171),
.A2(n_151),
.B1(n_120),
.B2(n_152),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_195),
.A2(n_206),
.B1(n_207),
.B2(n_156),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_154),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_197),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_174),
.Y(n_227)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_176),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_199),
.Y(n_233)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_200),
.A2(n_143),
.B1(n_145),
.B2(n_182),
.Y(n_232)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_157),
.A2(n_139),
.B1(n_142),
.B2(n_147),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_179),
.B1(n_178),
.B2(n_162),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_186),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_203),
.B(n_168),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_204),
.A2(n_213),
.B(n_175),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_159),
.B(n_144),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_205),
.B(n_212),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_171),
.A2(n_160),
.B1(n_183),
.B2(n_170),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_165),
.Y(n_216)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_175),
.A2(n_148),
.B1(n_155),
.B2(n_113),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_214),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_209),
.A2(n_160),
.B1(n_170),
.B2(n_157),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_215),
.A2(n_224),
.B1(n_208),
.B2(n_212),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_218),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_209),
.A2(n_161),
.B(n_157),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_217),
.A2(n_219),
.B(n_193),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_163),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_210),
.A2(n_175),
.B(n_178),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_220),
.B(n_227),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_223),
.A2(n_109),
.B1(n_96),
.B2(n_167),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_173),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_228),
.B(n_230),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_232),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_205),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_238),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_207),
.A2(n_162),
.B1(n_185),
.B2(n_179),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_236),
.A2(n_237),
.B1(n_198),
.B2(n_213),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_195),
.A2(n_185),
.B1(n_173),
.B2(n_181),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_192),
.B(n_181),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_189),
.B(n_137),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_239),
.B(n_229),
.Y(n_259)
);

OA21x2_ASAP7_75t_L g241 ( 
.A1(n_215),
.A2(n_204),
.B(n_202),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_241),
.A2(n_262),
.B1(n_266),
.B2(n_122),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_242),
.A2(n_254),
.B1(n_261),
.B2(n_265),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_243),
.A2(n_246),
.B1(n_235),
.B2(n_220),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_244),
.A2(n_263),
.B(n_219),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_224),
.A2(n_208),
.B1(n_206),
.B2(n_201),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_221),
.Y(n_248)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_249),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_199),
.Y(n_250)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_250),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_225),
.Y(n_252)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_252),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_188),
.Y(n_253)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

OAI21xp33_ASAP7_75t_SL g254 ( 
.A1(n_217),
.A2(n_189),
.B(n_143),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_255),
.Y(n_288)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_233),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_258),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_259),
.B(n_140),
.Y(n_276)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_225),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_260),
.Y(n_285)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_226),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_237),
.A2(n_236),
.B(n_214),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_222),
.B(n_197),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_267),
.Y(n_277)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_222),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_223),
.A2(n_200),
.B1(n_167),
.B2(n_145),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_218),
.B(n_191),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_268),
.A2(n_281),
.B(n_256),
.Y(n_304)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_271),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_260),
.A2(n_238),
.B1(n_216),
.B2(n_227),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_263),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_235),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_278),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_276),
.B(n_253),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_245),
.B(n_127),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_279),
.A2(n_283),
.B1(n_287),
.B2(n_246),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_251),
.A2(n_191),
.B(n_119),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_247),
.B(n_119),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_255),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_241),
.A2(n_266),
.B1(n_262),
.B2(n_242),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_119),
.C(n_108),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_286),
.C(n_290),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_240),
.B(n_108),
.C(n_66),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_241),
.A2(n_11),
.B1(n_19),
.B2(n_17),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_240),
.B(n_43),
.C(n_11),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_292),
.B(n_295),
.Y(n_326)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_288),
.Y(n_293)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_293),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_244),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_280),
.Y(n_296)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_296),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_297),
.B(n_303),
.Y(n_314)
);

INVx4_ASAP7_75t_SL g298 ( 
.A(n_289),
.Y(n_298)
);

INVx13_ASAP7_75t_L g328 ( 
.A(n_298),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_299),
.A2(n_279),
.B1(n_291),
.B2(n_269),
.Y(n_317)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_280),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_300),
.Y(n_330)
);

XOR2x2_ASAP7_75t_L g301 ( 
.A(n_273),
.B(n_243),
.Y(n_301)
);

AOI21xp33_ASAP7_75t_L g327 ( 
.A1(n_301),
.A2(n_8),
.B(n_17),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_271),
.B(n_257),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_302),
.B(n_257),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_241),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_304),
.A2(n_272),
.B1(n_283),
.B2(n_268),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_305),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_250),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_309),
.C(n_284),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_285),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_308),
.B(n_259),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_277),
.B(n_258),
.C(n_252),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_275),
.B(n_261),
.Y(n_310)
);

NOR2x1_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_311),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_270),
.B(n_264),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_313),
.B(n_297),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g338 ( 
.A(n_315),
.B(n_321),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_317),
.A2(n_304),
.B1(n_311),
.B2(n_298),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_294),
.B(n_277),
.C(n_272),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_318),
.B(n_325),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_312),
.A2(n_287),
.B1(n_248),
.B2(n_249),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_320),
.A2(n_323),
.B1(n_7),
.B2(n_15),
.Y(n_342)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_322),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_312),
.A2(n_265),
.B1(n_286),
.B2(n_290),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_294),
.B(n_281),
.C(n_11),
.Y(n_325)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_327),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_332),
.B(n_336),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_318),
.A2(n_292),
.B1(n_307),
.B2(n_310),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_333),
.B(n_328),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_313),
.B(n_303),
.C(n_301),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_324),
.B(n_309),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_337),
.B(n_314),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_319),
.B(n_307),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_339),
.B(n_344),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_326),
.B(n_306),
.C(n_295),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_340),
.B(n_343),
.C(n_345),
.Y(n_346)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_341),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_342),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_326),
.B(n_7),
.C(n_14),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_316),
.B(n_6),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_314),
.B(n_323),
.C(n_325),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_338),
.A2(n_324),
.B(n_329),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_347),
.A2(n_330),
.B(n_343),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_348),
.A2(n_356),
.B(n_345),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_340),
.B(n_317),
.Y(n_351)
);

NOR2xp67_ASAP7_75t_SL g360 ( 
.A(n_351),
.B(n_357),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_332),
.B(n_320),
.C(n_329),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_353),
.B(n_354),
.Y(n_359)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_334),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_338),
.A2(n_333),
.B(n_336),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_346),
.B(n_335),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_358),
.B(n_361),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_355),
.B(n_331),
.Y(n_361)
);

OAI221xp5_ASAP7_75t_L g374 ( 
.A1(n_362),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.C(n_4),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_363),
.A2(n_350),
.B(n_357),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_346),
.B(n_330),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_364),
.B(n_365),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_351),
.B(n_328),
.C(n_7),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_353),
.B(n_5),
.Y(n_366)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_366),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_349),
.B(n_5),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_367),
.B(n_368),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_352),
.A2(n_8),
.B(n_13),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_359),
.A2(n_347),
.B(n_356),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_369),
.B(n_374),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_370),
.Y(n_378)
);

AOI21xp33_ASAP7_75t_L g375 ( 
.A1(n_360),
.A2(n_4),
.B(n_19),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_375),
.B(n_4),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_376),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_379),
.B(n_380),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_373),
.B(n_365),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_371),
.B(n_363),
.Y(n_381)
);

OAI321xp33_ASAP7_75t_L g384 ( 
.A1(n_381),
.A2(n_382),
.A3(n_372),
.B1(n_370),
.B2(n_3),
.C(n_2),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_384),
.A2(n_385),
.B(n_378),
.Y(n_386)
);

AOI321xp33_ASAP7_75t_L g385 ( 
.A1(n_377),
.A2(n_0),
.A3(n_2),
.B1(n_3),
.B2(n_376),
.C(n_361),
.Y(n_385)
);

INVxp33_ASAP7_75t_L g388 ( 
.A(n_386),
.Y(n_388)
);

MAJx2_ASAP7_75t_L g387 ( 
.A(n_383),
.B(n_3),
.C(n_0),
.Y(n_387)
);

OR2x2_ASAP7_75t_L g389 ( 
.A(n_388),
.B(n_387),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_389),
.B(n_0),
.Y(n_390)
);


endmodule