module real_aes_1753_n_350 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_969, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_967, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_968, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_350);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_969;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_967;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_968;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_350;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_503;
wire n_357;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_364;
wire n_555;
wire n_766;
wire n_852;
wire n_919;
wire n_857;
wire n_461;
wire n_908;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_353;
wire n_431;
wire n_963;
wire n_865;
wire n_537;
wire n_884;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_550;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_356;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_746;
wire n_656;
wire n_532;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_725;
wire n_960;
wire n_455;
wire n_504;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_867;
wire n_722;
wire n_398;
wire n_688;
wire n_609;
wire n_425;
wire n_879;
wire n_449;
wire n_417;
wire n_754;
wire n_363;
wire n_607;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_617;
wire n_552;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_702;
wire n_954;
wire n_912;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_713;
wire n_598;
wire n_404;
wire n_728;
wire n_735;
wire n_756;
wire n_569;
wire n_785;
wire n_563;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_727;
wire n_649;
wire n_358;
wire n_385;
wire n_397;
wire n_663;
wire n_749;
wire n_588;
wire n_914;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_487;
wire n_831;
wire n_653;
wire n_365;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_922;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_959;
wire n_715;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_721;
wire n_446;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_575;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_587;
wire n_546;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_603;
wire n_854;
wire n_403;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_0), .A2(n_180), .B1(n_369), .B2(n_385), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_1), .A2(n_295), .B1(n_587), .B2(n_752), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_2), .A2(n_12), .B1(n_582), .B2(n_584), .Y(n_837) );
AOI22xp33_ASAP7_75t_SL g712 ( .A1(n_3), .A2(n_101), .B1(n_713), .B2(n_714), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_4), .A2(n_89), .B1(n_369), .B2(n_385), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_5), .A2(n_206), .B1(n_582), .B2(n_584), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_6), .A2(n_318), .B1(n_649), .B2(n_650), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g928 ( .A(n_7), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_8), .A2(n_78), .B1(n_440), .B2(n_522), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_9), .A2(n_144), .B1(n_477), .B2(n_478), .Y(n_476) );
AOI222xp33_ASAP7_75t_SL g791 ( .A1(n_10), .A2(n_34), .B1(n_122), .B2(n_583), .C1(n_792), .C2(n_793), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_11), .A2(n_298), .B1(n_506), .B2(n_544), .Y(n_738) );
AOI22xp33_ASAP7_75t_SL g715 ( .A1(n_13), .A2(n_106), .B1(n_458), .B2(n_580), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_14), .Y(n_492) );
AOI222xp33_ASAP7_75t_L g710 ( .A1(n_15), .A2(n_142), .B1(n_164), .B2(n_454), .C1(n_525), .C2(n_711), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_16), .A2(n_149), .B1(n_522), .B2(n_713), .Y(n_863) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_17), .A2(n_195), .B1(n_410), .B2(n_411), .Y(n_624) );
AOI222xp33_ASAP7_75t_L g865 ( .A1(n_18), .A2(n_100), .B1(n_259), .B2(n_553), .C1(n_731), .C2(n_866), .Y(n_865) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_19), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_20), .A2(n_66), .B1(n_390), .B2(n_395), .Y(n_389) );
AOI222xp33_ASAP7_75t_L g552 ( .A1(n_21), .A2(n_317), .B1(n_339), .B2(n_456), .C1(n_458), .C2(n_553), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_22), .A2(n_271), .B1(n_639), .B2(n_641), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_23), .B(n_762), .Y(n_761) );
AOI222xp33_ASAP7_75t_L g630 ( .A1(n_24), .A2(n_80), .B1(n_153), .B2(n_477), .C1(n_478), .C2(n_482), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_25), .A2(n_209), .B1(n_503), .B2(n_541), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_26), .A2(n_130), .B1(n_502), .B2(n_503), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_27), .A2(n_208), .B1(n_395), .B2(n_477), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g880 ( .A1(n_28), .A2(n_218), .B1(n_881), .B2(n_882), .Y(n_880) );
INVx1_ASAP7_75t_SL g380 ( .A(n_29), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g924 ( .A(n_29), .B(n_39), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_30), .A2(n_52), .B1(n_411), .B2(n_809), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_31), .B(n_762), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_32), .A2(n_82), .B1(n_458), .B2(n_653), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_33), .A2(n_335), .B1(n_470), .B2(n_543), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_35), .A2(n_269), .B1(n_438), .B2(n_440), .Y(n_567) );
AOI22xp33_ASAP7_75t_SL g498 ( .A1(n_36), .A2(n_74), .B1(n_469), .B2(n_499), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_37), .A2(n_53), .B1(n_447), .B2(n_806), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_38), .A2(n_236), .B1(n_598), .B2(n_842), .Y(n_841) );
AO22x2_ASAP7_75t_L g383 ( .A1(n_39), .A2(n_333), .B1(n_372), .B2(n_384), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_40), .A2(n_227), .B1(n_444), .B2(n_447), .Y(n_722) );
AOI22xp33_ASAP7_75t_SL g614 ( .A1(n_41), .A2(n_257), .B1(n_458), .B2(n_580), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_42), .A2(n_185), .B1(n_449), .B2(n_451), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_43), .A2(n_81), .B1(n_418), .B2(n_627), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_44), .A2(n_217), .B1(n_438), .B2(n_440), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_45), .A2(n_328), .B1(n_608), .B2(n_609), .Y(n_607) );
INVx1_ASAP7_75t_L g381 ( .A(n_46), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_47), .A2(n_205), .B1(n_449), .B2(n_547), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_48), .A2(n_224), .B1(n_421), .B2(n_424), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_49), .B(n_482), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_50), .A2(n_95), .B1(n_390), .B2(n_395), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_51), .A2(n_110), .B1(n_544), .B2(n_904), .Y(n_903) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_54), .A2(n_55), .B1(n_517), .B2(n_518), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_56), .A2(n_334), .B1(n_503), .B2(n_541), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_57), .A2(n_212), .B1(n_467), .B2(n_511), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_58), .B(n_565), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_59), .A2(n_121), .B1(n_598), .B2(n_599), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_60), .A2(n_138), .B1(n_670), .B2(n_671), .Y(n_669) );
AOI22xp33_ASAP7_75t_SL g613 ( .A1(n_61), .A2(n_230), .B1(n_435), .B2(n_584), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_62), .A2(n_102), .B1(n_462), .B2(n_718), .Y(n_717) );
AO22x2_ASAP7_75t_L g371 ( .A1(n_63), .A2(n_160), .B1(n_372), .B2(n_373), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_64), .A2(n_343), .B1(n_444), .B2(n_447), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_65), .A2(n_278), .B1(n_656), .B2(n_758), .Y(n_757) );
AOI22xp33_ASAP7_75t_SL g805 ( .A1(n_67), .A2(n_329), .B1(n_806), .B2(n_807), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_68), .A2(n_210), .B1(n_656), .B2(n_681), .Y(n_680) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_69), .A2(n_564), .B(n_566), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g939 ( .A1(n_70), .A2(n_246), .B1(n_506), .B2(n_544), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_71), .A2(n_148), .B1(n_414), .B2(n_415), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_72), .B(n_454), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_73), .A2(n_109), .B1(n_449), .B2(n_750), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_75), .A2(n_225), .B1(n_417), .B2(n_418), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_76), .A2(n_255), .B1(n_522), .B2(n_523), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_77), .A2(n_238), .B1(n_650), .B2(n_890), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_79), .A2(n_131), .B1(n_440), .B2(n_714), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_83), .A2(n_264), .B1(n_588), .B2(n_692), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_84), .A2(n_321), .B1(n_414), .B2(n_415), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g777 ( .A(n_85), .B(n_778), .Y(n_777) );
AOI22xp5_ASAP7_75t_L g849 ( .A1(n_86), .A2(n_266), .B1(n_564), .B2(n_670), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_87), .A2(n_173), .B1(n_418), .B2(n_627), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_88), .A2(n_305), .B1(n_451), .B2(n_813), .Y(n_812) );
OA22x2_ASAP7_75t_L g870 ( .A1(n_90), .A2(n_871), .B1(n_872), .B2(n_891), .Y(n_870) );
INVx1_ASAP7_75t_L g891 ( .A(n_90), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_91), .A2(n_248), .B1(n_398), .B2(n_399), .Y(n_483) );
AOI22x1_ASAP7_75t_L g494 ( .A1(n_92), .A2(n_495), .B1(n_526), .B2(n_527), .Y(n_494) );
CKINVDCx14_ASAP7_75t_R g527 ( .A(n_92), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_93), .A2(n_150), .B1(n_414), .B2(n_415), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_94), .A2(n_176), .B1(n_456), .B2(n_458), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_96), .A2(n_325), .B1(n_561), .B2(n_562), .Y(n_888) );
AOI22xp5_ASAP7_75t_L g759 ( .A1(n_97), .A2(n_289), .B1(n_670), .B2(n_760), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_98), .A2(n_182), .B1(n_462), .B2(n_842), .Y(n_952) );
AO22x2_ASAP7_75t_L g375 ( .A1(n_99), .A2(n_276), .B1(n_372), .B2(n_376), .Y(n_375) );
OA22x2_ASAP7_75t_L g852 ( .A1(n_103), .A2(n_853), .B1(n_854), .B2(n_867), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_103), .Y(n_853) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_104), .A2(n_242), .B1(n_467), .B2(n_469), .Y(n_466) );
AOI222xp33_ASAP7_75t_L g874 ( .A1(n_105), .A2(n_204), .B1(n_254), .B2(n_875), .C1(n_876), .C2(n_878), .Y(n_874) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_107), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_107), .B(n_571), .Y(n_570) );
OAI21xp5_ASAP7_75t_L g590 ( .A1(n_107), .A2(n_591), .B(n_592), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_108), .A2(n_241), .B1(n_398), .B2(n_731), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_111), .A2(n_275), .B1(n_506), .B2(n_718), .Y(n_814) );
AOI22xp5_ASAP7_75t_L g943 ( .A1(n_112), .A2(n_944), .B1(n_959), .B2(n_960), .Y(n_943) );
CKINVDCx20_ASAP7_75t_R g959 ( .A(n_112), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_113), .A2(n_285), .B1(n_414), .B2(n_415), .Y(n_938) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_114), .A2(n_231), .B1(n_456), .B2(n_458), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_115), .A2(n_340), .B1(n_678), .B2(n_771), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_116), .A2(n_168), .B1(n_369), .B2(n_385), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_117), .A2(n_197), .B1(n_587), .B2(n_588), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_118), .A2(n_265), .B1(n_561), .B2(n_562), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_119), .A2(n_184), .B1(n_369), .B2(n_385), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_120), .A2(n_221), .B1(n_417), .B2(n_418), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_123), .A2(n_253), .B1(n_646), .B2(n_695), .Y(n_840) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_124), .A2(n_296), .B1(n_573), .B2(n_574), .Y(n_572) );
BUFx2_ASAP7_75t_R g697 ( .A(n_125), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_126), .A2(n_223), .B1(n_458), .B2(n_580), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_127), .A2(n_261), .B1(n_601), .B2(n_602), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_128), .A2(n_250), .B1(n_643), .B2(n_644), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_129), .A2(n_309), .B1(n_410), .B2(n_411), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_132), .A2(n_181), .B1(n_601), .B2(n_775), .Y(n_843) );
AOI22xp33_ASAP7_75t_SL g687 ( .A1(n_133), .A2(n_213), .B1(n_650), .B2(n_688), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_134), .A2(n_314), .B1(n_562), .B2(n_695), .Y(n_694) );
AOI22xp5_ASAP7_75t_L g774 ( .A1(n_135), .A2(n_190), .B1(n_588), .B2(n_775), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_136), .A2(n_211), .B1(n_447), .B2(n_541), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_137), .A2(n_331), .B1(n_395), .B2(n_477), .Y(n_864) );
AOI22xp33_ASAP7_75t_SL g883 ( .A1(n_139), .A2(n_165), .B1(n_847), .B2(n_884), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_140), .A2(n_267), .B1(n_525), .B2(n_793), .Y(n_899) );
AOI22xp33_ASAP7_75t_SL g684 ( .A1(n_141), .A2(n_229), .B1(n_641), .B2(n_685), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_143), .A2(n_188), .B1(n_398), .B2(n_399), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_145), .A2(n_170), .B1(n_450), .B2(n_547), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_146), .A2(n_147), .B1(n_438), .B2(n_713), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_151), .A2(n_154), .B1(n_604), .B2(n_606), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_152), .A2(n_287), .B1(n_467), .B2(n_721), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_155), .A2(n_303), .B1(n_522), .B2(n_523), .Y(n_756) );
AOI22xp33_ASAP7_75t_SL g822 ( .A1(n_156), .A2(n_312), .B1(n_390), .B2(n_395), .Y(n_822) );
OA22x2_ASAP7_75t_L g724 ( .A1(n_157), .A2(n_725), .B1(n_726), .B2(n_727), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_157), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_158), .A2(n_308), .B1(n_721), .B2(n_861), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_159), .A2(n_171), .B1(n_506), .B2(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g923 ( .A(n_160), .Y(n_923) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_161), .A2(n_306), .B1(n_424), .B2(n_488), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_162), .A2(n_234), .B1(n_398), .B2(n_399), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_163), .A2(n_301), .B1(n_414), .B2(n_415), .Y(n_413) );
INVx1_ASAP7_75t_L g707 ( .A(n_166), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_167), .A2(n_349), .B1(n_444), .B2(n_574), .Y(n_859) );
OA22x2_ASAP7_75t_L g744 ( .A1(n_169), .A2(n_745), .B1(n_746), .B2(n_763), .Y(n_744) );
INVx1_ASAP7_75t_L g763 ( .A(n_169), .Y(n_763) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_172), .A2(n_260), .B1(n_509), .B2(n_511), .Y(n_508) );
INVx1_ASAP7_75t_L g776 ( .A(n_174), .Y(n_776) );
AOI21xp5_ASAP7_75t_L g784 ( .A1(n_174), .A2(n_175), .B(n_785), .Y(n_784) );
AOI22xp33_ASAP7_75t_SL g794 ( .A1(n_174), .A2(n_788), .B1(n_795), .B2(n_969), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_175), .Y(n_796) );
AOI22xp5_ASAP7_75t_L g789 ( .A1(n_177), .A2(n_252), .B1(n_447), .B2(n_790), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_178), .A2(n_228), .B1(n_949), .B2(n_950), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_179), .A2(n_244), .B1(n_721), .B2(n_861), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_183), .A2(n_191), .B1(n_541), .B2(n_754), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_186), .B(n_403), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_187), .A2(n_262), .B1(n_462), .B2(n_547), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_189), .A2(n_345), .B1(n_398), .B2(n_399), .Y(n_932) );
AOI22xp5_ASAP7_75t_L g780 ( .A1(n_192), .A2(n_288), .B1(n_561), .B2(n_562), .Y(n_780) );
INVx2_ASAP7_75t_L g357 ( .A(n_193), .Y(n_357) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_194), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_196), .A2(n_290), .B1(n_432), .B2(n_525), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_198), .A2(n_258), .B1(n_417), .B2(n_418), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_199), .A2(n_291), .B1(n_646), .B2(n_647), .Y(n_645) );
AOI211xp5_ASAP7_75t_L g350 ( .A1(n_200), .A2(n_351), .B(n_360), .C(n_925), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_201), .A2(n_347), .B1(n_438), .B2(n_440), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g936 ( .A1(n_202), .A2(n_237), .B1(n_410), .B2(n_411), .Y(n_936) );
INVx1_ASAP7_75t_L g668 ( .A(n_203), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_207), .A2(n_337), .B1(n_456), .B2(n_458), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_214), .A2(n_220), .B1(n_506), .B2(n_547), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_215), .A2(n_326), .B1(n_547), .B2(n_813), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_216), .A2(n_256), .B1(n_543), .B2(n_750), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_219), .A2(n_310), .B1(n_477), .B2(n_478), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_222), .A2(n_270), .B1(n_458), .B2(n_580), .Y(n_957) );
XNOR2x1_ASAP7_75t_L g428 ( .A(n_226), .B(n_429), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_232), .A2(n_292), .B1(n_424), .B2(n_488), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g958 ( .A(n_233), .B(n_454), .Y(n_958) );
AOI22xp33_ASAP7_75t_SL g631 ( .A1(n_235), .A2(n_307), .B1(n_369), .B2(n_385), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g832 ( .A1(n_239), .A2(n_833), .B1(n_834), .B2(n_850), .Y(n_832) );
INVx1_ASAP7_75t_L g850 ( .A(n_239), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_240), .A2(n_283), .B1(n_522), .B2(n_523), .Y(n_898) );
AOI22xp5_ASAP7_75t_L g770 ( .A1(n_243), .A2(n_346), .B1(n_771), .B2(n_773), .Y(n_770) );
AOI22xp33_ASAP7_75t_SL g431 ( .A1(n_245), .A2(n_319), .B1(n_432), .B2(n_435), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_247), .B(n_564), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_249), .A2(n_268), .B1(n_458), .B2(n_653), .Y(n_781) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_251), .Y(n_818) );
XNOR2x1_ASAP7_75t_L g635 ( .A(n_263), .B(n_636), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_272), .A2(n_322), .B1(n_410), .B2(n_411), .Y(n_737) );
AOI22xp5_ASAP7_75t_L g886 ( .A1(n_273), .A2(n_332), .B1(n_503), .B2(n_573), .Y(n_886) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_274), .A2(n_302), .B1(n_462), .B2(n_463), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g921 ( .A(n_276), .B(n_922), .Y(n_921) );
OA22x2_ASAP7_75t_L g895 ( .A1(n_277), .A2(n_896), .B1(n_908), .B2(n_909), .Y(n_895) );
INVx1_ASAP7_75t_L g908 ( .A(n_277), .Y(n_908) );
AOI22xp5_ASAP7_75t_L g934 ( .A1(n_279), .A2(n_342), .B1(n_369), .B2(n_385), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_280), .A2(n_344), .B1(n_582), .B2(n_656), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_281), .A2(n_327), .B1(n_449), .B2(n_599), .Y(n_856) );
CKINVDCx20_ASAP7_75t_R g845 ( .A(n_282), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_284), .A2(n_320), .B1(n_674), .B2(n_678), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_286), .A2(n_324), .B1(n_543), .B2(n_544), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_293), .A2(n_313), .B1(n_525), .B2(n_956), .Y(n_955) );
INVx3_ASAP7_75t_L g372 ( .A(n_294), .Y(n_372) );
XNOR2x2_ASAP7_75t_L g365 ( .A(n_297), .B(n_366), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_299), .A2(n_316), .B1(n_410), .B2(n_411), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_300), .B(n_564), .Y(n_615) );
CKINVDCx20_ASAP7_75t_R g633 ( .A(n_304), .Y(n_633) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_311), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_315), .B(n_565), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_323), .A2(n_348), .B1(n_410), .B2(n_411), .Y(n_409) );
XNOR2xp5_ASAP7_75t_L g594 ( .A(n_330), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_336), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g919 ( .A(n_336), .Y(n_919) );
INVx1_ASAP7_75t_L g354 ( .A(n_338), .Y(n_354) );
AND2x2_ASAP7_75t_R g962 ( .A(n_338), .B(n_919), .Y(n_962) );
INVxp67_ASAP7_75t_L g359 ( .A(n_341), .Y(n_359) );
BUFx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NOR2x1_ASAP7_75t_R g352 ( .A(n_353), .B(n_355), .Y(n_352) );
OR2x2_ASAP7_75t_L g965 ( .A(n_353), .B(n_356), .Y(n_965) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g918 ( .A(n_354), .B(n_919), .Y(n_918) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_700), .B1(n_914), .B2(n_915), .C(n_916), .Y(n_360) );
INVx1_ASAP7_75t_L g915 ( .A(n_361), .Y(n_915) );
OAI22xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_363), .B1(n_533), .B2(n_534), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AOI22xp33_ASAP7_75t_SL g363 ( .A1(n_364), .A2(n_425), .B1(n_426), .B2(n_532), .Y(n_363) );
INVx1_ASAP7_75t_SL g532 ( .A(n_364), .Y(n_532) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_408), .Y(n_366) );
NAND4xp25_ASAP7_75t_L g367 ( .A(n_368), .B(n_389), .C(n_397), .D(n_402), .Y(n_367) );
AND2x4_ASAP7_75t_L g369 ( .A(n_370), .B(n_377), .Y(n_369) );
AND2x6_ASAP7_75t_L g411 ( .A(n_370), .B(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g417 ( .A(n_370), .B(n_391), .Y(n_417) );
AND2x2_ASAP7_75t_L g439 ( .A(n_370), .B(n_377), .Y(n_439) );
AND2x2_ASAP7_75t_L g446 ( .A(n_370), .B(n_391), .Y(n_446) );
AND2x4_ASAP7_75t_L g465 ( .A(n_370), .B(n_412), .Y(n_465) );
AND2x2_ASAP7_75t_SL g627 ( .A(n_370), .B(n_391), .Y(n_627) );
AND2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_374), .Y(n_370) );
INVx2_ASAP7_75t_L g394 ( .A(n_371), .Y(n_394) );
AND2x2_ASAP7_75t_L g401 ( .A(n_371), .B(n_375), .Y(n_401) );
INVx1_ASAP7_75t_L g373 ( .A(n_372), .Y(n_373) );
INVx2_ASAP7_75t_L g376 ( .A(n_372), .Y(n_376) );
OAI22x1_ASAP7_75t_L g378 ( .A1(n_372), .A2(n_379), .B1(n_380), .B2(n_381), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_372), .Y(n_379) );
INVx1_ASAP7_75t_L g384 ( .A(n_372), .Y(n_384) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_374), .Y(n_387) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x4_ASAP7_75t_L g393 ( .A(n_375), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g407 ( .A(n_375), .Y(n_407) );
AND2x4_ASAP7_75t_L g398 ( .A(n_377), .B(n_393), .Y(n_398) );
AND2x2_ASAP7_75t_L g414 ( .A(n_377), .B(n_406), .Y(n_414) );
AND2x4_ASAP7_75t_L g450 ( .A(n_377), .B(n_406), .Y(n_450) );
AND2x2_ASAP7_75t_L g457 ( .A(n_377), .B(n_393), .Y(n_457) );
AND2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_382), .Y(n_377) );
AND2x2_ASAP7_75t_L g388 ( .A(n_378), .B(n_383), .Y(n_388) );
INVx2_ASAP7_75t_L g392 ( .A(n_378), .Y(n_392) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_378), .Y(n_400) );
AND2x4_ASAP7_75t_L g412 ( .A(n_382), .B(n_392), .Y(n_412) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g391 ( .A(n_383), .B(n_392), .Y(n_391) );
BUFx2_ASAP7_75t_L g419 ( .A(n_383), .Y(n_419) );
AND2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_388), .Y(n_385) );
AND2x4_ASAP7_75t_L g441 ( .A(n_386), .B(n_388), .Y(n_441) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g395 ( .A(n_388), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g405 ( .A(n_388), .B(n_406), .Y(n_405) );
AND2x4_ASAP7_75t_L g434 ( .A(n_388), .B(n_396), .Y(n_434) );
AND2x2_ASAP7_75t_L g478 ( .A(n_388), .B(n_396), .Y(n_478) );
AND2x4_ASAP7_75t_L g482 ( .A(n_388), .B(n_406), .Y(n_482) );
AND2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_393), .Y(n_390) );
AND2x6_ASAP7_75t_L g410 ( .A(n_391), .B(n_406), .Y(n_410) );
AND2x4_ASAP7_75t_L g436 ( .A(n_391), .B(n_393), .Y(n_436) );
AND2x2_ASAP7_75t_L g468 ( .A(n_391), .B(n_406), .Y(n_468) );
AND2x2_ASAP7_75t_L g477 ( .A(n_391), .B(n_393), .Y(n_477) );
AND2x2_ASAP7_75t_L g424 ( .A(n_393), .B(n_412), .Y(n_424) );
AND2x4_ASAP7_75t_L g470 ( .A(n_393), .B(n_412), .Y(n_470) );
INVxp67_ASAP7_75t_L g396 ( .A(n_394), .Y(n_396) );
AND2x4_ASAP7_75t_L g406 ( .A(n_394), .B(n_407), .Y(n_406) );
HB1xp67_ASAP7_75t_L g866 ( .A(n_398), .Y(n_866) );
AND2x2_ASAP7_75t_SL g399 ( .A(n_400), .B(n_401), .Y(n_399) );
AND2x2_ASAP7_75t_L g459 ( .A(n_400), .B(n_401), .Y(n_459) );
AND2x2_ASAP7_75t_SL g731 ( .A(n_400), .B(n_401), .Y(n_731) );
AND2x4_ASAP7_75t_L g415 ( .A(n_401), .B(n_412), .Y(n_415) );
AND2x4_ASAP7_75t_L g418 ( .A(n_401), .B(n_419), .Y(n_418) );
AND2x4_ASAP7_75t_L g447 ( .A(n_401), .B(n_419), .Y(n_447) );
AND2x4_ASAP7_75t_L g451 ( .A(n_401), .B(n_412), .Y(n_451) );
INVx4_ASAP7_75t_SL g403 ( .A(n_404), .Y(n_403) );
INVx3_ASAP7_75t_L g454 ( .A(n_404), .Y(n_454) );
BUFx2_ASAP7_75t_L g514 ( .A(n_404), .Y(n_514) );
INVx3_ASAP7_75t_SL g565 ( .A(n_404), .Y(n_565) );
INVx4_ASAP7_75t_SL g762 ( .A(n_404), .Y(n_762) );
INVx3_ASAP7_75t_L g792 ( .A(n_404), .Y(n_792) );
INVx6_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AND2x4_ASAP7_75t_L g423 ( .A(n_406), .B(n_412), .Y(n_423) );
AND2x2_ASAP7_75t_L g488 ( .A(n_406), .B(n_412), .Y(n_488) );
NAND4xp25_ASAP7_75t_L g408 ( .A(n_409), .B(n_413), .C(n_416), .D(n_420), .Y(n_408) );
INVx1_ASAP7_75t_L g810 ( .A(n_410), .Y(n_810) );
BUFx6f_ASAP7_75t_L g646 ( .A(n_421), .Y(n_646) );
INVx2_ASAP7_75t_L g689 ( .A(n_421), .Y(n_689) );
INVx4_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_SL g462 ( .A(n_422), .Y(n_462) );
INVx3_ASAP7_75t_L g506 ( .A(n_422), .Y(n_506) );
INVx3_ASAP7_75t_SL g543 ( .A(n_422), .Y(n_543) );
INVx2_ASAP7_75t_SL g608 ( .A(n_422), .Y(n_608) );
INVx2_ASAP7_75t_L g904 ( .A(n_422), .Y(n_904) );
INVx8_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AO22x2_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_471), .B1(n_530), .B2(n_531), .Y(n_426) );
INVx1_ASAP7_75t_L g530 ( .A(n_427), .Y(n_530) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NAND4xp75_ASAP7_75t_L g429 ( .A(n_430), .B(n_442), .C(n_452), .D(n_460), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_437), .Y(n_430) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_SL g584 ( .A(n_433), .Y(n_584) );
INVx2_ASAP7_75t_L g656 ( .A(n_433), .Y(n_656) );
INVx2_ASAP7_75t_SL g711 ( .A(n_433), .Y(n_711) );
INVx2_ASAP7_75t_L g793 ( .A(n_433), .Y(n_793) );
INVx2_ASAP7_75t_L g882 ( .A(n_433), .Y(n_882) );
INVx1_ASAP7_75t_L g956 ( .A(n_433), .Y(n_956) );
INVx6_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx3_ASAP7_75t_L g525 ( .A(n_436), .Y(n_525) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_436), .Y(n_583) );
BUFx2_ASAP7_75t_L g758 ( .A(n_436), .Y(n_758) );
BUFx6f_ASAP7_75t_SL g881 ( .A(n_438), .Y(n_881) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_439), .Y(n_522) );
INVx3_ASAP7_75t_L g677 ( .A(n_439), .Y(n_677) );
BUFx4f_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx3_ASAP7_75t_L g523 ( .A(n_441), .Y(n_523) );
INVx2_ASAP7_75t_L g679 ( .A(n_441), .Y(n_679) );
BUFx6f_ASAP7_75t_SL g713 ( .A(n_441), .Y(n_713) );
AND2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_448), .Y(n_442) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g605 ( .A(n_445), .Y(n_605) );
INVx1_ASAP7_75t_L g806 ( .A(n_445), .Y(n_806) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx3_ASAP7_75t_L g502 ( .A(n_446), .Y(n_502) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_446), .Y(n_541) );
BUFx3_ASAP7_75t_L g503 ( .A(n_447), .Y(n_503) );
INVx5_ASAP7_75t_SL g575 ( .A(n_447), .Y(n_575) );
BUFx2_ASAP7_75t_L g606 ( .A(n_447), .Y(n_606) );
BUFx2_ASAP7_75t_L g807 ( .A(n_447), .Y(n_807) );
BUFx3_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx6_ASAP7_75t_L g500 ( .A(n_450), .Y(n_500) );
BUFx3_ASAP7_75t_L g813 ( .A(n_450), .Y(n_813) );
BUFx3_ASAP7_75t_L g507 ( .A(n_451), .Y(n_507) );
BUFx3_ASAP7_75t_L g547 ( .A(n_451), .Y(n_547) );
INVx2_ASAP7_75t_L g610 ( .A(n_451), .Y(n_610) );
BUFx2_ASAP7_75t_SL g644 ( .A(n_451), .Y(n_644) );
BUFx2_ASAP7_75t_SL g695 ( .A(n_451), .Y(n_695) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_455), .Y(n_452) );
BUFx6f_ASAP7_75t_L g884 ( .A(n_456), .Y(n_884) );
BUFx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx3_ASAP7_75t_L g517 ( .A(n_457), .Y(n_517) );
BUFx5_ASAP7_75t_L g580 ( .A(n_457), .Y(n_580) );
INVx2_ASAP7_75t_L g654 ( .A(n_457), .Y(n_654) );
BUFx12f_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx3_ASAP7_75t_L g519 ( .A(n_459), .Y(n_519) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_466), .Y(n_460) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g511 ( .A(n_464), .Y(n_511) );
INVx2_ASAP7_75t_SL g587 ( .A(n_464), .Y(n_587) );
INVx1_ASAP7_75t_SL g602 ( .A(n_464), .Y(n_602) );
INVx2_ASAP7_75t_L g650 ( .A(n_464), .Y(n_650) );
INVx2_ASAP7_75t_L g721 ( .A(n_464), .Y(n_721) );
INVx2_ASAP7_75t_L g775 ( .A(n_464), .Y(n_775) );
INVx8_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g589 ( .A(n_467), .Y(n_589) );
BUFx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx3_ASAP7_75t_L g510 ( .A(n_468), .Y(n_510) );
BUFx2_ASAP7_75t_L g861 ( .A(n_468), .Y(n_861) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_470), .Y(n_544) );
BUFx3_ASAP7_75t_L g599 ( .A(n_470), .Y(n_599) );
INVx2_ASAP7_75t_L g719 ( .A(n_470), .Y(n_719) );
INVx2_ASAP7_75t_L g531 ( .A(n_471), .Y(n_531) );
OA22x2_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_493), .B1(n_494), .B2(n_528), .Y(n_471) );
XOR2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_492), .Y(n_472) );
XOR2x2_ASAP7_75t_L g529 ( .A(n_473), .B(n_492), .Y(n_529) );
NAND2x1_ASAP7_75t_SL g473 ( .A(n_474), .B(n_484), .Y(n_473) );
NOR2x1_ASAP7_75t_L g474 ( .A(n_475), .B(n_480), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_479), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_483), .Y(n_480) );
BUFx2_ASAP7_75t_L g553 ( .A(n_482), .Y(n_553) );
INVx2_ASAP7_75t_SL g817 ( .A(n_482), .Y(n_817) );
NOR2x1_ASAP7_75t_L g484 ( .A(n_485), .B(n_489), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g526 ( .A(n_495), .Y(n_526) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_512), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_497), .B(n_504), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_501), .Y(n_497) );
INVx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_SL g562 ( .A(n_500), .Y(n_562) );
INVx2_ASAP7_75t_L g598 ( .A(n_500), .Y(n_598) );
INVx2_ASAP7_75t_L g643 ( .A(n_500), .Y(n_643) );
INVx2_ASAP7_75t_L g949 ( .A(n_500), .Y(n_949) );
BUFx2_ASAP7_75t_L g573 ( .A(n_502), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_508), .Y(n_504) );
INVx3_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_SL g601 ( .A(n_510), .Y(n_601) );
INVx2_ASAP7_75t_SL g649 ( .A(n_510), .Y(n_649) );
INVx2_ASAP7_75t_L g752 ( .A(n_510), .Y(n_752) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_513), .B(n_520), .Y(n_512) );
OAI21xp5_ASAP7_75t_SL g513 ( .A1(n_514), .A2(n_515), .B(n_516), .Y(n_513) );
BUFx6f_ASAP7_75t_L g671 ( .A(n_518), .Y(n_671) );
INVx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g760 ( .A(n_519), .Y(n_760) );
INVx2_ASAP7_75t_L g848 ( .A(n_519), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_524), .Y(n_520) );
BUFx6f_ASAP7_75t_SL g773 ( .A(n_523), .Y(n_773) );
INVx1_ASAP7_75t_L g879 ( .A(n_525), .Y(n_879) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_617), .B1(n_618), .B2(n_699), .Y(n_534) );
INVx1_ASAP7_75t_L g699 ( .A(n_535), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_555), .B1(n_556), .B2(n_616), .Y(n_535) );
INVx2_ASAP7_75t_L g616 ( .A(n_536), .Y(n_616) );
BUFx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
XOR2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_554), .Y(n_537) );
NAND4xp75_ASAP7_75t_L g538 ( .A(n_539), .B(n_545), .C(n_549), .D(n_552), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_542), .Y(n_539) );
BUFx6f_ASAP7_75t_L g647 ( .A(n_544), .Y(n_647) );
INVx2_ASAP7_75t_L g693 ( .A(n_544), .Y(n_693) );
AND2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_548), .Y(n_545) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_547), .Y(n_561) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_558), .B1(n_593), .B2(n_594), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_576), .Y(n_558) );
A2O1A1Ixp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_563), .B(n_569), .C(n_570), .Y(n_559) );
NAND3xp33_ASAP7_75t_L g585 ( .A(n_560), .B(n_563), .C(n_586), .Y(n_585) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g667 ( .A(n_565), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
NAND3xp33_ASAP7_75t_L g577 ( .A(n_569), .B(n_572), .C(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g641 ( .A(n_575), .Y(n_641) );
INVx3_ASAP7_75t_L g754 ( .A(n_575), .Y(n_754) );
OAI21xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_585), .B(n_590), .Y(n_576) );
INVx1_ASAP7_75t_L g592 ( .A(n_578), .Y(n_592) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
BUFx4f_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
BUFx2_ASAP7_75t_L g681 ( .A(n_583), .Y(n_681) );
INVx1_ASAP7_75t_L g591 ( .A(n_586), .Y(n_591) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_611), .Y(n_595) );
NAND4xp25_ASAP7_75t_L g596 ( .A(n_597), .B(n_600), .C(n_603), .D(n_607), .Y(n_596) );
BUFx2_ASAP7_75t_L g778 ( .A(n_599), .Y(n_778) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g640 ( .A(n_605), .Y(n_640) );
INVx1_ASAP7_75t_L g686 ( .A(n_605), .Y(n_686) );
HB1xp67_ASAP7_75t_L g790 ( .A(n_605), .Y(n_790) );
BUFx2_ASAP7_75t_L g785 ( .A(n_608), .Y(n_785) );
INVx2_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_SL g950 ( .A(n_610), .Y(n_950) );
NAND4xp25_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .C(n_614), .D(n_615), .Y(n_611) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OA22x2_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_660), .B1(n_661), .B2(n_698), .Y(n_618) );
INVx2_ASAP7_75t_L g698 ( .A(n_619), .Y(n_698) );
AO22x2_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_634), .B1(n_635), .B2(n_659), .Y(n_619) );
BUFx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g659 ( .A(n_621), .Y(n_659) );
INVx1_ASAP7_75t_L g824 ( .A(n_621), .Y(n_824) );
XNOR2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_633), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_629), .Y(n_622) );
NAND4xp25_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .C(n_626), .D(n_628), .Y(n_623) );
NAND3xp33_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .C(n_632), .Y(n_629) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_651), .Y(n_636) );
NAND4xp25_ASAP7_75t_L g637 ( .A(n_638), .B(n_642), .C(n_645), .D(n_648), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND4xp25_ASAP7_75t_L g651 ( .A(n_652), .B(n_655), .C(n_657), .D(n_658), .Y(n_651) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g670 ( .A(n_654), .Y(n_670) );
OAI21xp5_ASAP7_75t_L g799 ( .A1(n_659), .A2(n_800), .B(n_823), .Y(n_799) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AOI22x1_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_664), .B1(n_696), .B2(n_697), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_682), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_666), .B(n_672), .Y(n_665) );
OAI21xp5_ASAP7_75t_SL g666 ( .A1(n_667), .A2(n_668), .B(n_669), .Y(n_666) );
INVx2_ASAP7_75t_L g875 ( .A(n_667), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_673), .B(n_680), .Y(n_672) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx2_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
INVx4_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g714 ( .A(n_677), .Y(n_714) );
INVx1_ASAP7_75t_L g772 ( .A(n_677), .Y(n_772) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
BUFx2_ASAP7_75t_L g877 ( .A(n_679), .Y(n_877) );
NOR2x1_ASAP7_75t_L g682 ( .A(n_683), .B(n_690), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_687), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_694), .Y(n_690) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g914 ( .A(n_700), .Y(n_914) );
XOR2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_828), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_766), .B1(n_826), .B2(n_827), .Y(n_701) );
INVx1_ASAP7_75t_L g827 ( .A(n_702), .Y(n_827) );
INVx4_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
OA22x2_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_705), .B1(n_742), .B2(n_764), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AOI22x1_ASAP7_75t_SL g705 ( .A1(n_706), .A2(n_724), .B1(n_740), .B2(n_741), .Y(n_705) );
INVx1_ASAP7_75t_SL g741 ( .A(n_706), .Y(n_741) );
XNOR2x1_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
OR2x2_ASAP7_75t_L g708 ( .A(n_709), .B(n_716), .Y(n_708) );
NAND3xp33_ASAP7_75t_L g709 ( .A(n_710), .B(n_712), .C(n_715), .Y(n_709) );
NAND4xp25_ASAP7_75t_L g716 ( .A(n_717), .B(n_720), .C(n_722), .D(n_723), .Y(n_716) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g750 ( .A(n_719), .Y(n_750) );
INVx1_ASAP7_75t_L g842 ( .A(n_719), .Y(n_842) );
INVx3_ASAP7_75t_L g740 ( .A(n_724), .Y(n_740) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
NOR2x1_ASAP7_75t_L g727 ( .A(n_728), .B(n_734), .Y(n_727) );
NAND4xp25_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .C(n_732), .D(n_733), .Y(n_728) );
NAND3xp33_ASAP7_75t_L g734 ( .A(n_735), .B(n_738), .C(n_739), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
BUFx2_ASAP7_75t_L g765 ( .A(n_744), .Y(n_765) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NOR2x1_ASAP7_75t_L g746 ( .A(n_747), .B(n_755), .Y(n_746) );
NAND4xp25_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .C(n_751), .D(n_753), .Y(n_747) );
NAND4xp25_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .C(n_759), .D(n_761), .Y(n_755) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx3_ASAP7_75t_L g826 ( .A(n_766), .Y(n_826) );
OA22x2_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_798), .B1(n_799), .B2(n_825), .Y(n_766) );
INVx2_ASAP7_75t_SL g825 ( .A(n_767), .Y(n_825) );
OR2x2_ASAP7_75t_L g767 ( .A(n_768), .B(n_782), .Y(n_767) );
OAI222xp33_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_776), .B1(n_777), .B2(n_779), .C1(n_967), .C2(n_968), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_769), .B(n_787), .Y(n_786) );
AND2x2_ASAP7_75t_L g769 ( .A(n_770), .B(n_774), .Y(n_769) );
BUFx3_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
NAND3xp33_ASAP7_75t_L g783 ( .A(n_777), .B(n_779), .C(n_784), .Y(n_783) );
AND2x2_ASAP7_75t_SL g779 ( .A(n_780), .B(n_781), .Y(n_779) );
OAI21xp5_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_786), .B(n_794), .Y(n_782) );
INVx1_ASAP7_75t_L g797 ( .A(n_785), .Y(n_797) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_789), .B(n_791), .Y(n_788) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .Y(n_795) );
INVx1_ASAP7_75t_SL g798 ( .A(n_799), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_800), .B(n_824), .Y(n_823) );
XNOR2x1_ASAP7_75t_L g800 ( .A(n_801), .B(n_802), .Y(n_800) );
NAND2x1p5_ASAP7_75t_L g802 ( .A(n_803), .B(n_815), .Y(n_802) );
NOR2x1_ASAP7_75t_L g803 ( .A(n_804), .B(n_811), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_805), .B(n_808), .Y(n_804) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_812), .B(n_814), .Y(n_811) );
NOR2x1_ASAP7_75t_L g815 ( .A(n_816), .B(n_820), .Y(n_815) );
OAI21xp5_ASAP7_75t_SL g816 ( .A1(n_817), .A2(n_818), .B(n_819), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_821), .B(n_822), .Y(n_820) );
AOI22xp5_ASAP7_75t_SL g828 ( .A1(n_829), .A2(n_869), .B1(n_912), .B2(n_913), .Y(n_828) );
INVx1_ASAP7_75t_L g912 ( .A(n_829), .Y(n_912) );
INVx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
AO22x1_ASAP7_75t_L g830 ( .A1(n_831), .A2(n_832), .B1(n_851), .B2(n_868), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
NOR3xp33_ASAP7_75t_SL g834 ( .A(n_835), .B(n_838), .C(n_844), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_836), .B(n_837), .Y(n_835) );
NAND4xp25_ASAP7_75t_SL g838 ( .A(n_839), .B(n_840), .C(n_841), .D(n_843), .Y(n_838) );
OAI21xp5_ASAP7_75t_SL g844 ( .A1(n_845), .A2(n_846), .B(n_849), .Y(n_844) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
BUFx2_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
BUFx2_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVxp67_ASAP7_75t_L g868 ( .A(n_852), .Y(n_868) );
AO22x1_ASAP7_75t_L g892 ( .A1(n_852), .A2(n_893), .B1(n_894), .B2(n_895), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_852), .Y(n_893) );
INVx2_ASAP7_75t_L g867 ( .A(n_854), .Y(n_867) );
NAND4xp75_ASAP7_75t_L g854 ( .A(n_855), .B(n_858), .C(n_862), .D(n_865), .Y(n_854) );
AND2x2_ASAP7_75t_L g855 ( .A(n_856), .B(n_857), .Y(n_855) );
AND2x2_ASAP7_75t_L g858 ( .A(n_859), .B(n_860), .Y(n_858) );
BUFx3_ASAP7_75t_L g890 ( .A(n_861), .Y(n_890) );
AND2x2_ASAP7_75t_L g862 ( .A(n_863), .B(n_864), .Y(n_862) );
INVx3_ASAP7_75t_L g913 ( .A(n_869), .Y(n_913) );
AO22x2_ASAP7_75t_L g869 ( .A1(n_870), .A2(n_892), .B1(n_910), .B2(n_911), .Y(n_869) );
INVx1_ASAP7_75t_L g910 ( .A(n_870), .Y(n_910) );
INVx2_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
OR2x2_ASAP7_75t_L g872 ( .A(n_873), .B(n_885), .Y(n_872) );
NAND3xp33_ASAP7_75t_L g873 ( .A(n_874), .B(n_880), .C(n_883), .Y(n_873) );
INVx3_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
NAND4xp25_ASAP7_75t_L g885 ( .A(n_886), .B(n_887), .C(n_888), .D(n_889), .Y(n_885) );
INVx1_ASAP7_75t_L g911 ( .A(n_892), .Y(n_911) );
INVx1_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
INVx1_ASAP7_75t_L g909 ( .A(n_896), .Y(n_909) );
NOR2x1_ASAP7_75t_L g896 ( .A(n_897), .B(n_902), .Y(n_896) );
NAND4xp25_ASAP7_75t_L g897 ( .A(n_898), .B(n_899), .C(n_900), .D(n_901), .Y(n_897) );
NAND4xp25_ASAP7_75t_L g902 ( .A(n_903), .B(n_905), .C(n_906), .D(n_907), .Y(n_902) );
CKINVDCx5p33_ASAP7_75t_R g916 ( .A(n_917), .Y(n_916) );
AND2x2_ASAP7_75t_L g917 ( .A(n_918), .B(n_920), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_918), .B(n_921), .Y(n_942) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_923), .B(n_924), .Y(n_922) );
OAI222xp33_ASAP7_75t_L g925 ( .A1(n_926), .A2(n_928), .B1(n_940), .B2(n_943), .C1(n_961), .C2(n_963), .Y(n_925) );
HB1xp67_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
XNOR2x1_ASAP7_75t_L g927 ( .A(n_928), .B(n_929), .Y(n_927) );
NOR2x1_ASAP7_75t_L g929 ( .A(n_930), .B(n_935), .Y(n_929) );
NAND4xp25_ASAP7_75t_L g930 ( .A(n_931), .B(n_932), .C(n_933), .D(n_934), .Y(n_930) );
NAND4xp25_ASAP7_75t_L g935 ( .A(n_936), .B(n_937), .C(n_938), .D(n_939), .Y(n_935) );
INVx1_ASAP7_75t_SL g940 ( .A(n_941), .Y(n_940) );
CKINVDCx6p67_ASAP7_75t_R g941 ( .A(n_942), .Y(n_941) );
CKINVDCx20_ASAP7_75t_R g960 ( .A(n_944), .Y(n_960) );
HB1xp67_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
NOR2xp67_ASAP7_75t_L g945 ( .A(n_946), .B(n_953), .Y(n_945) );
NAND4xp25_ASAP7_75t_L g946 ( .A(n_947), .B(n_948), .C(n_951), .D(n_952), .Y(n_946) );
NAND4xp25_ASAP7_75t_L g953 ( .A(n_954), .B(n_955), .C(n_957), .D(n_958), .Y(n_953) );
INVx2_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
CKINVDCx20_ASAP7_75t_R g963 ( .A(n_964), .Y(n_963) );
CKINVDCx20_ASAP7_75t_R g964 ( .A(n_965), .Y(n_964) );
endmodule