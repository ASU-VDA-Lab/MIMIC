module fake_ariane_2181_n_1975 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_172, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1975);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1975;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_181;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_177;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_118),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_77),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_45),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_48),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_68),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_149),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_139),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_85),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_78),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_49),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_4),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_2),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_0),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_62),
.Y(n_186)
);

BUFx10_ASAP7_75t_L g187 ( 
.A(n_25),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_163),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_26),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_129),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_146),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_43),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_26),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_87),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_58),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_1),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_25),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_8),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_10),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_71),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_66),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_37),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_135),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_137),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_96),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_58),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_140),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_142),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_21),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_131),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_54),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_84),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_172),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_136),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_106),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_101),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_3),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_168),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_23),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_124),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_62),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_22),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_104),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_6),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_133),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_117),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_166),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_45),
.Y(n_228)
);

BUFx10_ASAP7_75t_L g229 ( 
.A(n_55),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_68),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_114),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_64),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_141),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_30),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_88),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_2),
.Y(n_236)
);

BUFx5_ASAP7_75t_L g237 ( 
.A(n_162),
.Y(n_237)
);

BUFx5_ASAP7_75t_L g238 ( 
.A(n_120),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_156),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_43),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_126),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_11),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_159),
.Y(n_243)
);

BUFx5_ASAP7_75t_L g244 ( 
.A(n_12),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_155),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_92),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_8),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_60),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_145),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_54),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_3),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_1),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_134),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_169),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_41),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_79),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_12),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_105),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_112),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_4),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_63),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_11),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_154),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_150),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_69),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_81),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_63),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_23),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_158),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_46),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_76),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_143),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_61),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_160),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_46),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_49),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_70),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_95),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_47),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_24),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_116),
.Y(n_281)
);

INVxp67_ASAP7_75t_SL g282 ( 
.A(n_76),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_55),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_125),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_36),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_80),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_153),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_35),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_20),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_22),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_29),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_31),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_15),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_130),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_110),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_16),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_144),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_107),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_93),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_60),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_86),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_20),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_171),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_48),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_47),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_21),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_122),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_31),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_123),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_29),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_100),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_74),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_65),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_19),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_59),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_127),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_65),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_39),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_119),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_152),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_28),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_157),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_0),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_90),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_97),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_53),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_50),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_102),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_44),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_37),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_28),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_18),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_14),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_148),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_121),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_94),
.Y(n_336)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_18),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_67),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_27),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_91),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_64),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_164),
.Y(n_342)
);

BUFx10_ASAP7_75t_L g343 ( 
.A(n_108),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_14),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_337),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_244),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_176),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_244),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_244),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_244),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_244),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_191),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_185),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_247),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_176),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_337),
.B(n_5),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_337),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_218),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_319),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_340),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_283),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_244),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_336),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_244),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_192),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_192),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_182),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_186),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_337),
.B(n_244),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_244),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_193),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_179),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_195),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_197),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_179),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_190),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_190),
.B(n_5),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_210),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_210),
.B(n_6),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_181),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_213),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_277),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_198),
.Y(n_383)
);

NOR2xp67_ASAP7_75t_L g384 ( 
.A(n_175),
.B(n_7),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_213),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_200),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_220),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_220),
.B(n_7),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_226),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_226),
.B(n_9),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_201),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_209),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_211),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_231),
.Y(n_394)
);

INVxp33_ASAP7_75t_SL g395 ( 
.A(n_277),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_219),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_272),
.B(n_307),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_221),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_217),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_302),
.Y(n_400)
);

INVxp67_ASAP7_75t_SL g401 ( 
.A(n_177),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_231),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_230),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_302),
.B(n_9),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_339),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_340),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_233),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_236),
.Y(n_408)
);

NOR2xp67_ASAP7_75t_L g409 ( 
.A(n_175),
.B(n_10),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_242),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_233),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_259),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_339),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_252),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_177),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_255),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_259),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_261),
.Y(n_418)
);

INVxp67_ASAP7_75t_SL g419 ( 
.A(n_183),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_281),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_281),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_262),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_265),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_224),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_339),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_228),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_257),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_268),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_271),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_297),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_350),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_369),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_352),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_358),
.Y(n_434)
);

AND2x6_ASAP7_75t_L g435 ( 
.A(n_380),
.B(n_225),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_350),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_380),
.B(n_199),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_369),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_350),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_359),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_346),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_346),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_348),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_348),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g445 ( 
.A(n_367),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_363),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_R g447 ( 
.A(n_368),
.B(n_173),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_371),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_349),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_366),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_349),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_351),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_351),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_373),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_374),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_362),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_362),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_366),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_364),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_364),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_383),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_370),
.Y(n_462)
);

OA21x2_ASAP7_75t_L g463 ( 
.A1(n_372),
.A2(n_298),
.B(n_297),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_370),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_345),
.B(n_298),
.Y(n_465)
);

CKINVDCx14_ASAP7_75t_R g466 ( 
.A(n_353),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_391),
.Y(n_467)
);

BUFx8_ASAP7_75t_L g468 ( 
.A(n_404),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_392),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_372),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_345),
.B(n_311),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_375),
.Y(n_472)
);

BUFx8_ASAP7_75t_L g473 ( 
.A(n_404),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_375),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_380),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_393),
.Y(n_476)
);

NAND2x1_ASAP7_75t_L g477 ( 
.A(n_376),
.B(n_323),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_376),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_360),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_397),
.B(n_311),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_400),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_357),
.B(n_378),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_396),
.Y(n_483)
);

CKINVDCx11_ASAP7_75t_R g484 ( 
.A(n_386),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_378),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_381),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_398),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_381),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_385),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_385),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_387),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_387),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_403),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_R g494 ( 
.A(n_408),
.B(n_174),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_389),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_357),
.B(n_199),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_410),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_414),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_389),
.B(n_199),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_R g500 ( 
.A(n_416),
.B(n_178),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_394),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_394),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_402),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_402),
.Y(n_504)
);

AND3x2_ASAP7_75t_L g505 ( 
.A(n_347),
.B(n_365),
.C(n_355),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_407),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_418),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_478),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_478),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_447),
.B(n_360),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_478),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_478),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_436),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_478),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_482),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_436),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_482),
.B(n_401),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_436),
.Y(n_518)
);

AND2x6_ASAP7_75t_L g519 ( 
.A(n_432),
.B(n_316),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_484),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_432),
.B(n_406),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_478),
.Y(n_522)
);

INVx4_ASAP7_75t_L g523 ( 
.A(n_475),
.Y(n_523)
);

NAND2xp33_ASAP7_75t_SL g524 ( 
.A(n_448),
.B(n_422),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_438),
.B(n_406),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_494),
.B(n_423),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_482),
.B(n_405),
.Y(n_527)
);

AND2x4_ASAP7_75t_SL g528 ( 
.A(n_450),
.B(n_354),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_496),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_438),
.B(n_407),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_439),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_431),
.Y(n_532)
);

NOR3xp33_ASAP7_75t_L g533 ( 
.A(n_480),
.B(n_379),
.C(n_377),
.Y(n_533)
);

OAI22xp33_ASAP7_75t_SL g534 ( 
.A1(n_480),
.A2(n_397),
.B1(n_395),
.B2(n_465),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_475),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_491),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_491),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_445),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_465),
.B(n_428),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_491),
.Y(n_540)
);

CKINVDCx16_ASAP7_75t_R g541 ( 
.A(n_479),
.Y(n_541)
);

INVxp67_ASAP7_75t_SL g542 ( 
.A(n_475),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_431),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_491),
.Y(n_544)
);

AND2x2_ASAP7_75t_SL g545 ( 
.A(n_463),
.B(n_356),
.Y(n_545)
);

AND2x2_ASAP7_75t_SL g546 ( 
.A(n_463),
.B(n_225),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_496),
.B(n_411),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_491),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_496),
.B(n_401),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_491),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_500),
.B(n_429),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_437),
.B(n_411),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_492),
.Y(n_553)
);

BUFx10_ASAP7_75t_L g554 ( 
.A(n_454),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_492),
.Y(n_555)
);

AOI22x1_ASAP7_75t_L g556 ( 
.A1(n_456),
.A2(n_419),
.B1(n_282),
.B2(n_415),
.Y(n_556)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_475),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_475),
.Y(n_558)
);

AND2x6_ASAP7_75t_L g559 ( 
.A(n_506),
.B(n_316),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_475),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_471),
.B(n_347),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_439),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_431),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_471),
.B(n_355),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_470),
.B(n_365),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_492),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_455),
.B(n_382),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_431),
.Y(n_568)
);

BUFx10_ASAP7_75t_L g569 ( 
.A(n_461),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_492),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_443),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_439),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_431),
.Y(n_573)
);

INVxp67_ASAP7_75t_SL g574 ( 
.A(n_492),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_499),
.B(n_405),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_441),
.Y(n_576)
);

INVxp67_ASAP7_75t_SL g577 ( 
.A(n_492),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_441),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_441),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_503),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_443),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_503),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_437),
.B(n_412),
.Y(n_583)
);

INVx1_ASAP7_75t_SL g584 ( 
.A(n_445),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_503),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_437),
.B(n_412),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_463),
.A2(n_390),
.B1(n_388),
.B2(n_382),
.Y(n_587)
);

AO22x2_ASAP7_75t_L g588 ( 
.A1(n_468),
.A2(n_419),
.B1(n_417),
.B2(n_421),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_503),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_467),
.B(n_384),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_449),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_437),
.B(n_417),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_442),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_470),
.B(n_361),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_469),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_503),
.Y(n_596)
);

NAND2x1p5_ASAP7_75t_L g597 ( 
.A(n_463),
.B(n_420),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_503),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_442),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_476),
.B(n_384),
.Y(n_600)
);

NOR2x1p5_ASAP7_75t_L g601 ( 
.A(n_483),
.B(n_183),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_442),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_457),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_457),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_457),
.Y(n_605)
);

INVx4_ASAP7_75t_SL g606 ( 
.A(n_435),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_444),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_449),
.Y(n_608)
);

INVx4_ASAP7_75t_SL g609 ( 
.A(n_435),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_444),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_463),
.A2(n_400),
.B1(n_409),
.B2(n_421),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_499),
.B(n_413),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_506),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_456),
.Y(n_614)
);

NAND2x1p5_ASAP7_75t_L g615 ( 
.A(n_477),
.B(n_420),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_506),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_431),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_472),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_472),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_444),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_474),
.B(n_430),
.Y(n_621)
);

AND2x2_ASAP7_75t_SL g622 ( 
.A(n_479),
.B(n_245),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_474),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_499),
.B(n_415),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_468),
.A2(n_409),
.B1(n_260),
.B2(n_317),
.Y(n_625)
);

AND2x6_ASAP7_75t_L g626 ( 
.A(n_485),
.B(n_325),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_444),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_485),
.B(n_430),
.Y(n_628)
);

INVx4_ASAP7_75t_L g629 ( 
.A(n_444),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_499),
.A2(n_222),
.B1(n_314),
.B2(n_250),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_505),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_444),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_451),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_456),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_456),
.Y(n_635)
);

OR2x6_ASAP7_75t_L g636 ( 
.A(n_468),
.B(n_222),
.Y(n_636)
);

INVx5_ASAP7_75t_L g637 ( 
.A(n_435),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_486),
.B(n_413),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_486),
.B(n_425),
.Y(n_639)
);

OR2x6_ASAP7_75t_L g640 ( 
.A(n_468),
.B(n_425),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_488),
.B(n_334),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_488),
.B(n_489),
.Y(n_642)
);

BUFx8_ASAP7_75t_SL g643 ( 
.A(n_433),
.Y(n_643)
);

HB1xp67_ASAP7_75t_L g644 ( 
.A(n_434),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_489),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_490),
.B(n_305),
.Y(n_646)
);

INVx1_ASAP7_75t_SL g647 ( 
.A(n_440),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_487),
.B(n_187),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_SL g649 ( 
.A(n_493),
.B(n_497),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_490),
.B(n_334),
.Y(n_650)
);

OR2x2_ASAP7_75t_L g651 ( 
.A(n_450),
.B(n_240),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_452),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_452),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_495),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_498),
.B(n_187),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_495),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_501),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_459),
.Y(n_658)
);

INVx1_ASAP7_75t_SL g659 ( 
.A(n_446),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_501),
.B(n_305),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_539),
.B(n_502),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_561),
.B(n_502),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_549),
.B(n_507),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_549),
.B(n_473),
.Y(n_664)
);

INVxp67_ASAP7_75t_L g665 ( 
.A(n_584),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_564),
.B(n_504),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_529),
.B(n_504),
.Y(n_667)
);

O2A1O1Ixp33_ASAP7_75t_L g668 ( 
.A1(n_533),
.A2(n_451),
.B(n_453),
.C(n_464),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_513),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_549),
.B(n_473),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_549),
.B(n_529),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_515),
.B(n_459),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_515),
.B(n_459),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_517),
.B(n_459),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_613),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_517),
.B(n_505),
.Y(n_676)
);

NOR2xp67_ASAP7_75t_L g677 ( 
.A(n_637),
.B(n_453),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_513),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_517),
.B(n_547),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_517),
.B(n_460),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_613),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_643),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_574),
.A2(n_462),
.B(n_460),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_527),
.B(n_462),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_519),
.A2(n_473),
.B1(n_481),
.B2(n_458),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_527),
.B(n_464),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_616),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_639),
.B(n_473),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_554),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_519),
.A2(n_435),
.B1(n_321),
.B2(n_325),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_519),
.A2(n_481),
.B1(n_458),
.B2(n_435),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_530),
.B(n_452),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_651),
.B(n_399),
.Y(n_693)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_595),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_521),
.B(n_452),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_516),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_516),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_525),
.B(n_466),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_565),
.B(n_452),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_567),
.B(n_424),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_518),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_575),
.B(n_452),
.Y(n_702)
);

INVx8_ASAP7_75t_L g703 ( 
.A(n_640),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_649),
.B(n_187),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_575),
.B(n_612),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_624),
.B(n_187),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_612),
.B(n_435),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_587),
.B(n_435),
.Y(n_708)
);

AO22x1_ASAP7_75t_L g709 ( 
.A1(n_519),
.A2(n_626),
.B1(n_559),
.B2(n_624),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_556),
.B(n_435),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_616),
.Y(n_711)
);

NAND2x1p5_ASAP7_75t_L g712 ( 
.A(n_637),
.B(n_477),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_519),
.A2(n_343),
.B1(n_279),
.B2(n_229),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_519),
.A2(n_588),
.B1(n_611),
.B2(n_622),
.Y(n_714)
);

INVxp67_ASAP7_75t_SL g715 ( 
.A(n_571),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_556),
.B(n_250),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_552),
.B(n_251),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_624),
.B(n_229),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_538),
.B(n_594),
.Y(n_719)
);

INVx2_ASAP7_75t_SL g720 ( 
.A(n_622),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_624),
.B(n_229),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_631),
.B(n_622),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_519),
.A2(n_343),
.B1(n_229),
.B2(n_323),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_541),
.Y(n_724)
);

OR2x6_ASAP7_75t_L g725 ( 
.A(n_640),
.B(n_251),
.Y(n_725)
);

NOR2x2_ASAP7_75t_L g726 ( 
.A(n_636),
.B(n_314),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_583),
.B(n_305),
.Y(n_727)
);

OAI22x1_ASAP7_75t_SL g728 ( 
.A1(n_520),
.A2(n_427),
.B1(n_426),
.B2(n_344),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_586),
.B(n_308),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_592),
.B(n_308),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_588),
.A2(n_343),
.B1(n_323),
.B2(n_308),
.Y(n_731)
);

OR2x2_ASAP7_75t_SL g732 ( 
.A(n_541),
.B(n_184),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_554),
.Y(n_733)
);

NOR3xp33_ASAP7_75t_SL g734 ( 
.A(n_524),
.B(n_275),
.C(n_273),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_640),
.B(n_184),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_647),
.B(n_276),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_659),
.B(n_280),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_571),
.B(n_342),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_588),
.A2(n_343),
.B1(n_323),
.B2(n_294),
.Y(n_739)
);

INVx8_ASAP7_75t_L g740 ( 
.A(n_640),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_SL g741 ( 
.A(n_644),
.B(n_285),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_518),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_588),
.A2(n_323),
.B1(n_181),
.B2(n_258),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_545),
.A2(n_323),
.B1(n_181),
.B2(n_258),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_581),
.B(n_342),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_603),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_534),
.A2(n_212),
.B1(n_180),
.B2(n_335),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_581),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_626),
.A2(n_326),
.B1(n_338),
.B2(n_288),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_534),
.B(n_289),
.Y(n_750)
);

NOR2xp67_ASAP7_75t_L g751 ( 
.A(n_637),
.B(n_258),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_631),
.B(n_290),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_603),
.Y(n_753)
);

A2O1A1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_618),
.A2(n_206),
.B(n_333),
.C(n_331),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_604),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_577),
.A2(n_245),
.B(n_324),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_604),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_591),
.B(n_189),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_591),
.B(n_189),
.Y(n_759)
);

INVxp67_ASAP7_75t_SL g760 ( 
.A(n_608),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_608),
.B(n_633),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_633),
.B(n_196),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_626),
.A2(n_291),
.B1(n_292),
.B2(n_332),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_626),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_618),
.B(n_196),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_542),
.A2(n_204),
.B(n_328),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_531),
.Y(n_767)
);

O2A1O1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_642),
.A2(n_341),
.B(n_333),
.C(n_331),
.Y(n_768)
);

O2A1O1Ixp5_ASAP7_75t_L g769 ( 
.A1(n_570),
.A2(n_341),
.B(n_202),
.C(n_206),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_SL g770 ( 
.A(n_595),
.B(n_293),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_619),
.B(n_202),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_545),
.A2(n_294),
.B1(n_309),
.B2(n_320),
.Y(n_772)
);

O2A1O1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_619),
.A2(n_306),
.B(n_329),
.C(n_327),
.Y(n_773)
);

NOR3x1_ASAP7_75t_L g774 ( 
.A(n_651),
.B(n_306),
.C(n_329),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_531),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_562),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_623),
.B(n_232),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_554),
.B(n_300),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_638),
.B(n_232),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_510),
.B(n_310),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_569),
.B(n_312),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_526),
.B(n_315),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_562),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_614),
.A2(n_188),
.B(n_194),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_569),
.B(n_318),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_572),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_605),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_545),
.A2(n_203),
.B1(n_205),
.B2(n_322),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_626),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_605),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_SL g791 ( 
.A(n_569),
.B(n_330),
.Y(n_791)
);

BUFx4f_ASAP7_75t_L g792 ( 
.A(n_626),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_623),
.B(n_645),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_551),
.B(n_207),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_648),
.B(n_234),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_645),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_572),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_654),
.A2(n_327),
.B1(n_270),
.B2(n_313),
.Y(n_798)
);

OR2x2_ASAP7_75t_L g799 ( 
.A(n_528),
.B(n_234),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_655),
.B(n_248),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_590),
.B(n_248),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_625),
.B(n_208),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_654),
.B(n_267),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_576),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_614),
.A2(n_266),
.B(n_215),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_626),
.A2(n_214),
.B1(n_216),
.B2(n_223),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_656),
.Y(n_807)
);

AND2x6_ASAP7_75t_SL g808 ( 
.A(n_636),
.B(n_267),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_576),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_656),
.B(n_270),
.Y(n_810)
);

HB1xp67_ASAP7_75t_L g811 ( 
.A(n_528),
.Y(n_811)
);

OAI22xp33_ASAP7_75t_L g812 ( 
.A1(n_636),
.A2(n_313),
.B1(n_304),
.B2(n_296),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_625),
.B(n_227),
.Y(n_813)
);

NAND2xp33_ASAP7_75t_L g814 ( 
.A(n_597),
.B(n_237),
.Y(n_814)
);

NAND2xp33_ASAP7_75t_SL g815 ( 
.A(n_601),
.B(n_296),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_657),
.B(n_304),
.Y(n_816)
);

AND2x6_ASAP7_75t_SL g817 ( 
.A(n_636),
.B(n_13),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_657),
.B(n_235),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_600),
.B(n_239),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_614),
.B(n_241),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_636),
.B(n_294),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_634),
.B(n_243),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_L g823 ( 
.A1(n_634),
.A2(n_320),
.B1(n_309),
.B2(n_303),
.Y(n_823)
);

NOR2x2_ASAP7_75t_L g824 ( 
.A(n_601),
.B(n_13),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_634),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_646),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_635),
.B(n_246),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_635),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_578),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_635),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_658),
.B(n_249),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_658),
.B(n_254),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_621),
.B(n_256),
.Y(n_833)
);

INVxp67_ASAP7_75t_SL g834 ( 
.A(n_715),
.Y(n_834)
);

HB1xp67_ASAP7_75t_L g835 ( 
.A(n_665),
.Y(n_835)
);

INVxp67_ASAP7_75t_SL g836 ( 
.A(n_760),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_714),
.A2(n_546),
.B1(n_559),
.B2(n_630),
.Y(n_837)
);

BUFx8_ASAP7_75t_L g838 ( 
.A(n_733),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_662),
.B(n_666),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_719),
.B(n_628),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_792),
.B(n_658),
.Y(n_841)
);

BUFx2_ASAP7_75t_L g842 ( 
.A(n_724),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_671),
.B(n_606),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_671),
.B(n_606),
.Y(n_844)
);

AO22x1_ASAP7_75t_L g845 ( 
.A1(n_700),
.A2(n_559),
.B1(n_637),
.B2(n_641),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_669),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_733),
.B(n_606),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_703),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_796),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_661),
.B(n_650),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_R g851 ( 
.A(n_689),
.B(n_546),
.Y(n_851)
);

BUFx4f_ASAP7_75t_L g852 ( 
.A(n_725),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_R g853 ( 
.A(n_689),
.B(n_546),
.Y(n_853)
);

NAND3xp33_ASAP7_75t_L g854 ( 
.A(n_770),
.B(n_508),
.C(n_509),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_796),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_792),
.B(n_620),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_679),
.B(n_578),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_694),
.B(n_698),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_703),
.Y(n_859)
);

BUFx2_ASAP7_75t_R g860 ( 
.A(n_682),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_743),
.A2(n_559),
.B1(n_579),
.B2(n_593),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_722),
.B(n_610),
.Y(n_862)
);

BUFx4f_ASAP7_75t_L g863 ( 
.A(n_725),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_807),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_792),
.B(n_764),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_684),
.B(n_579),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_686),
.B(n_593),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_764),
.B(n_620),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_669),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_705),
.B(n_599),
.Y(n_870)
);

INVx4_ASAP7_75t_L g871 ( 
.A(n_703),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_693),
.B(n_615),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_811),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_674),
.B(n_599),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_748),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_720),
.B(n_610),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_720),
.B(n_606),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_678),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_725),
.B(n_609),
.Y(n_879)
);

AND3x1_ASAP7_75t_SL g880 ( 
.A(n_824),
.B(n_15),
.C(n_16),
.Y(n_880)
);

NOR3xp33_ASAP7_75t_SL g881 ( 
.A(n_682),
.B(n_660),
.C(n_274),
.Y(n_881)
);

NAND2xp33_ASAP7_75t_SL g882 ( 
.A(n_807),
.B(n_570),
.Y(n_882)
);

OR2x2_ASAP7_75t_L g883 ( 
.A(n_693),
.B(n_615),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_676),
.Y(n_884)
);

BUFx8_ASAP7_75t_L g885 ( 
.A(n_821),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_793),
.A2(n_629),
.B1(n_610),
.B2(n_597),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_703),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_748),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_678),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_696),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_725),
.B(n_609),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_724),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_664),
.B(n_609),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_744),
.A2(n_559),
.B1(n_602),
.B2(n_597),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_740),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_741),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_740),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_789),
.B(n_620),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_680),
.B(n_602),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_779),
.B(n_629),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_696),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_779),
.B(n_629),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_740),
.Y(n_903)
);

INVx1_ASAP7_75t_SL g904 ( 
.A(n_799),
.Y(n_904)
);

OR2x6_ASAP7_75t_L g905 ( 
.A(n_740),
.B(n_709),
.Y(n_905)
);

INVx1_ASAP7_75t_SL g906 ( 
.A(n_799),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_748),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_670),
.B(n_609),
.Y(n_908)
);

OR2x6_ASAP7_75t_SL g909 ( 
.A(n_791),
.B(n_264),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_735),
.Y(n_910)
);

BUFx3_ASAP7_75t_L g911 ( 
.A(n_825),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_735),
.Y(n_912)
);

AND2x6_ASAP7_75t_L g913 ( 
.A(n_690),
.B(n_607),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_697),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_789),
.B(n_620),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_825),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_735),
.B(n_637),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_663),
.B(n_750),
.Y(n_918)
);

BUFx2_ASAP7_75t_L g919 ( 
.A(n_732),
.Y(n_919)
);

BUFx10_ASAP7_75t_L g920 ( 
.A(n_780),
.Y(n_920)
);

BUFx3_ASAP7_75t_L g921 ( 
.A(n_828),
.Y(n_921)
);

INVx5_ASAP7_75t_L g922 ( 
.A(n_817),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_R g923 ( 
.A(n_815),
.B(n_585),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_675),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_688),
.B(n_620),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_695),
.B(n_585),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_728),
.Y(n_927)
);

AND3x1_ASAP7_75t_SL g928 ( 
.A(n_824),
.B(n_830),
.C(n_828),
.Y(n_928)
);

CKINVDCx20_ASAP7_75t_R g929 ( 
.A(n_732),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_667),
.B(n_585),
.Y(n_930)
);

CKINVDCx20_ASAP7_75t_R g931 ( 
.A(n_826),
.Y(n_931)
);

INVx5_ASAP7_75t_L g932 ( 
.A(n_808),
.Y(n_932)
);

INVxp67_ASAP7_75t_L g933 ( 
.A(n_815),
.Y(n_933)
);

INVxp67_ASAP7_75t_L g934 ( 
.A(n_801),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_702),
.B(n_589),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_758),
.B(n_589),
.Y(n_936)
);

NOR3xp33_ASAP7_75t_SL g937 ( 
.A(n_778),
.B(n_286),
.C(n_284),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_668),
.A2(n_589),
.B(n_598),
.C(n_509),
.Y(n_938)
);

OR2x2_ASAP7_75t_L g939 ( 
.A(n_802),
.B(n_615),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_821),
.B(n_637),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_R g941 ( 
.A(n_826),
.B(n_598),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_697),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_759),
.B(n_598),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_728),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_762),
.B(n_699),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_726),
.Y(n_946)
);

INVx2_ASAP7_75t_SL g947 ( 
.A(n_704),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_761),
.B(n_627),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_683),
.A2(n_653),
.B(n_607),
.Y(n_949)
);

AND2x6_ASAP7_75t_L g950 ( 
.A(n_690),
.B(n_632),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_691),
.B(n_570),
.Y(n_951)
);

BUFx2_ASAP7_75t_L g952 ( 
.A(n_726),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_706),
.B(n_558),
.Y(n_953)
);

INVx4_ASAP7_75t_L g954 ( 
.A(n_712),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_712),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_R g956 ( 
.A(n_814),
.B(n_508),
.Y(n_956)
);

NAND3xp33_ASAP7_75t_L g957 ( 
.A(n_749),
.B(n_566),
.C(n_550),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_672),
.B(n_511),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_701),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_681),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_774),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_749),
.B(n_627),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_712),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_763),
.B(n_627),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_734),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_673),
.B(n_511),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_SL g967 ( 
.A(n_812),
.B(n_559),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_687),
.Y(n_968)
);

NOR2xp67_ASAP7_75t_L g969 ( 
.A(n_782),
.B(n_512),
.Y(n_969)
);

HB1xp67_ASAP7_75t_L g970 ( 
.A(n_774),
.Y(n_970)
);

BUFx2_ASAP7_75t_L g971 ( 
.A(n_763),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_795),
.B(n_512),
.Y(n_972)
);

INVx6_ASAP7_75t_L g973 ( 
.A(n_709),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_687),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_713),
.A2(n_536),
.B1(n_553),
.B2(n_555),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_711),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_804),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_813),
.B(n_632),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_800),
.B(n_514),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_711),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_701),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_746),
.Y(n_982)
);

NOR3xp33_ASAP7_75t_SL g983 ( 
.A(n_781),
.B(n_785),
.C(n_737),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_717),
.B(n_746),
.Y(n_984)
);

HB1xp67_ASAP7_75t_L g985 ( 
.A(n_738),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_718),
.B(n_558),
.Y(n_986)
);

INVx3_ASAP7_75t_L g987 ( 
.A(n_830),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_753),
.B(n_514),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_753),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_742),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_755),
.B(n_522),
.Y(n_991)
);

AOI21xp33_ASAP7_75t_L g992 ( 
.A1(n_788),
.A2(n_540),
.B(n_522),
.Y(n_992)
);

BUFx4f_ASAP7_75t_L g993 ( 
.A(n_755),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_757),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_721),
.B(n_559),
.Y(n_995)
);

INVx2_ASAP7_75t_SL g996 ( 
.A(n_752),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_757),
.B(n_536),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_692),
.A2(n_653),
.B(n_557),
.Y(n_998)
);

INVx6_ASAP7_75t_L g999 ( 
.A(n_794),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_787),
.B(n_627),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_787),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_790),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_685),
.B(n_537),
.Y(n_1003)
);

INVx4_ASAP7_75t_L g1004 ( 
.A(n_804),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_790),
.Y(n_1005)
);

NAND3xp33_ASAP7_75t_SL g1006 ( 
.A(n_747),
.B(n_278),
.C(n_269),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_742),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_765),
.B(n_537),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_767),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_707),
.A2(n_544),
.B(n_548),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_771),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_777),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_819),
.A2(n_544),
.B1(n_540),
.B2(n_548),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_803),
.B(n_550),
.Y(n_1014)
);

INVx4_ASAP7_75t_L g1015 ( 
.A(n_809),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_R g1016 ( 
.A(n_814),
.B(n_553),
.Y(n_1016)
);

NOR2xp67_ASAP7_75t_L g1017 ( 
.A(n_745),
.B(n_555),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_810),
.B(n_566),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_708),
.A2(n_580),
.B(n_582),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_816),
.B(n_580),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_736),
.B(n_582),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_R g1022 ( 
.A(n_731),
.B(n_596),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_818),
.B(n_596),
.Y(n_1023)
);

AO21x1_ASAP7_75t_L g1024 ( 
.A1(n_710),
.A2(n_716),
.B(n_730),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_993),
.B(n_532),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_1019),
.A2(n_769),
.B(n_809),
.Y(n_1026)
);

OAI21x1_ASAP7_75t_L g1027 ( 
.A1(n_1024),
.A2(n_829),
.B(n_776),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_840),
.B(n_739),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_934),
.B(n_833),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_839),
.A2(n_773),
.B(n_768),
.C(n_772),
.Y(n_1030)
);

AOI21x1_ASAP7_75t_L g1031 ( 
.A1(n_925),
.A2(n_751),
.B(n_729),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_882),
.A2(n_832),
.B(n_831),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_859),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_993),
.A2(n_827),
.B1(n_822),
.B2(n_820),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_882),
.A2(n_850),
.B(n_866),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_867),
.A2(n_727),
.B(n_829),
.Y(n_1036)
);

BUFx3_ASAP7_75t_L g1037 ( 
.A(n_838),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1011),
.B(n_798),
.Y(n_1038)
);

AOI22xp33_ASAP7_75t_L g1039 ( 
.A1(n_971),
.A2(n_723),
.B1(n_786),
.B2(n_775),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_926),
.A2(n_783),
.B(n_767),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_973),
.A2(n_806),
.B1(n_823),
.B2(n_805),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_1012),
.A2(n_754),
.B(n_786),
.C(n_783),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_846),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_858),
.B(n_775),
.Y(n_1044)
);

NOR2x1_ASAP7_75t_SL g1045 ( 
.A(n_905),
.B(n_776),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_945),
.A2(n_797),
.B(n_784),
.Y(n_1046)
);

AOI21x1_ASAP7_75t_SL g1047 ( 
.A1(n_930),
.A2(n_756),
.B(n_523),
.Y(n_1047)
);

OA22x2_ASAP7_75t_L g1048 ( 
.A1(n_919),
.A2(n_797),
.B1(n_560),
.B2(n_557),
.Y(n_1048)
);

NAND2x1p5_ASAP7_75t_L g1049 ( 
.A(n_871),
.B(n_677),
.Y(n_1049)
);

O2A1O1Ixp5_ASAP7_75t_L g1050 ( 
.A1(n_925),
.A2(n_523),
.B(n_535),
.C(n_557),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_849),
.Y(n_1051)
);

AO21x2_ASAP7_75t_L g1052 ( 
.A1(n_948),
.A2(n_964),
.B(n_962),
.Y(n_1052)
);

OAI21x1_ASAP7_75t_L g1053 ( 
.A1(n_949),
.A2(n_751),
.B(n_677),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_938),
.A2(n_766),
.B(n_535),
.Y(n_1054)
);

CKINVDCx11_ASAP7_75t_R g1055 ( 
.A(n_931),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_846),
.Y(n_1056)
);

NAND3xp33_ASAP7_75t_L g1057 ( 
.A(n_967),
.B(n_652),
.C(n_627),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_1023),
.A2(n_886),
.B(n_984),
.Y(n_1058)
);

NOR2xp67_ASAP7_75t_L g1059 ( 
.A(n_896),
.B(n_835),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_985),
.B(n_652),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_973),
.A2(n_523),
.B1(n_535),
.B2(n_560),
.Y(n_1061)
);

AOI21xp33_ASAP7_75t_L g1062 ( 
.A1(n_883),
.A2(n_563),
.B(n_617),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_948),
.A2(n_532),
.B(n_617),
.Y(n_1063)
);

AOI21xp33_ASAP7_75t_L g1064 ( 
.A1(n_862),
.A2(n_902),
.B(n_900),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_973),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_869),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_998),
.A2(n_560),
.B(n_617),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_872),
.B(n_532),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_SL g1069 ( 
.A1(n_1010),
.A2(n_652),
.B(n_617),
.Y(n_1069)
);

AOI21xp33_ASAP7_75t_L g1070 ( 
.A1(n_862),
.A2(n_978),
.B(n_837),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_855),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_884),
.B(n_933),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_904),
.B(n_652),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_920),
.B(n_652),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_841),
.A2(n_617),
.B(n_573),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_938),
.A2(n_287),
.B(n_295),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_962),
.A2(n_573),
.B(n_568),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_941),
.Y(n_1078)
);

OR2x2_ASAP7_75t_L g1079 ( 
.A(n_906),
.B(n_532),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_841),
.A2(n_573),
.B(n_568),
.Y(n_1080)
);

CKINVDCx8_ASAP7_75t_R g1081 ( 
.A(n_892),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_964),
.A2(n_573),
.B(n_568),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_910),
.B(n_532),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_988),
.A2(n_573),
.B(n_568),
.Y(n_1084)
);

AO31x2_ASAP7_75t_L g1085 ( 
.A1(n_978),
.A2(n_568),
.A3(n_563),
.B(n_543),
.Y(n_1085)
);

AOI21x1_ASAP7_75t_L g1086 ( 
.A1(n_1000),
.A2(n_563),
.B(n_543),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_L g1087 ( 
.A1(n_1000),
.A2(n_563),
.B(n_543),
.Y(n_1087)
);

OA21x2_ASAP7_75t_L g1088 ( 
.A1(n_992),
.A2(n_299),
.B(n_301),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_912),
.B(n_563),
.Y(n_1089)
);

AOI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_931),
.A2(n_543),
.B1(n_320),
.B2(n_309),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_856),
.A2(n_543),
.B(n_238),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_1005),
.B(n_851),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_1005),
.A2(n_864),
.B1(n_837),
.B2(n_836),
.Y(n_1093)
);

BUFx4f_ASAP7_75t_L g1094 ( 
.A(n_905),
.Y(n_1094)
);

OAI22x1_ASAP7_75t_L g1095 ( 
.A1(n_918),
.A2(n_17),
.B1(n_19),
.B2(n_24),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_851),
.B(n_263),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_856),
.A2(n_238),
.B(n_237),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_991),
.A2(n_238),
.B(n_237),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_870),
.A2(n_17),
.B(n_27),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_834),
.B(n_30),
.Y(n_1100)
);

CKINVDCx16_ASAP7_75t_R g1101 ( 
.A(n_909),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_924),
.A2(n_974),
.B1(n_976),
.B2(n_980),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_SL g1103 ( 
.A1(n_905),
.A2(n_263),
.B(n_253),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_920),
.B(n_32),
.Y(n_1104)
);

OA21x2_ASAP7_75t_L g1105 ( 
.A1(n_894),
.A2(n_238),
.B(n_237),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_SL g1106 ( 
.A1(n_960),
.A2(n_32),
.B(n_33),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_968),
.A2(n_263),
.B1(n_253),
.B2(n_35),
.Y(n_1107)
);

INVxp67_ASAP7_75t_L g1108 ( 
.A(n_873),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_997),
.A2(n_238),
.B(n_237),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_894),
.A2(n_238),
.B(n_237),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_869),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_920),
.B(n_33),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_982),
.B(n_34),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_878),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_958),
.A2(n_966),
.B(n_1008),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_1014),
.A2(n_238),
.B(n_237),
.Y(n_1116)
);

BUFx3_ASAP7_75t_L g1117 ( 
.A(n_838),
.Y(n_1117)
);

INVx6_ASAP7_75t_SL g1118 ( 
.A(n_879),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_989),
.B(n_34),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_994),
.B(n_36),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1001),
.B(n_38),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1018),
.A2(n_1020),
.B(n_935),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_941),
.Y(n_1123)
);

NOR2xp67_ASAP7_75t_L g1124 ( 
.A(n_947),
.B(n_82),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_878),
.A2(n_238),
.B(n_237),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_SL g1126 ( 
.A(n_860),
.B(n_253),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_1002),
.A2(n_263),
.B(n_253),
.C(n_40),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_957),
.A2(n_38),
.B(n_39),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_853),
.Y(n_1129)
);

OA21x2_ASAP7_75t_L g1130 ( 
.A1(n_889),
.A2(n_238),
.B(n_237),
.Y(n_1130)
);

AOI21x1_ASAP7_75t_L g1131 ( 
.A1(n_845),
.A2(n_969),
.B(n_1017),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_889),
.A2(n_263),
.B(n_253),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_857),
.B(n_40),
.Y(n_1133)
);

OA21x2_ASAP7_75t_L g1134 ( 
.A1(n_890),
.A2(n_263),
.B(n_253),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_946),
.B(n_41),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_SL g1136 ( 
.A1(n_874),
.A2(n_42),
.B(n_44),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_890),
.A2(n_83),
.B(n_167),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_901),
.A2(n_170),
.B(n_165),
.Y(n_1138)
);

CKINVDCx11_ASAP7_75t_R g1139 ( 
.A(n_842),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_901),
.A2(n_161),
.B(n_151),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_SL g1141 ( 
.A1(n_951),
.A2(n_42),
.B(n_50),
.Y(n_1141)
);

OR2x2_ASAP7_75t_L g1142 ( 
.A(n_939),
.B(n_51),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_914),
.A2(n_959),
.B(n_990),
.Y(n_1143)
);

AOI21x1_ASAP7_75t_L g1144 ( 
.A1(n_936),
.A2(n_943),
.B(n_915),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_914),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_1021),
.A2(n_1006),
.B(n_979),
.C(n_972),
.Y(n_1146)
);

INVxp67_ASAP7_75t_L g1147 ( 
.A(n_961),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_996),
.B(n_51),
.Y(n_1148)
);

AO21x1_ASAP7_75t_L g1149 ( 
.A1(n_876),
.A2(n_915),
.B(n_898),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_871),
.B(n_848),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_942),
.A2(n_147),
.B(n_138),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_942),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_899),
.A2(n_132),
.B(n_128),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_868),
.A2(n_115),
.B(n_113),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_868),
.A2(n_111),
.B(n_109),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_959),
.A2(n_103),
.B(n_99),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_981),
.A2(n_98),
.B(n_89),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_848),
.B(n_75),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_981),
.A2(n_52),
.B(n_53),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_990),
.A2(n_52),
.B(n_56),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1021),
.A2(n_56),
.B(n_57),
.Y(n_1161)
);

AO22x2_ASAP7_75t_L g1162 ( 
.A1(n_927),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_1162)
);

INVxp67_ASAP7_75t_L g1163 ( 
.A(n_970),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1007),
.Y(n_1164)
);

BUFx3_ASAP7_75t_L g1165 ( 
.A(n_838),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1007),
.A2(n_66),
.B(n_67),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_898),
.A2(n_69),
.B(n_70),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1009),
.A2(n_71),
.B(n_72),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1009),
.A2(n_72),
.B(n_73),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_987),
.A2(n_73),
.B(n_74),
.Y(n_1170)
);

AOI21x1_ASAP7_75t_L g1171 ( 
.A1(n_854),
.A2(n_75),
.B(n_1003),
.Y(n_1171)
);

BUFx2_ASAP7_75t_SL g1172 ( 
.A(n_847),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1013),
.A2(n_975),
.B(n_876),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_859),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_987),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_859),
.Y(n_1176)
);

BUFx2_ASAP7_75t_L g1177 ( 
.A(n_853),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_865),
.A2(n_888),
.B(n_875),
.Y(n_1178)
);

AOI21xp33_ASAP7_75t_L g1179 ( 
.A1(n_953),
.A2(n_986),
.B(n_995),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_911),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_911),
.A2(n_921),
.B1(n_916),
.B2(n_907),
.Y(n_1181)
);

AO21x2_ASAP7_75t_L g1182 ( 
.A1(n_956),
.A2(n_1016),
.B(n_1022),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_875),
.A2(n_888),
.B(n_916),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1051),
.Y(n_1184)
);

OR2x6_ASAP7_75t_L g1185 ( 
.A(n_1172),
.B(n_897),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1132),
.A2(n_865),
.B(n_861),
.Y(n_1186)
);

AND2x6_ASAP7_75t_L g1187 ( 
.A(n_1033),
.B(n_891),
.Y(n_1187)
);

AO31x2_ASAP7_75t_L g1188 ( 
.A1(n_1149),
.A2(n_1015),
.A3(n_1004),
.B(n_954),
.Y(n_1188)
);

OA21x2_ASAP7_75t_L g1189 ( 
.A1(n_1116),
.A2(n_861),
.B(n_918),
.Y(n_1189)
);

AND2x6_ASAP7_75t_L g1190 ( 
.A(n_1033),
.B(n_891),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_SL g1191 ( 
.A1(n_1161),
.A2(n_954),
.B(n_1015),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1146),
.A2(n_983),
.B(n_937),
.Y(n_1192)
);

OR2x2_ASAP7_75t_L g1193 ( 
.A(n_1142),
.B(n_952),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1143),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1146),
.A2(n_918),
.B(n_913),
.Y(n_1195)
);

AO31x2_ASAP7_75t_L g1196 ( 
.A1(n_1149),
.A2(n_1004),
.A3(n_950),
.B(n_913),
.Y(n_1196)
);

NAND2x1p5_ASAP7_75t_L g1197 ( 
.A(n_1065),
.B(n_903),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1143),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1071),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1043),
.Y(n_1200)
);

NAND3xp33_ASAP7_75t_L g1201 ( 
.A(n_1128),
.B(n_1099),
.C(n_1127),
.Y(n_1201)
);

INVxp67_ASAP7_75t_SL g1202 ( 
.A(n_1065),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1132),
.A2(n_1016),
.B(n_956),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_1093),
.Y(n_1204)
);

AO31x2_ASAP7_75t_L g1205 ( 
.A1(n_1058),
.A2(n_913),
.A3(n_950),
.B(n_977),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1173),
.A2(n_1029),
.B1(n_1030),
.B2(n_1028),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1077),
.A2(n_977),
.B(n_921),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1098),
.A2(n_913),
.B(n_950),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1038),
.B(n_929),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1098),
.A2(n_913),
.B(n_950),
.Y(n_1210)
);

OAI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1035),
.A2(n_950),
.B(n_986),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_1070),
.B(n_907),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1109),
.A2(n_977),
.B(n_955),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_1064),
.B(n_923),
.Y(n_1214)
);

OA21x2_ASAP7_75t_L g1215 ( 
.A1(n_1116),
.A2(n_953),
.B(n_986),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1043),
.Y(n_1216)
);

O2A1O1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1030),
.A2(n_881),
.B(n_953),
.C(n_880),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1044),
.B(n_929),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1109),
.A2(n_1047),
.B(n_1125),
.Y(n_1219)
);

INVx4_ASAP7_75t_SL g1220 ( 
.A(n_1033),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1122),
.A2(n_852),
.B(n_863),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1100),
.A2(n_852),
.B(n_863),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1056),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1145),
.Y(n_1224)
);

OA21x2_ASAP7_75t_L g1225 ( 
.A1(n_1077),
.A2(n_908),
.B(n_893),
.Y(n_1225)
);

OAI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1095),
.A2(n_922),
.B1(n_932),
.B2(n_944),
.Y(n_1226)
);

CKINVDCx11_ASAP7_75t_R g1227 ( 
.A(n_1081),
.Y(n_1227)
);

AO21x2_ASAP7_75t_L g1228 ( 
.A1(n_1069),
.A2(n_1022),
.B(n_923),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1072),
.B(n_932),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1125),
.A2(n_977),
.B(n_963),
.Y(n_1230)
);

INVx6_ASAP7_75t_L g1231 ( 
.A(n_1150),
.Y(n_1231)
);

OR2x6_ASAP7_75t_L g1232 ( 
.A(n_1129),
.B(n_897),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1082),
.A2(n_963),
.B(n_955),
.Y(n_1233)
);

AND2x4_ASAP7_75t_L g1234 ( 
.A(n_1150),
.B(n_903),
.Y(n_1234)
);

INVx2_ASAP7_75t_SL g1235 ( 
.A(n_1037),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1082),
.A2(n_963),
.B(n_955),
.Y(n_1236)
);

INVx4_ASAP7_75t_L g1237 ( 
.A(n_1117),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1152),
.Y(n_1238)
);

AOI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1086),
.A2(n_893),
.B(n_908),
.Y(n_1239)
);

BUFx12f_ASAP7_75t_L g1240 ( 
.A(n_1055),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1097),
.A2(n_963),
.B(n_955),
.Y(n_1241)
);

NAND3x1_ASAP7_75t_L g1242 ( 
.A(n_1104),
.B(n_880),
.C(n_885),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1056),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1059),
.B(n_885),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_1150),
.B(n_895),
.Y(n_1245)
);

INVx4_ASAP7_75t_L g1246 ( 
.A(n_1117),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1102),
.A2(n_999),
.B1(n_965),
.B2(n_891),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1164),
.Y(n_1248)
);

A2O1A1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1127),
.A2(n_893),
.B(n_908),
.C(n_879),
.Y(n_1249)
);

BUFx3_ASAP7_75t_L g1250 ( 
.A(n_1078),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1097),
.A2(n_928),
.B(n_999),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1055),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_1078),
.Y(n_1253)
);

O2A1O1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1112),
.A2(n_928),
.B(n_847),
.C(n_844),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1066),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1066),
.Y(n_1256)
);

NAND3xp33_ASAP7_75t_L g1257 ( 
.A(n_1076),
.B(n_932),
.C(n_922),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1111),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1111),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1027),
.A2(n_1091),
.B(n_1063),
.Y(n_1260)
);

AND2x4_ASAP7_75t_L g1261 ( 
.A(n_1092),
.B(n_887),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1046),
.A2(n_843),
.B(n_844),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1027),
.A2(n_999),
.B(n_885),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1092),
.B(n_887),
.Y(n_1264)
);

OA21x2_ASAP7_75t_L g1265 ( 
.A1(n_1063),
.A2(n_940),
.B(n_877),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1114),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1091),
.A2(n_1053),
.B(n_1087),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1113),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1053),
.A2(n_887),
.B(n_895),
.Y(n_1269)
);

OA21x2_ASAP7_75t_L g1270 ( 
.A1(n_1087),
.A2(n_940),
.B(n_877),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1130),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1119),
.Y(n_1272)
);

OR2x2_ASAP7_75t_L g1273 ( 
.A(n_1142),
.B(n_887),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1108),
.B(n_932),
.Y(n_1274)
);

AOI221xp5_ASAP7_75t_L g1275 ( 
.A1(n_1135),
.A2(n_922),
.B1(n_844),
.B2(n_843),
.C(n_917),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1130),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1110),
.A2(n_895),
.B(n_859),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1120),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1110),
.A2(n_895),
.B(n_940),
.Y(n_1279)
);

OR2x6_ASAP7_75t_L g1280 ( 
.A(n_1129),
.B(n_879),
.Y(n_1280)
);

OR2x2_ASAP7_75t_L g1281 ( 
.A(n_1079),
.B(n_917),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1121),
.Y(n_1282)
);

O2A1O1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1148),
.A2(n_847),
.B(n_843),
.C(n_917),
.Y(n_1283)
);

NOR2x1_ASAP7_75t_R g1284 ( 
.A(n_1165),
.B(n_922),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1057),
.A2(n_877),
.B1(n_1177),
.B2(n_1123),
.Y(n_1285)
);

AO32x2_ASAP7_75t_L g1286 ( 
.A1(n_1107),
.A2(n_1181),
.A3(n_1034),
.B1(n_1041),
.B2(n_1052),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_1094),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1147),
.Y(n_1288)
);

OR2x2_ASAP7_75t_L g1289 ( 
.A(n_1079),
.B(n_1101),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1133),
.A2(n_1054),
.B(n_1115),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1032),
.A2(n_1084),
.B(n_1115),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1177),
.B(n_1073),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_1174),
.B(n_1068),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1069),
.A2(n_1140),
.B(n_1156),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1137),
.A2(n_1156),
.B(n_1140),
.Y(n_1295)
);

OR2x6_ASAP7_75t_L g1296 ( 
.A(n_1103),
.B(n_1165),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1162),
.A2(n_1095),
.B1(n_1182),
.B2(n_1179),
.Y(n_1297)
);

INVx8_ASAP7_75t_L g1298 ( 
.A(n_1033),
.Y(n_1298)
);

OR2x6_ASAP7_75t_L g1299 ( 
.A(n_1103),
.B(n_1068),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1060),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1175),
.A2(n_1094),
.B1(n_1096),
.B2(n_1158),
.Y(n_1301)
);

CKINVDCx20_ASAP7_75t_R g1302 ( 
.A(n_1081),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1137),
.A2(n_1157),
.B(n_1138),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1042),
.Y(n_1304)
);

BUFx3_ASAP7_75t_L g1305 ( 
.A(n_1174),
.Y(n_1305)
);

OA21x2_ASAP7_75t_L g1306 ( 
.A1(n_1159),
.A2(n_1160),
.B(n_1166),
.Y(n_1306)
);

OAI222xp33_ASAP7_75t_L g1307 ( 
.A1(n_1090),
.A2(n_1096),
.B1(n_1048),
.B2(n_1163),
.C1(n_1162),
.C2(n_1039),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1180),
.B(n_1182),
.Y(n_1308)
);

AO21x2_ASAP7_75t_L g1309 ( 
.A1(n_1052),
.A2(n_1036),
.B(n_1171),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1182),
.B(n_1126),
.Y(n_1310)
);

NAND2x1p5_ASAP7_75t_L g1311 ( 
.A(n_1094),
.B(n_1176),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1138),
.A2(n_1157),
.B(n_1151),
.Y(n_1312)
);

OAI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1061),
.A2(n_1042),
.B(n_1074),
.Y(n_1313)
);

OAI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1162),
.A2(n_1167),
.B1(n_1048),
.B2(n_1089),
.Y(n_1314)
);

NOR2x1_ASAP7_75t_SL g1315 ( 
.A(n_1025),
.B(n_1033),
.Y(n_1315)
);

OA21x2_ASAP7_75t_L g1316 ( 
.A1(n_1159),
.A2(n_1160),
.B(n_1168),
.Y(n_1316)
);

INVxp67_ASAP7_75t_SL g1317 ( 
.A(n_1083),
.Y(n_1317)
);

NAND3xp33_ASAP7_75t_L g1318 ( 
.A(n_1088),
.B(n_1183),
.C(n_1153),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_1045),
.B(n_1176),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1162),
.A2(n_1088),
.B1(n_1105),
.B2(n_1106),
.Y(n_1320)
);

BUFx2_ASAP7_75t_L g1321 ( 
.A(n_1118),
.Y(n_1321)
);

NOR4xp25_ASAP7_75t_L g1322 ( 
.A(n_1025),
.B(n_1062),
.C(n_1106),
.D(n_1141),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_SL g1323 ( 
.A1(n_1088),
.A2(n_1105),
.B1(n_1141),
.B2(n_1136),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1151),
.A2(n_1144),
.B(n_1026),
.Y(n_1324)
);

INVx3_ASAP7_75t_L g1325 ( 
.A(n_1176),
.Y(n_1325)
);

NAND3xp33_ASAP7_75t_L g1326 ( 
.A(n_1154),
.B(n_1155),
.C(n_1124),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1026),
.A2(n_1031),
.B(n_1067),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1176),
.Y(n_1328)
);

CKINVDCx6p67_ASAP7_75t_R g1329 ( 
.A(n_1139),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1118),
.A2(n_1049),
.B1(n_1176),
.B2(n_1105),
.Y(n_1330)
);

AO21x1_ASAP7_75t_L g1331 ( 
.A1(n_1131),
.A2(n_1040),
.B(n_1170),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1139),
.B(n_1118),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_SL g1333 ( 
.A1(n_1075),
.A2(n_1080),
.B(n_1130),
.Y(n_1333)
);

AO31x2_ASAP7_75t_L g1334 ( 
.A1(n_1052),
.A2(n_1085),
.A3(n_1134),
.B(n_1166),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1170),
.B(n_1168),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1134),
.Y(n_1336)
);

O2A1O1Ixp33_ASAP7_75t_SL g1337 ( 
.A1(n_1178),
.A2(n_1050),
.B(n_1085),
.C(n_1169),
.Y(n_1337)
);

BUFx3_ASAP7_75t_L g1338 ( 
.A(n_1178),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_1049),
.Y(n_1339)
);

NAND2xp33_ASAP7_75t_R g1340 ( 
.A(n_1134),
.B(n_1169),
.Y(n_1340)
);

NAND2x1p5_ASAP7_75t_L g1341 ( 
.A(n_1085),
.B(n_1065),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1085),
.A2(n_1132),
.B(n_1109),
.Y(n_1342)
);

INVx3_ASAP7_75t_L g1343 ( 
.A(n_1085),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1143),
.Y(n_1344)
);

AND2x4_ASAP7_75t_L g1345 ( 
.A(n_1065),
.B(n_848),
.Y(n_1345)
);

AND2x4_ASAP7_75t_L g1346 ( 
.A(n_1065),
.B(n_848),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1051),
.Y(n_1347)
);

INVx2_ASAP7_75t_SL g1348 ( 
.A(n_1037),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1200),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1206),
.A2(n_1201),
.B1(n_1297),
.B2(n_1226),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1200),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1295),
.A2(n_1312),
.B(n_1303),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1216),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1209),
.B(n_1193),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1293),
.B(n_1287),
.Y(n_1355)
);

AOI21xp33_ASAP7_75t_L g1356 ( 
.A1(n_1192),
.A2(n_1318),
.B(n_1217),
.Y(n_1356)
);

AND2x4_ASAP7_75t_L g1357 ( 
.A(n_1293),
.B(n_1287),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1293),
.B(n_1287),
.Y(n_1358)
);

INVx5_ASAP7_75t_L g1359 ( 
.A(n_1287),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_1227),
.Y(n_1360)
);

OR2x2_ASAP7_75t_L g1361 ( 
.A(n_1289),
.B(n_1218),
.Y(n_1361)
);

NOR2x1_ASAP7_75t_L g1362 ( 
.A(n_1257),
.B(n_1237),
.Y(n_1362)
);

OR2x6_ASAP7_75t_SL g1363 ( 
.A(n_1252),
.B(n_1244),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1297),
.A2(n_1226),
.B1(n_1204),
.B2(n_1195),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1184),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1199),
.Y(n_1366)
);

NAND2x1p5_ASAP7_75t_L g1367 ( 
.A(n_1345),
.B(n_1346),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1250),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1290),
.A2(n_1291),
.B(n_1326),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1295),
.A2(n_1312),
.B(n_1303),
.Y(n_1370)
);

NAND2xp33_ASAP7_75t_R g1371 ( 
.A(n_1296),
.B(n_1299),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1223),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1347),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1224),
.Y(n_1374)
);

BUFx2_ASAP7_75t_L g1375 ( 
.A(n_1250),
.Y(n_1375)
);

OAI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1204),
.A2(n_1268),
.B1(n_1278),
.B2(n_1272),
.Y(n_1376)
);

AO21x2_ASAP7_75t_L g1377 ( 
.A1(n_1333),
.A2(n_1310),
.B(n_1314),
.Y(n_1377)
);

OA21x2_ASAP7_75t_L g1378 ( 
.A1(n_1324),
.A2(n_1342),
.B(n_1219),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1229),
.B(n_1282),
.Y(n_1379)
);

INVx3_ASAP7_75t_SL g1380 ( 
.A(n_1252),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1211),
.A2(n_1337),
.B(n_1221),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1343),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1229),
.B(n_1202),
.Y(n_1383)
);

INVx2_ASAP7_75t_SL g1384 ( 
.A(n_1237),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1238),
.Y(n_1385)
);

BUFx4f_ASAP7_75t_SL g1386 ( 
.A(n_1302),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1248),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1214),
.A2(n_1212),
.B(n_1313),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1281),
.B(n_1273),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1275),
.A2(n_1320),
.B1(n_1214),
.B2(n_1247),
.Y(n_1390)
);

AOI221xp5_ASAP7_75t_SL g1391 ( 
.A1(n_1254),
.A2(n_1314),
.B1(n_1320),
.B2(n_1288),
.C(n_1274),
.Y(n_1391)
);

OR2x2_ASAP7_75t_L g1392 ( 
.A(n_1253),
.B(n_1300),
.Y(n_1392)
);

OR2x6_ASAP7_75t_L g1393 ( 
.A(n_1296),
.B(n_1299),
.Y(n_1393)
);

CKINVDCx16_ASAP7_75t_R g1394 ( 
.A(n_1240),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1223),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1292),
.B(n_1345),
.Y(n_1396)
);

BUFx2_ASAP7_75t_R g1397 ( 
.A(n_1339),
.Y(n_1397)
);

OAI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1212),
.A2(n_1292),
.B(n_1242),
.Y(n_1398)
);

INVx4_ASAP7_75t_L g1399 ( 
.A(n_1298),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1332),
.B(n_1235),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1332),
.B(n_1348),
.Y(n_1401)
);

AOI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1242),
.A2(n_1301),
.B1(n_1261),
.B2(n_1264),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1256),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_1240),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1258),
.Y(n_1405)
);

NAND2x1_ASAP7_75t_L g1406 ( 
.A(n_1191),
.B(n_1325),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_L g1407 ( 
.A(n_1187),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_SL g1408 ( 
.A1(n_1222),
.A2(n_1307),
.B1(n_1189),
.B2(n_1296),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1253),
.A2(n_1302),
.B1(n_1249),
.B2(n_1339),
.Y(n_1409)
);

O2A1O1Ixp33_ASAP7_75t_SL g1410 ( 
.A1(n_1249),
.A2(n_1262),
.B(n_1308),
.C(n_1304),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1243),
.Y(n_1411)
);

BUFx2_ASAP7_75t_L g1412 ( 
.A(n_1246),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1189),
.A2(n_1264),
.B1(n_1261),
.B2(n_1280),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1266),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1261),
.B(n_1264),
.Y(n_1415)
);

INVx2_ASAP7_75t_SL g1416 ( 
.A(n_1246),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1251),
.A2(n_1317),
.B(n_1322),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1243),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1255),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1329),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1255),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1259),
.Y(n_1422)
);

BUFx12f_ASAP7_75t_L g1423 ( 
.A(n_1321),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_SL g1424 ( 
.A1(n_1323),
.A2(n_1231),
.B1(n_1232),
.B2(n_1299),
.Y(n_1424)
);

BUFx3_ASAP7_75t_L g1425 ( 
.A(n_1305),
.Y(n_1425)
);

OR2x6_ASAP7_75t_L g1426 ( 
.A(n_1311),
.B(n_1280),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1219),
.A2(n_1294),
.B(n_1342),
.Y(n_1427)
);

BUFx2_ASAP7_75t_SL g1428 ( 
.A(n_1305),
.Y(n_1428)
);

OAI222xp33_ASAP7_75t_L g1429 ( 
.A1(n_1280),
.A2(n_1283),
.B1(n_1232),
.B2(n_1285),
.C1(n_1185),
.C2(n_1311),
.Y(n_1429)
);

AND2x4_ASAP7_75t_L g1430 ( 
.A(n_1319),
.B(n_1220),
.Y(n_1430)
);

BUFx12f_ASAP7_75t_L g1431 ( 
.A(n_1231),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1259),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1189),
.A2(n_1346),
.B1(n_1345),
.B2(n_1232),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1346),
.A2(n_1234),
.B1(n_1245),
.B2(n_1341),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1234),
.A2(n_1245),
.B1(n_1341),
.B2(n_1228),
.Y(n_1435)
);

OAI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1185),
.A2(n_1197),
.B1(n_1340),
.B2(n_1234),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1197),
.B(n_1196),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1294),
.A2(n_1324),
.B(n_1327),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1245),
.A2(n_1228),
.B1(n_1187),
.B2(n_1190),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1194),
.Y(n_1440)
);

AND2x4_ASAP7_75t_L g1441 ( 
.A(n_1319),
.B(n_1220),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1325),
.Y(n_1442)
);

OR2x6_ASAP7_75t_L g1443 ( 
.A(n_1185),
.B(n_1319),
.Y(n_1443)
);

INVxp67_ASAP7_75t_L g1444 ( 
.A(n_1284),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1328),
.A2(n_1335),
.B1(n_1330),
.B2(n_1343),
.Y(n_1445)
);

INVx4_ASAP7_75t_L g1446 ( 
.A(n_1298),
.Y(n_1446)
);

AND2x4_ASAP7_75t_L g1447 ( 
.A(n_1220),
.B(n_1263),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_SL g1448 ( 
.A1(n_1208),
.A2(n_1210),
.B1(n_1187),
.B2(n_1190),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1327),
.A2(n_1267),
.B(n_1213),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_SL g1450 ( 
.A1(n_1208),
.A2(n_1210),
.B1(n_1187),
.B2(n_1190),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_SL g1451 ( 
.A1(n_1315),
.A2(n_1225),
.B(n_1270),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1263),
.B(n_1187),
.Y(n_1452)
);

A2O1A1Ixp33_ASAP7_75t_L g1453 ( 
.A1(n_1203),
.A2(n_1251),
.B(n_1186),
.C(n_1286),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1188),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1188),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1338),
.A2(n_1298),
.B1(n_1270),
.B2(n_1306),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1194),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1196),
.B(n_1190),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_1190),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1198),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1196),
.B(n_1205),
.Y(n_1461)
);

INVx6_ASAP7_75t_L g1462 ( 
.A(n_1338),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1225),
.Y(n_1463)
);

CKINVDCx16_ASAP7_75t_R g1464 ( 
.A(n_1340),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1196),
.B(n_1205),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1198),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1205),
.Y(n_1467)
);

BUFx4f_ASAP7_75t_L g1468 ( 
.A(n_1225),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1337),
.A2(n_1203),
.B(n_1331),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_1344),
.Y(n_1470)
);

OR2x6_ASAP7_75t_SL g1471 ( 
.A(n_1344),
.B(n_1205),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1188),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1286),
.B(n_1188),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1271),
.Y(n_1474)
);

OAI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1186),
.A2(n_1269),
.B(n_1207),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1239),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_1271),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1306),
.Y(n_1478)
);

NAND3xp33_ASAP7_75t_L g1479 ( 
.A(n_1215),
.B(n_1270),
.C(n_1316),
.Y(n_1479)
);

CKINVDCx16_ASAP7_75t_R g1480 ( 
.A(n_1309),
.Y(n_1480)
);

INVx4_ASAP7_75t_L g1481 ( 
.A(n_1265),
.Y(n_1481)
);

AO31x2_ASAP7_75t_L g1482 ( 
.A1(n_1276),
.A2(n_1336),
.A3(n_1309),
.B(n_1334),
.Y(n_1482)
);

INVx2_ASAP7_75t_SL g1483 ( 
.A(n_1269),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1265),
.B(n_1334),
.Y(n_1484)
);

NAND2x1_ASAP7_75t_L g1485 ( 
.A(n_1265),
.B(n_1316),
.Y(n_1485)
);

AND2x4_ASAP7_75t_L g1486 ( 
.A(n_1233),
.B(n_1236),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1276),
.Y(n_1487)
);

INVx2_ASAP7_75t_SL g1488 ( 
.A(n_1233),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1334),
.B(n_1215),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1306),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1286),
.B(n_1334),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1316),
.A2(n_1215),
.B1(n_1286),
.B2(n_1336),
.Y(n_1492)
);

NAND2x1p5_ASAP7_75t_L g1493 ( 
.A(n_1279),
.B(n_1236),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1279),
.A2(n_1277),
.B1(n_1230),
.B2(n_1241),
.Y(n_1494)
);

NAND3xp33_ASAP7_75t_SL g1495 ( 
.A(n_1213),
.B(n_1260),
.C(n_1241),
.Y(n_1495)
);

AO21x2_ASAP7_75t_L g1496 ( 
.A1(n_1230),
.A2(n_1267),
.B(n_1260),
.Y(n_1496)
);

OAI222xp33_ASAP7_75t_L g1497 ( 
.A1(n_1277),
.A2(n_971),
.B1(n_625),
.B2(n_743),
.C1(n_731),
.C2(n_714),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1289),
.B(n_1209),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1209),
.B(n_919),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1379),
.B(n_1376),
.Y(n_1500)
);

OAI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1388),
.A2(n_1498),
.B1(n_1409),
.B2(n_1376),
.Y(n_1501)
);

INVx2_ASAP7_75t_SL g1502 ( 
.A(n_1386),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1383),
.B(n_1354),
.Y(n_1503)
);

BUFx12f_ASAP7_75t_L g1504 ( 
.A(n_1360),
.Y(n_1504)
);

AOI221xp5_ASAP7_75t_L g1505 ( 
.A1(n_1350),
.A2(n_1356),
.B1(n_1391),
.B2(n_1364),
.C(n_1473),
.Y(n_1505)
);

O2A1O1Ixp33_ASAP7_75t_L g1506 ( 
.A1(n_1350),
.A2(n_1398),
.B(n_1410),
.C(n_1497),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1385),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1396),
.B(n_1389),
.Y(n_1508)
);

AO21x1_ASAP7_75t_L g1509 ( 
.A1(n_1417),
.A2(n_1392),
.B(n_1456),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1364),
.A2(n_1390),
.B1(n_1402),
.B2(n_1424),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1387),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1365),
.Y(n_1512)
);

AOI21xp33_ASAP7_75t_L g1513 ( 
.A1(n_1390),
.A2(n_1377),
.B(n_1408),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1499),
.A2(n_1361),
.B1(n_1464),
.B2(n_1366),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1373),
.Y(n_1515)
);

INVx1_ASAP7_75t_SL g1516 ( 
.A(n_1386),
.Y(n_1516)
);

AOI222xp33_ASAP7_75t_L g1517 ( 
.A1(n_1491),
.A2(n_1465),
.B1(n_1429),
.B2(n_1467),
.C1(n_1436),
.C2(n_1405),
.Y(n_1517)
);

AOI21xp33_ASAP7_75t_L g1518 ( 
.A1(n_1377),
.A2(n_1437),
.B(n_1454),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1368),
.B(n_1375),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1403),
.Y(n_1520)
);

AOI221xp5_ASAP7_75t_L g1521 ( 
.A1(n_1492),
.A2(n_1410),
.B1(n_1453),
.B2(n_1479),
.C(n_1445),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_SL g1522 ( 
.A1(n_1458),
.A2(n_1461),
.B1(n_1407),
.B2(n_1393),
.Y(n_1522)
);

AOI222xp33_ASAP7_75t_L g1523 ( 
.A1(n_1436),
.A2(n_1414),
.B1(n_1413),
.B2(n_1444),
.C1(n_1415),
.C2(n_1433),
.Y(n_1523)
);

AOI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1369),
.A2(n_1469),
.B(n_1476),
.Y(n_1524)
);

INVx1_ASAP7_75t_SL g1525 ( 
.A(n_1397),
.Y(n_1525)
);

BUFx3_ASAP7_75t_L g1526 ( 
.A(n_1425),
.Y(n_1526)
);

INVx4_ASAP7_75t_SL g1527 ( 
.A(n_1393),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1421),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1428),
.B(n_1367),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_SL g1530 ( 
.A(n_1466),
.B(n_1470),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1400),
.B(n_1401),
.Y(n_1531)
);

OAI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1394),
.A2(n_1363),
.B1(n_1407),
.B2(n_1443),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1431),
.A2(n_1407),
.B1(n_1357),
.B2(n_1358),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1431),
.A2(n_1407),
.B1(n_1357),
.B2(n_1358),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1412),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1355),
.A2(n_1358),
.B1(n_1357),
.B2(n_1443),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1422),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1360),
.A2(n_1439),
.B1(n_1416),
.B2(n_1384),
.Y(n_1538)
);

AOI21xp5_ASAP7_75t_L g1539 ( 
.A1(n_1381),
.A2(n_1495),
.B(n_1468),
.Y(n_1539)
);

BUFx4f_ASAP7_75t_SL g1540 ( 
.A(n_1380),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1355),
.A2(n_1433),
.B1(n_1413),
.B2(n_1393),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1432),
.Y(n_1542)
);

INVx3_ASAP7_75t_L g1543 ( 
.A(n_1430),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1434),
.A2(n_1404),
.B1(n_1435),
.B2(n_1420),
.Y(n_1544)
);

CKINVDCx6p67_ASAP7_75t_R g1545 ( 
.A(n_1423),
.Y(n_1545)
);

AOI222xp33_ASAP7_75t_L g1546 ( 
.A1(n_1435),
.A2(n_1468),
.B1(n_1434),
.B2(n_1459),
.C1(n_1423),
.C2(n_1453),
.Y(n_1546)
);

AOI21xp33_ASAP7_75t_L g1547 ( 
.A1(n_1455),
.A2(n_1472),
.B(n_1489),
.Y(n_1547)
);

OAI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1371),
.A2(n_1426),
.B1(n_1404),
.B2(n_1359),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1349),
.Y(n_1549)
);

OAI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1371),
.A2(n_1426),
.B1(n_1359),
.B2(n_1420),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1442),
.B(n_1441),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1441),
.B(n_1470),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1441),
.B(n_1466),
.Y(n_1553)
);

AOI211xp5_ASAP7_75t_L g1554 ( 
.A1(n_1451),
.A2(n_1490),
.B(n_1478),
.C(n_1475),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1477),
.B(n_1480),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1426),
.A2(n_1452),
.B1(n_1477),
.B2(n_1447),
.Y(n_1556)
);

NAND3xp33_ASAP7_75t_L g1557 ( 
.A(n_1481),
.B(n_1406),
.C(n_1382),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1351),
.Y(n_1558)
);

OAI21xp5_ASAP7_75t_SL g1559 ( 
.A1(n_1448),
.A2(n_1450),
.B(n_1447),
.Y(n_1559)
);

OAI211xp5_ASAP7_75t_SL g1560 ( 
.A1(n_1382),
.A2(n_1494),
.B(n_1484),
.C(n_1483),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1452),
.A2(n_1447),
.B1(n_1351),
.B2(n_1353),
.Y(n_1561)
);

OAI221xp5_ASAP7_75t_L g1562 ( 
.A1(n_1481),
.A2(n_1485),
.B1(n_1462),
.B2(n_1494),
.C(n_1488),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1452),
.A2(n_1411),
.B1(n_1353),
.B2(n_1418),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1399),
.A2(n_1446),
.B1(n_1359),
.B2(n_1462),
.Y(n_1564)
);

OAI221xp5_ASAP7_75t_L g1565 ( 
.A1(n_1493),
.A2(n_1463),
.B1(n_1457),
.B2(n_1460),
.C(n_1440),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1471),
.A2(n_1463),
.B1(n_1486),
.B2(n_1378),
.Y(n_1566)
);

OAI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1463),
.A2(n_1460),
.B1(n_1457),
.B2(n_1440),
.Y(n_1567)
);

AOI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1496),
.A2(n_1449),
.B(n_1438),
.Y(n_1568)
);

OAI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1427),
.A2(n_1438),
.B(n_1449),
.Y(n_1569)
);

OAI21x1_ASAP7_75t_L g1570 ( 
.A1(n_1352),
.A2(n_1370),
.B(n_1378),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1372),
.A2(n_1419),
.B1(n_1395),
.B2(n_1411),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1395),
.A2(n_1487),
.B1(n_1474),
.B2(n_1486),
.Y(n_1572)
);

NAND4xp25_ASAP7_75t_L g1573 ( 
.A(n_1486),
.B(n_1474),
.C(n_1487),
.D(n_1352),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1378),
.A2(n_1496),
.B1(n_1370),
.B2(n_1482),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1482),
.Y(n_1575)
);

AOI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1482),
.A2(n_1206),
.B1(n_719),
.B2(n_971),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1482),
.A2(n_588),
.B1(n_622),
.B2(n_971),
.Y(n_1577)
);

INVx4_ASAP7_75t_L g1578 ( 
.A(n_1412),
.Y(n_1578)
);

BUFx12f_ASAP7_75t_L g1579 ( 
.A(n_1360),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1374),
.Y(n_1580)
);

BUFx6f_ASAP7_75t_L g1581 ( 
.A(n_1431),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1354),
.B(n_1396),
.Y(n_1582)
);

AOI222xp33_ASAP7_75t_L g1583 ( 
.A1(n_1350),
.A2(n_622),
.B1(n_815),
.B2(n_1095),
.C1(n_1226),
.C2(n_1206),
.Y(n_1583)
);

OAI21xp33_ASAP7_75t_L g1584 ( 
.A1(n_1356),
.A2(n_719),
.B(n_791),
.Y(n_1584)
);

CKINVDCx11_ASAP7_75t_R g1585 ( 
.A(n_1380),
.Y(n_1585)
);

OAI211xp5_ASAP7_75t_L g1586 ( 
.A1(n_1356),
.A2(n_1192),
.B(n_719),
.C(n_533),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1354),
.B(n_1396),
.Y(n_1587)
);

INVx3_ASAP7_75t_L g1588 ( 
.A(n_1425),
.Y(n_1588)
);

OAI221xp5_ASAP7_75t_L g1589 ( 
.A1(n_1350),
.A2(n_1192),
.B1(n_719),
.B2(n_770),
.C(n_533),
.Y(n_1589)
);

CKINVDCx20_ASAP7_75t_R g1590 ( 
.A(n_1386),
.Y(n_1590)
);

AOI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1350),
.A2(n_1206),
.B1(n_719),
.B2(n_971),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1379),
.B(n_1376),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_SL g1593 ( 
.A1(n_1464),
.A2(n_1162),
.B1(n_1204),
.B2(n_1206),
.Y(n_1593)
);

NAND2x1p5_ASAP7_75t_L g1594 ( 
.A(n_1362),
.B(n_1094),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1374),
.Y(n_1595)
);

CKINVDCx20_ASAP7_75t_R g1596 ( 
.A(n_1386),
.Y(n_1596)
);

AOI21xp5_ASAP7_75t_L g1597 ( 
.A1(n_1369),
.A2(n_1206),
.B(n_1058),
.Y(n_1597)
);

NAND4xp25_ASAP7_75t_L g1598 ( 
.A(n_1356),
.B(n_533),
.C(n_377),
.D(n_388),
.Y(n_1598)
);

OAI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1350),
.A2(n_1242),
.B1(n_1201),
.B2(n_1192),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1350),
.A2(n_1242),
.B1(n_1201),
.B2(n_1192),
.Y(n_1600)
);

INVx6_ASAP7_75t_L g1601 ( 
.A(n_1431),
.Y(n_1601)
);

NAND3xp33_ASAP7_75t_L g1602 ( 
.A(n_1356),
.B(n_1192),
.C(n_533),
.Y(n_1602)
);

AOI21x1_ASAP7_75t_L g1603 ( 
.A1(n_1369),
.A2(n_1206),
.B(n_1469),
.Y(n_1603)
);

OAI221xp5_ASAP7_75t_L g1604 ( 
.A1(n_1350),
.A2(n_1192),
.B1(n_719),
.B2(n_770),
.C(n_533),
.Y(n_1604)
);

BUFx5_ASAP7_75t_L g1605 ( 
.A(n_1486),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_L g1606 ( 
.A1(n_1350),
.A2(n_588),
.B1(n_622),
.B2(n_971),
.Y(n_1606)
);

AOI221xp5_ASAP7_75t_L g1607 ( 
.A1(n_1350),
.A2(n_533),
.B1(n_534),
.B2(n_1162),
.C(n_719),
.Y(n_1607)
);

OAI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1379),
.A2(n_1204),
.B1(n_971),
.B2(n_1206),
.Y(n_1608)
);

OA21x2_ASAP7_75t_L g1609 ( 
.A1(n_1570),
.A2(n_1568),
.B(n_1597),
.Y(n_1609)
);

INVxp67_ASAP7_75t_L g1610 ( 
.A(n_1573),
.Y(n_1610)
);

INVxp67_ASAP7_75t_L g1611 ( 
.A(n_1535),
.Y(n_1611)
);

AOI221xp5_ASAP7_75t_L g1612 ( 
.A1(n_1607),
.A2(n_1604),
.B1(n_1589),
.B2(n_1598),
.C(n_1501),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1549),
.Y(n_1613)
);

INVxp67_ASAP7_75t_L g1614 ( 
.A(n_1500),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1605),
.B(n_1582),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1558),
.Y(n_1616)
);

INVx3_ASAP7_75t_L g1617 ( 
.A(n_1605),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1605),
.B(n_1587),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1520),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1605),
.B(n_1507),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1503),
.B(n_1508),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1528),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1555),
.B(n_1592),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1605),
.B(n_1511),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1537),
.Y(n_1625)
);

INVx2_ASAP7_75t_SL g1626 ( 
.A(n_1526),
.Y(n_1626)
);

INVx1_ASAP7_75t_SL g1627 ( 
.A(n_1526),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1566),
.B(n_1574),
.Y(n_1628)
);

INVx3_ASAP7_75t_L g1629 ( 
.A(n_1569),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1524),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1608),
.B(n_1576),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1583),
.A2(n_1606),
.B1(n_1593),
.B2(n_1577),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1542),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1521),
.B(n_1554),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1512),
.B(n_1515),
.Y(n_1635)
);

AO31x2_ASAP7_75t_L g1636 ( 
.A1(n_1509),
.A2(n_1575),
.A3(n_1539),
.B(n_1600),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1527),
.B(n_1543),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1580),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1595),
.B(n_1603),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1572),
.B(n_1519),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1527),
.B(n_1543),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1572),
.B(n_1531),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1561),
.B(n_1563),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1514),
.B(n_1530),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1514),
.B(n_1530),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1552),
.B(n_1553),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1557),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1562),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1608),
.B(n_1501),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1565),
.Y(n_1650)
);

OA21x2_ASAP7_75t_L g1651 ( 
.A1(n_1518),
.A2(n_1505),
.B(n_1513),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1563),
.Y(n_1652)
);

INVxp67_ASAP7_75t_L g1653 ( 
.A(n_1588),
.Y(n_1653)
);

AO21x2_ASAP7_75t_L g1654 ( 
.A1(n_1567),
.A2(n_1547),
.B(n_1560),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1561),
.B(n_1551),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1571),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1522),
.B(n_1541),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1571),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1578),
.B(n_1591),
.Y(n_1659)
);

INVx4_ASAP7_75t_L g1660 ( 
.A(n_1601),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1522),
.B(n_1541),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1517),
.B(n_1556),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1567),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1606),
.A2(n_1599),
.B1(n_1602),
.B2(n_1593),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1556),
.B(n_1559),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1546),
.B(n_1523),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1532),
.B(n_1510),
.Y(n_1667)
);

NOR2x1_ASAP7_75t_SL g1668 ( 
.A(n_1564),
.B(n_1538),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1529),
.B(n_1544),
.Y(n_1669)
);

NOR2x1_ASAP7_75t_SL g1670 ( 
.A(n_1581),
.B(n_1586),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1536),
.B(n_1581),
.Y(n_1671)
);

A2O1A1Ixp33_ASAP7_75t_L g1672 ( 
.A1(n_1612),
.A2(n_1584),
.B(n_1506),
.C(n_1577),
.Y(n_1672)
);

OAI222xp33_ASAP7_75t_L g1673 ( 
.A1(n_1664),
.A2(n_1550),
.B1(n_1525),
.B2(n_1548),
.C1(n_1536),
.C2(n_1533),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1615),
.B(n_1502),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1615),
.B(n_1618),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1618),
.B(n_1516),
.Y(n_1676)
);

AOI211xp5_ASAP7_75t_L g1677 ( 
.A1(n_1612),
.A2(n_1560),
.B(n_1550),
.C(n_1548),
.Y(n_1677)
);

AOI221xp5_ASAP7_75t_L g1678 ( 
.A1(n_1664),
.A2(n_1581),
.B1(n_1596),
.B2(n_1590),
.C(n_1533),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1613),
.Y(n_1679)
);

AOI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1632),
.A2(n_1601),
.B1(n_1594),
.B2(n_1534),
.Y(n_1680)
);

AO21x2_ASAP7_75t_L g1681 ( 
.A1(n_1630),
.A2(n_1534),
.B(n_1601),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1614),
.B(n_1545),
.Y(n_1682)
);

OAI332xp33_ASAP7_75t_L g1683 ( 
.A1(n_1649),
.A2(n_1540),
.A3(n_1585),
.B1(n_1590),
.B2(n_1596),
.B3(n_1504),
.C1(n_1579),
.C2(n_1581),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_R g1684 ( 
.A(n_1634),
.B(n_1585),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1622),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1622),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1649),
.A2(n_1540),
.B1(n_1631),
.B2(n_1634),
.Y(n_1687)
);

OAI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1631),
.A2(n_1667),
.B1(n_1666),
.B2(n_1634),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1628),
.B(n_1620),
.Y(n_1689)
);

NAND3xp33_ASAP7_75t_L g1690 ( 
.A(n_1614),
.B(n_1610),
.C(n_1648),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1628),
.B(n_1620),
.Y(n_1691)
);

OAI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1667),
.A2(n_1666),
.B1(n_1644),
.B2(n_1645),
.Y(n_1692)
);

AOI221xp5_ASAP7_75t_L g1693 ( 
.A1(n_1662),
.A2(n_1610),
.B1(n_1665),
.B2(n_1648),
.C(n_1661),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1625),
.Y(n_1694)
);

INVxp67_ASAP7_75t_L g1695 ( 
.A(n_1647),
.Y(n_1695)
);

AO21x2_ASAP7_75t_L g1696 ( 
.A1(n_1630),
.A2(n_1654),
.B(n_1663),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1613),
.Y(n_1697)
);

AOI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1609),
.A2(n_1668),
.B(n_1654),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1623),
.B(n_1621),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1639),
.B(n_1647),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1623),
.B(n_1621),
.Y(n_1701)
);

OAI221xp5_ASAP7_75t_L g1702 ( 
.A1(n_1644),
.A2(n_1645),
.B1(n_1662),
.B2(n_1665),
.C(n_1651),
.Y(n_1702)
);

AND2x4_ASAP7_75t_SL g1703 ( 
.A(n_1637),
.B(n_1641),
.Y(n_1703)
);

INVx4_ASAP7_75t_L g1704 ( 
.A(n_1660),
.Y(n_1704)
);

AOI22xp33_ASAP7_75t_L g1705 ( 
.A1(n_1662),
.A2(n_1665),
.B1(n_1657),
.B2(n_1661),
.Y(n_1705)
);

AOI31xp33_ASAP7_75t_L g1706 ( 
.A1(n_1628),
.A2(n_1661),
.A3(n_1657),
.B(n_1659),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1640),
.B(n_1655),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1657),
.A2(n_1651),
.B1(n_1652),
.B2(n_1643),
.Y(n_1708)
);

OA21x2_ASAP7_75t_L g1709 ( 
.A1(n_1663),
.A2(n_1650),
.B(n_1639),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1639),
.B(n_1636),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1616),
.Y(n_1711)
);

OA21x2_ASAP7_75t_L g1712 ( 
.A1(n_1650),
.A2(n_1652),
.B(n_1658),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1624),
.B(n_1640),
.Y(n_1713)
);

INVxp67_ASAP7_75t_SL g1714 ( 
.A(n_1629),
.Y(n_1714)
);

OAI33xp33_ASAP7_75t_L g1715 ( 
.A1(n_1635),
.A2(n_1659),
.A3(n_1638),
.B1(n_1619),
.B2(n_1611),
.B3(n_1625),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1636),
.B(n_1638),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1624),
.B(n_1640),
.Y(n_1717)
);

INVxp67_ASAP7_75t_SL g1718 ( 
.A(n_1629),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1700),
.B(n_1636),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1695),
.B(n_1636),
.Y(n_1720)
);

BUFx2_ASAP7_75t_L g1721 ( 
.A(n_1714),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1713),
.B(n_1717),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1679),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1703),
.B(n_1617),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1695),
.B(n_1636),
.Y(n_1725)
);

INVx6_ASAP7_75t_L g1726 ( 
.A(n_1704),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_SL g1727 ( 
.A(n_1706),
.B(n_1626),
.Y(n_1727)
);

INVx6_ASAP7_75t_L g1728 ( 
.A(n_1704),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1700),
.B(n_1636),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1709),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1709),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1709),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1716),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1713),
.B(n_1609),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1713),
.B(n_1609),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1716),
.B(n_1636),
.Y(n_1736)
);

HB1xp67_ASAP7_75t_L g1737 ( 
.A(n_1710),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1703),
.B(n_1617),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1709),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1709),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1710),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1717),
.B(n_1609),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1706),
.B(n_1619),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1717),
.B(n_1609),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1707),
.B(n_1635),
.Y(n_1745)
);

NAND3xp33_ASAP7_75t_SL g1746 ( 
.A(n_1693),
.B(n_1627),
.C(n_1669),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_SL g1747 ( 
.A(n_1698),
.B(n_1690),
.Y(n_1747)
);

INVx3_ASAP7_75t_L g1748 ( 
.A(n_1703),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1689),
.B(n_1617),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1689),
.B(n_1617),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1689),
.B(n_1629),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1697),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1699),
.B(n_1633),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1697),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1711),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1711),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1707),
.B(n_1699),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1757),
.B(n_1701),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1757),
.B(n_1701),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1745),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1743),
.B(n_1690),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1722),
.B(n_1691),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_L g1763 ( 
.A(n_1743),
.B(n_1683),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1757),
.B(n_1745),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1722),
.B(n_1691),
.Y(n_1765)
);

OR2x6_ASAP7_75t_L g1766 ( 
.A(n_1747),
.B(n_1698),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1722),
.B(n_1691),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1745),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1753),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1753),
.B(n_1693),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1719),
.B(n_1702),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1736),
.B(n_1720),
.Y(n_1772)
);

AND3x2_ASAP7_75t_L g1773 ( 
.A(n_1737),
.B(n_1677),
.C(n_1678),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1722),
.B(n_1727),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1727),
.B(n_1675),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1736),
.B(n_1687),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1723),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1720),
.B(n_1687),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1737),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1723),
.Y(n_1780)
);

INVx3_ASAP7_75t_L g1781 ( 
.A(n_1748),
.Y(n_1781)
);

AOI211xp5_ASAP7_75t_SL g1782 ( 
.A1(n_1746),
.A2(n_1683),
.B(n_1702),
.C(n_1677),
.Y(n_1782)
);

AOI21xp5_ASAP7_75t_L g1783 ( 
.A1(n_1746),
.A2(n_1715),
.B(n_1668),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1719),
.B(n_1685),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1748),
.B(n_1675),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1719),
.B(n_1685),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1729),
.B(n_1686),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1725),
.B(n_1708),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1730),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1723),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1725),
.B(n_1686),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1748),
.B(n_1676),
.Y(n_1792)
);

INVx1_ASAP7_75t_SL g1793 ( 
.A(n_1747),
.Y(n_1793)
);

INVxp67_ASAP7_75t_L g1794 ( 
.A(n_1729),
.Y(n_1794)
);

AND2x4_ASAP7_75t_L g1795 ( 
.A(n_1748),
.B(n_1714),
.Y(n_1795)
);

CKINVDCx16_ASAP7_75t_R g1796 ( 
.A(n_1724),
.Y(n_1796)
);

AND2x4_ASAP7_75t_L g1797 ( 
.A(n_1762),
.B(n_1748),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1758),
.B(n_1729),
.Y(n_1798)
);

INVx1_ASAP7_75t_SL g1799 ( 
.A(n_1771),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1796),
.B(n_1762),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1758),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1782),
.B(n_1770),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1796),
.B(n_1748),
.Y(n_1803)
);

OAI211xp5_ASAP7_75t_L g1804 ( 
.A1(n_1793),
.A2(n_1684),
.B(n_1721),
.C(n_1705),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1759),
.Y(n_1805)
);

NAND5xp2_ASAP7_75t_L g1806 ( 
.A(n_1763),
.B(n_1678),
.C(n_1735),
.D(n_1734),
.E(n_1742),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1765),
.B(n_1751),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1793),
.B(n_1741),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1759),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1764),
.Y(n_1810)
);

NAND4xp25_ASAP7_75t_L g1811 ( 
.A(n_1783),
.B(n_1672),
.C(n_1721),
.D(n_1742),
.Y(n_1811)
);

AND2x4_ASAP7_75t_SL g1812 ( 
.A(n_1792),
.B(n_1724),
.Y(n_1812)
);

NAND2xp33_ASAP7_75t_R g1813 ( 
.A(n_1773),
.B(n_1651),
.Y(n_1813)
);

INVxp67_ASAP7_75t_L g1814 ( 
.A(n_1761),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1764),
.B(n_1760),
.Y(n_1815)
);

AOI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1788),
.A2(n_1715),
.B(n_1688),
.Y(n_1816)
);

OR2x6_ASAP7_75t_L g1817 ( 
.A(n_1766),
.B(n_1730),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1760),
.Y(n_1818)
);

INVxp67_ASAP7_75t_L g1819 ( 
.A(n_1771),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1768),
.B(n_1741),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1768),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1784),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1776),
.B(n_1733),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1784),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1765),
.B(n_1751),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1786),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1769),
.B(n_1778),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1786),
.Y(n_1828)
);

NOR2xp33_ASAP7_75t_L g1829 ( 
.A(n_1766),
.B(n_1682),
.Y(n_1829)
);

NOR2xp33_ASAP7_75t_SL g1830 ( 
.A(n_1774),
.B(n_1673),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1769),
.B(n_1733),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1779),
.B(n_1734),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1787),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1787),
.Y(n_1834)
);

NOR2xp33_ASAP7_75t_L g1835 ( 
.A(n_1766),
.B(n_1682),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1777),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1772),
.B(n_1611),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1789),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1789),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1810),
.Y(n_1840)
);

OAI22xp33_ASAP7_75t_L g1841 ( 
.A1(n_1830),
.A2(n_1766),
.B1(n_1692),
.B2(n_1740),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1801),
.Y(n_1842)
);

AOI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1802),
.A2(n_1766),
.B(n_1794),
.Y(n_1843)
);

OAI32xp33_ASAP7_75t_L g1844 ( 
.A1(n_1813),
.A2(n_1774),
.A3(n_1732),
.B1(n_1731),
.B2(n_1740),
.Y(n_1844)
);

AOI31xp33_ASAP7_75t_L g1845 ( 
.A1(n_1814),
.A2(n_1775),
.A3(n_1795),
.B(n_1785),
.Y(n_1845)
);

INVx1_ASAP7_75t_SL g1846 ( 
.A(n_1799),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1805),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1816),
.B(n_1767),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_SL g1849 ( 
.A1(n_1804),
.A2(n_1730),
.B1(n_1731),
.B2(n_1732),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1800),
.B(n_1767),
.Y(n_1850)
);

OAI21xp33_ASAP7_75t_L g1851 ( 
.A1(n_1806),
.A2(n_1791),
.B(n_1775),
.Y(n_1851)
);

OAI221xp5_ASAP7_75t_L g1852 ( 
.A1(n_1813),
.A2(n_1740),
.B1(n_1739),
.B2(n_1732),
.C(n_1731),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1809),
.Y(n_1853)
);

OR2x2_ASAP7_75t_L g1854 ( 
.A(n_1827),
.B(n_1777),
.Y(n_1854)
);

OAI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1811),
.A2(n_1732),
.B1(n_1730),
.B2(n_1739),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_L g1856 ( 
.A(n_1819),
.B(n_1781),
.Y(n_1856)
);

OAI31xp33_ASAP7_75t_L g1857 ( 
.A1(n_1829),
.A2(n_1731),
.A3(n_1739),
.B(n_1740),
.Y(n_1857)
);

INVx1_ASAP7_75t_SL g1858 ( 
.A(n_1803),
.Y(n_1858)
);

OAI21xp5_ASAP7_75t_L g1859 ( 
.A1(n_1829),
.A2(n_1835),
.B(n_1817),
.Y(n_1859)
);

NOR2xp33_ASAP7_75t_L g1860 ( 
.A(n_1835),
.B(n_1781),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1823),
.B(n_1734),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1815),
.B(n_1780),
.Y(n_1862)
);

OAI321xp33_ASAP7_75t_L g1863 ( 
.A1(n_1817),
.A2(n_1808),
.A3(n_1832),
.B1(n_1798),
.B2(n_1800),
.C(n_1739),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1837),
.B(n_1734),
.Y(n_1864)
);

OAI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1817),
.A2(n_1721),
.B(n_1744),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1817),
.Y(n_1866)
);

AOI322xp5_ASAP7_75t_L g1867 ( 
.A1(n_1838),
.A2(n_1735),
.A3(n_1744),
.B1(n_1742),
.B2(n_1839),
.C1(n_1828),
.C2(n_1826),
.Y(n_1867)
);

OAI21xp5_ASAP7_75t_L g1868 ( 
.A1(n_1803),
.A2(n_1744),
.B(n_1742),
.Y(n_1868)
);

OAI21xp33_ASAP7_75t_L g1869 ( 
.A1(n_1822),
.A2(n_1744),
.B(n_1735),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1818),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1812),
.B(n_1797),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_1812),
.B(n_1781),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1797),
.B(n_1785),
.Y(n_1873)
);

AOI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1821),
.A2(n_1696),
.B1(n_1651),
.B2(n_1712),
.Y(n_1874)
);

OAI22xp33_ASAP7_75t_L g1875 ( 
.A1(n_1820),
.A2(n_1669),
.B1(n_1651),
.B2(n_1680),
.Y(n_1875)
);

OAI21xp33_ASAP7_75t_SL g1876 ( 
.A1(n_1845),
.A2(n_1807),
.B(n_1825),
.Y(n_1876)
);

AOI322xp5_ASAP7_75t_L g1877 ( 
.A1(n_1848),
.A2(n_1735),
.A3(n_1839),
.B1(n_1838),
.B2(n_1834),
.C1(n_1833),
.C2(n_1824),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1870),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1850),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1850),
.B(n_1871),
.Y(n_1880)
);

NOR3xp33_ASAP7_75t_L g1881 ( 
.A(n_1863),
.B(n_1831),
.C(n_1673),
.Y(n_1881)
);

AOI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1875),
.A2(n_1841),
.B1(n_1855),
.B2(n_1851),
.Y(n_1882)
);

NOR2x1_ASAP7_75t_L g1883 ( 
.A(n_1846),
.B(n_1797),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1840),
.Y(n_1884)
);

AOI21xp33_ASAP7_75t_SL g1885 ( 
.A1(n_1859),
.A2(n_1795),
.B(n_1831),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1871),
.B(n_1807),
.Y(n_1886)
);

AOI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1849),
.A2(n_1696),
.B1(n_1712),
.B2(n_1680),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1858),
.B(n_1825),
.Y(n_1888)
);

NOR3xp33_ASAP7_75t_L g1889 ( 
.A(n_1844),
.B(n_1836),
.C(n_1718),
.Y(n_1889)
);

INVx1_ASAP7_75t_SL g1890 ( 
.A(n_1866),
.Y(n_1890)
);

AOI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1874),
.A2(n_1696),
.B1(n_1712),
.B2(n_1681),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1873),
.B(n_1792),
.Y(n_1892)
);

INVxp67_ASAP7_75t_L g1893 ( 
.A(n_1856),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1842),
.Y(n_1894)
);

AOI222xp33_ASAP7_75t_L g1895 ( 
.A1(n_1852),
.A2(n_1643),
.B1(n_1656),
.B2(n_1658),
.C1(n_1642),
.C2(n_1650),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_L g1896 ( 
.A(n_1847),
.B(n_1795),
.Y(n_1896)
);

XNOR2xp5_ASAP7_75t_L g1897 ( 
.A(n_1843),
.B(n_1671),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1873),
.A2(n_1795),
.B1(n_1728),
.B2(n_1726),
.Y(n_1898)
);

OAI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1865),
.A2(n_1728),
.B1(n_1726),
.B2(n_1751),
.Y(n_1899)
);

AOI22xp5_ASAP7_75t_SL g1900 ( 
.A1(n_1856),
.A2(n_1660),
.B1(n_1751),
.B2(n_1627),
.Y(n_1900)
);

AO22x1_ASAP7_75t_L g1901 ( 
.A1(n_1866),
.A2(n_1738),
.B1(n_1724),
.B2(n_1660),
.Y(n_1901)
);

NOR4xp25_ASAP7_75t_SL g1902 ( 
.A(n_1885),
.B(n_1853),
.C(n_1869),
.D(n_1867),
.Y(n_1902)
);

INVx1_ASAP7_75t_SL g1903 ( 
.A(n_1883),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1879),
.Y(n_1904)
);

AOI222xp33_ASAP7_75t_L g1905 ( 
.A1(n_1890),
.A2(n_1868),
.B1(n_1861),
.B2(n_1860),
.C1(n_1857),
.C2(n_1864),
.Y(n_1905)
);

NOR3xp33_ASAP7_75t_SL g1906 ( 
.A(n_1876),
.B(n_1860),
.C(n_1872),
.Y(n_1906)
);

NOR2x1_ASAP7_75t_L g1907 ( 
.A(n_1884),
.B(n_1872),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1879),
.Y(n_1908)
);

OAI21xp33_ASAP7_75t_L g1909 ( 
.A1(n_1882),
.A2(n_1854),
.B(n_1862),
.Y(n_1909)
);

INVx1_ASAP7_75t_SL g1910 ( 
.A(n_1880),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1888),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1886),
.B(n_1862),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1878),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1894),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1893),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1893),
.Y(n_1916)
);

OR2x2_ASAP7_75t_L g1917 ( 
.A(n_1881),
.B(n_1780),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1896),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1892),
.B(n_1896),
.Y(n_1919)
);

NAND2xp33_ASAP7_75t_SL g1920 ( 
.A(n_1898),
.B(n_1749),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1881),
.B(n_1790),
.Y(n_1921)
);

NOR2x1_ASAP7_75t_L g1922 ( 
.A(n_1899),
.B(n_1897),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1912),
.Y(n_1923)
);

OAI21xp33_ASAP7_75t_SL g1924 ( 
.A1(n_1905),
.A2(n_1877),
.B(n_1887),
.Y(n_1924)
);

INVx1_ASAP7_75t_SL g1925 ( 
.A(n_1910),
.Y(n_1925)
);

AOI211xp5_ASAP7_75t_L g1926 ( 
.A1(n_1909),
.A2(n_1889),
.B(n_1901),
.C(n_1891),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1912),
.Y(n_1927)
);

OAI21xp5_ASAP7_75t_L g1928 ( 
.A1(n_1906),
.A2(n_1889),
.B(n_1900),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1908),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_SL g1930 ( 
.A(n_1903),
.B(n_1660),
.Y(n_1930)
);

NOR2xp33_ASAP7_75t_L g1931 ( 
.A(n_1911),
.B(n_1726),
.Y(n_1931)
);

NOR2xp33_ASAP7_75t_L g1932 ( 
.A(n_1911),
.B(n_1790),
.Y(n_1932)
);

AOI22xp5_ASAP7_75t_L g1933 ( 
.A1(n_1921),
.A2(n_1895),
.B1(n_1696),
.B2(n_1712),
.Y(n_1933)
);

OAI22xp5_ASAP7_75t_L g1934 ( 
.A1(n_1902),
.A2(n_1728),
.B1(n_1726),
.B2(n_1738),
.Y(n_1934)
);

NOR4xp25_ASAP7_75t_L g1935 ( 
.A(n_1925),
.B(n_1915),
.C(n_1916),
.D(n_1908),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1923),
.Y(n_1936)
);

BUFx3_ASAP7_75t_L g1937 ( 
.A(n_1927),
.Y(n_1937)
);

AOI22xp5_ASAP7_75t_L g1938 ( 
.A1(n_1924),
.A2(n_1917),
.B1(n_1922),
.B2(n_1918),
.Y(n_1938)
);

AOI221xp5_ASAP7_75t_SL g1939 ( 
.A1(n_1928),
.A2(n_1918),
.B1(n_1904),
.B2(n_1914),
.C(n_1913),
.Y(n_1939)
);

AOI221xp5_ASAP7_75t_L g1940 ( 
.A1(n_1926),
.A2(n_1917),
.B1(n_1919),
.B2(n_1920),
.C(n_1907),
.Y(n_1940)
);

OAI21xp5_ASAP7_75t_L g1941 ( 
.A1(n_1929),
.A2(n_1919),
.B(n_1920),
.Y(n_1941)
);

INVx1_ASAP7_75t_SL g1942 ( 
.A(n_1930),
.Y(n_1942)
);

AOI311xp33_ASAP7_75t_L g1943 ( 
.A1(n_1934),
.A2(n_1718),
.A3(n_1694),
.B(n_1653),
.C(n_1728),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1932),
.B(n_1749),
.Y(n_1944)
);

AOI221xp5_ASAP7_75t_L g1945 ( 
.A1(n_1935),
.A2(n_1932),
.B1(n_1933),
.B2(n_1931),
.C(n_1654),
.Y(n_1945)
);

AO22x2_ASAP7_75t_L g1946 ( 
.A1(n_1936),
.A2(n_1754),
.B1(n_1755),
.B2(n_1756),
.Y(n_1946)
);

AOI21xp5_ASAP7_75t_L g1947 ( 
.A1(n_1938),
.A2(n_1670),
.B(n_1750),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1937),
.B(n_1750),
.Y(n_1948)
);

NAND3xp33_ASAP7_75t_SL g1949 ( 
.A(n_1940),
.B(n_1670),
.C(n_1676),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1942),
.B(n_1749),
.Y(n_1950)
);

NOR3xp33_ASAP7_75t_L g1951 ( 
.A(n_1949),
.B(n_1939),
.C(n_1945),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1950),
.B(n_1941),
.Y(n_1952)
);

NOR2xp33_ASAP7_75t_L g1953 ( 
.A(n_1948),
.B(n_1941),
.Y(n_1953)
);

AND3x2_ASAP7_75t_L g1954 ( 
.A(n_1947),
.B(n_1944),
.C(n_1943),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1946),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1946),
.B(n_1749),
.Y(n_1956)
);

NAND4xp25_ASAP7_75t_L g1957 ( 
.A(n_1953),
.B(n_1704),
.C(n_1724),
.D(n_1738),
.Y(n_1957)
);

XOR2x1_ASAP7_75t_L g1958 ( 
.A(n_1952),
.B(n_1955),
.Y(n_1958)
);

OR3x1_ASAP7_75t_L g1959 ( 
.A(n_1954),
.B(n_1728),
.C(n_1726),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1956),
.Y(n_1960)
);

AND4x1_ASAP7_75t_L g1961 ( 
.A(n_1951),
.B(n_1750),
.C(n_1676),
.D(n_1674),
.Y(n_1961)
);

XNOR2x1_ASAP7_75t_L g1962 ( 
.A(n_1958),
.B(n_1960),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1961),
.Y(n_1963)
);

XNOR2xp5_ASAP7_75t_L g1964 ( 
.A(n_1959),
.B(n_1671),
.Y(n_1964)
);

AO21x2_ASAP7_75t_L g1965 ( 
.A1(n_1962),
.A2(n_1957),
.B(n_1750),
.Y(n_1965)
);

OAI21xp5_ASAP7_75t_L g1966 ( 
.A1(n_1965),
.A2(n_1963),
.B(n_1964),
.Y(n_1966)
);

INVxp67_ASAP7_75t_L g1967 ( 
.A(n_1966),
.Y(n_1967)
);

BUFx6f_ASAP7_75t_L g1968 ( 
.A(n_1966),
.Y(n_1968)
);

AOI22xp33_ASAP7_75t_L g1969 ( 
.A1(n_1968),
.A2(n_1965),
.B1(n_1712),
.B2(n_1681),
.Y(n_1969)
);

OAI21xp5_ASAP7_75t_L g1970 ( 
.A1(n_1967),
.A2(n_1754),
.B(n_1755),
.Y(n_1970)
);

OA21x2_ASAP7_75t_L g1971 ( 
.A1(n_1969),
.A2(n_1968),
.B(n_1674),
.Y(n_1971)
);

AOI221xp5_ASAP7_75t_L g1972 ( 
.A1(n_1970),
.A2(n_1754),
.B1(n_1755),
.B2(n_1756),
.C(n_1752),
.Y(n_1972)
);

NOR3xp33_ASAP7_75t_SL g1973 ( 
.A(n_1971),
.B(n_1694),
.C(n_1752),
.Y(n_1973)
);

OAI221xp5_ASAP7_75t_L g1974 ( 
.A1(n_1973),
.A2(n_1972),
.B1(n_1726),
.B2(n_1728),
.C(n_1626),
.Y(n_1974)
);

AOI211xp5_ASAP7_75t_L g1975 ( 
.A1(n_1974),
.A2(n_1626),
.B(n_1646),
.C(n_1756),
.Y(n_1975)
);


endmodule