module fake_jpeg_8539_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx3_ASAP7_75t_SL g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

HB1xp67_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_28),
.A2(n_24),
.B1(n_30),
.B2(n_25),
.Y(n_48)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_30),
.Y(n_36)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_23),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_32),
.B(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_3),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_5),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_35),
.B(n_37),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_24),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_16),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_45),
.Y(n_54)
);

CKINVDCx6p67_ASAP7_75t_R g43 ( 
.A(n_26),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_19),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_20),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_28),
.C(n_21),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_48),
.A2(n_28),
.B1(n_31),
.B2(n_27),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_49),
.B(n_45),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_55),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_30),
.B1(n_25),
.B2(n_22),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_31),
.B1(n_44),
.B2(n_27),
.Y(n_69)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_35),
.B(n_30),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_60),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_31),
.B1(n_27),
.B2(n_29),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_42),
.B1(n_43),
.B2(n_29),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_59),
.A2(n_44),
.B1(n_31),
.B2(n_43),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_40),
.C(n_36),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_67),
.B1(n_50),
.B2(n_42),
.Y(n_83)
);

AO22x1_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_42),
.B1(n_27),
.B2(n_29),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_51),
.B(n_39),
.Y(n_81)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_68),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_57),
.B1(n_61),
.B2(n_62),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_68),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_70),
.B(n_77),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_62),
.A2(n_36),
.B(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_71),
.B(n_75),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_50),
.B1(n_55),
.B2(n_53),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_37),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_37),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_47),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_60),
.C(n_56),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_82),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_85),
.B(n_87),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_46),
.C(n_49),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_73),
.B1(n_78),
.B2(n_63),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_64),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_67),
.A2(n_47),
.B(n_18),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_17),
.B(n_20),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_88),
.A2(n_89),
.B1(n_55),
.B2(n_65),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_76),
.B(n_66),
.Y(n_89)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

NOR3xp33_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_71),
.C(n_63),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_93),
.Y(n_107)
);

OAI32xp33_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_84),
.A3(n_80),
.B1(n_82),
.B2(n_26),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_95),
.A2(n_98),
.B(n_74),
.C(n_15),
.Y(n_108)
);

A2O1A1O1Ixp25_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_65),
.B(n_26),
.C(n_17),
.D(n_13),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_17),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_81),
.A2(n_74),
.B1(n_26),
.B2(n_15),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_87),
.B(n_90),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_99),
.B1(n_94),
.B2(n_92),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_104),
.A2(n_108),
.B1(n_97),
.B2(n_7),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_105),
.B(n_110),
.Y(n_117)
);

INVxp33_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_74),
.C(n_13),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_111),
.C(n_92),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

XNOR2x1_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_5),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_112),
.A2(n_113),
.B(n_105),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_102),
.A2(n_110),
.B1(n_106),
.B2(n_111),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_115),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_10),
.C(n_11),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_6),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_108),
.A2(n_10),
.B1(n_11),
.B2(n_8),
.Y(n_119)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_121),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_118),
.B(n_116),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_125),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_117),
.B(n_107),
.Y(n_125)
);

BUFx24_ASAP7_75t_SL g127 ( 
.A(n_122),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_129),
.Y(n_133)
);

NOR3xp33_ASAP7_75t_SL g129 ( 
.A(n_124),
.B(n_114),
.C(n_113),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_6),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_7),
.C(n_8),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_132),
.C(n_9),
.Y(n_135)
);

XOR2x2_ASAP7_75t_SL g132 ( 
.A(n_126),
.B(n_9),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_133),
.A2(n_128),
.B(n_9),
.Y(n_134)
);

BUFx24_ASAP7_75t_SL g136 ( 
.A(n_134),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_135),
.Y(n_137)
);


endmodule