module real_jpeg_13369_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_300, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_300;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_288;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_249;
wire n_286;
wire n_292;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_197;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_216;
wire n_295;
wire n_244;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_213;
wire n_202;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

BUFx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_3),
.A2(n_35),
.B1(n_61),
.B2(n_63),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_5),
.A2(n_39),
.B1(n_40),
.B2(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_5),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_105),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_5),
.A2(n_61),
.B1(n_63),
.B2(n_105),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_105),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_6),
.A2(n_61),
.B1(n_63),
.B2(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_6),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_6),
.B(n_29),
.C(n_66),
.Y(n_144)
);

NAND2x1_ASAP7_75t_SL g148 ( 
.A(n_6),
.B(n_84),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_6),
.A2(n_96),
.B(n_156),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_6),
.A2(n_44),
.B(n_83),
.C(n_183),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_6),
.A2(n_44),
.B1(n_45),
.B2(n_140),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_6),
.B(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_6),
.B(n_39),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_7),
.A2(n_61),
.B1(n_63),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_7),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_71),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_7),
.A2(n_44),
.B1(n_45),
.B2(n_71),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_9),
.A2(n_44),
.B1(n_45),
.B2(n_86),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_9),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_9),
.A2(n_61),
.B1(n_63),
.B2(n_86),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_9),
.A2(n_39),
.B1(n_40),
.B2(n_86),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_86),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_10),
.A2(n_61),
.B1(n_63),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_10),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_152),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_152),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_10),
.A2(n_39),
.B1(n_40),
.B2(n_152),
.Y(n_255)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_11),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_12),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_12),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_41),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_12),
.A2(n_41),
.B1(n_61),
.B2(n_63),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_14),
.A2(n_39),
.B1(n_40),
.B2(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_14),
.A2(n_54),
.B1(n_61),
.B2(n_63),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_54),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_54),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_15),
.A2(n_60),
.B1(n_61),
.B2(n_63),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_15),
.A2(n_44),
.B1(n_45),
.B2(n_60),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_60),
.Y(n_245)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_127),
.B1(n_297),
.B2(n_298),
.Y(n_18)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_19),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_125),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_108),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_21),
.B(n_108),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_74),
.C(n_90),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_22),
.A2(n_23),
.B1(n_74),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_56),
.B2(n_73),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_36),
.B1(n_37),
.B2(n_55),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_26),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_26),
.A2(n_37),
.B(n_73),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_26),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_32),
.B(n_33),
.Y(n_26)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_27),
.A2(n_32),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_27),
.B(n_157),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_27),
.A2(n_32),
.B1(n_95),
.B2(n_245),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_28),
.A2(n_29),
.B1(n_66),
.B2(n_67),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_28),
.B(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_32),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_32),
.B(n_157),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_34),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_93)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_42),
.B(n_48),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_38),
.A2(n_42),
.B1(n_50),
.B2(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_40),
.B1(n_43),
.B2(n_47),
.Y(n_51)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

O2A1O1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_40),
.A2(n_50),
.B(n_140),
.C(n_227),
.Y(n_226)
);

AOI32xp33_ASAP7_75t_L g240 ( 
.A1(n_40),
.A2(n_44),
.A3(n_47),
.B1(n_228),
.B2(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_42),
.B(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_42),
.B(n_53),
.Y(n_107)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_42),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_42),
.A2(n_48),
.B(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_42),
.A2(n_50),
.B1(n_104),
.B2(n_255),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_42)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NAND2xp33_ASAP7_75t_SL g241 ( 
.A(n_43),
.B(n_45),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_44),
.A2(n_45),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_50),
.A2(n_104),
.B(n_106),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_64),
.B1(n_69),
.B2(n_72),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_59),
.A2(n_64),
.B1(n_72),
.B2(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_61),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_61),
.A2(n_63),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

AO22x1_ASAP7_75t_SL g84 ( 
.A1(n_61),
.A2(n_63),
.B1(n_82),
.B2(n_83),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_61),
.B(n_144),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_L g183 ( 
.A1(n_63),
.A2(n_82),
.B(n_140),
.Y(n_183)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_64),
.A2(n_72),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_64),
.B(n_142),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_64),
.A2(n_72),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_64),
.A2(n_72),
.B1(n_100),
.B2(n_234),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_68),
.A2(n_70),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_68),
.A2(n_151),
.B(n_153),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_68),
.B(n_140),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_68),
.A2(n_153),
.B(n_233),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_72),
.B(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_74),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_78),
.B(n_89),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_78),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_76),
.A2(n_139),
.B(n_141),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_76),
.A2(n_141),
.B(n_216),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_79),
.A2(n_85),
.B1(n_87),
.B2(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_79),
.A2(n_188),
.B(n_189),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_79),
.A2(n_87),
.B1(n_203),
.B2(n_231),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_79),
.A2(n_189),
.B(n_231),
.Y(n_253)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_80),
.A2(n_84),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_80),
.B(n_190),
.Y(n_204)
);

NOR2x1_ASAP7_75t_R g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_84),
.B(n_190),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_87),
.A2(n_203),
.B(n_204),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_87),
.A2(n_102),
.B(n_204),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_111),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_90),
.B(n_294),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_101),
.C(n_103),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_91),
.A2(n_92),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_98),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_93),
.A2(n_98),
.B1(n_99),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_93),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_96),
.A2(n_155),
.B(n_156),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_96),
.A2(n_97),
.B1(n_185),
.B2(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_96),
.A2(n_97),
.B1(n_211),
.B2(n_244),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_97),
.A2(n_162),
.B(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_97),
.B(n_140),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_97),
.A2(n_170),
.B(n_185),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_101),
.B(n_103),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_107),
.B(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_121),
.B1(n_122),
.B2(n_124),
.Y(n_111)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_117),
.B1(n_118),
.B2(n_120),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_113),
.Y(n_120)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_127),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_291),
.B(n_296),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_279),
.B(n_290),
.Y(n_129)
);

OAI321xp33_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_247),
.A3(n_272),
.B1(n_277),
.B2(n_278),
.C(n_300),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_220),
.B(n_246),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_197),
.B(n_219),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_178),
.B(n_196),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_158),
.B(n_177),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_145),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_136),
.B(n_145),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_143),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_137),
.A2(n_138),
.B1(n_143),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_154),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_150),
.C(n_154),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_166),
.B(n_176),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_160),
.B(n_164),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_171),
.B(n_175),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_168),
.B(n_169),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_179),
.B(n_180),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_186),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_191),
.C(n_195),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_184),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_191),
.B1(n_194),
.B2(n_195),
.Y(n_186)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_191),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_198),
.B(n_199),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_212),
.B2(n_213),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_215),
.C(n_217),
.Y(n_221)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_206),
.C(n_210),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_209),
.B2(n_210),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_217),
.B2(n_218),
.Y(n_213)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_214),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_221),
.B(n_222),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_236),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_223),
.B(n_237),
.C(n_238),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_229),
.B2(n_235),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_224),
.B(n_230),
.C(n_232),
.Y(n_261)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_229),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_232),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_242),
.B2(n_243),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_243),
.Y(n_257)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_262),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_262),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_258),
.C(n_261),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_249),
.A2(n_250),
.B1(n_275),
.B2(n_276),
.Y(n_274)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_257),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_256),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_256),
.C(n_257),
.Y(n_271)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_254),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_258),
.B(n_261),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_260),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_271),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_266),
.C(n_271),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_270),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_269),
.C(n_270),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_273),
.B(n_274),
.Y(n_277)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_289),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_289),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_284),
.C(n_285),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_293),
.Y(n_296)
);


endmodule