module fake_jpeg_28056_n_135 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_2),
.B(n_3),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_19),
.C(n_16),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_27),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_19),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_33),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_16),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_23),
.A2(n_15),
.B1(n_20),
.B2(n_14),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_15),
.B1(n_23),
.B2(n_22),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_37),
.B(n_22),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_50),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_33),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_54),
.Y(n_63)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_52),
.B1(n_39),
.B2(n_13),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_31),
.A2(n_30),
.B1(n_29),
.B2(n_11),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_49),
.A2(n_52),
.B1(n_39),
.B2(n_41),
.Y(n_57)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_27),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_30),
.B1(n_29),
.B2(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_25),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_27),
.Y(n_59)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_67),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_57),
.B(n_62),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_50),
.Y(n_77)
);

OAI22x1_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_68),
.B1(n_69),
.B2(n_38),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_49),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_65),
.B(n_66),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_13),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_43),
.B(n_11),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_14),
.B1(n_20),
.B2(n_17),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_45),
.A2(n_38),
.B1(n_41),
.B2(n_35),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_50),
.B(n_54),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_71),
.B(n_59),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_73),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

NOR2x1_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_75),
.Y(n_92)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_60),
.Y(n_94)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_78),
.B(n_80),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_51),
.Y(n_79)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_47),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_38),
.B1(n_58),
.B2(n_70),
.Y(n_95)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_93),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_88),
.B(n_79),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_L g88 ( 
.A1(n_77),
.A2(n_60),
.B(n_64),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_76),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_90),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_82),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_91),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_74),
.Y(n_93)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_95),
.A2(n_70),
.B1(n_58),
.B2(n_36),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_72),
.B1(n_73),
.B2(n_71),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_104),
.B1(n_88),
.B2(n_28),
.Y(n_113)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_102),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_100),
.B(n_101),
.Y(n_107)
);

AOI221xp5_ASAP7_75t_L g101 ( 
.A1(n_92),
.A2(n_83),
.B1(n_9),
.B2(n_10),
.C(n_8),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_89),
.B(n_9),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_87),
.C(n_94),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_109),
.C(n_112),
.Y(n_118)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_108),
.B(n_110),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_93),
.C(n_84),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_84),
.C(n_95),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_113),
.A2(n_99),
.B1(n_105),
.B2(n_103),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_114),
.A2(n_36),
.B1(n_28),
.B2(n_2),
.Y(n_120)
);

OA21x2_ASAP7_75t_SL g115 ( 
.A1(n_107),
.A2(n_10),
.B(n_8),
.Y(n_115)
);

NAND4xp25_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_4),
.C(n_5),
.D(n_6),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_27),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_119),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_27),
.C(n_28),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_120),
.A2(n_121),
.B(n_124),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_116),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_122),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_119),
.A2(n_5),
.B1(n_6),
.B2(n_36),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_118),
.C(n_117),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_128),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_118),
.C(n_36),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_120),
.C(n_36),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_129),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_5),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_131),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_130),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_133),
.Y(n_135)
);


endmodule