module real_aes_1539_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_505;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_733;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_0), .B(n_163), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_1), .A2(n_145), .B(n_196), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_2), .A2(n_468), .B1(n_473), .B2(n_818), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_3), .B(n_116), .Y(n_115) );
AOI22xp5_ASAP7_75t_L g129 ( .A1(n_4), .A2(n_11), .B1(n_130), .B2(n_131), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_4), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_5), .B(n_153), .Y(n_209) );
INVx1_ASAP7_75t_L g150 ( .A(n_6), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_7), .B(n_153), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g124 ( .A1(n_8), .A2(n_125), .B1(n_449), .B2(n_450), .Y(n_124) );
INVxp67_ASAP7_75t_L g450 ( .A(n_8), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_8), .B(n_140), .Y(n_509) );
INVx1_ASAP7_75t_L g537 ( .A(n_9), .Y(n_537) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_10), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_11), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g552 ( .A(n_12), .Y(n_552) );
NAND2xp33_ASAP7_75t_L g190 ( .A(n_13), .B(n_157), .Y(n_190) );
INVx2_ASAP7_75t_L g142 ( .A(n_14), .Y(n_142) );
AOI221x1_ASAP7_75t_L g232 ( .A1(n_15), .A2(n_28), .B1(n_145), .B2(n_163), .C(n_233), .Y(n_232) );
AND3x1_ASAP7_75t_L g113 ( .A(n_16), .B(n_40), .C(n_114), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g454 ( .A(n_16), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_17), .B(n_163), .Y(n_186) );
AO21x2_ASAP7_75t_L g183 ( .A1(n_18), .A2(n_184), .B(n_185), .Y(n_183) );
INVx1_ASAP7_75t_L g518 ( .A(n_19), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_20), .B(n_176), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_21), .B(n_153), .Y(n_152) );
AO21x1_ASAP7_75t_L g204 ( .A1(n_22), .A2(n_163), .B(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_SL g110 ( .A(n_23), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g458 ( .A(n_23), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_24), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g516 ( .A(n_25), .Y(n_516) );
INVx1_ASAP7_75t_SL g502 ( .A(n_26), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_27), .B(n_164), .Y(n_596) );
NAND2x1_ASAP7_75t_L g218 ( .A(n_29), .B(n_153), .Y(n_218) );
AOI33xp33_ASAP7_75t_L g564 ( .A1(n_30), .A2(n_55), .A3(n_492), .B1(n_499), .B2(n_565), .B3(n_566), .Y(n_564) );
NAND2x1_ASAP7_75t_L g172 ( .A(n_31), .B(n_157), .Y(n_172) );
INVx1_ASAP7_75t_L g546 ( .A(n_32), .Y(n_546) );
OR2x2_ASAP7_75t_L g141 ( .A(n_33), .B(n_90), .Y(n_141) );
OA21x2_ASAP7_75t_L g181 ( .A1(n_33), .A2(n_90), .B(n_142), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_34), .B(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_35), .B(n_157), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_36), .B(n_153), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_37), .B(n_157), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_38), .A2(n_145), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g146 ( .A(n_39), .B(n_147), .Y(n_146) );
AND2x2_ASAP7_75t_L g161 ( .A(n_39), .B(n_150), .Y(n_161) );
INVx1_ASAP7_75t_L g498 ( .A(n_39), .Y(n_498) );
OR2x6_ASAP7_75t_L g456 ( .A(n_40), .B(n_457), .Y(n_456) );
XNOR2xp5_ASAP7_75t_L g469 ( .A(n_41), .B(n_470), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_42), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_43), .B(n_163), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_44), .B(n_490), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_45), .A2(n_140), .B1(n_180), .B2(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_46), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_47), .B(n_164), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_48), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_49), .B(n_157), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_50), .B(n_184), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_51), .B(n_164), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_52), .A2(n_145), .B(n_171), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g593 ( .A(n_53), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_54), .B(n_157), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_56), .B(n_164), .Y(n_576) );
INVx1_ASAP7_75t_L g149 ( .A(n_57), .Y(n_149) );
INVx1_ASAP7_75t_L g159 ( .A(n_57), .Y(n_159) );
AND2x2_ASAP7_75t_L g577 ( .A(n_58), .B(n_176), .Y(n_577) );
AOI221xp5_ASAP7_75t_L g535 ( .A1(n_59), .A2(n_76), .B1(n_490), .B2(n_496), .C(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_60), .B(n_490), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_61), .B(n_153), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_62), .B(n_180), .Y(n_554) );
AOI21xp5_ASAP7_75t_SL g526 ( .A1(n_63), .A2(n_496), .B(n_527), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_64), .A2(n_145), .B(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g512 ( .A(n_65), .Y(n_512) );
AO21x1_ASAP7_75t_L g206 ( .A1(n_66), .A2(n_145), .B(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_67), .B(n_163), .Y(n_194) );
INVx1_ASAP7_75t_L g575 ( .A(n_68), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_69), .B(n_163), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_70), .A2(n_496), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g255 ( .A(n_71), .B(n_177), .Y(n_255) );
INVx1_ASAP7_75t_L g147 ( .A(n_72), .Y(n_147) );
INVx1_ASAP7_75t_L g155 ( .A(n_72), .Y(n_155) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_73), .A2(n_100), .B1(n_471), .B2(n_472), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_73), .Y(n_471) );
AND2x2_ASAP7_75t_L g178 ( .A(n_74), .B(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_75), .B(n_490), .Y(n_567) );
AND2x2_ASAP7_75t_L g505 ( .A(n_77), .B(n_179), .Y(n_505) );
INVx1_ASAP7_75t_L g513 ( .A(n_78), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_79), .A2(n_496), .B(n_501), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g594 ( .A1(n_80), .A2(n_496), .B(n_559), .C(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g111 ( .A(n_81), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_82), .B(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g192 ( .A(n_83), .B(n_179), .Y(n_192) );
AND2x2_ASAP7_75t_SL g524 ( .A(n_84), .B(n_179), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_85), .A2(n_496), .B1(n_562), .B2(n_563), .Y(n_561) );
CKINVDCx20_ASAP7_75t_R g827 ( .A(n_86), .Y(n_827) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_87), .A2(n_127), .B1(n_128), .B2(n_129), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_87), .Y(n_127) );
XNOR2xp5_ASAP7_75t_L g468 ( .A(n_88), .B(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g205 ( .A(n_89), .B(n_140), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_91), .B(n_157), .Y(n_156) );
AND2x2_ASAP7_75t_L g222 ( .A(n_92), .B(n_179), .Y(n_222) );
INVx1_ASAP7_75t_L g528 ( .A(n_93), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_94), .B(n_153), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_95), .A2(n_145), .B(n_151), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_96), .B(n_157), .Y(n_234) );
AND2x2_ASAP7_75t_L g568 ( .A(n_97), .B(n_179), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_98), .B(n_153), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_99), .A2(n_544), .B(n_545), .C(n_547), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_100), .Y(n_472) );
BUFx2_ASAP7_75t_L g122 ( .A(n_101), .Y(n_122) );
BUFx2_ASAP7_75t_SL g465 ( .A(n_101), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_102), .A2(n_145), .B(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_103), .B(n_164), .Y(n_529) );
AOI21xp33_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_117), .B(n_826), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_SL g828 ( .A(n_108), .Y(n_828) );
OR2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_112), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_111), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OA22x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_123), .B1(n_462), .B2(n_466), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
BUFx3_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_121), .Y(n_120) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OAI21xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_451), .B(n_459), .Y(n_123) );
INVx1_ASAP7_75t_L g449 ( .A(n_125), .Y(n_449) );
XNOR2x1_ASAP7_75t_L g125 ( .A(n_126), .B(n_132), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_129), .Y(n_128) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_132), .A2(n_474), .B1(n_478), .B2(n_481), .Y(n_473) );
INVx2_ASAP7_75t_L g823 ( .A(n_132), .Y(n_823) );
OR2x6_ASAP7_75t_L g132 ( .A(n_133), .B(n_347), .Y(n_132) );
NAND3xp33_ASAP7_75t_SL g133 ( .A(n_134), .B(n_259), .C(n_314), .Y(n_133) );
AOI221xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_199), .B1(n_223), .B2(n_227), .C(n_237), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_182), .Y(n_135) );
AND2x2_ASAP7_75t_SL g225 ( .A(n_136), .B(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g258 ( .A(n_136), .Y(n_258) );
AND2x2_ASAP7_75t_L g303 ( .A(n_136), .B(n_240), .Y(n_303) );
AND2x4_ASAP7_75t_L g136 ( .A(n_137), .B(n_167), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g291 ( .A(n_138), .Y(n_291) );
INVx1_ASAP7_75t_L g301 ( .A(n_138), .Y(n_301) );
AO21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_143), .B(n_165), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_139), .B(n_166), .Y(n_165) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_139), .A2(n_143), .B(n_165), .Y(n_265) );
INVx1_ASAP7_75t_SL g139 ( .A(n_140), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_140), .A2(n_186), .B(n_187), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_140), .B(n_211), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_140), .B(n_160), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_140), .A2(n_526), .B(n_530), .Y(n_525) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x2_ASAP7_75t_SL g177 ( .A(n_141), .B(n_142), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_162), .Y(n_143) );
AND2x6_ASAP7_75t_L g145 ( .A(n_146), .B(n_148), .Y(n_145) );
BUFx3_ASAP7_75t_L g494 ( .A(n_146), .Y(n_494) );
AND2x6_ASAP7_75t_L g157 ( .A(n_147), .B(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g500 ( .A(n_147), .Y(n_500) );
AND2x4_ASAP7_75t_L g496 ( .A(n_148), .B(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
AND2x4_ASAP7_75t_L g153 ( .A(n_149), .B(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g492 ( .A(n_149), .Y(n_492) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_150), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_156), .B(n_160), .Y(n_151) );
INVxp67_ASAP7_75t_L g519 ( .A(n_153), .Y(n_519) );
AND2x4_ASAP7_75t_L g164 ( .A(n_154), .B(n_158), .Y(n_164) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVxp67_ASAP7_75t_L g517 ( .A(n_157), .Y(n_517) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_160), .A2(n_172), .B(n_173), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_160), .A2(n_189), .B(n_190), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_160), .A2(n_197), .B(n_198), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_160), .A2(n_208), .B(n_209), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_160), .A2(n_218), .B(n_219), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_160), .A2(n_234), .B(n_235), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_160), .A2(n_252), .B(n_253), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_SL g501 ( .A1(n_160), .A2(n_502), .B(n_503), .C(n_504), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_160), .A2(n_503), .B(n_528), .C(n_529), .Y(n_527) );
O2A1O1Ixp33_ASAP7_75t_SL g536 ( .A1(n_160), .A2(n_503), .B(n_537), .C(n_538), .Y(n_536) );
INVx1_ASAP7_75t_L g562 ( .A(n_160), .Y(n_562) );
O2A1O1Ixp33_ASAP7_75t_L g574 ( .A1(n_160), .A2(n_503), .B(n_575), .C(n_576), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g595 ( .A1(n_160), .A2(n_596), .B(n_597), .Y(n_595) );
INVx5_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x4_ASAP7_75t_L g163 ( .A(n_161), .B(n_164), .Y(n_163) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_161), .Y(n_547) );
INVx1_ASAP7_75t_L g514 ( .A(n_164), .Y(n_514) );
OR2x2_ASAP7_75t_L g280 ( .A(n_167), .B(n_183), .Y(n_280) );
NAND2x1p5_ASAP7_75t_L g311 ( .A(n_167), .B(n_226), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_167), .B(n_191), .Y(n_324) );
INVx2_ASAP7_75t_L g333 ( .A(n_167), .Y(n_333) );
AND2x2_ASAP7_75t_L g354 ( .A(n_167), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g438 ( .A(n_167), .B(n_257), .Y(n_438) );
INVx4_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g266 ( .A(n_168), .B(n_191), .Y(n_266) );
AND2x2_ASAP7_75t_L g399 ( .A(n_168), .B(n_226), .Y(n_399) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_168), .Y(n_425) );
AO21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_175), .B(n_178), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_170), .B(n_174), .Y(n_169) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_175), .A2(n_488), .B(n_505), .Y(n_487) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_176), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_176), .A2(n_194), .B(n_195), .Y(n_193) );
OA21x2_ASAP7_75t_L g231 ( .A1(n_176), .A2(n_232), .B(n_236), .Y(n_231) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_176), .A2(n_232), .B(n_236), .Y(n_243) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx3_ASAP7_75t_L g221 ( .A(n_179), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_179), .A2(n_221), .B1(n_543), .B2(n_548), .Y(n_542) );
INVx4_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_180), .B(n_551), .Y(n_550) );
INVx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
BUFx4f_ASAP7_75t_L g184 ( .A(n_181), .Y(n_184) );
AND2x4_ASAP7_75t_L g353 ( .A(n_182), .B(n_354), .Y(n_353) );
AOI321xp33_ASAP7_75t_L g367 ( .A1(n_182), .A2(n_296), .A3(n_297), .B1(n_329), .B2(n_368), .C(n_371), .Y(n_367) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_191), .Y(n_182) );
BUFx3_ASAP7_75t_L g224 ( .A(n_183), .Y(n_224) );
INVx2_ASAP7_75t_L g257 ( .A(n_183), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_183), .B(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g290 ( .A(n_183), .B(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g323 ( .A(n_183), .Y(n_323) );
OA21x2_ASAP7_75t_L g534 ( .A1(n_184), .A2(n_535), .B(n_539), .Y(n_534) );
INVx2_ASAP7_75t_SL g559 ( .A(n_184), .Y(n_559) );
INVx5_ASAP7_75t_L g226 ( .A(n_191), .Y(n_226) );
NOR2x1_ASAP7_75t_SL g275 ( .A(n_191), .B(n_265), .Y(n_275) );
BUFx2_ASAP7_75t_L g370 ( .A(n_191), .Y(n_370) );
OR2x6_ASAP7_75t_L g191 ( .A(n_192), .B(n_193), .Y(n_191) );
INVxp67_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_201), .B(n_212), .Y(n_200) );
NOR2xp33_ASAP7_75t_SL g268 ( .A(n_201), .B(n_269), .Y(n_268) );
NOR4xp25_ASAP7_75t_L g371 ( .A(n_201), .B(n_365), .C(n_369), .D(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g409 ( .A(n_201), .Y(n_409) );
AND2x2_ASAP7_75t_L g443 ( .A(n_201), .B(n_383), .Y(n_443) );
BUFx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g244 ( .A(n_202), .Y(n_244) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g298 ( .A(n_203), .Y(n_298) );
OAI21x1_ASAP7_75t_SL g203 ( .A1(n_204), .A2(n_206), .B(n_210), .Y(n_203) );
INVx1_ASAP7_75t_L g211 ( .A(n_205), .Y(n_211) );
AOI33xp33_ASAP7_75t_L g439 ( .A1(n_212), .A2(n_241), .A3(n_272), .B1(n_288), .B2(n_394), .B3(n_440), .Y(n_439) );
INVx1_ASAP7_75t_SL g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g229 ( .A(n_213), .B(n_230), .Y(n_229) );
AND2x4_ASAP7_75t_L g239 ( .A(n_213), .B(n_240), .Y(n_239) );
BUFx3_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g246 ( .A(n_214), .Y(n_246) );
INVxp67_ASAP7_75t_L g327 ( .A(n_214), .Y(n_327) );
AND2x2_ASAP7_75t_L g383 ( .A(n_214), .B(n_248), .Y(n_383) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_221), .B(n_222), .Y(n_214) );
AO21x2_ASAP7_75t_L g287 ( .A1(n_215), .A2(n_221), .B(n_222), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_216), .B(n_220), .Y(n_215) );
AO21x2_ASAP7_75t_L g248 ( .A1(n_221), .A2(n_249), .B(n_255), .Y(n_248) );
AO21x2_ASAP7_75t_L g284 ( .A1(n_221), .A2(n_249), .B(n_255), .Y(n_284) );
AO21x2_ASAP7_75t_L g570 ( .A1(n_221), .A2(n_571), .B(n_577), .Y(n_570) );
AO21x2_ASAP7_75t_L g608 ( .A1(n_221), .A2(n_571), .B(n_577), .Y(n_608) );
AOI21xp5_ASAP7_75t_L g404 ( .A1(n_223), .A2(n_405), .B(n_406), .Y(n_404) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
AND2x2_ASAP7_75t_L g392 ( .A(n_224), .B(n_266), .Y(n_392) );
AND3x2_ASAP7_75t_L g394 ( .A(n_224), .B(n_278), .C(n_333), .Y(n_394) );
INVx3_ASAP7_75t_SL g346 ( .A(n_225), .Y(n_346) );
INVx4_ASAP7_75t_L g240 ( .A(n_226), .Y(n_240) );
AND2x2_ASAP7_75t_L g278 ( .A(n_226), .B(n_265), .Y(n_278) );
INVxp67_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
BUFx2_ASAP7_75t_L g272 ( .A(n_230), .Y(n_272) );
AND2x4_ASAP7_75t_L g297 ( .A(n_230), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g360 ( .A(n_230), .B(n_248), .Y(n_360) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g330 ( .A(n_231), .Y(n_330) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_231), .Y(n_352) );
O2A1O1Ixp33_ASAP7_75t_R g237 ( .A1(n_238), .A2(n_241), .B(n_245), .C(n_256), .Y(n_237) );
CKINVDCx16_ASAP7_75t_R g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g289 ( .A(n_240), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_240), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_240), .B(n_257), .Y(n_418) );
INVx1_ASAP7_75t_SL g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g400 ( .A(n_242), .B(n_390), .Y(n_400) );
AND2x2_ASAP7_75t_SL g242 ( .A(n_243), .B(n_244), .Y(n_242) );
AND2x2_ASAP7_75t_L g247 ( .A(n_243), .B(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g269 ( .A(n_243), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g285 ( .A(n_243), .B(n_286), .Y(n_285) );
AND2x4_ASAP7_75t_L g318 ( .A(n_243), .B(n_298), .Y(n_318) );
AND2x4_ASAP7_75t_L g283 ( .A(n_244), .B(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g307 ( .A(n_244), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g345 ( .A(n_244), .B(n_270), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
AND2x2_ASAP7_75t_L g273 ( .A(n_246), .B(n_270), .Y(n_273) );
AND2x2_ASAP7_75t_L g288 ( .A(n_246), .B(n_248), .Y(n_288) );
BUFx2_ASAP7_75t_L g344 ( .A(n_246), .Y(n_344) );
AND2x2_ASAP7_75t_L g358 ( .A(n_246), .B(n_269), .Y(n_358) );
INVx2_ASAP7_75t_L g270 ( .A(n_248), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_250), .B(n_254), .Y(n_249) );
OAI22xp33_ASAP7_75t_L g306 ( .A1(n_256), .A2(n_307), .B1(n_309), .B2(n_313), .Y(n_306) );
INVx2_ASAP7_75t_SL g337 ( .A(n_256), .Y(n_337) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
AND2x2_ASAP7_75t_L g312 ( .A(n_257), .B(n_265), .Y(n_312) );
INVx1_ASAP7_75t_L g419 ( .A(n_258), .Y(n_419) );
NOR3xp33_ASAP7_75t_L g259 ( .A(n_260), .B(n_292), .C(n_306), .Y(n_259) );
OAI221xp5_ASAP7_75t_SL g260 ( .A1(n_261), .A2(n_267), .B1(n_271), .B2(n_274), .C(n_276), .Y(n_260) );
INVx1_ASAP7_75t_SL g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_266), .Y(n_262) );
INVxp67_ASAP7_75t_SL g263 ( .A(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g320 ( .A(n_264), .Y(n_320) );
INVxp67_ASAP7_75t_SL g448 ( .A(n_264), .Y(n_448) );
INVx1_ASAP7_75t_L g411 ( .A(n_266), .Y(n_411) );
AND2x2_ASAP7_75t_SL g421 ( .A(n_266), .B(n_290), .Y(n_421) );
INVxp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_270), .B(n_298), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
OR2x2_ASAP7_75t_L g304 ( .A(n_272), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g382 ( .A(n_272), .Y(n_382) );
AND2x2_ASAP7_75t_L g317 ( .A(n_273), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g363 ( .A(n_275), .B(n_323), .Y(n_363) );
AND2x2_ASAP7_75t_L g440 ( .A(n_275), .B(n_438), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_281), .B1(n_288), .B2(n_289), .Y(n_276) );
AND2x4_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g299 ( .A(n_280), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
INVx2_ASAP7_75t_L g305 ( .A(n_283), .Y(n_305) );
AND2x4_ASAP7_75t_L g329 ( .A(n_283), .B(n_330), .Y(n_329) );
OAI21xp33_ASAP7_75t_SL g359 ( .A1(n_283), .A2(n_360), .B(n_361), .Y(n_359) );
AND2x2_ASAP7_75t_L g386 ( .A(n_283), .B(n_344), .Y(n_386) );
INVx2_ASAP7_75t_L g308 ( .A(n_284), .Y(n_308) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_284), .Y(n_341) );
INVx1_ASAP7_75t_SL g365 ( .A(n_285), .Y(n_365) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
BUFx2_ASAP7_75t_L g296 ( .A(n_287), .Y(n_296) );
AND2x4_ASAP7_75t_SL g390 ( .A(n_287), .B(n_308), .Y(n_390) );
AND2x2_ASAP7_75t_L g387 ( .A(n_290), .B(n_333), .Y(n_387) );
AND2x2_ASAP7_75t_L g413 ( .A(n_290), .B(n_399), .Y(n_413) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_291), .Y(n_335) );
INVx1_ASAP7_75t_L g355 ( .A(n_291), .Y(n_355) );
OAI22xp33_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_299), .B1(n_302), .B2(n_304), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_297), .B(n_308), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_297), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g436 ( .A(n_297), .Y(n_436) );
INVx2_ASAP7_75t_SL g361 ( .A(n_299), .Y(n_361) );
AND2x2_ASAP7_75t_L g373 ( .A(n_301), .B(n_333), .Y(n_373) );
INVx2_ASAP7_75t_L g379 ( .A(n_301), .Y(n_379) );
INVxp33_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g338 ( .A(n_304), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_307), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g429 ( .A(n_307), .Y(n_429) );
INVx1_ASAP7_75t_L g357 ( .A(n_309), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_310), .B(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g368 ( .A(n_312), .B(n_369), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_312), .A2(n_442), .B1(n_443), .B2(n_444), .Y(n_441) );
NOR3xp33_ASAP7_75t_L g314 ( .A(n_315), .B(n_336), .C(n_339), .Y(n_314) );
OAI221xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_319), .B1(n_321), .B2(n_325), .C(n_328), .Y(n_315) );
INVx1_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_SL g434 ( .A(n_319), .Y(n_434) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g403 ( .A(n_320), .B(n_369), .Y(n_403) );
OR2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g334 ( .A(n_323), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g405 ( .A(n_325), .Y(n_405) );
OR2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
INVx1_ASAP7_75t_L g402 ( .A(n_326), .Y(n_402) );
INVx1_ASAP7_75t_L g408 ( .A(n_327), .Y(n_408) );
OR2x2_ASAP7_75t_L g431 ( .A(n_327), .B(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_331), .Y(n_328) );
INVx1_ASAP7_75t_SL g340 ( .A(n_330), .Y(n_340) );
AND2x2_ASAP7_75t_L g410 ( .A(n_330), .B(n_390), .Y(n_410) );
AND2x2_ASAP7_75t_SL g442 ( .A(n_330), .B(n_343), .Y(n_442) );
INVx1_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx1_ASAP7_75t_L g447 ( .A(n_333), .Y(n_447) );
INVx1_ASAP7_75t_L g397 ( .A(n_335), .Y(n_397) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
O2A1O1Ixp33_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_341), .B(n_342), .C(n_346), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_340), .B(n_390), .Y(n_414) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_343), .B(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
AND2x2_ASAP7_75t_L g351 ( .A(n_345), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g432 ( .A(n_345), .Y(n_432) );
NAND4xp75_ASAP7_75t_L g347 ( .A(n_348), .B(n_404), .C(n_420), .D(n_441), .Y(n_347) );
NOR3x1_ASAP7_75t_L g348 ( .A(n_349), .B(n_366), .C(n_388), .Y(n_348) );
NAND4xp75_ASAP7_75t_L g349 ( .A(n_350), .B(n_356), .C(n_359), .D(n_362), .Y(n_349) );
NAND2xp5_ASAP7_75t_SL g350 ( .A(n_351), .B(n_353), .Y(n_350) );
AND2x2_ASAP7_75t_L g401 ( .A(n_352), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g426 ( .A(n_353), .Y(n_426) );
NAND2xp5_ASAP7_75t_SL g356 ( .A(n_357), .B(n_358), .Y(n_356) );
INVx1_ASAP7_75t_SL g415 ( .A(n_358), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_374), .Y(n_366) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_370), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
AOI21xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_380), .B(n_384), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OAI322xp33_ASAP7_75t_L g406 ( .A1(n_378), .A2(n_407), .A3(n_411), .B1(n_412), .B2(n_414), .C1(n_415), .C2(n_416), .Y(n_406) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_379), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_382), .B(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_383), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
OAI211xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_391), .B(n_393), .C(n_395), .Y(n_388) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_400), .B1(n_401), .B2(n_403), .Y(n_395) );
NOR2xp33_ASAP7_75t_SL g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx2_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_409), .B(n_410), .Y(n_407) );
INVxp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_413), .B(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_417), .B(n_419), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g423 ( .A(n_418), .B(n_424), .Y(n_423) );
O2A1O1Ixp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_422), .B(n_427), .C(n_430), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g422 ( .A(n_423), .B(n_426), .Y(n_422) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OAI221xp5_ASAP7_75t_SL g430 ( .A1(n_431), .A2(n_433), .B1(n_435), .B2(n_437), .C(n_439), .Y(n_430) );
INVxp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx2_ASAP7_75t_L g461 ( .A(n_453), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
AND2x6_ASAP7_75t_SL g477 ( .A(n_454), .B(n_456), .Y(n_477) );
OR2x6_ASAP7_75t_SL g480 ( .A(n_454), .B(n_455), .Y(n_480) );
OR2x2_ASAP7_75t_L g819 ( .A(n_454), .B(n_456), .Y(n_819) );
CKINVDCx5p33_ASAP7_75t_R g455 ( .A(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_459), .B(n_463), .Y(n_462) );
INVx1_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
CKINVDCx11_ASAP7_75t_R g463 ( .A(n_464), .Y(n_463) );
CKINVDCx8_ASAP7_75t_R g464 ( .A(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_467), .B(n_820), .Y(n_466) );
INVx1_ASAP7_75t_L g821 ( .A(n_468), .Y(n_821) );
CKINVDCx6p67_ASAP7_75t_R g474 ( .A(n_475), .Y(n_474) );
INVx4_ASAP7_75t_SL g824 ( .A(n_475), .Y(n_824) );
INVx3_ASAP7_75t_SL g475 ( .A(n_476), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
CKINVDCx11_ASAP7_75t_R g479 ( .A(n_480), .Y(n_479) );
OAI22x1_ASAP7_75t_L g822 ( .A1(n_480), .A2(n_823), .B1(n_824), .B2(n_825), .Y(n_822) );
INVx1_ASAP7_75t_L g825 ( .A(n_481), .Y(n_825) );
OR3x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_683), .C(n_754), .Y(n_481) );
NAND3x1_ASAP7_75t_SL g482 ( .A(n_483), .B(n_610), .C(n_632), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_600), .Y(n_483) );
AOI22xp33_ASAP7_75t_SL g484 ( .A1(n_485), .A2(n_531), .B1(n_578), .B2(n_582), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_485), .A2(n_786), .B1(n_787), .B2(n_789), .Y(n_785) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_506), .Y(n_485) );
AND2x2_ASAP7_75t_L g601 ( .A(n_486), .B(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_486), .B(n_648), .Y(n_667) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g585 ( .A(n_487), .Y(n_585) );
AND2x2_ASAP7_75t_L g635 ( .A(n_487), .B(n_508), .Y(n_635) );
INVx1_ASAP7_75t_L g674 ( .A(n_487), .Y(n_674) );
OR2x2_ASAP7_75t_L g711 ( .A(n_487), .B(n_523), .Y(n_711) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_487), .Y(n_723) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_487), .Y(n_747) );
AND2x2_ASAP7_75t_L g804 ( .A(n_487), .B(n_631), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_495), .Y(n_488) );
INVx1_ASAP7_75t_L g555 ( .A(n_490), .Y(n_555) );
AND2x4_ASAP7_75t_L g490 ( .A(n_491), .B(n_494), .Y(n_490) );
INVx1_ASAP7_75t_L g591 ( .A(n_491), .Y(n_591) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .Y(n_491) );
OR2x6_ASAP7_75t_L g503 ( .A(n_492), .B(n_500), .Y(n_503) );
INVxp33_ASAP7_75t_L g565 ( .A(n_492), .Y(n_565) );
INVx1_ASAP7_75t_L g592 ( .A(n_494), .Y(n_592) );
INVxp67_ASAP7_75t_L g553 ( .A(n_496), .Y(n_553) );
NOR2x1p5_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
INVx1_ASAP7_75t_L g566 ( .A(n_499), .Y(n_566) );
INVx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_503), .A2(n_512), .B1(n_513), .B2(n_514), .Y(n_511) );
INVxp67_ASAP7_75t_L g544 ( .A(n_503), .Y(n_544) );
INVx2_ASAP7_75t_L g598 ( .A(n_503), .Y(n_598) );
NOR2x1_ASAP7_75t_L g506 ( .A(n_507), .B(n_521), .Y(n_506) );
INVx1_ASAP7_75t_L g679 ( .A(n_507), .Y(n_679) );
AND2x2_ASAP7_75t_L g705 ( .A(n_507), .B(n_523), .Y(n_705) );
NAND2x1_ASAP7_75t_L g721 ( .A(n_507), .B(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g602 ( .A(n_508), .B(n_588), .Y(n_602) );
INVx3_ASAP7_75t_L g631 ( .A(n_508), .Y(n_631) );
NOR2x1_ASAP7_75t_SL g750 ( .A(n_508), .B(n_523), .Y(n_750) );
AND2x4_ASAP7_75t_L g508 ( .A(n_509), .B(n_510), .Y(n_508) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_515), .B(n_520), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_514), .B(n_546), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_517), .B1(n_518), .B2(n_519), .Y(n_515) );
NOR2x1_ASAP7_75t_L g658 ( .A(n_521), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g629 ( .A(n_522), .B(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx4_ASAP7_75t_L g599 ( .A(n_523), .Y(n_599) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_523), .Y(n_644) );
AND2x2_ASAP7_75t_L g716 ( .A(n_523), .B(n_588), .Y(n_716) );
AND2x4_ASAP7_75t_L g733 ( .A(n_523), .B(n_677), .Y(n_733) );
NAND2xp5_ASAP7_75t_SL g780 ( .A(n_523), .B(n_675), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_523), .B(n_584), .Y(n_809) );
OR2x6_ASAP7_75t_L g523 ( .A(n_524), .B(n_525), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g738 ( .A1(n_531), .A2(n_626), .B1(n_697), .B2(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_556), .Y(n_531) );
INVx2_ASAP7_75t_L g699 ( .A(n_532), .Y(n_699) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_540), .Y(n_532) );
BUFx3_ASAP7_75t_L g689 ( .A(n_533), .Y(n_689) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_534), .B(n_558), .Y(n_581) );
INVx2_ASAP7_75t_L g605 ( .A(n_534), .Y(n_605) );
INVx1_ASAP7_75t_L g617 ( .A(n_534), .Y(n_617) );
AND2x4_ASAP7_75t_L g624 ( .A(n_534), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g641 ( .A(n_534), .B(n_541), .Y(n_641) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_534), .Y(n_655) );
INVxp67_ASAP7_75t_L g663 ( .A(n_534), .Y(n_663) );
AND2x2_ASAP7_75t_L g692 ( .A(n_540), .B(n_608), .Y(n_692) );
AND2x2_ASAP7_75t_L g708 ( .A(n_540), .B(n_609), .Y(n_708) );
NOR2xp67_ASAP7_75t_L g795 ( .A(n_540), .B(n_608), .Y(n_795) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x4_ASAP7_75t_L g604 ( .A(n_541), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g615 ( .A(n_541), .Y(n_615) );
INVx1_ASAP7_75t_L g628 ( .A(n_541), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_541), .B(n_570), .Y(n_665) );
OR2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_549), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_553), .B1(n_554), .B2(n_555), .Y(n_549) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g788 ( .A(n_556), .Y(n_788) );
AND2x4_ASAP7_75t_L g556 ( .A(n_557), .B(n_569), .Y(n_556) );
AND2x2_ASAP7_75t_L g662 ( .A(n_557), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g691 ( .A(n_557), .Y(n_691) );
AND2x2_ASAP7_75t_L g793 ( .A(n_557), .B(n_608), .Y(n_793) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_558), .B(n_570), .Y(n_653) );
AO21x2_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_560), .B(n_568), .Y(n_558) );
AO21x2_ASAP7_75t_L g609 ( .A1(n_559), .A2(n_560), .B(n_568), .Y(n_609) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_561), .B(n_567), .Y(n_560) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx3_ASAP7_75t_L g579 ( .A(n_569), .Y(n_579) );
NAND2x1p5_ASAP7_75t_L g768 ( .A(n_569), .B(n_689), .Y(n_768) );
INVx3_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_570), .Y(n_682) );
AND2x2_ASAP7_75t_L g709 ( .A(n_570), .B(n_655), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
AND2x2_ASAP7_75t_L g623 ( .A(n_579), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g639 ( .A(n_579), .Y(n_639) );
AND2x2_ASAP7_75t_L g727 ( .A(n_579), .B(n_604), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_579), .B(n_747), .Y(n_752) );
AND2x2_ASAP7_75t_L g762 ( .A(n_579), .B(n_641), .Y(n_762) );
OR2x2_ASAP7_75t_L g799 ( .A(n_579), .B(n_699), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_580), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g759 ( .A(n_580), .B(n_615), .Y(n_759) );
AND2x2_ASAP7_75t_L g775 ( .A(n_580), .B(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g769 ( .A(n_581), .B(n_665), .Y(n_769) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_586), .Y(n_582) );
INVx1_ASAP7_75t_L g651 ( .A(n_583), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_583), .B(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g749 ( .A(n_583), .B(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_583), .B(n_630), .Y(n_774) );
INVx3_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_584), .Y(n_621) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_585), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_586), .A2(n_619), .B1(n_637), .B2(n_640), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_586), .B(n_721), .Y(n_720) );
INVx2_ASAP7_75t_SL g753 ( .A(n_586), .Y(n_753) );
AND2x4_ASAP7_75t_SL g586 ( .A(n_587), .B(n_599), .Y(n_586) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x4_ASAP7_75t_L g630 ( .A(n_588), .B(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g650 ( .A(n_588), .Y(n_650) );
INVx1_ASAP7_75t_L g677 ( .A(n_588), .Y(n_677) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_594), .Y(n_588) );
NOR3xp33_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .C(n_593), .Y(n_590) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_599), .Y(n_619) );
AND2x4_ASAP7_75t_L g676 ( .A(n_599), .B(n_677), .Y(n_676) );
NOR2x1_ASAP7_75t_L g737 ( .A(n_599), .B(n_706), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
AND2x2_ASAP7_75t_L g701 ( .A(n_601), .B(n_644), .Y(n_701) );
OAI21xp5_ASAP7_75t_L g781 ( .A1(n_601), .A2(n_782), .B(n_783), .Y(n_781) );
INVx2_ASAP7_75t_L g659 ( .A(n_602), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g712 ( .A1(n_603), .A2(n_713), .B1(n_717), .B2(n_720), .Y(n_712) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_606), .Y(n_603) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_604), .Y(n_670) );
AND2x2_ASAP7_75t_L g680 ( .A(n_604), .B(n_681), .Y(n_680) );
INVx3_ASAP7_75t_L g719 ( .A(n_604), .Y(n_719) );
NAND2x1_ASAP7_75t_SL g744 ( .A(n_604), .B(n_613), .Y(n_744) );
AND2x2_ASAP7_75t_L g640 ( .A(n_606), .B(n_641), .Y(n_640) );
AND2x4_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NOR2x1_ASAP7_75t_L g616 ( .A(n_608), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g613 ( .A(n_609), .Y(n_613) );
INVx2_ASAP7_75t_L g625 ( .A(n_609), .Y(n_625) );
AOI21xp5_ASAP7_75t_SL g610 ( .A1(n_611), .A2(n_618), .B(n_622), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_613), .B(n_807), .Y(n_806) );
AOI22xp5_ASAP7_75t_L g702 ( .A1(n_614), .A2(n_703), .B1(n_707), .B2(n_710), .Y(n_702) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
BUFx2_ASAP7_75t_L g807 ( .A(n_615), .Y(n_807) );
INVx1_ASAP7_75t_SL g814 ( .A(n_615), .Y(n_814) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_616), .Y(n_777) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OA21x2_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_626), .B(n_629), .Y(n_622) );
AND2x2_ASAP7_75t_L g626 ( .A(n_624), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g668 ( .A(n_624), .B(n_664), .Y(n_668) );
AND2x2_ASAP7_75t_L g783 ( .A(n_624), .B(n_681), .Y(n_783) );
AND2x2_ASAP7_75t_L g786 ( .A(n_624), .B(n_692), .Y(n_786) );
AND2x4_ASAP7_75t_L g794 ( .A(n_624), .B(n_795), .Y(n_794) );
OAI21xp33_ASAP7_75t_L g748 ( .A1(n_626), .A2(n_749), .B(n_751), .Y(n_748) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g776 ( .A(n_628), .Y(n_776) );
AND2x2_ASAP7_75t_L g792 ( .A(n_628), .B(n_793), .Y(n_792) );
INVx4_ASAP7_75t_L g706 ( .A(n_630), .Y(n_706) );
INVx1_ASAP7_75t_L g675 ( .A(n_631), .Y(n_675) );
AND2x2_ASAP7_75t_L g697 ( .A(n_631), .B(n_650), .Y(n_697) );
NOR2x1_ASAP7_75t_L g632 ( .A(n_633), .B(n_656), .Y(n_632) );
OAI21xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_636), .B(n_642), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g643 ( .A(n_635), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_SL g796 ( .A(n_635), .B(n_648), .Y(n_796) );
AND2x2_ASAP7_75t_L g817 ( .A(n_635), .B(n_733), .Y(n_817) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g743 ( .A(n_640), .Y(n_743) );
OAI21xp5_ASAP7_75t_SL g642 ( .A1(n_643), .A2(n_645), .B(n_652), .Y(n_642) );
OR2x6_ASAP7_75t_L g695 ( .A(n_644), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_651), .Y(n_646) );
INVx2_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
OR2x2_ASAP7_75t_L g718 ( .A(n_653), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g815 ( .A(n_653), .Y(n_815) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_654), .B(n_788), .Y(n_787) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_669), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_660), .B1(n_666), .B2(n_668), .Y(n_657) );
OR2x2_ASAP7_75t_L g729 ( .A(n_659), .B(n_730), .Y(n_729) );
INVx3_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_661), .Y(n_686) );
NAND2x1p5_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .Y(n_661) );
INVx1_ASAP7_75t_L g735 ( .A(n_664), .Y(n_735) );
INVx2_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
INVxp67_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_671), .B1(n_678), .B2(n_680), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_673), .B(n_676), .Y(n_672) );
AND2x4_ASAP7_75t_SL g673 ( .A(n_674), .B(n_675), .Y(n_673) );
AND2x2_ASAP7_75t_L g678 ( .A(n_676), .B(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g739 ( .A(n_679), .B(n_733), .Y(n_739) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_684), .B(n_724), .Y(n_683) );
NOR2xp67_ASAP7_75t_L g684 ( .A(n_685), .B(n_698), .Y(n_684) );
AOI21xp33_ASAP7_75t_SL g685 ( .A1(n_686), .A2(n_687), .B(n_693), .Y(n_685) );
OR2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_690), .Y(n_687) );
INVx3_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND2x1p5_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OAI22xp33_ASAP7_75t_SL g763 ( .A1(n_695), .A2(n_764), .B1(n_766), .B2(n_769), .Y(n_763) );
NOR2x1_ASAP7_75t_L g710 ( .A(n_696), .B(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g746 ( .A(n_697), .B(n_747), .Y(n_746) );
OAI211xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_700), .B(n_702), .C(n_712), .Y(n_698) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND2xp33_ASAP7_75t_SL g703 ( .A(n_704), .B(n_706), .Y(n_703) );
INVxp33_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g715 ( .A(n_706), .Y(n_715) );
AOI221xp5_ASAP7_75t_L g726 ( .A1(n_707), .A2(n_727), .B1(n_728), .B2(n_731), .C(n_734), .Y(n_726) );
AND2x4_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
INVx1_ASAP7_75t_L g767 ( .A(n_708), .Y(n_767) );
INVx2_ASAP7_75t_SL g765 ( .A(n_711), .Y(n_765) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
NAND2x1_ASAP7_75t_L g764 ( .A(n_715), .B(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g761 ( .A(n_721), .Y(n_761) );
INVx1_ASAP7_75t_L g790 ( .A(n_722), .Y(n_790) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
NOR2x1_ASAP7_75t_L g724 ( .A(n_725), .B(n_740), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_726), .B(n_738), .Y(n_725) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g779 ( .A(n_730), .Y(n_779) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AND2x2_ASAP7_75t_L g800 ( .A(n_733), .B(n_801), .Y(n_800) );
INVx2_ASAP7_75t_L g805 ( .A(n_733), .Y(n_805) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
INVxp33_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
BUFx2_ASAP7_75t_L g758 ( .A(n_737), .Y(n_758) );
OAI21xp5_ASAP7_75t_SL g740 ( .A1(n_741), .A2(n_745), .B(n_748), .Y(n_740) );
INVxp67_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
BUFx2_ASAP7_75t_L g801 ( .A(n_747), .Y(n_801) );
AND2x2_ASAP7_75t_L g789 ( .A(n_750), .B(n_790), .Y(n_789) );
NOR2xp33_ASAP7_75t_R g751 ( .A(n_752), .B(n_753), .Y(n_751) );
NAND3xp33_ASAP7_75t_L g754 ( .A(n_755), .B(n_770), .C(n_797), .Y(n_754) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_756), .B(n_763), .Y(n_755) );
NAND2xp5_ASAP7_75t_SL g756 ( .A(n_757), .B(n_760), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
OR2x2_ASAP7_75t_L g766 ( .A(n_767), .B(n_768), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g770 ( .A(n_771), .B(n_784), .Y(n_770) );
NAND2xp5_ASAP7_75t_SL g771 ( .A(n_772), .B(n_781), .Y(n_771) );
AOI22xp33_ASAP7_75t_SL g772 ( .A1(n_773), .A2(n_775), .B1(n_777), .B2(n_778), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
NOR2x1_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
INVxp67_ASAP7_75t_SL g782 ( .A(n_780), .Y(n_782) );
NAND2xp5_ASAP7_75t_SL g784 ( .A(n_785), .B(n_791), .Y(n_784) );
OAI21xp5_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_794), .B(n_796), .Y(n_791) );
INVx1_ASAP7_75t_L g810 ( .A(n_794), .Y(n_810) );
AOI211xp5_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_800), .B(n_802), .C(n_811), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g802 ( .A1(n_803), .A2(n_806), .B1(n_808), .B2(n_810), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .Y(n_803) );
HB1xp67_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
NOR2xp33_ASAP7_75t_L g811 ( .A(n_812), .B(n_816), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
AND2x2_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .Y(n_813) );
INVxp67_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx2_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_821), .B(n_822), .Y(n_820) );
NOR2xp33_ASAP7_75t_L g826 ( .A(n_827), .B(n_828), .Y(n_826) );
endmodule