module fake_jpeg_30034_n_407 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_407);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_407;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx4f_ASAP7_75t_SL g41 ( 
.A(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_2),
.B(n_12),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_51),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_15),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_44),
.B(n_47),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_14),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_20),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_50),
.B(n_52),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_13),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_20),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_20),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_56),
.B(n_58),
.Y(n_116)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_27),
.B(n_40),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_63),
.Y(n_119)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_17),
.B(n_0),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_68),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_27),
.B(n_13),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_12),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_70),
.B(n_71),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_10),
.Y(n_71)
);

BUFx16f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_72),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_79),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_40),
.B(n_10),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_80),
.Y(n_101)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_43),
.A2(n_31),
.B1(n_38),
.B2(n_17),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_82),
.B(n_122),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_31),
.B1(n_38),
.B2(n_29),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_84),
.A2(n_118),
.B1(n_124),
.B2(n_127),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_76),
.A2(n_34),
.B1(n_35),
.B2(n_21),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_98),
.A2(n_105),
.B1(n_121),
.B2(n_125),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g104 ( 
.A(n_66),
.B(n_18),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_37),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_57),
.A2(n_35),
.B1(n_34),
.B2(n_28),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_72),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_123),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_65),
.A2(n_29),
.B1(n_24),
.B2(n_19),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_77),
.A2(n_35),
.B1(n_34),
.B2(n_28),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_43),
.A2(n_24),
.B1(n_19),
.B2(n_16),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_72),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_67),
.A2(n_16),
.B1(n_28),
.B2(n_32),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_59),
.A2(n_28),
.B1(n_32),
.B2(n_18),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_L g127 ( 
.A1(n_45),
.A2(n_28),
.B1(n_37),
.B2(n_32),
.Y(n_127)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_129),
.Y(n_184)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_132),
.Y(n_174)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_134),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_82),
.A2(n_54),
.B1(n_48),
.B2(n_49),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_136),
.A2(n_163),
.B1(n_103),
.B2(n_119),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_137),
.Y(n_202)
);

BUFx8_ASAP7_75t_L g138 ( 
.A(n_86),
.Y(n_138)
);

BUFx10_ASAP7_75t_L g185 ( 
.A(n_138),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_106),
.A2(n_64),
.B1(n_62),
.B2(n_74),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_139),
.Y(n_203)
);

INVx11_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_140),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_46),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_141),
.B(n_149),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_94),
.A2(n_53),
.B1(n_81),
.B2(n_69),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_142),
.A2(n_173),
.B1(n_88),
.B2(n_109),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_143),
.B(n_148),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_85),
.A2(n_60),
.B1(n_55),
.B2(n_73),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_144),
.A2(n_153),
.B1(n_7),
.B2(n_9),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_145),
.Y(n_214)
);

OR2x2_ASAP7_75t_SL g146 ( 
.A(n_122),
.B(n_37),
.Y(n_146)
);

NAND3xp33_ASAP7_75t_L g196 ( 
.A(n_146),
.B(n_4),
.C(n_5),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_83),
.B(n_37),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_151),
.Y(n_183)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_104),
.B(n_92),
.Y(n_149)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_95),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_152),
.Y(n_179)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_114),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_85),
.A2(n_75),
.B1(n_78),
.B2(n_4),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

BUFx12_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_101),
.B(n_116),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_158),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_78),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_157),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_99),
.B(n_1),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_113),
.Y(n_158)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_100),
.B(n_3),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_159),
.B(n_109),
.C(n_6),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_79),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_168),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_95),
.B(n_61),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_162),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_117),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_112),
.A2(n_102),
.B1(n_94),
.B2(n_110),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_100),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_164),
.B(n_169),
.Y(n_177)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_167),
.Y(n_206)
);

INVx11_ASAP7_75t_L g166 ( 
.A(n_119),
.Y(n_166)
);

BUFx12_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_86),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_87),
.B(n_61),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_102),
.B(n_3),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_86),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_171),
.Y(n_210)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_87),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_111),
.B(n_3),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_167),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_103),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_180),
.B(n_190),
.Y(n_226)
);

OAI22x1_ASAP7_75t_SL g182 ( 
.A1(n_131),
.A2(n_111),
.B1(n_120),
.B2(n_110),
.Y(n_182)
);

AO22x1_ASAP7_75t_SL g248 ( 
.A1(n_182),
.A2(n_190),
.B1(n_188),
.B2(n_176),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_128),
.A2(n_93),
.B(n_90),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_188),
.A2(n_194),
.B(n_205),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_128),
.A2(n_96),
.B1(n_93),
.B2(n_90),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_149),
.B(n_120),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_191),
.B(n_209),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_160),
.A2(n_4),
.B(n_5),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_151),
.B(n_88),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_208),
.C(n_212),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_196),
.A2(n_157),
.B(n_143),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_200),
.B(n_212),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_160),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_128),
.A2(n_141),
.B1(n_156),
.B2(n_169),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_204),
.A2(n_207),
.B1(n_135),
.B2(n_163),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_168),
.A2(n_7),
.B(n_9),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_147),
.B(n_7),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_147),
.B(n_159),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_167),
.Y(n_231)
);

XOR2x2_ASAP7_75t_L g212 ( 
.A(n_146),
.B(n_159),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_132),
.B(n_168),
.C(n_164),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_154),
.C(n_145),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_215),
.Y(n_271)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_174),
.Y(n_216)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_216),
.Y(n_258)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_174),
.Y(n_217)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_217),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_198),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_218),
.B(n_231),
.Y(n_259)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_186),
.Y(n_220)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_220),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_182),
.A2(n_135),
.B1(n_152),
.B2(n_133),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_221),
.A2(n_240),
.B1(n_248),
.B2(n_189),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_192),
.B(n_130),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_228),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_227),
.A2(n_213),
.B1(n_200),
.B2(n_183),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_187),
.B(n_148),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_150),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_229),
.B(n_236),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_203),
.A2(n_162),
.B(n_137),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_230),
.A2(n_234),
.B(n_247),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_210),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_239),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_209),
.A2(n_165),
.B(n_129),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_235),
.B(n_242),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_181),
.B(n_134),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_177),
.B(n_167),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_237),
.B(n_241),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_203),
.A2(n_166),
.B1(n_140),
.B2(n_138),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_238),
.B(n_245),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_206),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_180),
.A2(n_138),
.B1(n_191),
.B2(n_177),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_184),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_195),
.B(n_192),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_186),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_243),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_199),
.B(n_204),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_244),
.Y(n_264)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_179),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_193),
.C(n_202),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_212),
.A2(n_183),
.B(n_194),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_185),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_249),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_183),
.B(n_208),
.Y(n_250)
);

OAI21xp33_ASAP7_75t_SL g266 ( 
.A1(n_250),
.A2(n_178),
.B(n_185),
.Y(n_266)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_193),
.Y(n_251)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_251),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_253),
.A2(n_256),
.B1(n_216),
.B2(n_217),
.Y(n_310)
);

XOR2x1_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_176),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_254),
.A2(n_257),
.B(n_276),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_227),
.A2(n_199),
.B1(n_205),
.B2(n_207),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_222),
.A2(n_175),
.B1(n_202),
.B2(n_184),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_265),
.C(n_235),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_219),
.A2(n_214),
.B(n_175),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_261),
.A2(n_277),
.B(n_215),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_225),
.B(n_214),
.C(n_178),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_237),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_232),
.A2(n_189),
.B1(n_178),
.B2(n_185),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_272),
.Y(n_286)
);

AO22x1_ASAP7_75t_L g269 ( 
.A1(n_248),
.A2(n_189),
.B1(n_178),
.B2(n_185),
.Y(n_269)
);

OA21x2_ASAP7_75t_L g304 ( 
.A1(n_269),
.A2(n_229),
.B(n_251),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_230),
.A2(n_189),
.B(n_234),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_219),
.A2(n_224),
.B(n_225),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_236),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_233),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_226),
.A2(n_231),
.B(n_248),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_280),
.A2(n_226),
.B(n_238),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_221),
.A2(n_226),
.B1(n_240),
.B2(n_248),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_282),
.B(n_272),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_284),
.A2(n_282),
.B1(n_283),
.B2(n_259),
.Y(n_321)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_258),
.Y(n_285)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_285),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_287),
.B(n_291),
.C(n_300),
.Y(n_312)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_270),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_290),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_289),
.A2(n_304),
.B(n_307),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_268),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_242),
.C(n_246),
.Y(n_291)
);

NOR2x1_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_223),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_292),
.B(n_296),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_293),
.A2(n_280),
.B(n_274),
.Y(n_320)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_258),
.Y(n_294)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_294),
.Y(n_327)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_267),
.Y(n_295)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_295),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_262),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_267),
.Y(n_297)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_297),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_298),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_250),
.C(n_224),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_255),
.B(n_228),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_308),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_263),
.B(n_218),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_302),
.Y(n_326)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_281),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_303),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_264),
.B(n_245),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_305),
.B(n_306),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_273),
.A2(n_276),
.B(n_261),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_263),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_255),
.B(n_278),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_270),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_310),
.B(n_254),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_287),
.B(n_265),
.C(n_260),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_315),
.B(n_319),
.C(n_325),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_316),
.B(n_321),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_286),
.A2(n_269),
.B1(n_273),
.B2(n_274),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_317),
.A2(n_284),
.B1(n_288),
.B2(n_286),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_291),
.B(n_300),
.C(n_277),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_320),
.B(n_322),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_306),
.B(n_283),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_310),
.B(n_271),
.C(n_274),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_331),
.C(n_286),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_293),
.B(n_299),
.C(n_307),
.Y(n_331)
);

AO21x2_ASAP7_75t_L g336 ( 
.A1(n_328),
.A2(n_304),
.B(n_299),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_336),
.A2(n_304),
.B1(n_321),
.B2(n_301),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_328),
.A2(n_292),
.B(n_289),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_337),
.B(n_341),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_338),
.B(n_340),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_339),
.B(n_315),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_313),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_326),
.B(n_302),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_314),
.Y(n_342)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_342),
.Y(n_353)
);

BUFx12_ASAP7_75t_L g344 ( 
.A(n_317),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_344),
.B(n_350),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_333),
.B(n_298),
.Y(n_345)
);

CKINVDCx14_ASAP7_75t_R g365 ( 
.A(n_345),
.Y(n_365)
);

CKINVDCx14_ASAP7_75t_R g346 ( 
.A(n_311),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_346),
.B(n_348),
.Y(n_356)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_324),
.Y(n_347)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_347),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_316),
.B(n_309),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_331),
.A2(n_286),
.B(n_292),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_349),
.A2(n_352),
.B(n_329),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_325),
.B(n_296),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_318),
.B(n_305),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_351),
.B(n_318),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_323),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_355),
.B(n_358),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_357),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_343),
.B(n_322),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_336),
.A2(n_304),
.B(n_308),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_359),
.B(n_366),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_360),
.B(n_338),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_363),
.B(n_335),
.C(n_312),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_336),
.A2(n_271),
.B(n_319),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_340),
.A2(n_312),
.B1(n_330),
.B2(n_327),
.Y(n_367)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_367),
.Y(n_373)
);

BUFx4f_ASAP7_75t_SL g368 ( 
.A(n_365),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_368),
.B(n_374),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_364),
.B(n_342),
.Y(n_371)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_371),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_372),
.B(n_363),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_361),
.B(n_345),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_375),
.B(n_334),
.Y(n_388)
);

NOR2x1_ASAP7_75t_L g377 ( 
.A(n_360),
.B(n_348),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_377),
.A2(n_378),
.B1(n_356),
.B2(n_367),
.Y(n_382)
);

INVx5_ASAP7_75t_L g378 ( 
.A(n_353),
.Y(n_378)
);

A2O1A1Ixp33_ASAP7_75t_L g379 ( 
.A1(n_370),
.A2(n_359),
.B(n_337),
.C(n_362),
.Y(n_379)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_379),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_376),
.A2(n_336),
.B1(n_352),
.B2(n_354),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_381),
.A2(n_384),
.B1(n_385),
.B2(n_386),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_382),
.B(n_383),
.Y(n_394)
);

OAI321xp33_ASAP7_75t_L g384 ( 
.A1(n_368),
.A2(n_362),
.A3(n_334),
.B1(n_336),
.B2(n_366),
.C(n_344),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_373),
.A2(n_357),
.B(n_349),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_372),
.A2(n_339),
.B(n_335),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_388),
.B(n_369),
.C(n_355),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_390),
.B(n_392),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_380),
.B(n_368),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_391),
.A2(n_395),
.B(n_378),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_387),
.B(n_388),
.C(n_379),
.Y(n_392)
);

NAND3xp33_ASAP7_75t_L g395 ( 
.A(n_381),
.B(n_377),
.C(n_347),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_387),
.Y(n_396)
);

AOI322xp5_ASAP7_75t_L g398 ( 
.A1(n_396),
.A2(n_393),
.A3(n_389),
.B1(n_323),
.B2(n_303),
.C1(n_332),
.C2(n_391),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_397),
.B(n_398),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_394),
.B(n_249),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_400),
.B(n_275),
.C(n_252),
.Y(n_402)
);

AOI322xp5_ASAP7_75t_L g401 ( 
.A1(n_395),
.A2(n_294),
.A3(n_297),
.B1(n_285),
.B2(n_295),
.C1(n_344),
.C2(n_281),
.Y(n_401)
);

A2O1A1O1Ixp25_ASAP7_75t_L g403 ( 
.A1(n_401),
.A2(n_275),
.B(n_220),
.C(n_252),
.D(n_243),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_402),
.B(n_403),
.C(n_399),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_405),
.B(n_404),
.C(n_369),
.Y(n_406)
);

FAx1_ASAP7_75t_SL g407 ( 
.A(n_406),
.B(n_358),
.CI(n_343),
.CON(n_407),
.SN(n_407)
);


endmodule