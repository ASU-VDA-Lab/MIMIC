module fake_jpeg_1825_n_721 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_721);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_721;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_716;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_717;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_718;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_713;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_701;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_704;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_715;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_539;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_720;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_710;
wire n_610;
wire n_174;
wire n_714;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_709;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_708;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_703;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_702;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_719;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_707;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_705;
wire n_665;
wire n_706;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_700;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_712;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_711;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_19),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_4),
.B(n_19),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_1),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_11),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_1),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_31),
.B(n_8),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_62),
.B(n_70),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_63),
.Y(n_149)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_31),
.B(n_9),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_65),
.B(n_74),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_66),
.Y(n_157)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g180 ( 
.A(n_67),
.Y(n_180)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_68),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_69),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_22),
.B(n_9),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_35),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_71),
.B(n_75),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_72),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_73),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_22),
.B(n_9),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_35),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_76),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_77),
.Y(n_172)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_45),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g146 ( 
.A(n_78),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_79),
.Y(n_190)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_80),
.Y(n_182)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_82),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_36),
.B(n_9),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_83),
.B(n_96),
.Y(n_143)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_85),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_86),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_87),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_88),
.Y(n_218)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_89),
.Y(n_176)
);

BUFx12_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx6_ASAP7_75t_SL g223 ( 
.A(n_90),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_23),
.Y(n_91)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_91),
.Y(n_177)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_92),
.Y(n_166)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_93),
.Y(n_174)
);

BUFx4f_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_94),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_95),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_7),
.Y(n_96)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

INVx3_ASAP7_75t_SL g153 ( 
.A(n_97),
.Y(n_153)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_27),
.Y(n_98)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_98),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_100),
.Y(n_184)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_101),
.Y(n_178)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_103),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_41),
.Y(n_104)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_106),
.Y(n_175)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_21),
.Y(n_107)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_107),
.Y(n_194)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_108),
.Y(n_162)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_21),
.Y(n_109)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_109),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_110),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_111),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_112),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_25),
.Y(n_113)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_40),
.Y(n_114)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_114),
.Y(n_173)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_25),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_115),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_61),
.B(n_7),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_116),
.B(n_117),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_50),
.B(n_17),
.Y(n_117)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_118),
.Y(n_206)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_25),
.Y(n_119)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_119),
.Y(n_221)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_50),
.Y(n_120)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_120),
.Y(n_210)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_40),
.Y(n_121)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_121),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_40),
.Y(n_122)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_42),
.Y(n_123)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_42),
.Y(n_124)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_124),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_42),
.B(n_7),
.C(n_16),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_128),
.Y(n_152)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_40),
.Y(n_126)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_126),
.Y(n_227)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_39),
.Y(n_127)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_127),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_20),
.B(n_10),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_39),
.Y(n_129)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_129),
.Y(n_224)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_39),
.Y(n_130)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_130),
.Y(n_181)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_39),
.Y(n_131)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_131),
.Y(n_189)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_39),
.Y(n_132)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_132),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_20),
.B(n_10),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_133),
.B(n_134),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_24),
.B(n_10),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_70),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_136),
.A2(n_154),
.B1(n_159),
.B2(n_167),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_100),
.A2(n_59),
.B1(n_26),
.B2(n_57),
.Y(n_151)
);

OA22x2_ASAP7_75t_L g292 ( 
.A1(n_151),
.A2(n_158),
.B1(n_202),
.B2(n_203),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_97),
.A2(n_59),
.B1(n_26),
.B2(n_57),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_78),
.B(n_79),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_156),
.B(n_183),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_94),
.A2(n_53),
.B1(n_37),
.B2(n_44),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_103),
.A2(n_24),
.B1(n_30),
.B2(n_52),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_88),
.A2(n_52),
.B1(n_30),
.B2(n_58),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_110),
.A2(n_53),
.B1(n_34),
.B2(n_58),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_169),
.A2(n_195),
.B1(n_208),
.B2(n_131),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_79),
.B(n_34),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_108),
.B(n_29),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_188),
.B(n_193),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_104),
.A2(n_44),
.B1(n_29),
.B2(n_43),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_192),
.A2(n_209),
.B1(n_219),
.B2(n_222),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_122),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_105),
.A2(n_37),
.B1(n_43),
.B2(n_46),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_124),
.B(n_46),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_199),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_90),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_114),
.Y(n_200)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_200),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_123),
.A2(n_37),
.B1(n_44),
.B2(n_54),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_95),
.A2(n_44),
.B1(n_54),
.B2(n_55),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_111),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_204),
.B(n_205),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_72),
.B(n_12),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_73),
.A2(n_48),
.B1(n_54),
.B2(n_51),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_207),
.A2(n_219),
.B1(n_222),
.B2(n_228),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_112),
.A2(n_48),
.B1(n_54),
.B2(n_55),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_99),
.A2(n_66),
.B1(n_63),
.B2(n_76),
.Y(n_209)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_118),
.Y(n_215)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_215),
.Y(n_250)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_129),
.Y(n_217)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_217),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_77),
.A2(n_54),
.B1(n_48),
.B2(n_2),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_95),
.A2(n_54),
.B1(n_48),
.B2(n_51),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_90),
.A2(n_48),
.B1(n_51),
.B2(n_11),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_228),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_91),
.B(n_48),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_229),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_230),
.Y(n_348)
);

INVx8_ASAP7_75t_L g231 ( 
.A(n_138),
.Y(n_231)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_231),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_223),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_232),
.B(n_240),
.Y(n_315)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

INVx4_ASAP7_75t_L g341 ( 
.A(n_233),
.Y(n_341)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_235),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_198),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_236),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_237),
.A2(n_249),
.B1(n_262),
.B2(n_270),
.Y(n_343)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_227),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g329 ( 
.A(n_238),
.Y(n_329)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_198),
.Y(n_239)
);

INVx8_ASAP7_75t_L g352 ( 
.A(n_239),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_226),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_147),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_241),
.B(n_252),
.Y(n_317)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_161),
.Y(n_243)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_243),
.Y(n_314)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_192),
.Y(n_244)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_244),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_126),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_246),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_143),
.B(n_113),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_247),
.Y(n_342)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_153),
.Y(n_248)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_248),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_209),
.A2(n_64),
.B1(n_51),
.B2(n_2),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_201),
.Y(n_251)
);

INVx6_ASAP7_75t_L g312 ( 
.A(n_251),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_11),
.Y(n_252)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_153),
.Y(n_254)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_254),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_201),
.Y(n_255)
);

INVx6_ASAP7_75t_L g354 ( 
.A(n_255),
.Y(n_354)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_216),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_256),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_179),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_258),
.B(n_261),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_213),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g374 ( 
.A(n_259),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_213),
.Y(n_260)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_260),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_135),
.B(n_144),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_152),
.A2(n_64),
.B1(n_51),
.B2(n_2),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_195),
.A2(n_17),
.B1(n_16),
.B2(n_15),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_263),
.A2(n_279),
.B1(n_137),
.B2(n_142),
.Y(n_327)
);

O2A1O1Ixp33_ASAP7_75t_L g264 ( 
.A1(n_203),
.A2(n_202),
.B(n_145),
.C(n_148),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_264),
.A2(n_172),
.B(n_137),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_265),
.B(n_280),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_146),
.B(n_0),
.Y(n_266)
);

AND2x2_ASAP7_75t_SL g367 ( 
.A(n_266),
.B(n_286),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_179),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_267),
.B(n_277),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_182),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_268),
.A2(n_274),
.B1(n_281),
.B2(n_290),
.Y(n_323)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_190),
.Y(n_269)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_269),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_185),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_182),
.A2(n_14),
.B1(n_12),
.B2(n_3),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_166),
.B(n_0),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_275),
.B(n_168),
.Y(n_320)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_227),
.Y(n_276)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_276),
.Y(n_361)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_206),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_218),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_278),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_174),
.A2(n_12),
.B1(n_1),
.B2(n_3),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_178),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_146),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_282),
.B(n_284),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_194),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_283),
.A2(n_302),
.B1(n_303),
.B2(n_248),
.Y(n_369)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_221),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_181),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_285),
.B(n_287),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_196),
.B(n_210),
.Y(n_286)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_171),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_221),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_288),
.B(n_289),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_211),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_171),
.A2(n_4),
.B1(n_6),
.B2(n_184),
.Y(n_290)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_218),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_291),
.Y(n_336)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_177),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_293),
.B(n_295),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_211),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_294),
.B(n_305),
.Y(n_350)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_150),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_176),
.A2(n_141),
.B1(n_162),
.B2(n_173),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_296),
.A2(n_180),
.B1(n_138),
.B2(n_173),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_186),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_297),
.B(n_298),
.Y(n_357)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_177),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_189),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_299),
.B(n_300),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_149),
.Y(n_300)
);

INVx4_ASAP7_75t_SL g301 ( 
.A(n_138),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_301),
.B(n_306),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_155),
.A2(n_225),
.B1(n_163),
.B2(n_158),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_155),
.A2(n_225),
.B1(n_163),
.B2(n_139),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_141),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_186),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_190),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_307),
.B(n_308),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_140),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_224),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_309),
.B(n_310),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_170),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_162),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_311),
.B(n_310),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_244),
.A2(n_170),
.B1(n_157),
.B2(n_160),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_313),
.A2(n_356),
.B1(n_364),
.B2(n_369),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_242),
.B(n_165),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_319),
.B(n_305),
.C(n_233),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_320),
.B(n_345),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_275),
.B(n_175),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_325),
.B(n_332),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_L g389 ( 
.A1(n_327),
.A2(n_251),
.B1(n_278),
.B2(n_236),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_270),
.B(n_212),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_335),
.Y(n_379)
);

NAND2xp33_ASAP7_75t_SL g337 ( 
.A(n_273),
.B(n_191),
.Y(n_337)
);

OAI21xp33_ASAP7_75t_L g402 ( 
.A1(n_337),
.A2(n_360),
.B(n_350),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_262),
.B(n_214),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_338),
.B(n_339),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_304),
.B(n_140),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_272),
.A2(n_180),
.B1(n_164),
.B2(n_149),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_340),
.A2(n_344),
.B1(n_358),
.B2(n_301),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_246),
.A2(n_164),
.B1(n_157),
.B2(n_160),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_257),
.B(n_142),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_346),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_266),
.B(n_172),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_353),
.B(n_360),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_L g356 ( 
.A1(n_271),
.A2(n_237),
.B1(n_263),
.B2(n_264),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_246),
.A2(n_234),
.B1(n_249),
.B2(n_292),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_286),
.B(n_266),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_292),
.A2(n_280),
.B1(n_286),
.B2(n_291),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_253),
.B(n_250),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_371),
.B(n_317),
.Y(n_410)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_372),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_L g373 ( 
.A1(n_292),
.A2(n_295),
.B1(n_288),
.B2(n_284),
.Y(n_373)
);

OAI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_373),
.A2(n_254),
.B1(n_298),
.B2(n_293),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_292),
.A2(n_239),
.B1(n_277),
.B2(n_259),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_375),
.A2(n_346),
.B1(n_364),
.B2(n_327),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_376),
.B(n_407),
.Y(n_457)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_318),
.Y(n_378)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_378),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_380),
.B(n_424),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_365),
.B(n_245),
.C(n_243),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_381),
.B(n_391),
.C(n_393),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_349),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_382),
.Y(n_463)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_318),
.Y(n_383)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_383),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_342),
.B(n_240),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_385),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_386),
.A2(n_420),
.B(n_347),
.Y(n_442)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_333),
.Y(n_387)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_387),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_343),
.A2(n_303),
.B1(n_283),
.B2(n_309),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_388),
.A2(n_415),
.B1(n_336),
.B2(n_326),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_L g427 ( 
.A1(n_389),
.A2(n_392),
.B1(n_374),
.B2(n_331),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_328),
.A2(n_307),
.B1(n_276),
.B2(n_238),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_SL g429 ( 
.A1(n_390),
.A2(n_408),
.B1(n_374),
.B2(n_331),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_365),
.B(n_311),
.C(n_287),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_319),
.B(n_294),
.Y(n_393)
);

OAI321xp33_ASAP7_75t_L g394 ( 
.A1(n_328),
.A2(n_255),
.A3(n_260),
.B1(n_269),
.B2(n_300),
.C(n_256),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_394),
.B(n_406),
.Y(n_433)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_333),
.Y(n_395)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_395),
.Y(n_439)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_314),
.Y(n_397)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_397),
.Y(n_448)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_314),
.Y(n_399)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_399),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_367),
.B(n_231),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_400),
.B(n_403),
.C(n_413),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_316),
.B(n_235),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_401),
.B(n_404),
.Y(n_435)
);

CKINVDCx14_ASAP7_75t_R g455 ( 
.A(n_402),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_367),
.B(n_320),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_371),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_368),
.Y(n_405)
);

INVx2_ASAP7_75t_SL g430 ( 
.A(n_405),
.Y(n_430)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_368),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_L g408 ( 
.A1(n_351),
.A2(n_375),
.B1(n_338),
.B2(n_339),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_325),
.B(n_332),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_409),
.B(n_421),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_410),
.B(n_412),
.Y(n_450)
);

BUFx5_ASAP7_75t_L g411 ( 
.A(n_321),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_411),
.Y(n_444)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_329),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_367),
.B(n_360),
.Y(n_413)
);

INVx13_ASAP7_75t_L g414 ( 
.A(n_363),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_414),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_343),
.A2(n_328),
.B1(n_369),
.B2(n_351),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_350),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_416),
.B(n_422),
.Y(n_459)
);

NAND2x1p5_ASAP7_75t_L g417 ( 
.A(n_367),
.B(n_337),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_417),
.A2(n_423),
.B(n_420),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_316),
.B(n_345),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_418),
.B(n_425),
.Y(n_440)
);

FAx1_ASAP7_75t_L g420 ( 
.A(n_353),
.B(n_357),
.CI(n_366),
.CON(n_420),
.SN(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_357),
.B(n_362),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_350),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_315),
.B(n_330),
.C(n_366),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_315),
.B(n_330),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_420),
.A2(n_323),
.B(n_347),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_426),
.A2(n_437),
.B(n_442),
.Y(n_471)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_427),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_428),
.A2(n_441),
.B1(n_456),
.B2(n_468),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_429),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_421),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_431),
.B(n_438),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_414),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_376),
.A2(n_336),
.B1(n_362),
.B2(n_374),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_405),
.B(n_326),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_445),
.B(n_465),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_407),
.A2(n_372),
.B(n_370),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_449),
.A2(n_464),
.B(n_416),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_419),
.A2(n_334),
.B1(n_370),
.B2(n_355),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_451),
.A2(n_422),
.B1(n_399),
.B2(n_397),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_415),
.A2(n_334),
.B1(n_355),
.B2(n_352),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_398),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_458),
.B(n_396),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_398),
.B(n_329),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_460),
.B(n_462),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_384),
.B(n_329),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_387),
.A2(n_361),
.B(n_363),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_378),
.B(n_361),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_403),
.B(n_321),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_466),
.B(n_393),
.C(n_380),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_395),
.B(n_324),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_467),
.B(n_377),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_388),
.A2(n_352),
.B1(n_354),
.B2(n_312),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_457),
.A2(n_426),
.B1(n_433),
.B2(n_437),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_469),
.A2(n_490),
.B1(n_495),
.B2(n_466),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_437),
.A2(n_379),
.B(n_417),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_473),
.A2(n_455),
.B(n_430),
.Y(n_508)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_465),
.Y(n_475)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_475),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_477),
.B(n_485),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_454),
.B(n_383),
.Y(n_478)
);

INVxp33_ASAP7_75t_L g517 ( 
.A(n_478),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_467),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_479),
.A2(n_484),
.B1(n_486),
.B2(n_487),
.Y(n_528)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_448),
.Y(n_480)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_480),
.Y(n_521)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_448),
.Y(n_481)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_481),
.Y(n_536)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_452),
.Y(n_482)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_482),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_483),
.A2(n_498),
.B(n_459),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_431),
.B(n_377),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_457),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_452),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_449),
.B(n_404),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_488),
.B(n_489),
.Y(n_531)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_430),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_457),
.A2(n_396),
.B1(n_409),
.B2(n_379),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_445),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_491),
.B(n_499),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_492),
.B(n_504),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_494),
.B(n_506),
.C(n_443),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_458),
.A2(n_400),
.B1(n_406),
.B2(n_424),
.Y(n_495)
);

AOI21xp33_ASAP7_75t_L g497 ( 
.A1(n_442),
.A2(n_417),
.B(n_413),
.Y(n_497)
);

AOI21xp33_ASAP7_75t_L g546 ( 
.A1(n_497),
.A2(n_503),
.B(n_447),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_457),
.A2(n_391),
.B(n_412),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_430),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_432),
.B(n_381),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_500),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_432),
.B(n_382),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_501),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_460),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_502),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_434),
.B(n_324),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_430),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_434),
.B(n_436),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_505),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_461),
.B(n_348),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_435),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_507),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_508),
.B(n_519),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_473),
.A2(n_455),
.B(n_459),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_511),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_512),
.B(n_523),
.C(n_527),
.Y(n_554)
);

CKINVDCx14_ASAP7_75t_R g563 ( 
.A(n_514),
.Y(n_563)
);

FAx1_ASAP7_75t_SL g516 ( 
.A(n_469),
.B(n_461),
.CI(n_446),
.CON(n_516),
.SN(n_516)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_516),
.B(n_546),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_SL g518 ( 
.A(n_506),
.B(n_453),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_SL g573 ( 
.A(n_518),
.B(n_483),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_470),
.A2(n_441),
.B1(n_433),
.B2(n_428),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_522),
.B(n_530),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_506),
.B(n_453),
.C(n_494),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_471),
.A2(n_464),
.B(n_429),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_524),
.B(n_525),
.Y(n_553)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_471),
.A2(n_441),
.B(n_439),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_496),
.A2(n_446),
.B1(n_451),
.B2(n_439),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_526),
.A2(n_529),
.B1(n_532),
.B2(n_538),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_494),
.B(n_453),
.C(n_443),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_496),
.A2(n_436),
.B1(n_435),
.B2(n_462),
.Y(n_529)
);

CKINVDCx16_ASAP7_75t_R g530 ( 
.A(n_472),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_496),
.A2(n_456),
.B1(n_468),
.B2(n_440),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_495),
.B(n_443),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_535),
.B(n_537),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_488),
.B(n_461),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_469),
.A2(n_490),
.B1(n_486),
.B2(n_502),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_477),
.A2(n_440),
.B1(n_427),
.B2(n_450),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_539),
.A2(n_541),
.B1(n_475),
.B2(n_479),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_500),
.B(n_466),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_540),
.B(n_484),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_490),
.A2(n_456),
.B1(n_450),
.B2(n_438),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_498),
.B(n_348),
.C(n_359),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_543),
.B(n_473),
.C(n_498),
.Y(n_572)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_534),
.Y(n_547)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_547),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_542),
.B(n_472),
.Y(n_549)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_549),
.Y(n_612)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_534),
.Y(n_550)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_550),
.Y(n_598)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_515),
.Y(n_552)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_552),
.Y(n_602)
);

XOR2xp5_ASAP7_75t_L g583 ( 
.A(n_556),
.B(n_573),
.Y(n_583)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_521),
.Y(n_557)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_557),
.Y(n_606)
);

FAx1_ASAP7_75t_L g558 ( 
.A(n_516),
.B(n_471),
.CI(n_497),
.CON(n_558),
.SN(n_558)
);

OAI21xp5_ASAP7_75t_SL g590 ( 
.A1(n_558),
.A2(n_574),
.B(n_514),
.Y(n_590)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_515),
.Y(n_559)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_559),
.Y(n_608)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_521),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_561),
.B(n_562),
.Y(n_596)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_536),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_531),
.Y(n_564)
);

CKINVDCx14_ASAP7_75t_R g587 ( 
.A(n_564),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_508),
.B(n_504),
.Y(n_565)
);

INVxp67_ASAP7_75t_L g592 ( 
.A(n_565),
.Y(n_592)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_539),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_566),
.B(n_567),
.Y(n_610)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_536),
.Y(n_567)
);

CKINVDCx14_ASAP7_75t_R g568 ( 
.A(n_531),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_568),
.A2(n_570),
.B(n_581),
.Y(n_605)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_545),
.Y(n_569)
);

BUFx24_ASAP7_75t_SL g603 ( 
.A(n_569),
.Y(n_603)
);

INVx13_ASAP7_75t_L g570 ( 
.A(n_544),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_572),
.B(n_575),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_509),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_545),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_517),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_576),
.A2(n_578),
.B1(n_513),
.B2(n_533),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_523),
.B(n_507),
.C(n_478),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_577),
.B(n_579),
.C(n_560),
.Y(n_586)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_528),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_527),
.B(n_491),
.C(n_483),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g581 ( 
.A(n_513),
.B(n_493),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_SL g584 ( 
.A1(n_582),
.A2(n_541),
.B1(n_520),
.B2(n_538),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_584),
.A2(n_600),
.B1(n_563),
.B2(n_551),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_585),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_586),
.B(n_593),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_571),
.A2(n_529),
.B1(n_526),
.B2(n_520),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_588),
.A2(n_599),
.B1(n_601),
.B2(n_547),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_SL g631 ( 
.A1(n_590),
.A2(n_604),
.B(n_555),
.Y(n_631)
);

XOR2xp5_ASAP7_75t_L g591 ( 
.A(n_560),
.B(n_512),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_591),
.B(n_595),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_554),
.B(n_535),
.C(n_518),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g595 ( 
.A(n_577),
.B(n_579),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g597 ( 
.A(n_554),
.B(n_537),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g632 ( 
.A(n_597),
.B(n_591),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_571),
.A2(n_510),
.B1(n_532),
.B2(n_524),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_SL g600 ( 
.A1(n_582),
.A2(n_519),
.B1(n_525),
.B2(n_522),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_578),
.A2(n_544),
.B1(n_533),
.B2(n_511),
.Y(n_601)
);

OAI21xp5_ASAP7_75t_L g604 ( 
.A1(n_555),
.A2(n_533),
.B(n_476),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_572),
.B(n_540),
.C(n_543),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_607),
.B(n_609),
.C(n_611),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_580),
.B(n_499),
.C(n_489),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_580),
.B(n_516),
.C(n_505),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_SL g613 ( 
.A(n_603),
.B(n_493),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_613),
.B(n_619),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_SL g650 ( 
.A1(n_614),
.A2(n_626),
.B1(n_629),
.B2(n_633),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_616),
.A2(n_618),
.B1(n_620),
.B2(n_623),
.Y(n_643)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_596),
.Y(n_617)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_617),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_612),
.A2(n_581),
.B1(n_549),
.B2(n_548),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_605),
.Y(n_619)
);

CKINVDCx14_ASAP7_75t_R g620 ( 
.A(n_590),
.Y(n_620)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_605),
.Y(n_622)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_622),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_SL g623 ( 
.A1(n_599),
.A2(n_551),
.B1(n_558),
.B2(n_564),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_606),
.Y(n_624)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_624),
.Y(n_657)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_589),
.Y(n_625)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_625),
.Y(n_652)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_585),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_SL g627 ( 
.A1(n_588),
.A2(n_601),
.B1(n_610),
.B2(n_551),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_627),
.A2(n_636),
.B1(n_638),
.B2(n_592),
.Y(n_644)
);

XNOR2x2_ASAP7_75t_SL g628 ( 
.A(n_604),
.B(n_558),
.Y(n_628)
);

XNOR2xp5_ASAP7_75t_L g646 ( 
.A(n_628),
.B(n_600),
.Y(n_646)
);

CKINVDCx14_ASAP7_75t_R g629 ( 
.A(n_609),
.Y(n_629)
);

OAI21xp5_ASAP7_75t_L g649 ( 
.A1(n_631),
.A2(n_637),
.B(n_583),
.Y(n_649)
);

NOR2xp67_ASAP7_75t_SL g654 ( 
.A(n_632),
.B(n_573),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_584),
.A2(n_553),
.B1(n_565),
.B2(n_476),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_587),
.B(n_557),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_635),
.A2(n_562),
.B(n_501),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_SL g636 ( 
.A1(n_598),
.A2(n_553),
.B1(n_565),
.B2(n_570),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_592),
.A2(n_553),
.B(n_556),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_SL g638 ( 
.A1(n_602),
.A2(n_474),
.B1(n_485),
.B2(n_561),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g639 ( 
.A(n_621),
.B(n_595),
.C(n_597),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_639),
.B(n_642),
.Y(n_674)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_621),
.B(n_586),
.C(n_593),
.Y(n_642)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_644),
.Y(n_668)
);

XOR2xp5_ASAP7_75t_L g645 ( 
.A(n_614),
.B(n_594),
.Y(n_645)
);

XNOR2xp5_ASAP7_75t_L g670 ( 
.A(n_645),
.B(n_646),
.Y(n_670)
);

XNOR2xp5_ASAP7_75t_L g647 ( 
.A(n_628),
.B(n_594),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_647),
.B(n_655),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_622),
.A2(n_608),
.B1(n_611),
.B2(n_607),
.Y(n_648)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_648),
.Y(n_673)
);

XOR2xp5_ASAP7_75t_L g662 ( 
.A(n_649),
.B(n_654),
.Y(n_662)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_651),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_627),
.A2(n_474),
.B1(n_583),
.B2(n_492),
.Y(n_653)
);

INVxp67_ASAP7_75t_L g664 ( 
.A(n_653),
.Y(n_664)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_632),
.B(n_487),
.C(n_482),
.Y(n_655)
);

MAJIxp5_ASAP7_75t_L g658 ( 
.A(n_634),
.B(n_480),
.C(n_481),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_658),
.B(n_659),
.Y(n_666)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_630),
.B(n_615),
.C(n_626),
.Y(n_659)
);

MAJIxp5_ASAP7_75t_L g660 ( 
.A(n_630),
.B(n_444),
.C(n_503),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_660),
.B(n_447),
.Y(n_676)
);

AOI22x1_ASAP7_75t_SL g661 ( 
.A1(n_650),
.A2(n_623),
.B1(n_615),
.B2(n_636),
.Y(n_661)
);

MAJx2_ASAP7_75t_L g693 ( 
.A(n_661),
.B(n_354),
.C(n_341),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_SL g663 ( 
.A1(n_641),
.A2(n_617),
.B1(n_625),
.B2(n_635),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_663),
.A2(n_677),
.B(n_660),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_SL g665 ( 
.A(n_640),
.B(n_648),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_665),
.B(n_675),
.Y(n_686)
);

MAJIxp5_ASAP7_75t_L g667 ( 
.A(n_659),
.B(n_633),
.C(n_631),
.Y(n_667)
);

MAJIxp5_ASAP7_75t_L g680 ( 
.A(n_667),
.B(n_669),
.C(n_672),
.Y(n_680)
);

MAJIxp5_ASAP7_75t_L g669 ( 
.A(n_639),
.B(n_637),
.C(n_638),
.Y(n_669)
);

XOR2xp5_ASAP7_75t_L g671 ( 
.A(n_655),
.B(n_624),
.Y(n_671)
);

XNOR2xp5_ASAP7_75t_L g683 ( 
.A(n_671),
.B(n_653),
.Y(n_683)
);

MAJIxp5_ASAP7_75t_L g672 ( 
.A(n_642),
.B(n_444),
.C(n_463),
.Y(n_672)
);

XNOR2xp5_ASAP7_75t_L g675 ( 
.A(n_658),
.B(n_349),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_676),
.A2(n_657),
.B1(n_652),
.B2(n_647),
.Y(n_684)
);

MAJIxp5_ASAP7_75t_L g677 ( 
.A(n_645),
.B(n_463),
.C(n_322),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_SL g681 ( 
.A1(n_674),
.A2(n_643),
.B(n_656),
.Y(n_681)
);

OAI21xp5_ASAP7_75t_SL g694 ( 
.A1(n_681),
.A2(n_689),
.B(n_664),
.Y(n_694)
);

OAI21xp5_ASAP7_75t_L g682 ( 
.A1(n_673),
.A2(n_644),
.B(n_649),
.Y(n_682)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_682),
.Y(n_697)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_683),
.Y(n_702)
);

XNOR2xp5_ASAP7_75t_L g701 ( 
.A(n_684),
.B(n_687),
.Y(n_701)
);

XOR2xp5_ASAP7_75t_L g695 ( 
.A(n_685),
.B(n_691),
.Y(n_695)
);

XOR2xp5_ASAP7_75t_L g687 ( 
.A(n_670),
.B(n_646),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_667),
.B(n_463),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_SL g698 ( 
.A(n_688),
.B(n_692),
.Y(n_698)
);

OAI21xp5_ASAP7_75t_SL g689 ( 
.A1(n_666),
.A2(n_349),
.B(n_411),
.Y(n_689)
);

AO21x1_ASAP7_75t_L g690 ( 
.A1(n_668),
.A2(n_322),
.B(n_359),
.Y(n_690)
);

OAI21xp33_ASAP7_75t_L g700 ( 
.A1(n_690),
.A2(n_672),
.B(n_664),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_678),
.A2(n_352),
.B1(n_341),
.B2(n_312),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_679),
.B(n_312),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_693),
.B(n_677),
.Y(n_699)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_694),
.Y(n_710)
);

MAJIxp5_ASAP7_75t_L g696 ( 
.A(n_680),
.B(n_671),
.C(n_669),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_696),
.B(n_699),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_700),
.B(n_662),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_680),
.B(n_670),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_703),
.B(n_686),
.Y(n_707)
);

OAI21x1_ASAP7_75t_L g704 ( 
.A1(n_697),
.A2(n_682),
.B(n_661),
.Y(n_704)
);

AOI21x1_ASAP7_75t_L g713 ( 
.A1(n_704),
.A2(n_709),
.B(n_693),
.Y(n_713)
);

XNOR2xp5_ASAP7_75t_L g706 ( 
.A(n_696),
.B(n_687),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_706),
.B(n_707),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_701),
.B(n_683),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_708),
.A2(n_695),
.B(n_700),
.Y(n_714)
);

OAI21xp5_ASAP7_75t_SL g712 ( 
.A1(n_710),
.A2(n_702),
.B(n_701),
.Y(n_712)
);

NOR3xp33_ASAP7_75t_L g716 ( 
.A(n_712),
.B(n_713),
.C(n_714),
.Y(n_716)
);

A2O1A1Ixp33_ASAP7_75t_L g715 ( 
.A1(n_711),
.A2(n_705),
.B(n_709),
.C(n_690),
.Y(n_715)
);

INVxp33_ASAP7_75t_L g717 ( 
.A(n_715),
.Y(n_717)
);

MAJIxp5_ASAP7_75t_L g718 ( 
.A(n_717),
.B(n_716),
.C(n_695),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_718),
.Y(n_719)
);

MAJIxp5_ASAP7_75t_L g720 ( 
.A(n_719),
.B(n_662),
.C(n_698),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_720),
.A2(n_691),
.B(n_354),
.Y(n_721)
);


endmodule