module fake_jpeg_812_n_540 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_540);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_540;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_16),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_53),
.B(n_70),
.Y(n_134)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx5_ASAP7_75t_SL g159 ( 
.A(n_55),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_21),
.B(n_52),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_66),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_58),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_59),
.B(n_85),
.Y(n_113)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_61),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_62),
.Y(n_155)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_63),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_64),
.Y(n_136)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g109 ( 
.A(n_65),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_1),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_1),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_67),
.B(n_78),
.Y(n_131)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_47),
.Y(n_68)
);

INVx5_ASAP7_75t_SL g161 ( 
.A(n_68),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_42),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_72),
.Y(n_140)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_75),
.Y(n_156)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_76),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_48),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_77),
.B(n_83),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_21),
.B(n_17),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

BUFx24_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_80),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_23),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_84),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_23),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_52),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_87),
.B(n_88),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_47),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_34),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_90),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_39),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_47),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_20),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_24),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_96),
.B(n_33),
.Y(n_138)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_99),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_39),
.B(n_44),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_101),
.B(n_102),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_45),
.B(n_17),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_28),
.Y(n_103)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_28),
.B(n_17),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_104),
.B(n_32),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_55),
.A2(n_20),
.B1(n_37),
.B2(n_36),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_111),
.A2(n_112),
.B1(n_114),
.B2(n_120),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_55),
.A2(n_20),
.B1(n_37),
.B2(n_36),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_66),
.A2(n_33),
.B1(n_43),
.B2(n_41),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_83),
.B(n_24),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_118),
.B(n_147),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_119),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_67),
.A2(n_35),
.B1(n_50),
.B2(n_31),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_35),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_121),
.B(n_150),
.Y(n_209)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_123),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_54),
.B(n_50),
.C(n_31),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_133),
.B(n_19),
.Y(n_231)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_137),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_138),
.B(n_160),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_77),
.A2(n_40),
.B1(n_43),
.B2(n_41),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_141),
.A2(n_143),
.B1(n_158),
.B2(n_80),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_53),
.A2(n_26),
.B1(n_40),
.B2(n_32),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_70),
.A2(n_26),
.B1(n_22),
.B2(n_46),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_149),
.A2(n_95),
.B1(n_99),
.B2(n_100),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_87),
.B(n_16),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_65),
.A2(n_22),
.B1(n_34),
.B2(n_46),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_151),
.A2(n_164),
.B1(n_80),
.B2(n_64),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_75),
.A2(n_81),
.B1(n_69),
.B2(n_56),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_68),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_76),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_79),
.A2(n_46),
.B1(n_19),
.B2(n_18),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_60),
.Y(n_165)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_165),
.Y(n_199)
);

AOI21xp33_ASAP7_75t_L g168 ( 
.A1(n_96),
.A2(n_15),
.B(n_14),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_168),
.B(n_170),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_88),
.B(n_15),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_94),
.Y(n_198)
);

AOI21xp33_ASAP7_75t_L g170 ( 
.A1(n_98),
.A2(n_46),
.B(n_19),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_163),
.Y(n_171)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_171),
.Y(n_238)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_117),
.Y(n_172)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_172),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_173),
.A2(n_210),
.B1(n_136),
.B2(n_115),
.Y(n_250)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_174),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_131),
.B(n_86),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_175),
.B(n_182),
.Y(n_240)
);

OAI21x1_ASAP7_75t_SL g262 ( 
.A1(n_177),
.A2(n_181),
.B(n_183),
.Y(n_262)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_178),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_127),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_179),
.B(n_196),
.Y(n_236)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_180),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_119),
.B(n_97),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_105),
.B(n_71),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_121),
.B(n_63),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_62),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_184),
.B(n_185),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_141),
.B(n_61),
.Y(n_185)
);

INVx6_ASAP7_75t_SL g186 ( 
.A(n_161),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_186),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_58),
.Y(n_187)
);

NAND2x1_ASAP7_75t_L g282 ( 
.A(n_187),
.B(n_195),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_116),
.B(n_58),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_190),
.B(n_191),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_130),
.B(n_93),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_120),
.B(n_113),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_192),
.B(n_126),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_193),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_153),
.B(n_93),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_129),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_198),
.B(n_224),
.Y(n_263)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_109),
.Y(n_201)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_110),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_202),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_203),
.Y(n_285)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_109),
.Y(n_204)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_204),
.Y(n_253)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_142),
.Y(n_205)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_205),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_161),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_206),
.B(n_208),
.Y(n_247)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_117),
.Y(n_207)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_207),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_167),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_149),
.A2(n_82),
.B1(n_84),
.B2(n_46),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_148),
.Y(n_211)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_164),
.A2(n_151),
.B1(n_112),
.B2(n_111),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_212),
.A2(n_232),
.B1(n_5),
.B2(n_6),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_144),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_213),
.Y(n_271)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_108),
.Y(n_214)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_214),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_132),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_216),
.B(n_223),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_128),
.Y(n_217)
);

INVx11_ASAP7_75t_L g291 ( 
.A(n_217),
.Y(n_291)
);

INVx13_ASAP7_75t_L g218 ( 
.A(n_159),
.Y(n_218)
);

INVx11_ASAP7_75t_L g249 ( 
.A(n_218),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_128),
.Y(n_219)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_219),
.Y(n_273)
);

BUFx12_ASAP7_75t_L g220 ( 
.A(n_159),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_108),
.Y(n_222)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_222),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_144),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_132),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_126),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_225),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_157),
.A2(n_91),
.B1(n_74),
.B2(n_73),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_226),
.Y(n_270)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_107),
.Y(n_227)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_227),
.Y(n_286)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_107),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_229),
.Y(n_255)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_157),
.Y(n_229)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_110),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_230),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_152),
.C(n_155),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_156),
.A2(n_94),
.B1(n_18),
.B2(n_49),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_124),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_122),
.Y(n_246)
);

MAJx2_ASAP7_75t_L g235 ( 
.A(n_175),
.B(n_156),
.C(n_145),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_235),
.B(n_244),
.Y(n_320)
);

BUFx24_ASAP7_75t_SL g242 ( 
.A(n_194),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_242),
.B(n_266),
.Y(n_305)
);

INVxp33_ASAP7_75t_L g314 ( 
.A(n_246),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_188),
.A2(n_136),
.B(n_122),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_248),
.A2(n_261),
.B(n_207),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_250),
.A2(n_269),
.B1(n_222),
.B2(n_214),
.Y(n_304)
);

NOR2x1_ASAP7_75t_R g252 ( 
.A(n_174),
.B(n_215),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_252),
.Y(n_296)
);

OAI211xp5_ASAP7_75t_L g338 ( 
.A1(n_259),
.A2(n_287),
.B(n_6),
.C(n_7),
.Y(n_338)
);

OR2x2_ASAP7_75t_SL g260 ( 
.A(n_231),
.B(n_106),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_260),
.Y(n_301)
);

O2A1O1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_185),
.A2(n_155),
.B(n_115),
.C(n_106),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_197),
.B(n_154),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_182),
.B(n_135),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_267),
.B(n_275),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_173),
.A2(n_135),
.B1(n_125),
.B2(n_166),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_184),
.B(n_125),
.C(n_154),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_277),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_215),
.B(n_166),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_180),
.B(n_1),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_276),
.B(n_280),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_221),
.B(n_18),
.C(n_2),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g278 ( 
.A(n_192),
.B(n_186),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_278),
.B(n_218),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_183),
.B(n_1),
.C(n_2),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_279),
.B(n_195),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_209),
.B(n_2),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_190),
.B(n_3),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_281),
.B(n_283),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_191),
.B(n_4),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_171),
.B(n_176),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_284),
.B(n_211),
.Y(n_328)
);

OAI21xp33_ASAP7_75t_SL g337 ( 
.A1(n_288),
.A2(n_258),
.B(n_270),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_255),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_293),
.B(n_303),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_278),
.A2(n_209),
.B(n_183),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_295),
.A2(n_298),
.B(n_299),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_181),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_297),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_275),
.A2(n_181),
.B(n_200),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_240),
.A2(n_187),
.B(n_195),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_284),
.Y(n_300)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_300),
.Y(n_366)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_238),
.Y(n_302)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_302),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_304),
.A2(n_324),
.B1(n_326),
.B2(n_268),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_240),
.B(n_178),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_306),
.B(n_328),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_263),
.B(n_236),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_308),
.B(n_317),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_282),
.B(n_187),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_310),
.Y(n_346)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_238),
.Y(n_311)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_311),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_255),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_313),
.B(n_318),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_315),
.A2(n_325),
.B(n_338),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_316),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_265),
.B(n_189),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_255),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_247),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_319),
.B(n_327),
.Y(n_379)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_289),
.Y(n_321)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_321),
.Y(n_376)
);

AND2x2_ASAP7_75t_SL g322 ( 
.A(n_243),
.B(n_199),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_322),
.B(n_277),
.Y(n_364)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_289),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_323),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_241),
.A2(n_228),
.B1(n_227),
.B2(n_199),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_259),
.A2(n_229),
.B(n_233),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_241),
.A2(n_230),
.B1(n_202),
.B2(n_225),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_271),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_248),
.A2(n_172),
.B1(n_203),
.B2(n_213),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_329),
.A2(n_337),
.B1(n_270),
.B2(n_256),
.Y(n_343)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_286),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_330),
.B(n_331),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_267),
.B(n_219),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_235),
.B(n_217),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_332),
.B(n_334),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_244),
.B(n_220),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_333),
.B(n_260),
.C(n_282),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_243),
.B(n_5),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_251),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_335),
.B(n_339),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_265),
.B(n_220),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_336),
.B(n_340),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_272),
.B(n_7),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_258),
.B(n_7),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_273),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_341),
.Y(n_349)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_274),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_251),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_343),
.A2(n_360),
.B(n_310),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_347),
.B(n_355),
.C(n_363),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_L g412 ( 
.A1(n_353),
.A2(n_356),
.B1(n_359),
.B2(n_249),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_320),
.B(n_252),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_319),
.A2(n_287),
.B1(n_288),
.B2(n_262),
.Y(n_356)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_357),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_325),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_358),
.B(n_378),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_300),
.A2(n_316),
.B1(n_296),
.B2(n_304),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_332),
.A2(n_254),
.B(n_237),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_309),
.A2(n_283),
.B1(n_281),
.B2(n_261),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_361),
.A2(n_380),
.B1(n_377),
.B2(n_354),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_320),
.B(n_253),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_364),
.B(n_330),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_333),
.B(n_294),
.C(n_301),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_365),
.B(n_381),
.C(n_382),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_306),
.B(n_279),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_369),
.B(n_372),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_309),
.B(n_245),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_301),
.A2(n_245),
.B1(n_264),
.B2(n_292),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_373),
.A2(n_313),
.B1(n_318),
.B2(n_293),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_299),
.A2(n_237),
.B(n_264),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_375),
.A2(n_346),
.B(n_367),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_341),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_322),
.A2(n_290),
.B1(n_292),
.B2(n_257),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_294),
.B(n_239),
.C(n_234),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_296),
.B(n_297),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_312),
.B(n_234),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_384),
.B(n_303),
.C(n_302),
.Y(n_403)
);

INVxp33_ASAP7_75t_L g429 ( 
.A(n_385),
.Y(n_429)
);

NAND2x1_ASAP7_75t_SL g387 ( 
.A(n_350),
.B(n_346),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_387),
.A2(n_411),
.B(n_416),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_366),
.A2(n_324),
.B1(n_326),
.B2(n_331),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_388),
.A2(n_390),
.B1(n_392),
.B2(n_395),
.Y(n_434)
);

CKINVDCx14_ASAP7_75t_R g389 ( 
.A(n_348),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_389),
.B(n_391),
.Y(n_449)
);

AOI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_350),
.A2(n_329),
.B1(n_327),
.B2(n_310),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_357),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_366),
.A2(n_334),
.B1(n_298),
.B2(n_339),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_372),
.A2(n_322),
.B1(n_314),
.B2(n_295),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_393),
.A2(n_402),
.B1(n_361),
.B2(n_367),
.Y(n_425)
);

AO21x1_ASAP7_75t_L g440 ( 
.A1(n_394),
.A2(n_419),
.B(n_348),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_351),
.A2(n_328),
.B1(n_297),
.B2(n_312),
.Y(n_395)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_371),
.Y(n_397)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_397),
.Y(n_420)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_371),
.Y(n_401)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_401),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_351),
.A2(n_323),
.B1(n_321),
.B2(n_311),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_403),
.B(n_399),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_370),
.B(n_307),
.Y(n_404)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_404),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_383),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_405),
.B(n_417),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_383),
.Y(n_406)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_406),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_407),
.B(n_368),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_365),
.B(n_305),
.C(n_342),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_408),
.B(n_410),
.C(n_347),
.Y(n_427)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_374),
.Y(n_409)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_409),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_363),
.B(n_335),
.C(n_285),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_412),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_362),
.B(n_285),
.Y(n_413)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_413),
.Y(n_431)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_374),
.Y(n_414)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_414),
.Y(n_433)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_376),
.Y(n_415)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_415),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_375),
.A2(n_249),
.B(n_291),
.Y(n_416)
);

OA21x2_ASAP7_75t_L g417 ( 
.A1(n_343),
.A2(n_291),
.B(n_290),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_379),
.B(n_9),
.Y(n_418)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_418),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_387),
.A2(n_344),
.B(n_360),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_421),
.A2(n_440),
.B(n_447),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_425),
.A2(n_432),
.B1(n_436),
.B2(n_443),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_427),
.B(n_438),
.C(n_442),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_430),
.B(n_439),
.Y(n_453)
);

AOI22x1_ASAP7_75t_L g432 ( 
.A1(n_385),
.A2(n_380),
.B1(n_345),
.B2(n_344),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_419),
.A2(n_345),
.B1(n_352),
.B2(n_382),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_400),
.B(n_381),
.C(n_355),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_400),
.B(n_364),
.C(n_384),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_391),
.A2(n_352),
.B1(n_354),
.B2(n_376),
.Y(n_443)
);

AOI21xp33_ASAP7_75t_L g444 ( 
.A1(n_411),
.A2(n_369),
.B(n_373),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_444),
.B(n_394),
.Y(n_452)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_398),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_445),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_399),
.B(n_349),
.C(n_10),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_446),
.B(n_392),
.C(n_395),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_386),
.A2(n_10),
.B1(n_12),
.B2(n_393),
.Y(n_447)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_445),
.Y(n_450)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_450),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_452),
.B(n_455),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_431),
.B(n_398),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_454),
.B(n_473),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_423),
.B(n_408),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_430),
.B(n_407),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_SL g478 ( 
.A(n_458),
.B(n_461),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_443),
.B(n_402),
.Y(n_459)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_459),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_449),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_460),
.B(n_470),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_442),
.B(n_438),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_439),
.B(n_403),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_462),
.B(n_467),
.C(n_469),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_435),
.A2(n_421),
.B(n_429),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_464),
.A2(n_448),
.B(n_432),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_465),
.B(n_466),
.Y(n_485)
);

XNOR2x1_ASAP7_75t_L g466 ( 
.A(n_434),
.B(n_410),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_427),
.B(n_387),
.C(n_396),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_429),
.B(n_396),
.Y(n_468)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_468),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_436),
.B(n_416),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_424),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_425),
.A2(n_417),
.B1(n_405),
.B2(n_409),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_471),
.A2(n_448),
.B1(n_428),
.B2(n_388),
.Y(n_489)
);

NAND2xp33_ASAP7_75t_SL g472 ( 
.A(n_435),
.B(n_401),
.Y(n_472)
);

OAI221xp5_ASAP7_75t_L g476 ( 
.A1(n_472),
.A2(n_440),
.B1(n_417),
.B2(n_428),
.C(n_432),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_441),
.B(n_397),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_476),
.A2(n_482),
.B(n_491),
.Y(n_497)
);

INVx13_ASAP7_75t_L g479 ( 
.A(n_457),
.Y(n_479)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_479),
.Y(n_501)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_468),
.Y(n_484)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_484),
.Y(n_507)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_450),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_486),
.B(n_471),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_461),
.B(n_446),
.C(n_448),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_488),
.B(n_492),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_489),
.A2(n_490),
.B1(n_459),
.B2(n_463),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_451),
.A2(n_420),
.B1(n_433),
.B2(n_426),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_464),
.A2(n_422),
.B(n_437),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_456),
.B(n_414),
.C(n_415),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_467),
.B(n_10),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_487),
.B(n_465),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_494),
.B(n_495),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_480),
.B(n_487),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_482),
.A2(n_463),
.B(n_469),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_496),
.A2(n_474),
.B(n_486),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_492),
.B(n_460),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_499),
.B(n_500),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_493),
.B(n_470),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_488),
.B(n_456),
.C(n_458),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_502),
.B(n_503),
.C(n_478),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_481),
.B(n_466),
.C(n_453),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_504),
.B(n_505),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_SL g505 ( 
.A(n_481),
.B(n_453),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_506),
.A2(n_475),
.B1(n_483),
.B2(n_491),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_497),
.A2(n_489),
.B1(n_483),
.B2(n_484),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_508),
.B(n_510),
.Y(n_519)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_509),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_497),
.A2(n_475),
.B1(n_477),
.B2(n_490),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_511),
.A2(n_496),
.B(n_501),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_503),
.B(n_485),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_512),
.B(n_514),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_507),
.A2(n_474),
.B1(n_479),
.B2(n_462),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_513),
.B(n_514),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_498),
.B(n_478),
.C(n_502),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_516),
.B(n_505),
.C(n_506),
.Y(n_521)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_520),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_521),
.B(n_523),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_517),
.B(n_504),
.Y(n_523)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_524),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_515),
.B(n_518),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_525),
.B(n_516),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_530),
.B(n_524),
.Y(n_532)
);

NOR2xp67_ASAP7_75t_SL g531 ( 
.A(n_521),
.B(n_512),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_531),
.B(n_526),
.C(n_519),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_532),
.B(n_533),
.C(n_534),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_528),
.B(n_522),
.C(n_513),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_532),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_536),
.A2(n_529),
.B(n_527),
.Y(n_537)
);

AO21x1_ASAP7_75t_L g538 ( 
.A1(n_537),
.A2(n_509),
.B(n_518),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_538),
.B(n_535),
.C(n_508),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_539),
.B(n_510),
.Y(n_540)
);


endmodule