module fake_netlist_6_4305_n_1217 (n_52, n_1, n_91, n_326, n_256, n_209, n_63, n_223, n_278, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_56, n_119, n_235, n_147, n_191, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_53, n_44, n_232, n_16, n_163, n_46, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_323, n_152, n_92, n_321, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_325, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_231, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_215, n_178, n_247, n_225, n_308, n_309, n_317, n_149, n_90, n_24, n_54, n_328, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_315, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1217);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_323;
input n_152;
input n_92;
input n_321;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_325;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_231;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_317;
input n_149;
input n_90;
input n_24;
input n_54;
input n_328;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1217;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_801;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_881;
wire n_1199;
wire n_875;
wire n_465;
wire n_367;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_1189;
wire n_1079;
wire n_341;
wire n_362;
wire n_1212;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1052;
wire n_419;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_595;
wire n_627;
wire n_1203;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_1208;
wire n_798;
wire n_1164;
wire n_509;
wire n_1209;
wire n_575;
wire n_368;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_1151;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_1214;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_1204;
wire n_1160;
wire n_883;
wire n_557;
wire n_823;
wire n_1132;
wire n_643;
wire n_349;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_807;
wire n_1036;
wire n_739;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_1138;
wire n_893;
wire n_925;
wire n_485;
wire n_1101;
wire n_1026;
wire n_443;
wire n_1099;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_935;
wire n_1192;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_1127;
wire n_1095;
wire n_573;
wire n_769;
wire n_639;
wire n_676;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_597;
wire n_685;
wire n_832;
wire n_353;
wire n_1187;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_1139;
wire n_718;
wire n_517;
wire n_1018;
wire n_1172;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_1206;
wire n_621;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_544;
wire n_372;
wire n_468;
wire n_901;
wire n_504;
wire n_923;
wire n_1140;
wire n_378;
wire n_413;
wire n_1196;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_601;
wire n_375;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_1147;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_1143;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_1182;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_761;
wire n_428;
wire n_785;
wire n_746;
wire n_1205;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_1163;
wire n_1173;
wire n_1180;
wire n_1116;
wire n_611;
wire n_943;
wire n_1168;
wire n_491;
wire n_1216;
wire n_878;
wire n_656;
wire n_843;
wire n_772;
wire n_989;
wire n_1174;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_1094;
wire n_1176;
wire n_1190;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_1213;
wire n_638;
wire n_1181;
wire n_910;
wire n_1211;
wire n_486;
wire n_947;
wire n_381;
wire n_911;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_809;
wire n_1043;
wire n_1011;
wire n_926;
wire n_927;
wire n_1215;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_1084;
wire n_1171;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_526;
wire n_1109;
wire n_921;
wire n_712;
wire n_1183;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_1193;
wire n_1148;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_1161;
wire n_458;
wire n_1070;
wire n_1085;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_1145;
wire n_330;
wire n_771;
wire n_1121;
wire n_1152;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_492;
wire n_972;
wire n_699;
wire n_551;
wire n_456;
wire n_1149;
wire n_564;
wire n_1178;
wire n_451;
wire n_624;
wire n_1184;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_686;
wire n_796;
wire n_1041;
wire n_757;
wire n_594;
wire n_565;
wire n_719;
wire n_1195;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1186;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_829;
wire n_1156;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_1142;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_1201;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_645;
wire n_331;
wire n_916;
wire n_1078;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_608;
wire n_474;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_543;
wire n_1144;
wire n_889;
wire n_357;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_1162;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_600;
wire n_464;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_959;
wire n_879;
wire n_1198;
wire n_584;
wire n_1110;
wire n_399;
wire n_979;
wire n_548;
wire n_905;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_993;
wire n_345;
wire n_409;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_1155;
wire n_756;
wire n_547;
wire n_537;
wire n_558;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_1194;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_1146;
wire n_1141;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_1158;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_1125;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_1159;
wire n_569;
wire n_1092;
wire n_441;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_1207;
wire n_1111;
wire n_511;
wire n_715;
wire n_467;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1106;
wire n_790;
wire n_1055;
wire n_582;
wire n_1167;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_651;
wire n_404;
wire n_439;
wire n_1153;
wire n_518;
wire n_1210;
wire n_679;
wire n_1069;
wire n_1185;
wire n_612;
wire n_453;
wire n_633;
wire n_1170;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_1165;
wire n_426;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_1166;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1131;
wire n_1033;
wire n_502;
wire n_1175;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_834;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1179;
wire n_1169;
wire n_1135;
wire n_1089;
wire n_401;
wire n_743;
wire n_766;
wire n_816;
wire n_1157;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_1188;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_1019;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_438;
wire n_1124;
wire n_339;
wire n_784;
wire n_434;
wire n_515;
wire n_983;
wire n_427;
wire n_1200;
wire n_1059;
wire n_1197;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1154;
wire n_1082;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_457;
wire n_391;
wire n_1098;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_1134;
wire n_1177;
wire n_332;
wire n_891;
wire n_336;
wire n_1150;
wire n_410;
wire n_398;
wire n_1129;
wire n_1191;
wire n_566;
wire n_554;
wire n_602;
wire n_1023;
wire n_1013;
wire n_1076;
wire n_1118;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_12),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_215),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_245),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_269),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_121),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_164),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_248),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_296),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_142),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_187),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_298),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_199),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_249),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_211),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_102),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_326),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_325),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_186),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_231),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_143),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_224),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_144),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_288),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_27),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_127),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_192),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_221),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_317),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_179),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_140),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_181),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_103),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_83),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_307),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_275),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_51),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_290),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_162),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_262),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_312),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_327),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_225),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_66),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_283),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_209),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_226),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_161),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g376 ( 
.A(n_114),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_217),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_126),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_253),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_295),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_158),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_174),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_87),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_223),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_235),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_202),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_282),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_229),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_273),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_255),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_280),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_303),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_292),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_101),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_328),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_203),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_277),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_89),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_299),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_267),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_208),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_155),
.Y(n_402)
);

INVx2_ASAP7_75t_SL g403 ( 
.A(n_210),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_39),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g405 ( 
.A(n_220),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_185),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_10),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_252),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_194),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_15),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_50),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_56),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_149),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_191),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_236),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_131),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_109),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_251),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_132),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_138),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_234),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_243),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_63),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_47),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_133),
.B(n_148),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_261),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_214),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_29),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_169),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_70),
.B(n_117),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_232),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_98),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_313),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_38),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_176),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_287),
.Y(n_436)
);

BUFx10_ASAP7_75t_L g437 ( 
.A(n_154),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_108),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_141),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_159),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_206),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_157),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_81),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_118),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_6),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_38),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_135),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_19),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_59),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_218),
.Y(n_450)
);

NOR2xp67_ASAP7_75t_L g451 ( 
.A(n_30),
.B(n_40),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_319),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_145),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_321),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_247),
.Y(n_455)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_284),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_233),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_304),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_89),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_160),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_52),
.Y(n_461)
);

BUFx8_ASAP7_75t_SL g462 ( 
.A(n_258),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_204),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_198),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g465 ( 
.A(n_30),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_134),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_23),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_173),
.Y(n_468)
);

BUFx10_ASAP7_75t_L g469 ( 
.A(n_83),
.Y(n_469)
);

BUFx10_ASAP7_75t_L g470 ( 
.A(n_266),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_33),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_324),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_182),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_256),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_55),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_34),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_264),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_88),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_289),
.Y(n_479)
);

NOR2xp67_ASAP7_75t_L g480 ( 
.A(n_167),
.B(n_291),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_54),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_115),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_86),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_265),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_90),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_175),
.Y(n_486)
);

BUFx2_ASAP7_75t_L g487 ( 
.A(n_222),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_97),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_124),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_103),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_139),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_136),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_178),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_123),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_240),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_449),
.Y(n_496)
);

AND2x2_ASAP7_75t_SL g497 ( 
.A(n_422),
.B(n_0),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_421),
.Y(n_498)
);

AND2x6_ASAP7_75t_L g499 ( 
.A(n_397),
.B(n_116),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_397),
.A2(n_120),
.B(n_119),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_456),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_386),
.B(n_1),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_332),
.B(n_2),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_421),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_449),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_487),
.B(n_3),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_330),
.B(n_3),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_421),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_386),
.B(n_4),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_364),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_421),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_436),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_436),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_434),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_364),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_436),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_361),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_376),
.B(n_4),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_402),
.B(n_444),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_437),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_371),
.Y(n_521)
);

INVx5_ASAP7_75t_L g522 ( 
.A(n_460),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_469),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_445),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_460),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_445),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_404),
.Y(n_527)
);

OAI22x1_ASAP7_75t_SL g528 ( 
.A1(n_412),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_437),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_402),
.B(n_5),
.Y(n_530)
);

INVx6_ASAP7_75t_L g531 ( 
.A(n_470),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_331),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_424),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_467),
.A2(n_343),
.B1(n_352),
.B2(n_329),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_403),
.B(n_405),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_479),
.B(n_7),
.Y(n_536)
);

NOR2x1_ASAP7_75t_L g537 ( 
.A(n_444),
.B(n_122),
.Y(n_537)
);

OAI21x1_ASAP7_75t_L g538 ( 
.A1(n_333),
.A2(n_128),
.B(n_125),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_428),
.Y(n_539)
);

AOI22x1_ASAP7_75t_SL g540 ( 
.A1(n_412),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_490),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_333),
.B(n_8),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_341),
.B(n_11),
.Y(n_543)
);

OAI22x1_ASAP7_75t_SL g544 ( 
.A1(n_360),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_544)
);

AOI22x1_ASAP7_75t_SL g545 ( 
.A1(n_383),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_341),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_366),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_470),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_366),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_378),
.B(n_14),
.Y(n_550)
);

AOI22x1_ASAP7_75t_SL g551 ( 
.A1(n_394),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_410),
.A2(n_465),
.B1(n_477),
.B2(n_407),
.Y(n_552)
);

INVx5_ASAP7_75t_L g553 ( 
.A(n_462),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_378),
.A2(n_130),
.B(n_129),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_337),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_395),
.B(n_16),
.Y(n_556)
);

AND2x6_ASAP7_75t_L g557 ( 
.A(n_395),
.B(n_408),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_398),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_461),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_478),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_481),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_408),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_411),
.B(n_417),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_418),
.B(n_17),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_423),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_418),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_496),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_531),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_502),
.B(n_435),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_498),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_498),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_496),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_498),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_505),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_505),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_519),
.B(n_358),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_519),
.B(n_389),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_553),
.B(n_477),
.Y(n_578)
);

AO21x2_ASAP7_75t_L g579 ( 
.A1(n_550),
.A2(n_480),
.B(n_451),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_504),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_546),
.Y(n_581)
);

AND2x2_ASAP7_75t_SL g582 ( 
.A(n_497),
.B(n_430),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_508),
.Y(n_583)
);

INVx1_ASAP7_75t_SL g584 ( 
.A(n_531),
.Y(n_584)
);

NAND2xp33_ASAP7_75t_SL g585 ( 
.A(n_542),
.B(n_432),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_508),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_508),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_553),
.B(n_390),
.Y(n_588)
);

AND2x6_ASAP7_75t_L g589 ( 
.A(n_542),
.B(n_439),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_511),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_546),
.Y(n_591)
);

NAND2xp33_ASAP7_75t_L g592 ( 
.A(n_499),
.B(n_438),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_511),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_502),
.B(n_509),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_529),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_535),
.B(n_439),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_511),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_512),
.Y(n_598)
);

INVx8_ASAP7_75t_L g599 ( 
.A(n_499),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_512),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_509),
.B(n_452),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_563),
.B(n_452),
.Y(n_602)
);

BUFx10_ASAP7_75t_L g603 ( 
.A(n_532),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_513),
.Y(n_604)
);

BUFx10_ASAP7_75t_L g605 ( 
.A(n_555),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_558),
.B(n_443),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_513),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_547),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_516),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_516),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_547),
.Y(n_611)
);

NOR2xp67_ASAP7_75t_L g612 ( 
.A(n_568),
.B(n_548),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_595),
.B(n_565),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_594),
.B(n_557),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_595),
.B(n_534),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_576),
.B(n_520),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_587),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_584),
.B(n_503),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_576),
.B(n_506),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_577),
.B(n_523),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_587),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_SL g622 ( 
.A(n_582),
.B(n_462),
.Y(n_622)
);

NAND3xp33_ASAP7_75t_L g623 ( 
.A(n_596),
.B(n_536),
.C(n_541),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_606),
.B(n_602),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_606),
.B(n_507),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_602),
.B(n_522),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_577),
.B(n_603),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_569),
.B(n_530),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_569),
.B(n_601),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_604),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_L g631 ( 
.A1(n_582),
.A2(n_501),
.B1(n_552),
.B2(n_514),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_578),
.B(n_518),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_580),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_585),
.B(n_530),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_580),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_603),
.Y(n_636)
);

NOR2x1p5_ASAP7_75t_L g637 ( 
.A(n_567),
.B(n_446),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_597),
.Y(n_638)
);

O2A1O1Ixp33_ASAP7_75t_L g639 ( 
.A1(n_592),
.A2(n_564),
.B(n_561),
.C(n_521),
.Y(n_639)
);

BUFx8_ASAP7_75t_L g640 ( 
.A(n_567),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_588),
.B(n_543),
.Y(n_641)
);

NAND2xp33_ASAP7_75t_SL g642 ( 
.A(n_579),
.B(n_336),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_605),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_607),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_589),
.A2(n_556),
.B1(n_579),
.B2(n_592),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_589),
.B(n_525),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_605),
.B(n_526),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_609),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_605),
.B(n_556),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_589),
.B(n_557),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_599),
.B(n_345),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_581),
.B(n_517),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_591),
.B(n_527),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_589),
.B(n_557),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_579),
.B(n_557),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_608),
.B(n_499),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_L g657 ( 
.A1(n_572),
.A2(n_459),
.B1(n_471),
.B2(n_448),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_611),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_572),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_610),
.B(n_499),
.Y(n_660)
);

OR2x6_ASAP7_75t_L g661 ( 
.A(n_599),
.B(n_533),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_610),
.B(n_547),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_599),
.B(n_351),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_574),
.B(n_539),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_600),
.B(n_549),
.Y(n_665)
);

OA21x2_ASAP7_75t_L g666 ( 
.A1(n_574),
.A2(n_500),
.B(n_538),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_625),
.B(n_354),
.Y(n_667)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_616),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_629),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_628),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_614),
.A2(n_571),
.B(n_570),
.Y(n_671)
);

BUFx12f_ASAP7_75t_L g672 ( 
.A(n_640),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_637),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_645),
.B(n_562),
.Y(n_674)
);

OAI21xp5_ASAP7_75t_L g675 ( 
.A1(n_655),
.A2(n_554),
.B(n_537),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_624),
.B(n_562),
.Y(n_676)
);

INVx4_ASAP7_75t_L g677 ( 
.A(n_661),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_634),
.B(n_356),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_SL g679 ( 
.A(n_636),
.B(n_359),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_632),
.B(n_566),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_655),
.A2(n_642),
.B1(n_623),
.B2(n_631),
.Y(n_681)
);

OAI21xp5_ASAP7_75t_L g682 ( 
.A1(n_660),
.A2(n_656),
.B(n_619),
.Y(n_682)
);

OAI22xp5_ASAP7_75t_L g683 ( 
.A1(n_651),
.A2(n_385),
.B1(n_400),
.B2(n_384),
.Y(n_683)
);

A2O1A1Ixp33_ASAP7_75t_L g684 ( 
.A1(n_639),
.A2(n_335),
.B(n_340),
.C(n_334),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_626),
.B(n_566),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_641),
.B(n_659),
.Y(n_686)
);

BUFx2_ASAP7_75t_L g687 ( 
.A(n_640),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_633),
.B(n_573),
.Y(n_688)
);

AND2x2_ASAP7_75t_SL g689 ( 
.A(n_622),
.B(n_528),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_635),
.B(n_583),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_643),
.Y(n_691)
);

AOI21x1_ASAP7_75t_L g692 ( 
.A1(n_646),
.A2(n_575),
.B(n_586),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_631),
.A2(n_441),
.B1(n_473),
.B2(n_454),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_615),
.A2(n_415),
.B1(n_425),
.B2(n_339),
.Y(n_694)
);

O2A1O1Ixp5_ASAP7_75t_L g695 ( 
.A1(n_613),
.A2(n_593),
.B(n_598),
.C(n_590),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_620),
.B(n_559),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_665),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_644),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_649),
.B(n_475),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_648),
.B(n_590),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_627),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_650),
.A2(n_350),
.B1(n_353),
.B2(n_349),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_662),
.Y(n_703)
);

AOI22xp5_ASAP7_75t_L g704 ( 
.A1(n_663),
.A2(n_342),
.B1(n_344),
.B2(n_338),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_617),
.B(n_575),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_621),
.B(n_638),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_612),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_658),
.Y(n_708)
);

AND2x6_ASAP7_75t_L g709 ( 
.A(n_654),
.B(n_362),
.Y(n_709)
);

O2A1O1Ixp33_ASAP7_75t_L g710 ( 
.A1(n_654),
.A2(n_560),
.B(n_370),
.C(n_375),
.Y(n_710)
);

OAI21xp5_ASAP7_75t_L g711 ( 
.A1(n_666),
.A2(n_379),
.B(n_367),
.Y(n_711)
);

OAI21xp5_ASAP7_75t_L g712 ( 
.A1(n_666),
.A2(n_381),
.B(n_380),
.Y(n_712)
);

OAI21xp5_ASAP7_75t_L g713 ( 
.A1(n_618),
.A2(n_388),
.B(n_387),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_652),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_SL g715 ( 
.A(n_657),
.B(n_476),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_622),
.B(n_483),
.Y(n_716)
);

A2O1A1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_664),
.A2(n_409),
.B(n_414),
.C(n_406),
.Y(n_717)
);

OAI21xp5_ASAP7_75t_L g718 ( 
.A1(n_653),
.A2(n_427),
.B(n_426),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_657),
.B(n_526),
.Y(n_719)
);

OAI21xp5_ASAP7_75t_L g720 ( 
.A1(n_630),
.A2(n_447),
.B(n_433),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_630),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_628),
.B(n_450),
.Y(n_722)
);

A2O1A1Ixp33_ASAP7_75t_L g723 ( 
.A1(n_625),
.A2(n_455),
.B(n_457),
.C(n_453),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_625),
.B(n_485),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_625),
.B(n_488),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_628),
.B(n_458),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_628),
.B(n_463),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_628),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_629),
.Y(n_729)
);

HB1xp67_ASAP7_75t_L g730 ( 
.A(n_616),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_647),
.B(n_346),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_629),
.A2(n_482),
.B(n_474),
.Y(n_732)
);

HB1xp67_ASAP7_75t_L g733 ( 
.A(n_616),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_647),
.B(n_347),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_628),
.B(n_348),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_628),
.B(n_355),
.Y(n_736)
);

NOR3xp33_ASAP7_75t_L g737 ( 
.A(n_625),
.B(n_363),
.C(n_357),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_SL g738 ( 
.A(n_636),
.B(n_365),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_616),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_629),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_629),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_625),
.B(n_368),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_629),
.A2(n_372),
.B(n_369),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_628),
.B(n_373),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_629),
.A2(n_377),
.B(n_374),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_628),
.B(n_382),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_629),
.A2(n_392),
.B(n_391),
.Y(n_747)
);

OAI21xp5_ASAP7_75t_L g748 ( 
.A1(n_655),
.A2(n_396),
.B(n_393),
.Y(n_748)
);

INVxp67_ASAP7_75t_L g749 ( 
.A(n_668),
.Y(n_749)
);

OAI22x1_ASAP7_75t_L g750 ( 
.A1(n_693),
.A2(n_667),
.B1(n_694),
.B2(n_716),
.Y(n_750)
);

A2O1A1Ixp33_ASAP7_75t_L g751 ( 
.A1(n_724),
.A2(n_401),
.B(n_413),
.C(n_399),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_674),
.A2(n_419),
.B(n_416),
.Y(n_752)
);

A2O1A1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_725),
.A2(n_429),
.B(n_431),
.C(n_420),
.Y(n_753)
);

OAI21x1_ASAP7_75t_SL g754 ( 
.A1(n_682),
.A2(n_712),
.B(n_711),
.Y(n_754)
);

NAND3xp33_ASAP7_75t_L g755 ( 
.A(n_742),
.B(n_540),
.C(n_545),
.Y(n_755)
);

OAI21x1_ASAP7_75t_L g756 ( 
.A1(n_692),
.A2(n_515),
.B(n_510),
.Y(n_756)
);

AOI21x1_ASAP7_75t_L g757 ( 
.A1(n_671),
.A2(n_524),
.B(n_515),
.Y(n_757)
);

BUFx8_ASAP7_75t_L g758 ( 
.A(n_687),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_688),
.Y(n_759)
);

OAI21xp5_ASAP7_75t_L g760 ( 
.A1(n_675),
.A2(n_442),
.B(n_440),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_730),
.Y(n_761)
);

OAI21x1_ASAP7_75t_SL g762 ( 
.A1(n_720),
.A2(n_544),
.B(n_528),
.Y(n_762)
);

AO22x1_ASAP7_75t_L g763 ( 
.A1(n_678),
.A2(n_544),
.B1(n_540),
.B2(n_545),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_729),
.B(n_740),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_733),
.Y(n_765)
);

INVx1_ASAP7_75t_SL g766 ( 
.A(n_739),
.Y(n_766)
);

INVxp67_ASAP7_75t_L g767 ( 
.A(n_699),
.Y(n_767)
);

AOI221xp5_ASAP7_75t_L g768 ( 
.A1(n_715),
.A2(n_468),
.B1(n_472),
.B2(n_466),
.C(n_464),
.Y(n_768)
);

AO31x2_ASAP7_75t_L g769 ( 
.A1(n_684),
.A2(n_20),
.A3(n_18),
.B(n_19),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_696),
.Y(n_770)
);

OAI21xp5_ASAP7_75t_L g771 ( 
.A1(n_748),
.A2(n_486),
.B(n_484),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_741),
.B(n_489),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_701),
.Y(n_773)
);

OAI21xp5_ASAP7_75t_L g774 ( 
.A1(n_676),
.A2(n_680),
.B(n_695),
.Y(n_774)
);

AO21x1_ASAP7_75t_L g775 ( 
.A1(n_718),
.A2(n_551),
.B(n_20),
.Y(n_775)
);

OAI21xp5_ASAP7_75t_L g776 ( 
.A1(n_686),
.A2(n_492),
.B(n_491),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_714),
.B(n_493),
.Y(n_777)
);

OA22x2_ASAP7_75t_L g778 ( 
.A1(n_693),
.A2(n_551),
.B1(n_495),
.B2(n_494),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_703),
.B(n_21),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_690),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_672),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_700),
.Y(n_782)
);

NAND2xp33_ASAP7_75t_L g783 ( 
.A(n_670),
.B(n_137),
.Y(n_783)
);

INVxp67_ASAP7_75t_L g784 ( 
.A(n_708),
.Y(n_784)
);

BUFx3_ASAP7_75t_L g785 ( 
.A(n_673),
.Y(n_785)
);

O2A1O1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_723),
.A2(n_24),
.B(n_22),
.C(n_23),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_685),
.A2(n_706),
.B(n_697),
.Y(n_787)
);

AND3x4_ASAP7_75t_L g788 ( 
.A(n_737),
.B(n_25),
.C(n_26),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_722),
.A2(n_147),
.B(n_146),
.Y(n_789)
);

INVx3_ASAP7_75t_SL g790 ( 
.A(n_691),
.Y(n_790)
);

OAI21x1_ASAP7_75t_SL g791 ( 
.A1(n_732),
.A2(n_151),
.B(n_150),
.Y(n_791)
);

AO31x2_ASAP7_75t_L g792 ( 
.A1(n_717),
.A2(n_29),
.A3(n_27),
.B(n_28),
.Y(n_792)
);

AO31x2_ASAP7_75t_L g793 ( 
.A1(n_726),
.A2(n_32),
.A3(n_28),
.B(n_31),
.Y(n_793)
);

O2A1O1Ixp5_ASAP7_75t_L g794 ( 
.A1(n_727),
.A2(n_153),
.B(n_156),
.C(n_152),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_719),
.B(n_31),
.Y(n_795)
);

BUFx4f_ASAP7_75t_L g796 ( 
.A(n_728),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_705),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_728),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_683),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_728),
.B(n_163),
.Y(n_800)
);

NOR2xp67_ASAP7_75t_L g801 ( 
.A(n_707),
.B(n_165),
.Y(n_801)
);

AND2x6_ASAP7_75t_SL g802 ( 
.A(n_735),
.B(n_736),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_SL g803 ( 
.A(n_679),
.B(n_166),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_738),
.B(n_35),
.Y(n_804)
);

AO21x1_ASAP7_75t_L g805 ( 
.A1(n_710),
.A2(n_36),
.B(n_37),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_698),
.B(n_36),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_677),
.B(n_168),
.Y(n_807)
);

NOR2xp67_ASAP7_75t_L g808 ( 
.A(n_677),
.B(n_170),
.Y(n_808)
);

OAI21xp5_ASAP7_75t_L g809 ( 
.A1(n_743),
.A2(n_172),
.B(n_171),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_744),
.B(n_37),
.Y(n_810)
);

A2O1A1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_746),
.A2(n_42),
.B(n_40),
.C(n_41),
.Y(n_811)
);

AO21x2_ASAP7_75t_L g812 ( 
.A1(n_721),
.A2(n_180),
.B(n_177),
.Y(n_812)
);

OAI21x1_ASAP7_75t_L g813 ( 
.A1(n_745),
.A2(n_184),
.B(n_183),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_731),
.A2(n_734),
.B(n_747),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_702),
.A2(n_704),
.B(n_709),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_709),
.A2(n_189),
.B(n_188),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_709),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_689),
.B(n_41),
.Y(n_818)
);

AOI211x1_ASAP7_75t_L g819 ( 
.A1(n_713),
.A2(n_44),
.B(n_42),
.C(n_43),
.Y(n_819)
);

AO31x2_ASAP7_75t_L g820 ( 
.A1(n_684),
.A2(n_45),
.A3(n_43),
.B(n_44),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_691),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_742),
.B(n_45),
.Y(n_822)
);

OAI21x1_ASAP7_75t_SL g823 ( 
.A1(n_682),
.A2(n_193),
.B(n_190),
.Y(n_823)
);

O2A1O1Ixp5_ASAP7_75t_L g824 ( 
.A1(n_748),
.A2(n_196),
.B(n_197),
.C(n_195),
.Y(n_824)
);

NAND2xp33_ASAP7_75t_L g825 ( 
.A(n_674),
.B(n_200),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_670),
.B(n_201),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_742),
.B(n_46),
.Y(n_827)
);

OR2x2_ASAP7_75t_L g828 ( 
.A(n_667),
.B(n_46),
.Y(n_828)
);

OR2x2_ASAP7_75t_L g829 ( 
.A(n_667),
.B(n_48),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_742),
.B(n_48),
.Y(n_830)
);

INVx5_ASAP7_75t_L g831 ( 
.A(n_670),
.Y(n_831)
);

AOI221x1_ASAP7_75t_L g832 ( 
.A1(n_684),
.A2(n_230),
.B1(n_323),
.B2(n_322),
.C(n_320),
.Y(n_832)
);

OAI21xp5_ASAP7_75t_L g833 ( 
.A1(n_711),
.A2(n_207),
.B(n_205),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_691),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_742),
.B(n_49),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_711),
.A2(n_213),
.B(n_212),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_742),
.B(n_49),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_674),
.A2(n_219),
.B(n_216),
.Y(n_838)
);

BUFx2_ASAP7_75t_L g839 ( 
.A(n_668),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_668),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_742),
.B(n_50),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_742),
.B(n_51),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_742),
.B(n_52),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_742),
.B(n_53),
.Y(n_844)
);

NAND3x1_ASAP7_75t_L g845 ( 
.A(n_693),
.B(n_53),
.C(n_54),
.Y(n_845)
);

AO31x2_ASAP7_75t_L g846 ( 
.A1(n_684),
.A2(n_55),
.A3(n_56),
.B(n_57),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_742),
.B(n_57),
.Y(n_847)
);

NAND2xp33_ASAP7_75t_SL g848 ( 
.A(n_681),
.B(n_58),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_742),
.B(n_58),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_L g850 ( 
.A1(n_711),
.A2(n_228),
.B(n_227),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_742),
.B(n_59),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_667),
.B(n_60),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_667),
.B(n_60),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_667),
.B(n_61),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_667),
.B(n_62),
.Y(n_855)
);

OA22x2_ASAP7_75t_L g856 ( 
.A1(n_693),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_691),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_742),
.B(n_64),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_L g859 ( 
.A1(n_711),
.A2(n_238),
.B(n_237),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_839),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_785),
.Y(n_861)
);

BUFx2_ASAP7_75t_R g862 ( 
.A(n_834),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_840),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_764),
.B(n_239),
.Y(n_864)
);

AOI21x1_ASAP7_75t_L g865 ( 
.A1(n_757),
.A2(n_787),
.B(n_814),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_761),
.Y(n_866)
);

INVx1_ASAP7_75t_SL g867 ( 
.A(n_765),
.Y(n_867)
);

OAI21xp5_ASAP7_75t_L g868 ( 
.A1(n_774),
.A2(n_318),
.B(n_260),
.Y(n_868)
);

AO21x2_ASAP7_75t_L g869 ( 
.A1(n_754),
.A2(n_259),
.B(n_315),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_750),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_848),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_797),
.B(n_241),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_831),
.B(n_242),
.Y(n_873)
);

INVx6_ASAP7_75t_L g874 ( 
.A(n_758),
.Y(n_874)
);

AO21x1_ASAP7_75t_L g875 ( 
.A1(n_822),
.A2(n_69),
.B(n_70),
.Y(n_875)
);

AO21x2_ASAP7_75t_L g876 ( 
.A1(n_833),
.A2(n_268),
.B(n_314),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_790),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_777),
.B(n_71),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_767),
.B(n_72),
.Y(n_879)
);

AO21x2_ASAP7_75t_L g880 ( 
.A1(n_836),
.A2(n_270),
.B(n_311),
.Y(n_880)
);

NOR2xp67_ASAP7_75t_L g881 ( 
.A(n_831),
.B(n_244),
.Y(n_881)
);

AO21x2_ASAP7_75t_L g882 ( 
.A1(n_850),
.A2(n_263),
.B(n_310),
.Y(n_882)
);

AOI221xp5_ASAP7_75t_L g883 ( 
.A1(n_854),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.C(n_75),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_759),
.B(n_780),
.Y(n_884)
);

AOI221xp5_ASAP7_75t_L g885 ( 
.A1(n_755),
.A2(n_763),
.B1(n_855),
.B2(n_799),
.C(n_818),
.Y(n_885)
);

NAND2x1p5_ASAP7_75t_L g886 ( 
.A(n_831),
.B(n_246),
.Y(n_886)
);

AO31x2_ASAP7_75t_L g887 ( 
.A1(n_832),
.A2(n_73),
.A3(n_74),
.B(n_75),
.Y(n_887)
);

AO21x2_ASAP7_75t_L g888 ( 
.A1(n_859),
.A2(n_271),
.B(n_309),
.Y(n_888)
);

INVx8_ASAP7_75t_L g889 ( 
.A(n_826),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_766),
.Y(n_890)
);

NAND2x1p5_ASAP7_75t_L g891 ( 
.A(n_796),
.B(n_250),
.Y(n_891)
);

CKINVDCx6p67_ASAP7_75t_R g892 ( 
.A(n_781),
.Y(n_892)
);

CKINVDCx20_ASAP7_75t_R g893 ( 
.A(n_857),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_749),
.Y(n_894)
);

INVx1_ASAP7_75t_SL g895 ( 
.A(n_795),
.Y(n_895)
);

INVx1_ASAP7_75t_SL g896 ( 
.A(n_806),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_758),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_782),
.B(n_254),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_824),
.A2(n_272),
.B(n_308),
.Y(n_899)
);

AO21x2_ASAP7_75t_L g900 ( 
.A1(n_823),
.A2(n_257),
.B(n_306),
.Y(n_900)
);

CKINVDCx6p67_ASAP7_75t_R g901 ( 
.A(n_804),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_773),
.Y(n_902)
);

OAI21xp5_ASAP7_75t_L g903 ( 
.A1(n_815),
.A2(n_316),
.B(n_305),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_852),
.B(n_274),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_853),
.B(n_302),
.Y(n_905)
);

OA21x2_ASAP7_75t_L g906 ( 
.A1(n_789),
.A2(n_301),
.B(n_300),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_796),
.B(n_297),
.Y(n_907)
);

OAI21x1_ASAP7_75t_L g908 ( 
.A1(n_813),
.A2(n_294),
.B(n_293),
.Y(n_908)
);

OA21x2_ASAP7_75t_L g909 ( 
.A1(n_809),
.A2(n_286),
.B(n_285),
.Y(n_909)
);

A2O1A1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_827),
.A2(n_76),
.B(n_77),
.C(n_78),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_830),
.A2(n_281),
.B(n_279),
.Y(n_911)
);

AO21x1_ASAP7_75t_L g912 ( 
.A1(n_835),
.A2(n_76),
.B(n_77),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_784),
.B(n_78),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_770),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_828),
.B(n_79),
.Y(n_915)
);

AO21x2_ASAP7_75t_L g916 ( 
.A1(n_760),
.A2(n_858),
.B(n_837),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_807),
.Y(n_917)
);

OA21x2_ASAP7_75t_L g918 ( 
.A1(n_794),
.A2(n_278),
.B(n_276),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_829),
.B(n_79),
.Y(n_919)
);

OAI21x1_ASAP7_75t_L g920 ( 
.A1(n_817),
.A2(n_80),
.B(n_82),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_779),
.Y(n_921)
);

OAI21x1_ASAP7_75t_SL g922 ( 
.A1(n_791),
.A2(n_84),
.B(n_85),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_802),
.Y(n_923)
);

OR2x6_ASAP7_75t_L g924 ( 
.A(n_798),
.B(n_85),
.Y(n_924)
);

NAND3xp33_ASAP7_75t_L g925 ( 
.A(n_841),
.B(n_86),
.C(n_87),
.Y(n_925)
);

AO21x2_ASAP7_75t_L g926 ( 
.A1(n_842),
.A2(n_851),
.B(n_843),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_810),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_825),
.A2(n_91),
.B(n_92),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_844),
.B(n_847),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_849),
.B(n_93),
.Y(n_930)
);

AO21x2_ASAP7_75t_L g931 ( 
.A1(n_771),
.A2(n_113),
.B(n_95),
.Y(n_931)
);

OAI21x1_ASAP7_75t_L g932 ( 
.A1(n_838),
.A2(n_94),
.B(n_96),
.Y(n_932)
);

AO21x2_ASAP7_75t_L g933 ( 
.A1(n_816),
.A2(n_97),
.B(n_98),
.Y(n_933)
);

NAND2x1p5_ASAP7_75t_L g934 ( 
.A(n_807),
.B(n_99),
.Y(n_934)
);

INVx8_ASAP7_75t_L g935 ( 
.A(n_808),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_772),
.B(n_99),
.Y(n_936)
);

AO31x2_ASAP7_75t_L g937 ( 
.A1(n_805),
.A2(n_100),
.A3(n_101),
.B(n_102),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_778),
.B(n_100),
.Y(n_938)
);

NOR4xp25_ASAP7_75t_L g939 ( 
.A(n_845),
.B(n_104),
.C(n_105),
.D(n_106),
.Y(n_939)
);

AOI22x1_ASAP7_75t_L g940 ( 
.A1(n_752),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_940)
);

INVx1_ASAP7_75t_SL g941 ( 
.A(n_856),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_776),
.B(n_107),
.Y(n_942)
);

BUFx4f_ASAP7_75t_L g943 ( 
.A(n_788),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_801),
.B(n_107),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_811),
.Y(n_945)
);

OAI21x1_ASAP7_75t_SL g946 ( 
.A1(n_786),
.A2(n_110),
.B(n_111),
.Y(n_946)
);

CKINVDCx8_ASAP7_75t_R g947 ( 
.A(n_803),
.Y(n_947)
);

AO21x2_ASAP7_75t_L g948 ( 
.A1(n_751),
.A2(n_112),
.B(n_113),
.Y(n_948)
);

INVx3_ASAP7_75t_SL g949 ( 
.A(n_800),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_769),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_819),
.B(n_753),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_769),
.Y(n_952)
);

INVx4_ASAP7_75t_L g953 ( 
.A(n_812),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_768),
.A2(n_775),
.B1(n_762),
.B2(n_783),
.Y(n_954)
);

NAND3xp33_ASAP7_75t_L g955 ( 
.A(n_820),
.B(n_846),
.C(n_792),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_820),
.Y(n_956)
);

BUFx8_ASAP7_75t_SL g957 ( 
.A(n_793),
.Y(n_957)
);

CKINVDCx6p67_ASAP7_75t_R g958 ( 
.A(n_846),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_846),
.B(n_792),
.Y(n_959)
);

OA21x2_ASAP7_75t_L g960 ( 
.A1(n_792),
.A2(n_774),
.B(n_756),
.Y(n_960)
);

INVx4_ASAP7_75t_L g961 ( 
.A(n_831),
.Y(n_961)
);

BUFx2_ASAP7_75t_SL g962 ( 
.A(n_821),
.Y(n_962)
);

CKINVDCx20_ASAP7_75t_R g963 ( 
.A(n_821),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_767),
.B(n_667),
.Y(n_964)
);

AO21x2_ASAP7_75t_L g965 ( 
.A1(n_754),
.A2(n_774),
.B(n_712),
.Y(n_965)
);

INVx6_ASAP7_75t_L g966 ( 
.A(n_758),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_764),
.B(n_669),
.Y(n_967)
);

AO21x1_ASAP7_75t_L g968 ( 
.A1(n_822),
.A2(n_830),
.B(n_827),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_764),
.B(n_669),
.Y(n_969)
);

OAI21xp33_ASAP7_75t_SL g970 ( 
.A1(n_764),
.A2(n_645),
.B(n_674),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_831),
.B(n_826),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_866),
.Y(n_972)
);

NAND2x1p5_ASAP7_75t_L g973 ( 
.A(n_971),
.B(n_961),
.Y(n_973)
);

AOI22xp33_ASAP7_75t_L g974 ( 
.A1(n_883),
.A2(n_942),
.B1(n_945),
.B2(n_925),
.Y(n_974)
);

BUFx4f_ASAP7_75t_SL g975 ( 
.A(n_893),
.Y(n_975)
);

HB1xp67_ASAP7_75t_L g976 ( 
.A(n_860),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_L g977 ( 
.A1(n_967),
.A2(n_969),
.B1(n_884),
.B2(n_947),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_961),
.Y(n_978)
);

HB1xp67_ASAP7_75t_L g979 ( 
.A(n_867),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_867),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_964),
.B(n_895),
.Y(n_981)
);

HB1xp67_ASAP7_75t_L g982 ( 
.A(n_863),
.Y(n_982)
);

BUFx3_ASAP7_75t_L g983 ( 
.A(n_861),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_890),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_877),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_894),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_963),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_873),
.Y(n_988)
);

AOI21x1_ASAP7_75t_L g989 ( 
.A1(n_865),
.A2(n_959),
.B(n_950),
.Y(n_989)
);

AO31x2_ASAP7_75t_L g990 ( 
.A1(n_952),
.A2(n_956),
.A3(n_959),
.B(n_968),
.Y(n_990)
);

INVx8_ASAP7_75t_L g991 ( 
.A(n_889),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_862),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_921),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_896),
.B(n_919),
.Y(n_994)
);

INVx4_ASAP7_75t_L g995 ( 
.A(n_889),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_941),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_929),
.B(n_927),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_941),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_862),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_914),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_896),
.B(n_878),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_873),
.Y(n_1002)
);

BUFx12f_ASAP7_75t_L g1003 ( 
.A(n_874),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_920),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_929),
.B(n_926),
.Y(n_1005)
);

OR2x6_ASAP7_75t_L g1006 ( 
.A(n_962),
.B(n_917),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_883),
.A2(n_925),
.B1(n_870),
.B2(n_915),
.Y(n_1007)
);

OA21x2_ASAP7_75t_L g1008 ( 
.A1(n_955),
.A2(n_899),
.B(n_903),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_936),
.Y(n_1009)
);

AOI21x1_ASAP7_75t_L g1010 ( 
.A1(n_960),
.A2(n_905),
.B(n_904),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_936),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_902),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_935),
.Y(n_1013)
);

NOR2x1_ASAP7_75t_L g1014 ( 
.A(n_897),
.B(n_872),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_898),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_898),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_901),
.Y(n_1017)
);

AO21x2_ASAP7_75t_L g1018 ( 
.A1(n_955),
.A2(n_899),
.B(n_916),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_872),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_924),
.Y(n_1020)
);

AOI21x1_ASAP7_75t_L g1021 ( 
.A1(n_904),
.A2(n_905),
.B(n_930),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_970),
.A2(n_951),
.B(n_868),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_SL g1023 ( 
.A1(n_943),
.A2(n_924),
.B1(n_954),
.B2(n_933),
.Y(n_1023)
);

AO21x2_ASAP7_75t_L g1024 ( 
.A1(n_916),
.A2(n_965),
.B(n_868),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_970),
.A2(n_951),
.B(n_930),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_944),
.Y(n_1026)
);

CKINVDCx11_ASAP7_75t_R g1027 ( 
.A(n_892),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_879),
.B(n_885),
.Y(n_1028)
);

CKINVDCx16_ASAP7_75t_R g1029 ( 
.A(n_924),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_874),
.Y(n_1030)
);

BUFx2_ASAP7_75t_SL g1031 ( 
.A(n_881),
.Y(n_1031)
);

INVx1_ASAP7_75t_SL g1032 ( 
.A(n_949),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_966),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_864),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_875),
.A2(n_912),
.B1(n_871),
.B2(n_933),
.Y(n_1035)
);

INVx3_ASAP7_75t_L g1036 ( 
.A(n_935),
.Y(n_1036)
);

NAND3xp33_ASAP7_75t_L g1037 ( 
.A(n_911),
.B(n_910),
.C(n_954),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_932),
.Y(n_1038)
);

OAI22xp33_ASAP7_75t_L g1039 ( 
.A1(n_943),
.A2(n_934),
.B1(n_923),
.B2(n_913),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_946),
.Y(n_1040)
);

INVx6_ASAP7_75t_L g1041 ( 
.A(n_966),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_937),
.Y(n_1042)
);

AOI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_940),
.A2(n_931),
.B1(n_911),
.B2(n_948),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_957),
.Y(n_1044)
);

INVx3_ASAP7_75t_L g1045 ( 
.A(n_935),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_958),
.Y(n_1046)
);

AOI22xp33_ASAP7_75t_L g1047 ( 
.A1(n_931),
.A2(n_948),
.B1(n_938),
.B2(n_876),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_965),
.B(n_882),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_887),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_886),
.Y(n_1050)
);

INVx1_ASAP7_75t_SL g1051 ( 
.A(n_907),
.Y(n_1051)
);

OR2x6_ASAP7_75t_L g1052 ( 
.A(n_891),
.B(n_928),
.Y(n_1052)
);

AO21x1_ASAP7_75t_SL g1053 ( 
.A1(n_939),
.A2(n_888),
.B(n_880),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_922),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_939),
.B(n_900),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_908),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_900),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_994),
.B(n_869),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_1001),
.B(n_1028),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_995),
.B(n_953),
.Y(n_1060)
);

INVxp67_ASAP7_75t_L g1061 ( 
.A(n_979),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_995),
.B(n_953),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_981),
.B(n_909),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_1007),
.A2(n_906),
.B1(n_918),
.B2(n_974),
.Y(n_1064)
);

HB1xp67_ASAP7_75t_L g1065 ( 
.A(n_979),
.Y(n_1065)
);

HB1xp67_ASAP7_75t_L g1066 ( 
.A(n_980),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_974),
.A2(n_1037),
.B1(n_1023),
.B2(n_977),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_981),
.B(n_977),
.Y(n_1068)
);

HB1xp67_ASAP7_75t_L g1069 ( 
.A(n_980),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_1000),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_983),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_996),
.B(n_998),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_993),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_1009),
.B(n_1011),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_997),
.B(n_1026),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1005),
.B(n_1015),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_972),
.B(n_986),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_976),
.B(n_1012),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_985),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_1037),
.A2(n_1023),
.B1(n_1035),
.B2(n_1039),
.Y(n_1080)
);

AND2x4_ASAP7_75t_SL g1081 ( 
.A(n_982),
.B(n_978),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_991),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_988),
.B(n_1002),
.Y(n_1083)
);

INVxp67_ASAP7_75t_L g1084 ( 
.A(n_982),
.Y(n_1084)
);

INVx3_ASAP7_75t_SL g1085 ( 
.A(n_1030),
.Y(n_1085)
);

OR2x2_ASAP7_75t_L g1086 ( 
.A(n_987),
.B(n_1029),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_1035),
.A2(n_1039),
.B1(n_1022),
.B2(n_1025),
.Y(n_1087)
);

INVx4_ASAP7_75t_L g1088 ( 
.A(n_978),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_978),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1005),
.B(n_1016),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_1041),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_984),
.B(n_1020),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_1050),
.Y(n_1093)
);

NOR2x1_ASAP7_75t_SL g1094 ( 
.A(n_1052),
.B(n_1031),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_SL g1095 ( 
.A1(n_1032),
.A2(n_1043),
.B(n_1044),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1019),
.B(n_1034),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_1006),
.B(n_1032),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_1050),
.Y(n_1098)
);

INVx2_ASAP7_75t_SL g1099 ( 
.A(n_1003),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1042),
.Y(n_1100)
);

OR2x2_ASAP7_75t_L g1101 ( 
.A(n_987),
.B(n_1006),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_990),
.Y(n_1102)
);

INVxp67_ASAP7_75t_L g1103 ( 
.A(n_1014),
.Y(n_1103)
);

HB1xp67_ASAP7_75t_L g1104 ( 
.A(n_989),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1004),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1049),
.Y(n_1106)
);

AND2x4_ASAP7_75t_SL g1107 ( 
.A(n_1013),
.B(n_1045),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_1051),
.B(n_1044),
.Y(n_1108)
);

OR2x2_ASAP7_75t_L g1109 ( 
.A(n_1017),
.B(n_1025),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1022),
.B(n_1021),
.Y(n_1110)
);

AND2x4_ASAP7_75t_SL g1111 ( 
.A(n_1036),
.B(n_1045),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_973),
.B(n_1036),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1106),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1058),
.B(n_1055),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_1059),
.B(n_1046),
.Y(n_1115)
);

OR2x2_ASAP7_75t_L g1116 ( 
.A(n_1065),
.B(n_1047),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1100),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1068),
.B(n_1040),
.Y(n_1118)
);

AO22x1_ASAP7_75t_L g1119 ( 
.A1(n_1103),
.A2(n_992),
.B1(n_999),
.B2(n_1030),
.Y(n_1119)
);

OR2x2_ASAP7_75t_L g1120 ( 
.A(n_1066),
.B(n_1054),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1075),
.B(n_975),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_1063),
.B(n_1053),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1074),
.B(n_1052),
.Y(n_1123)
);

HB1xp67_ASAP7_75t_L g1124 ( 
.A(n_1104),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1105),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1078),
.B(n_1024),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1096),
.B(n_1008),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_1070),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_1077),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1069),
.B(n_1018),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1072),
.B(n_1010),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_1109),
.B(n_1057),
.Y(n_1132)
);

INVx2_ASAP7_75t_SL g1133 ( 
.A(n_1081),
.Y(n_1133)
);

INVxp67_ASAP7_75t_L g1134 ( 
.A(n_1073),
.Y(n_1134)
);

BUFx2_ASAP7_75t_SL g1135 ( 
.A(n_1079),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_1094),
.B(n_1060),
.Y(n_1136)
);

OR2x2_ASAP7_75t_L g1137 ( 
.A(n_1061),
.B(n_1048),
.Y(n_1137)
);

AOI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_1067),
.A2(n_1108),
.B1(n_1080),
.B2(n_1095),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1097),
.B(n_1038),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_1067),
.A2(n_1080),
.B1(n_1087),
.B2(n_1064),
.Y(n_1140)
);

INVx4_ASAP7_75t_R g1141 ( 
.A(n_1079),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_1108),
.B(n_1057),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1061),
.B(n_1033),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_1062),
.B(n_1056),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_1086),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1142),
.B(n_1076),
.Y(n_1146)
);

NAND3xp33_ASAP7_75t_L g1147 ( 
.A(n_1138),
.B(n_1064),
.C(n_1103),
.Y(n_1147)
);

OR2x2_ASAP7_75t_L g1148 ( 
.A(n_1114),
.B(n_1110),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1114),
.B(n_1102),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1142),
.B(n_1090),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1126),
.B(n_1122),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1113),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1139),
.B(n_1090),
.Y(n_1153)
);

OR2x2_ASAP7_75t_L g1154 ( 
.A(n_1130),
.B(n_1110),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1117),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1125),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_1121),
.B(n_1101),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_1129),
.B(n_1071),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_1136),
.B(n_1083),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1124),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1118),
.B(n_1084),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1120),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1145),
.B(n_1084),
.Y(n_1163)
);

HB1xp67_ASAP7_75t_L g1164 ( 
.A(n_1131),
.Y(n_1164)
);

INVxp67_ASAP7_75t_L g1165 ( 
.A(n_1128),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1155),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1156),
.Y(n_1167)
);

NAND3xp33_ASAP7_75t_L g1168 ( 
.A(n_1147),
.B(n_1140),
.C(n_1132),
.Y(n_1168)
);

OR2x2_ASAP7_75t_L g1169 ( 
.A(n_1148),
.B(n_1116),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1151),
.B(n_1132),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1156),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1146),
.B(n_1134),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1150),
.B(n_1162),
.Y(n_1173)
);

INVxp67_ASAP7_75t_L g1174 ( 
.A(n_1163),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1164),
.B(n_1134),
.Y(n_1175)
);

NAND4xp25_ASAP7_75t_L g1176 ( 
.A(n_1157),
.B(n_1140),
.C(n_1115),
.D(n_1143),
.Y(n_1176)
);

OR2x2_ASAP7_75t_L g1177 ( 
.A(n_1148),
.B(n_1137),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1152),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1149),
.B(n_1127),
.Y(n_1179)
);

INVx3_ASAP7_75t_R g1180 ( 
.A(n_1177),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1166),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1167),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1179),
.B(n_1154),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_SL g1184 ( 
.A(n_1168),
.B(n_1158),
.Y(n_1184)
);

OR2x2_ASAP7_75t_L g1185 ( 
.A(n_1169),
.B(n_1154),
.Y(n_1185)
);

NAND2x1_ASAP7_75t_L g1186 ( 
.A(n_1171),
.B(n_1141),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1179),
.B(n_1160),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1184),
.A2(n_1159),
.B(n_1176),
.Y(n_1188)
);

OAI21xp33_ASAP7_75t_L g1189 ( 
.A1(n_1183),
.A2(n_1172),
.B(n_1173),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_1185),
.A2(n_1174),
.B1(n_1136),
.B2(n_1144),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1181),
.Y(n_1191)
);

NOR3xp33_ASAP7_75t_L g1192 ( 
.A(n_1186),
.B(n_1119),
.C(n_1165),
.Y(n_1192)
);

OAI21xp33_ASAP7_75t_L g1193 ( 
.A1(n_1183),
.A2(n_1175),
.B(n_1153),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1191),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1189),
.B(n_1085),
.Y(n_1195)
);

OAI211xp5_ASAP7_75t_L g1196 ( 
.A1(n_1188),
.A2(n_1161),
.B(n_1187),
.C(n_1178),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1192),
.A2(n_1136),
.B(n_1123),
.Y(n_1197)
);

OAI211xp5_ASAP7_75t_SL g1198 ( 
.A1(n_1196),
.A2(n_1193),
.B(n_1190),
.C(n_1027),
.Y(n_1198)
);

NOR3xp33_ASAP7_75t_L g1199 ( 
.A(n_1195),
.B(n_1099),
.C(n_1091),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1194),
.B(n_1170),
.Y(n_1200)
);

AOI211xp5_ASAP7_75t_L g1201 ( 
.A1(n_1197),
.A2(n_1085),
.B(n_1180),
.C(n_1092),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1194),
.Y(n_1202)
);

NAND4xp75_ASAP7_75t_L g1203 ( 
.A(n_1202),
.B(n_1133),
.C(n_1027),
.D(n_1112),
.Y(n_1203)
);

NOR2x1_ASAP7_75t_L g1204 ( 
.A(n_1198),
.B(n_1135),
.Y(n_1204)
);

NOR3xp33_ASAP7_75t_L g1205 ( 
.A(n_1199),
.B(n_1093),
.C(n_1098),
.Y(n_1205)
);

NOR2x1_ASAP7_75t_L g1206 ( 
.A(n_1203),
.B(n_1071),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1204),
.B(n_1200),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1206),
.Y(n_1208)
);

XNOR2xp5_ASAP7_75t_L g1209 ( 
.A(n_1208),
.B(n_1201),
.Y(n_1209)
);

NAND3xp33_ASAP7_75t_L g1210 ( 
.A(n_1209),
.B(n_1207),
.C(n_1205),
.Y(n_1210)
);

NAND3xp33_ASAP7_75t_L g1211 ( 
.A(n_1210),
.B(n_1088),
.C(n_1089),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1211),
.Y(n_1212)
);

OA22x2_ASAP7_75t_L g1213 ( 
.A1(n_1212),
.A2(n_1081),
.B1(n_1111),
.B2(n_1107),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1213),
.B(n_1182),
.Y(n_1214)
);

OR2x6_ASAP7_75t_L g1215 ( 
.A(n_1214),
.B(n_1082),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1215),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1216),
.A2(n_1089),
.B1(n_1088),
.B2(n_1082),
.Y(n_1217)
);


endmodule