module real_jpeg_12015_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_215;
wire n_221;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_202;
wire n_179;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_1),
.A2(n_33),
.B1(n_57),
.B2(n_59),
.Y(n_88)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g93 ( 
.A(n_3),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_4),
.A2(n_37),
.B(n_38),
.C(n_44),
.Y(n_36)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_4),
.A2(n_40),
.B1(n_44),
.B2(n_45),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_4),
.B(n_116),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_4),
.A2(n_40),
.B1(n_57),
.B2(n_59),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_4),
.A2(n_101),
.B1(n_105),
.B2(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_4),
.B(n_62),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_6),
.A2(n_44),
.B1(n_45),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_6),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_6),
.A2(n_41),
.B1(n_42),
.B2(n_72),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_6),
.A2(n_57),
.B1(n_59),
.B2(n_72),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_72),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_10),
.A2(n_41),
.B1(n_42),
.B2(n_75),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_10),
.A2(n_57),
.B1(n_59),
.B2(n_75),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_75),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_11),
.A2(n_35),
.B1(n_57),
.B2(n_59),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_12),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_12),
.A2(n_57),
.B1(n_59),
.B2(n_85),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_12),
.A2(n_41),
.B1(n_42),
.B2(n_85),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_13),
.A2(n_41),
.B1(n_42),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_13),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_64),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_13),
.A2(n_57),
.B1(n_59),
.B2(n_64),
.Y(n_123)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_15),
.A2(n_41),
.B1(n_42),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_15),
.A2(n_44),
.B1(n_45),
.B2(n_51),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_15),
.A2(n_51),
.B1(n_57),
.B2(n_59),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_51),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_132),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_130),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_117),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_19),
.B(n_117),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_76),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_48),
.C(n_65),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_21),
.A2(n_22),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_23),
.A2(n_24),
.B1(n_36),
.B2(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_25),
.B(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_25),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_25),
.A2(n_81),
.B(n_104),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_25),
.A2(n_30),
.B1(n_188),
.B2(n_190),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_26),
.A2(n_27),
.B1(n_91),
.B2(n_92),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_26),
.B(n_40),
.C(n_92),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_26),
.B(n_195),
.Y(n_194)
);

CKINVDCx6p67_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_30),
.B(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_30),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_32),
.A2(n_82),
.B(n_105),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_34),
.Y(n_102)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_36),
.Y(n_142)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_37),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_37),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_69)
);

OAI21xp33_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B(n_41),
.Y(n_38)
);

HAxp5_ASAP7_75t_SL g159 ( 
.A(n_40),
.B(n_42),
.CON(n_159),
.SN(n_159)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_40),
.B(n_105),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_40),
.B(n_94),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_42),
.B1(n_55),
.B2(n_56),
.Y(n_60)
);

NOR3xp33_ASAP7_75t_L g160 ( 
.A(n_41),
.B(n_56),
.C(n_57),
.Y(n_160)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_48),
.B(n_65),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_52),
.B(n_61),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_50),
.A2(n_53),
.B1(n_62),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_52),
.A2(n_54),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_53),
.A2(n_63),
.B(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_53),
.A2(n_62),
.B1(n_149),
.B2(n_159),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_60),
.Y(n_53)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_54),
.B(n_113),
.Y(n_112)
);

OA22x2_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_SL g157 ( 
.A1(n_55),
.A2(n_59),
.B(n_158),
.C(n_160),
.Y(n_157)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_57),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_57),
.A2(n_59),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_59),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_69),
.B1(n_70),
.B2(n_73),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_67),
.A2(n_74),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_67),
.A2(n_71),
.B1(n_116),
.B2(n_128),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_98),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_86),
.B2(n_97),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_80),
.A2(n_101),
.B(n_191),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_105),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_86),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_89),
.B1(n_95),
.B2(n_96),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_94),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_108),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_123),
.B(n_124),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_89),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_89),
.A2(n_95),
.B1(n_165),
.B2(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_89),
.A2(n_95),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_89),
.A2(n_95),
.B1(n_174),
.B2(n_184),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_94),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_94),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_109),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_95),
.B(n_123),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_110),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_106),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_106),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B(n_103),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_101),
.A2(n_105),
.B1(n_189),
.B2(n_197),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_114),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_121),
.C(n_129),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_129),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_125),
.C(n_127),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_125),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_126),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_140),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_224),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_151),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_136),
.B(n_138),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.C(n_143),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_139),
.B(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_141),
.B(n_143),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.C(n_147),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_147),
.B(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_219),
.B(n_223),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_175),
.B(n_218),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_170),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_154),
.B(n_170),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_167),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_162),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_156),
.B(n_162),
.C(n_167),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_161),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_157),
.B(n_161),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_164),
.B(n_166),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.C(n_173),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_171),
.B(n_215),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_172),
.B(n_173),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_213),
.B(n_217),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_203),
.B(n_212),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_192),
.B(n_202),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_187),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_187),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_182),
.B1(n_185),
.B2(n_186),
.Y(n_179)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_180),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_182),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_185),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_198),
.B(n_201),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_199),
.B(n_200),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_205),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_208),
.C(n_211),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_210),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_216),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_222),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);


endmodule