module real_jpeg_29033_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx11_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_1),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_2),
.A2(n_25),
.B1(n_28),
.B2(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_4),
.A2(n_25),
.B1(n_28),
.B2(n_33),
.Y(n_102)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_5),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_6),
.A2(n_63),
.B1(n_64),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_6),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_71),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_6),
.A2(n_25),
.B1(n_28),
.B2(n_71),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_7),
.A2(n_25),
.B1(n_28),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_8),
.A2(n_74),
.B1(n_75),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_8),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_8),
.A2(n_63),
.B1(n_64),
.B2(n_83),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_83),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_8),
.A2(n_25),
.B1(n_28),
.B2(n_83),
.Y(n_183)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_10),
.A2(n_56),
.B1(n_63),
.B2(n_64),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_10),
.A2(n_25),
.B1(n_28),
.B2(n_56),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_11),
.A2(n_63),
.B1(n_64),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_11),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_11),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_69),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_11),
.A2(n_25),
.B1(n_28),
.B2(n_69),
.Y(n_175)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_13),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_62)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_66),
.Y(n_67)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_13),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_14),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_14),
.B(n_81),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_14),
.B(n_63),
.Y(n_132)
);

AOI21xp33_ASAP7_75t_L g136 ( 
.A1(n_14),
.A2(n_63),
.B(n_132),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_76),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_14),
.A2(n_25),
.B(n_29),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_14),
.B(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_14),
.A2(n_41),
.B1(n_49),
.B2(n_183),
.Y(n_185)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_15),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_120),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_118),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_103),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_20),
.B(n_103),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_84),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_51),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_34),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_24),
.A2(n_36),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_24),
.A2(n_36),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_24),
.A2(n_36),
.B1(n_139),
.B2(n_158),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_24),
.B(n_76),
.Y(n_181)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_24)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_27),
.A2(n_32),
.B(n_76),
.C(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_28),
.B(n_187),
.Y(n_186)
);

AOI32xp33_ASAP7_75t_L g128 ( 
.A1(n_31),
.A2(n_64),
.A3(n_129),
.B1(n_132),
.B2(n_133),
.Y(n_128)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp33_ASAP7_75t_SL g133 ( 
.A(n_32),
.B(n_130),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_54),
.B(n_57),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_36),
.A2(n_140),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_38),
.B(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_45),
.B(n_47),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_41),
.A2(n_44),
.B1(n_45),
.B2(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_41),
.A2(n_169),
.B(n_170),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_41),
.A2(n_49),
.B1(n_175),
.B2(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_42),
.B(n_117),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_42),
.A2(n_48),
.B(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_42),
.A2(n_43),
.B1(n_174),
.B2(n_176),
.Y(n_173)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_43),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_43),
.B(n_127),
.Y(n_170)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_49),
.B(n_76),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_50),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_59),
.C(n_72),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_52),
.A2(n_53),
.B1(n_59),
.B2(n_60),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_55),
.B(n_58),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_60)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_61),
.A2(n_67),
.B1(n_68),
.B2(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_61),
.A2(n_67),
.B1(n_111),
.B2(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_67),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_64),
.B1(n_78),
.B2(n_79),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_78),
.Y(n_100)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_64),
.A2(n_73),
.B1(n_80),
.B2(n_100),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_67),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_72),
.B(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_77),
.B1(n_81),
.B2(n_82),
.Y(n_72)
);

HAxp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_76),
.CON(n_73),
.SN(n_73)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_74),
.A2(n_78),
.B(n_80),
.C(n_81),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_78),
.Y(n_80)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_82),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_98),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_92),
.B2(n_93),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B(n_96),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_101),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_102),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.C(n_109),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_104),
.A2(n_105),
.B1(n_201),
.B2(n_203),
.Y(n_200)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_109),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.C(n_114),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_114),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_198),
.B(n_204),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_151),
.B(n_197),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_141),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_123),
.B(n_141),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_134),
.C(n_137),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_124),
.A2(n_125),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_128),
.Y(n_148)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_134),
.A2(n_135),
.B1(n_137),
.B2(n_138),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_146),
.B2(n_147),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_142),
.B(n_148),
.C(n_149),
.Y(n_199)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_191),
.B(n_196),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_171),
.B(n_190),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_161),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_154),
.B(n_161),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_159),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_155),
.A2(n_156),
.B1(n_159),
.B2(n_178),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_159),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_168),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_166),
.B2(n_167),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_167),
.C(n_168),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_169),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_179),
.B(n_189),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_177),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_173),
.B(n_177),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_184),
.B(n_188),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_181),
.B(n_182),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_192),
.B(n_193),
.Y(n_196)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_199),
.B(n_200),
.Y(n_204)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_201),
.Y(n_203)
);


endmodule