module fake_jpeg_9959_n_199 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_199);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_36),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_26),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_28),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_43),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_46),
.B(n_40),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_38),
.A2(n_30),
.B1(n_19),
.B2(n_20),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_47),
.A2(n_48),
.B1(n_51),
.B2(n_58),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_29),
.B1(n_22),
.B2(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_53),
.B(n_56),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_31),
.B1(n_32),
.B2(n_17),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_29),
.B1(n_22),
.B2(n_17),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_31),
.B1(n_16),
.B2(n_27),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_23),
.B1(n_25),
.B2(n_24),
.Y(n_67)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_61),
.B(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_40),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_81),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_23),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_70),
.Y(n_94)
);

OA21x2_ASAP7_75t_L g100 ( 
.A1(n_67),
.A2(n_27),
.B(n_16),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVxp33_ASAP7_75t_SL g91 ( 
.A(n_68),
.Y(n_91)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_25),
.Y(n_70)
);

INVx5_ASAP7_75t_SL g71 ( 
.A(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_76),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_72),
.Y(n_87)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_74),
.B(n_75),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_46),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_77),
.B(n_56),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_34),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_80),
.B(n_45),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_61),
.B(n_50),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_36),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_73),
.A2(n_54),
.B1(n_36),
.B2(n_52),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_82),
.A2(n_85),
.B1(n_99),
.B2(n_69),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_63),
.B1(n_52),
.B2(n_49),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_100),
.B1(n_71),
.B2(n_64),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_79),
.A2(n_45),
.B1(n_63),
.B2(n_34),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_88),
.B(n_92),
.Y(n_107)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_98),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_57),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_35),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_68),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_57),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_96),
.B(n_97),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_53),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_78),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_81),
.A2(n_67),
.B1(n_72),
.B2(n_77),
.Y(n_99)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_78),
.B(n_33),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_80),
.C(n_64),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_114),
.B1(n_85),
.B2(n_93),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_109),
.C(n_102),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_98),
.A2(n_35),
.B(n_74),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_87),
.B(n_100),
.Y(n_122)
);

A2O1A1O1Ixp25_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_67),
.B(n_80),
.C(n_42),
.D(n_33),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_110),
.B(n_113),
.Y(n_127)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_111),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_112),
.A2(n_99),
.B1(n_82),
.B2(n_100),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_49),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_87),
.A2(n_49),
.B1(n_18),
.B2(n_67),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_115),
.B(n_116),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_93),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_102),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_120),
.B(n_121),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_42),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_122),
.A2(n_107),
.B(n_108),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_123),
.B(n_125),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_120),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_135),
.C(n_35),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_128),
.A2(n_132),
.B1(n_133),
.B2(n_90),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_130),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_121),
.A2(n_118),
.B1(n_109),
.B2(n_112),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_116),
.A2(n_83),
.B1(n_95),
.B2(n_94),
.Y(n_133)
);

NAND2x1_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_95),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_108),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_94),
.C(n_37),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_137),
.B(n_115),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_127),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_139),
.B(n_140),
.Y(n_158)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_145),
.Y(n_159)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_124),
.B(n_117),
.Y(n_145)
);

A2O1A1O1Ixp25_ASAP7_75t_L g164 ( 
.A1(n_146),
.A2(n_147),
.B(n_149),
.C(n_150),
.D(n_129),
.Y(n_164)
);

A2O1A1O1Ixp25_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_111),
.B(n_37),
.C(n_28),
.D(n_35),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

OAI32xp33_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_28),
.A3(n_24),
.B1(n_37),
.B2(n_18),
.Y(n_149)
);

A2O1A1O1Ixp25_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_35),
.B(n_110),
.C(n_4),
.D(n_5),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_152),
.C(n_122),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_136),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_153),
.A2(n_143),
.B1(n_130),
.B2(n_149),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_126),
.C(n_135),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_155),
.C(n_160),
.Y(n_168)
);

BUFx12_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_157),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_133),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_129),
.C(n_124),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_163),
.C(n_4),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_128),
.Y(n_163)
);

AO21x1_ASAP7_75t_L g167 ( 
.A1(n_164),
.A2(n_150),
.B(n_141),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_165),
.B(n_146),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_166),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_167),
.B(n_164),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_162),
.B(n_158),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_172),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_161),
.A2(n_138),
.B1(n_8),
.B2(n_9),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_156),
.B1(n_163),
.B2(n_12),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_160),
.A2(n_138),
.B(n_3),
.Y(n_171)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_171),
.Y(n_177)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_159),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_157),
.A2(n_2),
.B(n_3),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_175),
.C(n_154),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_179),
.A2(n_180),
.B1(n_182),
.B2(n_4),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_168),
.C(n_170),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_174),
.A2(n_156),
.B1(n_157),
.B2(n_11),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_168),
.C(n_175),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_184),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_180),
.A2(n_171),
.B1(n_167),
.B2(n_12),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_185),
.B(n_186),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_176),
.A2(n_9),
.B(n_13),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_15),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_187),
.B(n_188),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_183),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_5),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_192),
.A2(n_187),
.B(n_182),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_195),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_181),
.Y(n_194)
);

AOI322xp5_ASAP7_75t_L g196 ( 
.A1(n_194),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_189),
.C1(n_195),
.C2(n_187),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_196),
.A2(n_6),
.B(n_7),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_197),
.Y(n_199)
);


endmodule